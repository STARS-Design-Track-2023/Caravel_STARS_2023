magic
tech sky130A
magscale 1 2
timestamp 1691545468
<< viali >>
rect 1501 39049 1535 39083
rect 2145 39049 2179 39083
rect 5365 39049 5399 39083
rect 9873 39049 9907 39083
rect 14565 39049 14599 39083
rect 17601 39049 17635 39083
rect 23489 39049 23523 39083
rect 25421 39049 25455 39083
rect 27353 39049 27387 39083
rect 32321 39049 32355 39083
rect 34897 39049 34931 39083
rect 36369 39049 36403 39083
rect 20913 38981 20947 39015
rect 37841 38981 37875 39015
rect 1777 38913 1811 38947
rect 2053 38913 2087 38947
rect 5641 38913 5675 38947
rect 10149 38913 10183 38947
rect 14749 38913 14783 38947
rect 17785 38913 17819 38947
rect 23397 38913 23431 38947
rect 25237 38913 25271 38947
rect 27261 38913 27295 38947
rect 32229 38913 32263 38947
rect 34805 38913 34839 38947
rect 36185 38913 36219 38947
rect 37657 38913 37691 38947
rect 20729 38777 20763 38811
rect 1961 38505 1995 38539
rect 11437 38505 11471 38539
rect 24225 38437 24259 38471
rect 17325 38369 17359 38403
rect 19717 38369 19751 38403
rect 21833 38369 21867 38403
rect 24409 38369 24443 38403
rect 24685 38369 24719 38403
rect 1777 38301 1811 38335
rect 11621 38301 11655 38335
rect 15025 38301 15059 38335
rect 24041 38301 24075 38335
rect 15301 38233 15335 38267
rect 17601 38233 17635 38267
rect 19993 38233 20027 38267
rect 22109 38233 22143 38267
rect 16773 38165 16807 38199
rect 19073 38165 19107 38199
rect 21465 38165 21499 38199
rect 23581 38165 23615 38199
rect 26157 38165 26191 38199
rect 10241 37961 10275 37995
rect 12817 37961 12851 37995
rect 15577 37961 15611 37995
rect 16681 37961 16715 37995
rect 17049 37961 17083 37995
rect 17601 37961 17635 37995
rect 17969 37961 18003 37995
rect 20085 37961 20119 37995
rect 20729 37961 20763 37995
rect 22293 37961 22327 37995
rect 22569 37961 22603 37995
rect 22937 37961 22971 37995
rect 24409 37961 24443 37995
rect 24777 37961 24811 37995
rect 25237 37961 25271 37995
rect 26617 37961 26651 37995
rect 1777 37825 1811 37859
rect 10425 37825 10459 37859
rect 13001 37825 13035 37859
rect 15761 37825 15795 37859
rect 16129 37825 16163 37859
rect 16221 37825 16255 37859
rect 16313 37825 16347 37859
rect 16497 37825 16531 37859
rect 20269 37825 20303 37859
rect 22477 37825 22511 37859
rect 25513 37825 25547 37859
rect 25605 37825 25639 37859
rect 25697 37825 25731 37859
rect 25881 37825 25915 37859
rect 25973 37825 26007 37859
rect 26157 37825 26191 37859
rect 26249 37825 26283 37859
rect 26341 37825 26375 37859
rect 37657 37825 37691 37859
rect 13185 37757 13219 37791
rect 17141 37757 17175 37791
rect 17325 37757 17359 37791
rect 18061 37757 18095 37791
rect 18153 37757 18187 37791
rect 20821 37757 20855 37791
rect 20913 37757 20947 37791
rect 23029 37757 23063 37791
rect 23213 37757 23247 37791
rect 24869 37757 24903 37791
rect 24961 37757 24995 37791
rect 20361 37689 20395 37723
rect 1501 37621 1535 37655
rect 15853 37621 15887 37655
rect 37841 37621 37875 37655
rect 11621 37417 11655 37451
rect 12081 37417 12115 37451
rect 16405 37417 16439 37451
rect 19993 37417 20027 37451
rect 25421 37417 25455 37451
rect 25881 37417 25915 37451
rect 11989 37281 12023 37315
rect 11805 37213 11839 37247
rect 12265 37213 12299 37247
rect 12449 37213 12483 37247
rect 12725 37213 12759 37247
rect 16221 37213 16255 37247
rect 20269 37213 20303 37247
rect 20361 37213 20395 37247
rect 20453 37213 20487 37247
rect 20637 37213 20671 37247
rect 20913 37213 20947 37247
rect 25513 37213 25547 37247
rect 16037 37145 16071 37179
rect 20729 37145 20763 37179
rect 21097 37145 21131 37179
rect 25053 37145 25087 37179
rect 25237 37145 25271 37179
rect 25697 37145 25731 37179
rect 12909 37077 12943 37111
rect 12725 36873 12759 36907
rect 20729 36873 20763 36907
rect 23305 36873 23339 36907
rect 33609 36873 33643 36907
rect 37565 36873 37599 36907
rect 13093 36805 13127 36839
rect 22169 36805 22203 36839
rect 22385 36805 22419 36839
rect 12357 36737 12391 36771
rect 18153 36737 18187 36771
rect 21097 36737 21131 36771
rect 22753 36737 22787 36771
rect 23673 36737 23707 36771
rect 25145 36737 25179 36771
rect 25329 36737 25363 36771
rect 33425 36737 33459 36771
rect 37381 36737 37415 36771
rect 12081 36669 12115 36703
rect 12265 36669 12299 36703
rect 12817 36669 12851 36703
rect 18429 36669 18463 36703
rect 21189 36669 21223 36703
rect 21281 36669 21315 36703
rect 22661 36669 22695 36703
rect 23121 36669 23155 36703
rect 23765 36669 23799 36703
rect 23857 36669 23891 36703
rect 14565 36533 14599 36567
rect 19901 36533 19935 36567
rect 22017 36533 22051 36567
rect 22201 36533 22235 36567
rect 25329 36533 25363 36567
rect 14841 36329 14875 36363
rect 16773 36329 16807 36363
rect 18521 36329 18555 36363
rect 21741 36329 21775 36363
rect 24869 36329 24903 36363
rect 25973 36329 26007 36363
rect 28457 36329 28491 36363
rect 29009 36329 29043 36363
rect 19257 36261 19291 36295
rect 21465 36261 21499 36295
rect 13921 36193 13955 36227
rect 15393 36193 15427 36227
rect 15485 36193 15519 36227
rect 16405 36193 16439 36227
rect 16681 36193 16715 36227
rect 17233 36193 17267 36227
rect 17417 36193 17451 36227
rect 19809 36193 19843 36227
rect 25329 36193 25363 36227
rect 25421 36193 25455 36227
rect 9505 36125 9539 36159
rect 14197 36125 14231 36159
rect 14381 36125 14415 36159
rect 14473 36125 14507 36159
rect 14565 36125 14599 36159
rect 15301 36125 15335 36159
rect 16313 36125 16347 36159
rect 18705 36125 18739 36159
rect 19625 36125 19659 36159
rect 21189 36125 21223 36159
rect 21557 36125 21591 36159
rect 21741 36125 21775 36159
rect 22937 36125 22971 36159
rect 25697 36125 25731 36159
rect 25973 36125 26007 36159
rect 28089 36125 28123 36159
rect 28273 36125 28307 36159
rect 28641 36125 28675 36159
rect 28825 36125 28859 36159
rect 9781 36057 9815 36091
rect 13553 36057 13587 36091
rect 13737 36057 13771 36091
rect 21281 36057 21315 36091
rect 21465 36057 21499 36091
rect 22753 36057 22787 36091
rect 11253 35989 11287 36023
rect 14933 35989 14967 36023
rect 17141 35989 17175 36023
rect 19717 35989 19751 36023
rect 23121 35989 23155 36023
rect 25237 35989 25271 36023
rect 25789 35989 25823 36023
rect 10057 35785 10091 35819
rect 10609 35785 10643 35819
rect 10977 35785 11011 35819
rect 17325 35785 17359 35819
rect 18153 35785 18187 35819
rect 25605 35785 25639 35819
rect 12909 35717 12943 35751
rect 16297 35717 16331 35751
rect 16497 35717 16531 35751
rect 25757 35717 25791 35751
rect 25973 35717 26007 35751
rect 8217 35649 8251 35683
rect 10241 35649 10275 35683
rect 11989 35649 12023 35683
rect 12265 35649 12299 35683
rect 12449 35649 12483 35683
rect 12725 35649 12759 35683
rect 13093 35649 13127 35683
rect 13287 35649 13321 35683
rect 16957 35649 16991 35683
rect 17049 35649 17083 35683
rect 17509 35649 17543 35683
rect 17877 35649 17911 35683
rect 18061 35649 18095 35683
rect 18521 35649 18555 35683
rect 19717 35649 19751 35683
rect 22661 35649 22695 35683
rect 25145 35649 25179 35683
rect 37657 35649 37691 35683
rect 8493 35581 8527 35615
rect 9965 35581 9999 35615
rect 11069 35581 11103 35615
rect 11161 35581 11195 35615
rect 12541 35581 12575 35615
rect 14197 35581 14231 35615
rect 14473 35581 14507 35615
rect 16865 35581 16899 35615
rect 17141 35581 17175 35615
rect 17693 35581 17727 35615
rect 17969 35581 18003 35615
rect 18613 35581 18647 35615
rect 18797 35581 18831 35615
rect 22477 35581 22511 35615
rect 25053 35581 25087 35615
rect 12081 35513 12115 35547
rect 11897 35445 11931 35479
rect 13185 35445 13219 35479
rect 15945 35445 15979 35479
rect 16129 35445 16163 35479
rect 16313 35445 16347 35479
rect 16681 35445 16715 35479
rect 19625 35445 19659 35479
rect 22845 35445 22879 35479
rect 25513 35445 25547 35479
rect 25789 35445 25823 35479
rect 37841 35445 37875 35479
rect 8953 35241 8987 35275
rect 11345 35241 11379 35275
rect 13369 35241 13403 35275
rect 14657 35241 14691 35275
rect 16405 35241 16439 35275
rect 17969 35241 18003 35275
rect 19993 35241 20027 35275
rect 20729 35241 20763 35275
rect 37565 35241 37599 35275
rect 10057 35105 10091 35139
rect 12265 35105 12299 35139
rect 12541 35105 12575 35139
rect 16129 35105 16163 35139
rect 19441 35105 19475 35139
rect 19533 35105 19567 35139
rect 21741 35105 21775 35139
rect 22845 35105 22879 35139
rect 24961 35105 24995 35139
rect 25697 35105 25731 35139
rect 25789 35105 25823 35139
rect 9137 35037 9171 35071
rect 9781 35037 9815 35071
rect 11529 35037 11563 35071
rect 11621 35037 11655 35071
rect 11989 35037 12023 35071
rect 12357 35037 12391 35071
rect 12449 35037 12483 35071
rect 12725 35037 12759 35071
rect 13001 35037 13035 35071
rect 13093 35037 13127 35071
rect 13185 35037 13219 35071
rect 13461 35037 13495 35071
rect 13829 35037 13863 35071
rect 14841 35037 14875 35071
rect 16589 35037 16623 35071
rect 16773 35037 16807 35071
rect 17049 35037 17083 35071
rect 17969 35037 18003 35071
rect 18153 35037 18187 35071
rect 18889 35037 18923 35071
rect 19073 35037 19107 35071
rect 20085 35037 20119 35071
rect 20269 35037 20303 35071
rect 20361 35037 20395 35071
rect 20453 35037 20487 35071
rect 21189 35037 21223 35071
rect 22477 35037 22511 35071
rect 22661 35037 22695 35071
rect 22753 35037 22787 35071
rect 22937 35037 22971 35071
rect 24777 35037 24811 35071
rect 37381 35037 37415 35071
rect 1501 34969 1535 35003
rect 1685 34969 1719 35003
rect 11713 34969 11747 35003
rect 11851 34969 11885 35003
rect 12883 34969 12917 35003
rect 13645 34969 13679 35003
rect 15393 34969 15427 35003
rect 16681 34969 16715 35003
rect 16891 34969 16925 35003
rect 21925 34969 21959 35003
rect 22569 34969 22603 35003
rect 9413 34901 9447 34935
rect 9873 34901 9907 34935
rect 12081 34901 12115 34935
rect 19073 34901 19107 34935
rect 19625 34901 19659 34935
rect 21005 34901 21039 34935
rect 22017 34901 22051 34935
rect 22385 34901 22419 34935
rect 24409 34901 24443 34935
rect 24869 34901 24903 34935
rect 25237 34901 25271 34935
rect 25605 34901 25639 34935
rect 11529 34697 11563 34731
rect 12985 34697 13019 34731
rect 16221 34697 16255 34731
rect 20085 34697 20119 34731
rect 21833 34697 21867 34731
rect 22293 34697 22327 34731
rect 25053 34697 25087 34731
rect 29745 34697 29779 34731
rect 11253 34629 11287 34663
rect 11805 34629 11839 34663
rect 11897 34629 11931 34663
rect 12449 34629 12483 34663
rect 13185 34629 13219 34663
rect 22201 34629 22235 34663
rect 29561 34629 29595 34663
rect 11345 34561 11379 34595
rect 11713 34561 11747 34595
rect 12035 34561 12069 34595
rect 12173 34561 12207 34595
rect 12725 34561 12759 34595
rect 16129 34561 16163 34595
rect 19901 34561 19935 34595
rect 20085 34561 20119 34595
rect 29377 34561 29411 34595
rect 29653 34561 29687 34595
rect 29837 34561 29871 34595
rect 29929 34561 29963 34595
rect 30113 34561 30147 34595
rect 22477 34493 22511 34527
rect 23305 34493 23339 34527
rect 23581 34493 23615 34527
rect 29193 34493 29227 34527
rect 12817 34357 12851 34391
rect 13001 34357 13035 34391
rect 30113 34357 30147 34391
rect 14749 34153 14783 34187
rect 22477 34153 22511 34187
rect 23765 34153 23799 34187
rect 26893 34153 26927 34187
rect 27537 34153 27571 34187
rect 6929 34085 6963 34119
rect 26525 34085 26559 34119
rect 20729 34017 20763 34051
rect 26341 34017 26375 34051
rect 30205 34017 30239 34051
rect 30573 34017 30607 34051
rect 5181 33949 5215 33983
rect 14105 33949 14139 33983
rect 14289 33949 14323 33983
rect 14381 33949 14415 33983
rect 14473 33949 14507 33983
rect 15393 33949 15427 33983
rect 15577 33949 15611 33983
rect 17785 33949 17819 33983
rect 17969 33949 18003 33983
rect 23121 33949 23155 33983
rect 23949 33949 23983 33983
rect 25237 33949 25271 33983
rect 25421 33949 25455 33983
rect 26617 33949 26651 33983
rect 27353 33949 27387 33983
rect 27537 33949 27571 33983
rect 29837 33949 29871 33983
rect 30021 33949 30055 33983
rect 30297 33949 30331 33983
rect 30389 33949 30423 33983
rect 5457 33881 5491 33915
rect 15761 33881 15795 33915
rect 21005 33881 21039 33915
rect 22937 33881 22971 33915
rect 26709 33881 26743 33915
rect 17785 33813 17819 33847
rect 23305 33813 23339 33847
rect 25053 33813 25087 33847
rect 26341 33813 26375 33847
rect 26909 33813 26943 33847
rect 27077 33813 27111 33847
rect 27169 33813 27203 33847
rect 30573 33813 30607 33847
rect 5917 33609 5951 33643
rect 6929 33609 6963 33643
rect 8769 33609 8803 33643
rect 12909 33609 12943 33643
rect 14289 33609 14323 33643
rect 15025 33609 15059 33643
rect 15669 33609 15703 33643
rect 26341 33609 26375 33643
rect 28273 33609 28307 33643
rect 29101 33609 29135 33643
rect 31769 33609 31803 33643
rect 4353 33541 4387 33575
rect 7297 33541 7331 33575
rect 9505 33541 9539 33575
rect 12015 33541 12049 33575
rect 12541 33541 12575 33575
rect 15485 33541 15519 33575
rect 27721 33541 27755 33575
rect 6101 33473 6135 33507
rect 6745 33473 6779 33507
rect 11713 33473 11747 33507
rect 11805 33473 11839 33507
rect 11897 33473 11931 33507
rect 12725 33473 12759 33507
rect 13001 33473 13035 33507
rect 14841 33473 14875 33507
rect 15025 33473 15059 33507
rect 15117 33473 15151 33507
rect 15301 33473 15335 33507
rect 15393 33473 15427 33507
rect 15577 33473 15611 33507
rect 15945 33473 15979 33507
rect 16037 33473 16071 33507
rect 16129 33473 16163 33507
rect 16313 33473 16347 33507
rect 18153 33473 18187 33507
rect 18521 33473 18555 33507
rect 18705 33473 18739 33507
rect 18797 33473 18831 33507
rect 19809 33473 19843 33507
rect 19993 33473 20027 33507
rect 25881 33473 25915 33507
rect 26065 33473 26099 33507
rect 26157 33473 26191 33507
rect 26525 33473 26559 33507
rect 26985 33473 27019 33507
rect 27261 33473 27295 33507
rect 27353 33473 27387 33507
rect 27537 33473 27571 33507
rect 28181 33473 28215 33507
rect 28457 33473 28491 33507
rect 28641 33473 28675 33507
rect 28733 33473 28767 33507
rect 28917 33473 28951 33507
rect 29285 33473 29319 33507
rect 29837 33473 29871 33507
rect 29929 33473 29963 33507
rect 31125 33473 31159 33507
rect 31401 33473 31435 33507
rect 31493 33473 31527 33507
rect 31644 33473 31678 33507
rect 32597 33473 32631 33507
rect 4077 33405 4111 33439
rect 7021 33405 7055 33439
rect 9229 33405 9263 33439
rect 12173 33405 12207 33439
rect 17417 33405 17451 33439
rect 18061 33405 18095 33439
rect 18889 33405 18923 33439
rect 26709 33405 26743 33439
rect 27905 33405 27939 33439
rect 28549 33405 28583 33439
rect 30205 33405 30239 33439
rect 30297 33405 30331 33439
rect 32505 33405 32539 33439
rect 27445 33337 27479 33371
rect 28089 33337 28123 33371
rect 28917 33337 28951 33371
rect 31125 33337 31159 33371
rect 31953 33337 31987 33371
rect 5825 33269 5859 33303
rect 10977 33269 11011 33303
rect 11529 33269 11563 33303
rect 15209 33269 15243 33303
rect 18521 33269 18555 33303
rect 19809 33269 19843 33303
rect 25697 33269 25731 33303
rect 27997 33269 28031 33303
rect 29653 33269 29687 33303
rect 32873 33269 32907 33303
rect 4445 33065 4479 33099
rect 5825 33065 5859 33099
rect 6837 33065 6871 33099
rect 9781 33065 9815 33099
rect 11805 33065 11839 33099
rect 14381 33065 14415 33099
rect 16037 33065 16071 33099
rect 18337 33065 18371 33099
rect 20085 33065 20119 33099
rect 26525 33065 26559 33099
rect 26709 33065 26743 33099
rect 29561 33065 29595 33099
rect 30021 33065 30055 33099
rect 33149 33065 33183 33099
rect 8401 32997 8435 33031
rect 12265 32997 12299 33031
rect 13737 32997 13771 33031
rect 17233 32997 17267 33031
rect 19441 32997 19475 33031
rect 28089 32997 28123 33031
rect 31401 32997 31435 33031
rect 32597 32997 32631 33031
rect 34161 32997 34195 33031
rect 5273 32929 5307 32963
rect 6469 32929 6503 32963
rect 7481 32929 7515 32963
rect 7757 32929 7791 32963
rect 10977 32929 11011 32963
rect 16589 32929 16623 32963
rect 18245 32929 18279 32963
rect 18889 32929 18923 32963
rect 20637 32929 20671 32963
rect 27629 32929 27663 32963
rect 29285 32929 29319 32963
rect 29837 32929 29871 32963
rect 34713 32929 34747 32963
rect 34897 32929 34931 32963
rect 4629 32861 4663 32895
rect 5089 32861 5123 32895
rect 6285 32861 6319 32895
rect 8033 32861 8067 32895
rect 8677 32861 8711 32895
rect 9965 32861 9999 32895
rect 10793 32861 10827 32895
rect 10885 32861 10919 32895
rect 11713 32861 11747 32895
rect 11897 32861 11931 32895
rect 12449 32861 12483 32895
rect 13185 32861 13219 32895
rect 13461 32861 13495 32895
rect 13553 32861 13587 32895
rect 14105 32861 14139 32895
rect 14841 32861 14875 32895
rect 14933 32861 14967 32895
rect 15117 32861 15151 32895
rect 15485 32861 15519 32895
rect 15761 32861 15795 32895
rect 16405 32861 16439 32895
rect 17509 32861 17543 32895
rect 17601 32861 17635 32895
rect 17785 32861 17819 32895
rect 17877 32861 17911 32895
rect 17970 32861 18004 32895
rect 18797 32861 18831 32895
rect 19625 32861 19659 32895
rect 19717 32861 19751 32895
rect 19901 32861 19935 32895
rect 19993 32861 20027 32895
rect 21741 32861 21775 32895
rect 22063 32861 22097 32895
rect 22193 32871 22227 32905
rect 25513 32861 25547 32895
rect 25697 32861 25731 32895
rect 26157 32861 26191 32895
rect 26617 32861 26651 32895
rect 26801 32861 26835 32895
rect 27721 32861 27755 32895
rect 29193 32861 29227 32895
rect 29377 32861 29411 32895
rect 30113 32861 30147 32895
rect 31401 32861 31435 32895
rect 31585 32861 31619 32895
rect 31953 32861 31987 32895
rect 32137 32861 32171 32895
rect 32229 32861 32263 32895
rect 33057 32861 33091 32895
rect 33333 32861 33367 32895
rect 33425 32861 33459 32895
rect 34161 32861 34195 32895
rect 34437 32861 34471 32895
rect 34989 32861 35023 32895
rect 35081 32861 35115 32895
rect 35173 32861 35207 32895
rect 37933 32861 37967 32895
rect 5181 32793 5215 32827
rect 7941 32793 7975 32827
rect 12633 32793 12667 32827
rect 13369 32793 13403 32827
rect 14749 32793 14783 32827
rect 15025 32793 15059 32827
rect 15577 32793 15611 32827
rect 17233 32793 17267 32827
rect 18705 32793 18739 32827
rect 21833 32793 21867 32827
rect 21925 32793 21959 32827
rect 26341 32793 26375 32827
rect 30389 32793 30423 32827
rect 30573 32793 30607 32827
rect 32413 32793 32447 32827
rect 4721 32725 4755 32759
rect 6193 32725 6227 32759
rect 7205 32725 7239 32759
rect 7297 32725 7331 32759
rect 8493 32725 8527 32759
rect 10425 32725 10459 32759
rect 14565 32725 14599 32759
rect 15945 32725 15979 32759
rect 16497 32725 16531 32759
rect 17417 32725 17451 32759
rect 20453 32725 20487 32759
rect 20545 32725 20579 32759
rect 21557 32725 21591 32759
rect 22293 32725 22327 32759
rect 25513 32725 25547 32759
rect 30205 32725 30239 32759
rect 31861 32725 31895 32759
rect 33609 32725 33643 32759
rect 34345 32725 34379 32759
rect 37749 32725 37783 32759
rect 18889 32521 18923 32555
rect 20453 32521 20487 32555
rect 21833 32521 21867 32555
rect 29853 32521 29887 32555
rect 30021 32521 30055 32555
rect 7941 32453 7975 32487
rect 12541 32453 12575 32487
rect 21557 32453 21591 32487
rect 22661 32453 22695 32487
rect 23673 32453 23707 32487
rect 24133 32453 24167 32487
rect 24225 32453 24259 32487
rect 25053 32453 25087 32487
rect 29653 32453 29687 32487
rect 32321 32453 32355 32487
rect 12265 32385 12299 32419
rect 12449 32385 12483 32419
rect 12685 32385 12719 32419
rect 18153 32385 18187 32419
rect 18705 32385 18739 32419
rect 18797 32385 18831 32419
rect 19809 32385 19843 32419
rect 20361 32385 20395 32419
rect 20545 32385 20579 32419
rect 20637 32385 20671 32419
rect 21189 32385 21223 32419
rect 21373 32385 21407 32419
rect 21465 32385 21499 32419
rect 21649 32385 21683 32419
rect 22385 32385 22419 32419
rect 22569 32385 22603 32419
rect 22845 32385 22879 32419
rect 22937 32385 22971 32419
rect 23121 32385 23155 32419
rect 23213 32385 23247 32419
rect 23581 32385 23615 32419
rect 23765 32385 23799 32419
rect 24041 32385 24075 32419
rect 24409 32385 24443 32419
rect 24501 32385 24535 32419
rect 24685 32385 24719 32419
rect 24961 32385 24995 32419
rect 32137 32385 32171 32419
rect 33241 32385 33275 32419
rect 33701 32385 33735 32419
rect 33977 32385 34011 32419
rect 34437 32385 34471 32419
rect 7665 32317 7699 32351
rect 9413 32317 9447 32351
rect 19165 32317 19199 32351
rect 19625 32317 19659 32351
rect 19901 32317 19935 32351
rect 19993 32317 20027 32351
rect 20085 32317 20119 32351
rect 22293 32317 22327 32351
rect 33425 32317 33459 32351
rect 34621 32317 34655 32351
rect 34713 32317 34747 32351
rect 35081 32317 35115 32351
rect 20729 32249 20763 32283
rect 21373 32249 21407 32283
rect 21925 32249 21959 32283
rect 32873 32249 32907 32283
rect 12817 32181 12851 32215
rect 18245 32181 18279 32215
rect 22477 32181 22511 32215
rect 23857 32181 23891 32215
rect 24869 32181 24903 32215
rect 29837 32181 29871 32215
rect 32505 32181 32539 32215
rect 3801 31977 3835 32011
rect 21465 31977 21499 32011
rect 24409 31977 24443 32011
rect 25789 31977 25823 32011
rect 32321 31977 32355 32011
rect 27813 31909 27847 31943
rect 5549 31841 5583 31875
rect 6377 31841 6411 31875
rect 14933 31841 14967 31875
rect 17969 31841 18003 31875
rect 18153 31841 18187 31875
rect 18337 31841 18371 31875
rect 22753 31841 22787 31875
rect 24593 31841 24627 31875
rect 27721 31841 27755 31875
rect 31585 31841 31619 31875
rect 34161 31841 34195 31875
rect 34345 31841 34379 31875
rect 11621 31773 11655 31807
rect 11805 31773 11839 31807
rect 11989 31773 12023 31807
rect 12081 31773 12115 31807
rect 14841 31773 14875 31807
rect 15853 31773 15887 31807
rect 15945 31773 15979 31807
rect 16129 31773 16163 31807
rect 16221 31773 16255 31807
rect 18245 31773 18279 31807
rect 18429 31773 18463 31807
rect 21649 31773 21683 31807
rect 21925 31773 21959 31807
rect 22661 31773 22695 31807
rect 23121 31773 23155 31807
rect 23397 31773 23431 31807
rect 23581 31773 23615 31807
rect 23673 31773 23707 31807
rect 23857 31773 23891 31807
rect 24041 31773 24075 31807
rect 24225 31773 24259 31807
rect 24685 31773 24719 31807
rect 25697 31773 25731 31807
rect 25881 31773 25915 31807
rect 27905 31773 27939 31807
rect 27997 31773 28031 31807
rect 31493 31773 31527 31807
rect 32137 31773 32171 31807
rect 32413 31773 32447 31807
rect 33793 31773 33827 31807
rect 34069 31773 34103 31807
rect 5273 31705 5307 31739
rect 6653 31705 6687 31739
rect 21833 31705 21867 31739
rect 8125 31637 8159 31671
rect 16405 31637 16439 31671
rect 22201 31637 22235 31671
rect 22569 31637 22603 31671
rect 23219 31637 23253 31671
rect 23305 31637 23339 31671
rect 25053 31637 25087 31671
rect 4905 31433 4939 31467
rect 6561 31433 6595 31467
rect 8769 31433 8803 31467
rect 13645 31433 13679 31467
rect 15025 31433 15059 31467
rect 15761 31433 15795 31467
rect 19073 31433 19107 31467
rect 19993 31433 20027 31467
rect 21557 31433 21591 31467
rect 24317 31433 24351 31467
rect 27721 31433 27755 31467
rect 29101 31433 29135 31467
rect 31493 31433 31527 31467
rect 32873 31433 32907 31467
rect 33977 31433 34011 31467
rect 35909 31433 35943 31467
rect 7021 31365 7055 31399
rect 7481 31365 7515 31399
rect 11253 31365 11287 31399
rect 11805 31365 11839 31399
rect 11897 31365 11931 31399
rect 14105 31365 14139 31399
rect 15393 31365 15427 31399
rect 18153 31365 18187 31399
rect 19165 31365 19199 31399
rect 21373 31365 21407 31399
rect 27353 31365 27387 31399
rect 34069 31365 34103 31399
rect 36461 31365 36495 31399
rect 3341 31297 3375 31331
rect 6377 31297 6411 31331
rect 7113 31297 7147 31331
rect 9321 31297 9355 31331
rect 11161 31297 11195 31331
rect 11713 31297 11747 31331
rect 12035 31297 12069 31331
rect 12357 31297 12391 31331
rect 12541 31297 12575 31331
rect 12633 31297 12667 31331
rect 12725 31297 12759 31331
rect 13461 31297 13495 31331
rect 13645 31297 13679 31331
rect 13737 31297 13771 31331
rect 13921 31297 13955 31331
rect 14013 31297 14047 31331
rect 14197 31297 14231 31331
rect 14336 31297 14370 31331
rect 14565 31297 14599 31331
rect 14674 31297 14708 31331
rect 14933 31297 14967 31331
rect 15212 31297 15246 31331
rect 15485 31297 15519 31331
rect 15577 31297 15611 31331
rect 15853 31297 15887 31331
rect 16129 31297 16163 31331
rect 16221 31297 16255 31331
rect 16405 31297 16439 31331
rect 16773 31297 16807 31331
rect 17049 31297 17083 31331
rect 17969 31297 18003 31331
rect 18245 31297 18279 31331
rect 18337 31297 18371 31331
rect 18705 31297 18739 31331
rect 18889 31297 18923 31331
rect 19349 31297 19383 31331
rect 19533 31297 19567 31331
rect 19809 31297 19843 31331
rect 21649 31297 21683 31331
rect 21833 31297 21867 31331
rect 22164 31297 22198 31331
rect 22385 31297 22419 31331
rect 24133 31297 24167 31331
rect 24317 31297 24351 31331
rect 24961 31297 24995 31331
rect 25145 31297 25179 31331
rect 25237 31297 25271 31331
rect 25329 31297 25363 31331
rect 27169 31297 27203 31331
rect 27997 31297 28031 31331
rect 28365 31297 28399 31331
rect 28549 31297 28583 31331
rect 28917 31297 28951 31331
rect 29837 31297 29871 31331
rect 29929 31297 29963 31331
rect 30113 31297 30147 31331
rect 30389 31297 30423 31331
rect 30665 31297 30699 31331
rect 30849 31297 30883 31331
rect 31125 31297 31159 31331
rect 32137 31297 32171 31331
rect 32321 31297 32355 31331
rect 32689 31297 32723 31331
rect 33241 31297 33275 31331
rect 33333 31297 33367 31331
rect 33425 31297 33459 31331
rect 33609 31297 33643 31331
rect 33701 31297 33735 31331
rect 34161 31297 34195 31331
rect 34529 31297 34563 31331
rect 34621 31297 34655 31331
rect 34805 31297 34839 31331
rect 34897 31297 34931 31331
rect 35449 31297 35483 31331
rect 35541 31297 35575 31331
rect 35633 31297 35667 31331
rect 35817 31297 35851 31331
rect 36093 31297 36127 31331
rect 36277 31297 36311 31331
rect 36369 31297 36403 31331
rect 36553 31297 36587 31331
rect 3065 31229 3099 31263
rect 3433 31229 3467 31263
rect 4353 31229 4387 31263
rect 5641 31229 5675 31263
rect 7205 31229 7239 31263
rect 9597 31229 9631 31263
rect 12173 31229 12207 31263
rect 15136 31229 15170 31263
rect 16313 31229 16347 31263
rect 16957 31229 16991 31263
rect 18613 31229 18647 31263
rect 19625 31229 19659 31263
rect 26985 31229 27019 31263
rect 27721 31229 27755 31263
rect 28641 31229 28675 31263
rect 28733 31229 28767 31263
rect 31033 31229 31067 31263
rect 32413 31229 32447 31263
rect 32505 31229 32539 31263
rect 35173 31229 35207 31263
rect 6653 31161 6687 31195
rect 12909 31161 12943 31195
rect 13921 31161 13955 31195
rect 14841 31161 14875 31195
rect 15577 31161 15611 31195
rect 16865 31161 16899 31195
rect 18521 31161 18555 31195
rect 21373 31161 21407 31195
rect 21925 31161 21959 31195
rect 27905 31161 27939 31195
rect 34345 31161 34379 31195
rect 1593 31093 1627 31127
rect 4077 31093 4111 31127
rect 5089 31093 5123 31127
rect 11069 31093 11103 31127
rect 11529 31093 11563 31127
rect 14381 31093 14415 31127
rect 15945 31093 15979 31127
rect 17233 31093 17267 31127
rect 25605 31093 25639 31127
rect 30205 31093 30239 31127
rect 32965 31093 32999 31127
rect 3157 30889 3191 30923
rect 4445 30889 4479 30923
rect 5089 30889 5123 30923
rect 9781 30889 9815 30923
rect 11621 30889 11655 30923
rect 14197 30889 14231 30923
rect 18613 30889 18647 30923
rect 19441 30889 19475 30923
rect 25605 30889 25639 30923
rect 34713 30889 34747 30923
rect 36185 30889 36219 30923
rect 4537 30821 4571 30855
rect 11437 30821 11471 30855
rect 16865 30821 16899 30855
rect 32505 30821 32539 30855
rect 6837 30753 6871 30787
rect 7021 30753 7055 30787
rect 8769 30753 8803 30787
rect 9413 30753 9447 30787
rect 9505 30753 9539 30787
rect 10793 30753 10827 30787
rect 10885 30753 10919 30787
rect 15945 30753 15979 30787
rect 16129 30753 16163 30787
rect 16313 30753 16347 30787
rect 29285 30753 29319 30787
rect 36001 30753 36035 30787
rect 3341 30685 3375 30719
rect 3525 30685 3559 30719
rect 3617 30685 3651 30719
rect 3801 30685 3835 30719
rect 3949 30685 3983 30719
rect 4307 30685 4341 30719
rect 4905 30685 4939 30719
rect 9965 30685 9999 30719
rect 10701 30685 10735 30719
rect 12449 30685 12483 30719
rect 12633 30685 12667 30719
rect 12725 30685 12759 30719
rect 12817 30685 12851 30719
rect 13266 30685 13300 30719
rect 14289 30685 14323 30719
rect 16221 30685 16255 30719
rect 16405 30685 16439 30719
rect 16589 30685 16623 30719
rect 16773 30685 16807 30719
rect 18521 30685 18555 30719
rect 18705 30685 18739 30719
rect 18889 30685 18923 30719
rect 18981 30685 19015 30719
rect 19257 30685 19291 30719
rect 19441 30685 19475 30719
rect 25237 30685 25271 30719
rect 26249 30685 26283 30719
rect 26801 30685 26835 30719
rect 27721 30685 27755 30719
rect 27905 30685 27939 30719
rect 27997 30685 28031 30719
rect 28549 30685 28583 30719
rect 28917 30685 28951 30719
rect 32229 30685 32263 30719
rect 32505 30685 32539 30719
rect 35081 30685 35115 30719
rect 35909 30685 35943 30719
rect 4077 30617 4111 30651
rect 4169 30617 4203 30651
rect 4721 30617 4755 30651
rect 6561 30617 6595 30651
rect 7297 30617 7331 30651
rect 11589 30617 11623 30651
rect 11805 30617 11839 30651
rect 13093 30617 13127 30651
rect 25421 30617 25455 30651
rect 27629 30617 27663 30651
rect 34897 30617 34931 30651
rect 8953 30549 8987 30583
rect 9321 30549 9355 30583
rect 10333 30549 10367 30583
rect 13001 30549 13035 30583
rect 13461 30549 13495 30583
rect 32321 30549 32355 30583
rect 3525 30345 3559 30379
rect 4445 30345 4479 30379
rect 8125 30345 8159 30379
rect 20545 30345 20579 30379
rect 27997 30345 28031 30379
rect 4905 30277 4939 30311
rect 4997 30277 5031 30311
rect 19993 30277 20027 30311
rect 20209 30277 20243 30311
rect 20729 30277 20763 30311
rect 23305 30277 23339 30311
rect 27629 30277 27663 30311
rect 29653 30277 29687 30311
rect 3433 30209 3467 30243
rect 3525 30209 3559 30243
rect 4537 30209 4571 30243
rect 4629 30209 4663 30243
rect 4777 30209 4811 30243
rect 5133 30209 5167 30243
rect 8309 30209 8343 30243
rect 13277 30209 13311 30243
rect 13369 30209 13403 30243
rect 13461 30209 13495 30243
rect 13645 30209 13679 30243
rect 20453 30209 20487 30243
rect 23121 30209 23155 30243
rect 23765 30209 23799 30243
rect 24225 30209 24259 30243
rect 24409 30209 24443 30243
rect 27813 30209 27847 30243
rect 28089 30209 28123 30243
rect 28273 30209 28307 30243
rect 29561 30209 29595 30243
rect 29745 30209 29779 30243
rect 30021 30209 30055 30243
rect 30297 30209 30331 30243
rect 30481 30209 30515 30243
rect 30757 30209 30791 30243
rect 32781 30209 32815 30243
rect 3249 30141 3283 30175
rect 3617 30141 3651 30175
rect 23673 30141 23707 30175
rect 23857 30141 23891 30175
rect 23949 30141 23983 30175
rect 24133 30141 24167 30175
rect 28181 30141 28215 30175
rect 30573 30141 30607 30175
rect 30941 30141 30975 30175
rect 32689 30141 32723 30175
rect 33609 30141 33643 30175
rect 5273 30073 5307 30107
rect 23489 30073 23523 30107
rect 24501 30073 24535 30107
rect 4261 30005 4295 30039
rect 13001 30005 13035 30039
rect 20177 30005 20211 30039
rect 20361 30005 20395 30039
rect 20729 30005 20763 30039
rect 29837 30005 29871 30039
rect 14565 29801 14599 29835
rect 20269 29801 20303 29835
rect 20637 29801 20671 29835
rect 23765 29801 23799 29835
rect 31033 29801 31067 29835
rect 34161 29801 34195 29835
rect 3157 29733 3191 29767
rect 5089 29733 5123 29767
rect 10149 29733 10183 29767
rect 15577 29733 15611 29767
rect 16589 29733 16623 29767
rect 21465 29733 21499 29767
rect 28365 29733 28399 29767
rect 34253 29733 34287 29767
rect 36737 29733 36771 29767
rect 1409 29665 1443 29699
rect 7021 29665 7055 29699
rect 10701 29665 10735 29699
rect 12817 29665 12851 29699
rect 14381 29665 14415 29699
rect 15209 29665 15243 29699
rect 15485 29665 15519 29699
rect 16037 29665 16071 29699
rect 16129 29665 16163 29699
rect 20085 29665 20119 29699
rect 20545 29665 20579 29699
rect 28831 29665 28865 29699
rect 36461 29665 36495 29699
rect 4997 29597 5031 29631
rect 5181 29597 5215 29631
rect 9873 29597 9907 29631
rect 11437 29597 11471 29631
rect 13093 29597 13127 29631
rect 14289 29597 14323 29631
rect 15117 29597 15151 29631
rect 16405 29597 16439 29631
rect 16589 29597 16623 29631
rect 20361 29597 20395 29631
rect 20453 29597 20487 29631
rect 21097 29597 21131 29631
rect 21189 29597 21223 29631
rect 21465 29597 21499 29631
rect 23489 29597 23523 29631
rect 23765 29597 23799 29631
rect 24409 29597 24443 29631
rect 24586 29597 24620 29631
rect 26433 29597 26467 29631
rect 26617 29597 26651 29631
rect 26709 29597 26743 29631
rect 26893 29597 26927 29631
rect 26985 29597 27019 29631
rect 28112 29597 28146 29631
rect 28273 29597 28307 29631
rect 28549 29597 28583 29631
rect 28733 29597 28767 29631
rect 28917 29597 28951 29631
rect 29101 29597 29135 29631
rect 30849 29597 30883 29631
rect 31033 29597 31067 29631
rect 31769 29597 31803 29631
rect 32045 29597 32079 29631
rect 33793 29597 33827 29631
rect 33977 29597 34011 29631
rect 34069 29597 34103 29631
rect 34345 29597 34379 29631
rect 36369 29597 36403 29631
rect 37197 29597 37231 29631
rect 37473 29597 37507 29631
rect 1685 29529 1719 29563
rect 7297 29529 7331 29563
rect 10517 29529 10551 29563
rect 11621 29529 11655 29563
rect 13001 29529 13035 29563
rect 15945 29529 15979 29563
rect 21281 29529 21315 29563
rect 8769 29461 8803 29495
rect 9689 29461 9723 29495
rect 10609 29461 10643 29495
rect 11805 29461 11839 29495
rect 13461 29461 13495 29495
rect 20085 29461 20119 29495
rect 20821 29461 20855 29495
rect 21005 29461 21039 29495
rect 23581 29461 23615 29495
rect 24501 29461 24535 29495
rect 26249 29461 26283 29495
rect 28273 29461 28307 29495
rect 32045 29461 32079 29495
rect 36829 29461 36863 29495
rect 1869 29257 1903 29291
rect 3617 29257 3651 29291
rect 5181 29257 5215 29291
rect 8033 29257 8067 29291
rect 10885 29257 10919 29291
rect 11529 29257 11563 29291
rect 13093 29257 13127 29291
rect 21189 29257 21223 29291
rect 24409 29257 24443 29291
rect 26341 29257 26375 29291
rect 27813 29257 27847 29291
rect 28273 29257 28307 29291
rect 28365 29257 28399 29291
rect 34713 29257 34747 29291
rect 7481 29189 7515 29223
rect 9413 29189 9447 29223
rect 11897 29189 11931 29223
rect 12725 29189 12759 29223
rect 18521 29189 18555 29223
rect 21281 29189 21315 29223
rect 21481 29189 21515 29223
rect 31401 29189 31435 29223
rect 33425 29189 33459 29223
rect 34989 29189 35023 29223
rect 35357 29189 35391 29223
rect 36277 29189 36311 29223
rect 2053 29121 2087 29155
rect 3709 29121 3743 29155
rect 4537 29121 4571 29155
rect 4837 29121 4871 29155
rect 4997 29121 5031 29155
rect 5089 29121 5123 29155
rect 5273 29121 5307 29155
rect 7573 29121 7607 29155
rect 8217 29121 8251 29155
rect 11161 29121 11195 29155
rect 11345 29121 11379 29155
rect 11713 29121 11747 29155
rect 11805 29121 11839 29155
rect 12035 29121 12069 29155
rect 12449 29121 12483 29155
rect 12633 29121 12667 29155
rect 12817 29121 12851 29155
rect 13277 29121 13311 29155
rect 15853 29121 15887 29155
rect 15945 29121 15979 29155
rect 16129 29121 16163 29155
rect 17877 29121 17911 29155
rect 17969 29121 18003 29155
rect 18153 29121 18187 29155
rect 20821 29121 20855 29155
rect 22017 29121 22051 29155
rect 23949 29121 23983 29155
rect 24777 29121 24811 29155
rect 25973 29121 26007 29155
rect 27169 29121 27203 29155
rect 27445 29121 27479 29155
rect 27537 29121 27571 29155
rect 27721 29121 27755 29155
rect 28457 29121 28491 29155
rect 28549 29121 28583 29155
rect 28733 29121 28767 29155
rect 29009 29121 29043 29155
rect 29469 29121 29503 29155
rect 30021 29121 30055 29155
rect 30113 29121 30147 29155
rect 31309 29121 31343 29155
rect 31493 29121 31527 29155
rect 32137 29121 32171 29155
rect 32873 29121 32907 29155
rect 33149 29121 33183 29155
rect 33333 29121 33367 29155
rect 33517 29121 33551 29155
rect 33977 29121 34011 29155
rect 34161 29121 34195 29155
rect 34262 29121 34296 29155
rect 34529 29121 34563 29155
rect 35173 29121 35207 29155
rect 35633 29121 35667 29155
rect 36185 29121 36219 29155
rect 36369 29121 36403 29155
rect 3893 29053 3927 29087
rect 4353 29053 4387 29087
rect 7297 29053 7331 29087
rect 9137 29053 9171 29087
rect 11253 29053 11287 29087
rect 12173 29053 12207 29087
rect 13461 29053 13495 29087
rect 20913 29053 20947 29087
rect 21925 29053 21959 29087
rect 24041 29053 24075 29087
rect 24685 29053 24719 29087
rect 26065 29053 26099 29087
rect 27353 29053 27387 29087
rect 27997 29053 28031 29087
rect 28089 29053 28123 29087
rect 29377 29053 29411 29087
rect 29929 29053 29963 29087
rect 30205 29053 30239 29087
rect 32229 29053 32263 29087
rect 33241 29053 33275 29087
rect 34345 29053 34379 29087
rect 36093 29053 36127 29087
rect 3249 28985 3283 29019
rect 4997 28985 5031 29019
rect 7941 28985 7975 29019
rect 13001 28985 13035 29019
rect 16129 28985 16163 29019
rect 21649 28985 21683 29019
rect 24317 28985 24351 29019
rect 26985 28985 27019 29019
rect 28733 28985 28767 29019
rect 29653 28985 29687 29019
rect 32505 28985 32539 29019
rect 4721 28917 4755 28951
rect 18521 28917 18555 28951
rect 21465 28917 21499 28951
rect 22293 28917 22327 28951
rect 29745 28917 29779 28951
rect 32137 28917 32171 28951
rect 35725 28917 35759 28951
rect 3617 28713 3651 28747
rect 4629 28713 4663 28747
rect 5273 28713 5307 28747
rect 6837 28713 6871 28747
rect 15945 28713 15979 28747
rect 17601 28713 17635 28747
rect 22201 28713 22235 28747
rect 27169 28713 27203 28747
rect 27905 28713 27939 28747
rect 29561 28713 29595 28747
rect 29929 28713 29963 28747
rect 31677 28713 31711 28747
rect 32781 28713 32815 28747
rect 33057 28713 33091 28747
rect 35633 28713 35667 28747
rect 36461 28713 36495 28747
rect 6745 28645 6779 28679
rect 17693 28645 17727 28679
rect 22661 28645 22695 28679
rect 31493 28645 31527 28679
rect 32597 28645 32631 28679
rect 35449 28645 35483 28679
rect 35725 28645 35759 28679
rect 36093 28645 36127 28679
rect 1869 28577 1903 28611
rect 3801 28577 3835 28611
rect 5733 28577 5767 28611
rect 5917 28577 5951 28611
rect 7113 28577 7147 28611
rect 7297 28577 7331 28611
rect 15577 28577 15611 28611
rect 17325 28577 17359 28611
rect 17785 28577 17819 28611
rect 22201 28577 22235 28611
rect 22845 28577 22879 28611
rect 27261 28577 27295 28611
rect 30021 28577 30055 28611
rect 30849 28577 30883 28611
rect 32873 28577 32907 28611
rect 36737 28577 36771 28611
rect 4445 28509 4479 28543
rect 4537 28509 4571 28543
rect 4813 28509 4847 28543
rect 5273 28509 5307 28543
rect 5365 28509 5399 28543
rect 5549 28509 5583 28543
rect 5641 28509 5675 28543
rect 6009 28509 6043 28543
rect 6101 28509 6135 28543
rect 7021 28509 7055 28543
rect 7205 28509 7239 28543
rect 13001 28509 13035 28543
rect 15301 28509 15335 28543
rect 15485 28509 15519 28543
rect 15761 28509 15795 28543
rect 16037 28509 16071 28543
rect 16129 28509 16163 28543
rect 16313 28509 16347 28543
rect 16497 28509 16531 28543
rect 17233 28509 17267 28543
rect 18061 28509 18095 28543
rect 18521 28509 18555 28543
rect 18889 28509 18923 28543
rect 19441 28509 19475 28543
rect 19533 28509 19567 28543
rect 19717 28509 19751 28543
rect 19809 28509 19843 28543
rect 19901 28509 19935 28543
rect 20085 28509 20119 28543
rect 22114 28509 22148 28543
rect 22569 28509 22603 28543
rect 24685 28509 24719 28543
rect 24777 28509 24811 28543
rect 24869 28509 24903 28543
rect 25053 28509 25087 28543
rect 26709 28509 26743 28543
rect 26801 28509 26835 28543
rect 26985 28509 27019 28543
rect 27537 28509 27571 28543
rect 27721 28509 27755 28543
rect 27997 28509 28031 28543
rect 29745 28509 29779 28543
rect 30757 28509 30791 28543
rect 30941 28509 30975 28543
rect 31125 28509 31159 28543
rect 31309 28509 31343 28543
rect 31585 28509 31619 28543
rect 31769 28509 31803 28543
rect 32965 28509 32999 28543
rect 33057 28509 33091 28543
rect 33241 28509 33275 28543
rect 35909 28509 35943 28543
rect 36001 28509 36035 28543
rect 36185 28509 36219 28543
rect 36369 28509 36403 28543
rect 36645 28509 36679 28543
rect 36829 28509 36863 28543
rect 36921 28509 36955 28543
rect 2145 28441 2179 28475
rect 6586 28441 6620 28475
rect 12817 28441 12851 28475
rect 35173 28441 35207 28475
rect 4997 28373 5031 28407
rect 5733 28373 5767 28407
rect 6377 28373 6411 28407
rect 6469 28373 6503 28407
rect 13185 28373 13219 28407
rect 15393 28373 15427 28407
rect 16405 28373 16439 28407
rect 19257 28373 19291 28407
rect 19993 28373 20027 28407
rect 22477 28373 22511 28407
rect 22845 28373 22879 28407
rect 24409 28373 24443 28407
rect 27629 28373 27663 28407
rect 6469 28169 6503 28203
rect 15761 28169 15795 28203
rect 17601 28169 17635 28203
rect 19901 28169 19935 28203
rect 24133 28169 24167 28203
rect 26065 28169 26099 28203
rect 32781 28169 32815 28203
rect 35909 28169 35943 28203
rect 4721 28101 4755 28135
rect 22385 28101 22419 28135
rect 23121 28101 23155 28135
rect 27077 28101 27111 28135
rect 22615 28067 22649 28101
rect 1961 28033 1995 28067
rect 6377 28033 6411 28067
rect 6561 28033 6595 28067
rect 11713 28033 11747 28067
rect 13553 28033 13587 28067
rect 13645 28033 13679 28067
rect 13737 28033 13771 28067
rect 13921 28033 13955 28067
rect 15669 28033 15703 28067
rect 15853 28033 15887 28067
rect 17233 28033 17267 28067
rect 17877 28033 17911 28067
rect 18153 28033 18187 28067
rect 19073 28033 19107 28067
rect 19257 28033 19291 28067
rect 19533 28033 19567 28067
rect 19809 28033 19843 28067
rect 22848 28033 22882 28067
rect 22937 28033 22971 28067
rect 23949 28033 23983 28067
rect 24225 28033 24259 28067
rect 24777 28033 24811 28067
rect 24869 28033 24903 28067
rect 25605 28033 25639 28067
rect 25881 28033 25915 28067
rect 26985 28033 27019 28067
rect 27169 28033 27203 28067
rect 32137 28033 32171 28067
rect 32321 28033 32355 28067
rect 32413 28033 32447 28067
rect 32505 28033 32539 28067
rect 32873 28033 32907 28067
rect 33057 28033 33091 28067
rect 33517 28033 33551 28067
rect 33885 28033 33919 28067
rect 34437 28033 34471 28067
rect 34529 28033 34563 28067
rect 35081 28033 35115 28067
rect 36001 28033 36035 28067
rect 36185 28033 36219 28067
rect 8033 27965 8067 27999
rect 8309 27965 8343 27999
rect 11805 27965 11839 27999
rect 17141 27965 17175 27999
rect 18337 27965 18371 27999
rect 19441 27965 19475 27999
rect 35449 27965 35483 27999
rect 12081 27897 12115 27931
rect 17969 27897 18003 27931
rect 19349 27897 19383 27931
rect 19717 27897 19751 27931
rect 24869 27897 24903 27931
rect 25697 27897 25731 27931
rect 25789 27897 25823 27931
rect 33885 27897 33919 27931
rect 35725 27897 35759 27931
rect 36277 27897 36311 27931
rect 1777 27829 1811 27863
rect 4997 27829 5031 27863
rect 9781 27829 9815 27863
rect 13277 27829 13311 27863
rect 22569 27829 22603 27863
rect 22753 27829 22787 27863
rect 23121 27829 23155 27863
rect 23949 27829 23983 27863
rect 32873 27829 32907 27863
rect 4905 27625 4939 27659
rect 6377 27625 6411 27659
rect 7205 27625 7239 27659
rect 8309 27625 8343 27659
rect 19441 27625 19475 27659
rect 19993 27625 20027 27659
rect 20361 27625 20395 27659
rect 36645 27625 36679 27659
rect 6745 27557 6779 27591
rect 13277 27557 13311 27591
rect 15761 27557 15795 27591
rect 27353 27557 27387 27591
rect 29285 27557 29319 27591
rect 6653 27489 6687 27523
rect 9413 27489 9447 27523
rect 9505 27489 9539 27523
rect 11897 27489 11931 27523
rect 13461 27489 13495 27523
rect 30113 27489 30147 27523
rect 37289 27489 37323 27523
rect 4905 27421 4939 27455
rect 5089 27421 5123 27455
rect 6561 27421 6595 27455
rect 6837 27421 6871 27455
rect 7113 27421 7147 27455
rect 8493 27421 8527 27455
rect 11069 27421 11103 27455
rect 12357 27421 12391 27455
rect 12449 27421 12483 27455
rect 12541 27421 12575 27455
rect 12705 27421 12739 27455
rect 13001 27421 13035 27455
rect 13553 27421 13587 27455
rect 14381 27421 14415 27455
rect 14841 27421 14875 27455
rect 15945 27421 15979 27455
rect 16129 27421 16163 27455
rect 19441 27421 19475 27455
rect 19625 27421 19659 27455
rect 19809 27421 19843 27455
rect 19901 27421 19935 27455
rect 19993 27421 20027 27455
rect 20177 27421 20211 27455
rect 20269 27421 20303 27455
rect 20453 27421 20487 27455
rect 22385 27421 22419 27455
rect 22569 27421 22603 27455
rect 22753 27421 22787 27455
rect 27261 27421 27295 27455
rect 27445 27421 27479 27455
rect 29193 27421 29227 27455
rect 29377 27421 29411 27455
rect 29561 27421 29595 27455
rect 29837 27421 29871 27455
rect 30297 27421 30331 27455
rect 30573 27421 30607 27455
rect 34713 27421 34747 27455
rect 34897 27421 34931 27455
rect 36461 27421 36495 27455
rect 36645 27421 36679 27455
rect 37381 27421 37415 27455
rect 11713 27353 11747 27387
rect 12817 27353 12851 27387
rect 13829 27353 13863 27387
rect 13921 27353 13955 27387
rect 22937 27353 22971 27387
rect 23029 27353 23063 27387
rect 29653 27353 29687 27387
rect 30021 27353 30055 27387
rect 30481 27353 30515 27387
rect 36737 27353 36771 27387
rect 4721 27285 4755 27319
rect 7573 27285 7607 27319
rect 8953 27285 8987 27319
rect 9321 27285 9355 27319
rect 11253 27285 11287 27319
rect 11345 27285 11379 27319
rect 11805 27285 11839 27319
rect 12173 27285 12207 27319
rect 13185 27285 13219 27319
rect 14197 27285 14231 27319
rect 34805 27285 34839 27319
rect 5641 27081 5675 27115
rect 7113 27081 7147 27115
rect 8217 27081 8251 27115
rect 8861 27081 8895 27115
rect 14289 27081 14323 27115
rect 15301 27081 15335 27115
rect 17509 27081 17543 27115
rect 19257 27081 19291 27115
rect 25237 27081 25271 27115
rect 26157 27081 26191 27115
rect 27629 27081 27663 27115
rect 28365 27081 28399 27115
rect 30849 27081 30883 27115
rect 31769 27081 31803 27115
rect 36277 27081 36311 27115
rect 9229 27013 9263 27047
rect 13001 27013 13035 27047
rect 25697 27013 25731 27047
rect 30113 27013 30147 27047
rect 32965 27013 32999 27047
rect 33977 27013 34011 27047
rect 35081 27013 35115 27047
rect 36093 27013 36127 27047
rect 36737 27013 36771 27047
rect 2145 26945 2179 26979
rect 3985 26945 4019 26979
rect 4721 26945 4755 26979
rect 4997 26945 5031 26979
rect 5365 26945 5399 26979
rect 5825 26945 5859 26979
rect 5917 26945 5951 26979
rect 6101 26945 6135 26979
rect 6193 26945 6227 26979
rect 6564 26945 6598 26979
rect 7021 26945 7055 26979
rect 7665 26945 7699 26979
rect 7757 26945 7791 26979
rect 7849 26945 7883 26979
rect 8033 26945 8067 26979
rect 8677 26945 8711 26979
rect 15393 26945 15427 26979
rect 16405 26945 16439 26979
rect 17233 26945 17267 26979
rect 17417 26945 17451 26979
rect 17509 26945 17543 26979
rect 17693 26945 17727 26979
rect 19441 26945 19475 26979
rect 19533 26945 19567 26979
rect 19625 26945 19659 26979
rect 19809 26945 19843 26979
rect 20729 26945 20763 26979
rect 22937 26945 22971 26979
rect 23121 26945 23155 26979
rect 24501 26945 24535 26979
rect 24593 26945 24627 26979
rect 24869 26945 24903 26979
rect 25053 26945 25087 26979
rect 25237 26945 25271 26979
rect 25513 26945 25547 26979
rect 25789 26945 25823 26979
rect 25973 26945 26007 26979
rect 26617 26945 26651 26979
rect 26801 26945 26835 26979
rect 27077 26945 27111 26979
rect 27169 26945 27203 26979
rect 27353 26945 27387 26979
rect 27445 26945 27479 26979
rect 27721 26945 27755 26979
rect 27905 26945 27939 26979
rect 27997 26945 28031 26979
rect 28089 26945 28123 26979
rect 29377 26945 29411 26979
rect 29561 26945 29595 26979
rect 29745 26945 29779 26979
rect 29929 26945 29963 26979
rect 30205 26945 30239 26979
rect 30389 26945 30423 26979
rect 30481 26945 30515 26979
rect 30573 26945 30607 26979
rect 31125 26945 31159 26979
rect 31309 26945 31343 26979
rect 31585 26945 31619 26979
rect 33149 26945 33183 26979
rect 33241 26945 33275 26979
rect 33701 26945 33735 26979
rect 33794 26945 33828 26979
rect 34069 26945 34103 26979
rect 34207 26945 34241 26979
rect 34713 26945 34747 26979
rect 34989 26945 35023 26979
rect 35265 26945 35299 26979
rect 35449 26945 35483 26979
rect 35633 26945 35667 26979
rect 35817 26945 35851 26979
rect 36369 26945 36403 26979
rect 36553 26945 36587 26979
rect 36921 26945 36955 26979
rect 2421 26877 2455 26911
rect 3893 26877 3927 26911
rect 6653 26877 6687 26911
rect 7389 26877 7423 26911
rect 8953 26877 8987 26911
rect 15485 26877 15519 26911
rect 20821 26877 20855 26911
rect 25329 26877 25363 26911
rect 26709 26877 26743 26911
rect 29653 26877 29687 26911
rect 32965 26877 32999 26911
rect 35541 26877 35575 26911
rect 10701 26809 10735 26843
rect 23029 26809 23063 26843
rect 34345 26809 34379 26843
rect 34897 26809 34931 26843
rect 36093 26809 36127 26843
rect 4077 26741 4111 26775
rect 4813 26741 4847 26775
rect 5273 26741 5307 26775
rect 6377 26741 6411 26775
rect 6837 26741 6871 26775
rect 7297 26741 7331 26775
rect 14933 26741 14967 26775
rect 16313 26741 16347 26775
rect 17325 26741 17359 26775
rect 21005 26741 21039 26775
rect 34529 26741 34563 26775
rect 35725 26741 35759 26775
rect 5549 26537 5583 26571
rect 7205 26537 7239 26571
rect 7573 26537 7607 26571
rect 9045 26537 9079 26571
rect 13277 26537 13311 26571
rect 15853 26537 15887 26571
rect 22569 26537 22603 26571
rect 24961 26537 24995 26571
rect 27813 26537 27847 26571
rect 29009 26537 29043 26571
rect 29745 26537 29779 26571
rect 29929 26537 29963 26571
rect 32965 26537 32999 26571
rect 35173 26537 35207 26571
rect 36829 26537 36863 26571
rect 37013 26537 37047 26571
rect 3617 26469 3651 26503
rect 16313 26469 16347 26503
rect 17049 26469 17083 26503
rect 18245 26469 18279 26503
rect 21741 26469 21775 26503
rect 28089 26469 28123 26503
rect 34437 26469 34471 26503
rect 1409 26401 1443 26435
rect 1685 26401 1719 26435
rect 3157 26401 3191 26435
rect 4353 26401 4387 26435
rect 9505 26401 9539 26435
rect 9689 26401 9723 26435
rect 11805 26401 11839 26435
rect 14381 26401 14415 26435
rect 15945 26401 15979 26435
rect 17233 26401 17267 26435
rect 18337 26401 18371 26435
rect 21281 26401 21315 26435
rect 22201 26401 22235 26435
rect 25513 26401 25547 26435
rect 26709 26401 26743 26435
rect 28641 26401 28675 26435
rect 32505 26401 32539 26435
rect 32597 26401 32631 26435
rect 34805 26401 34839 26435
rect 36185 26401 36219 26435
rect 36553 26401 36587 26435
rect 3433 26333 3467 26367
rect 3617 26333 3651 26367
rect 4905 26333 4939 26367
rect 7113 26333 7147 26367
rect 11529 26333 11563 26367
rect 14105 26333 14139 26367
rect 16129 26333 16163 26367
rect 16957 26333 16991 26367
rect 17141 26333 17175 26367
rect 17601 26333 17635 26367
rect 17693 26333 17727 26367
rect 18153 26333 18187 26367
rect 18429 26333 18463 26367
rect 21373 26333 21407 26367
rect 22371 26333 22405 26367
rect 23581 26333 23615 26367
rect 23765 26333 23799 26367
rect 23857 26333 23891 26367
rect 23949 26333 23983 26367
rect 25329 26333 25363 26367
rect 25973 26333 26007 26367
rect 26157 26333 26191 26367
rect 26617 26333 26651 26367
rect 26801 26333 26835 26367
rect 27077 26333 27111 26367
rect 27261 26333 27295 26367
rect 27353 26333 27387 26367
rect 27445 26333 27479 26367
rect 27629 26333 27663 26367
rect 28917 26335 28951 26369
rect 29101 26333 29135 26367
rect 32229 26333 32263 26367
rect 32413 26333 32447 26367
rect 32781 26333 32815 26367
rect 34529 26333 34563 26367
rect 34897 26333 34931 26367
rect 36645 26333 36679 26367
rect 36921 26333 36955 26367
rect 37105 26333 37139 26367
rect 3801 26265 3835 26299
rect 4537 26265 4571 26299
rect 7021 26265 7055 26299
rect 15853 26265 15887 26299
rect 24225 26265 24259 26299
rect 25421 26265 25455 26299
rect 26065 26265 26099 26299
rect 28457 26265 28491 26299
rect 29561 26265 29595 26299
rect 29761 26265 29795 26299
rect 9413 26197 9447 26231
rect 17877 26197 17911 26231
rect 17969 26197 18003 26231
rect 28549 26197 28583 26231
rect 3433 25993 3467 26027
rect 5641 25993 5675 26027
rect 6653 25993 6687 26027
rect 14105 25993 14139 26027
rect 30113 25993 30147 26027
rect 31861 25993 31895 26027
rect 33057 25993 33091 26027
rect 1777 25925 1811 25959
rect 7113 25925 7147 25959
rect 13369 25925 13403 25959
rect 14841 25925 14875 25959
rect 16037 25925 16071 25959
rect 16129 25925 16163 25959
rect 29653 25925 29687 25959
rect 30757 25925 30791 25959
rect 30941 25925 30975 25959
rect 31125 25925 31159 25959
rect 32873 25925 32907 25959
rect 1409 25857 1443 25891
rect 3341 25857 3375 25891
rect 3525 25857 3559 25891
rect 4629 25857 4663 25891
rect 5641 25857 5675 25891
rect 6377 25857 6411 25891
rect 13180 25857 13214 25891
rect 13277 25857 13311 25891
rect 13553 25857 13587 25891
rect 13829 25857 13863 25891
rect 14381 25857 14415 25891
rect 14744 25857 14778 25891
rect 14933 25857 14967 25891
rect 15117 25857 15151 25891
rect 15940 25857 15974 25891
rect 16313 25857 16347 25891
rect 19257 25857 19291 25891
rect 19349 25857 19383 25891
rect 19462 25863 19496 25897
rect 19625 25857 19659 25891
rect 19901 25857 19935 25891
rect 19993 25857 20027 25891
rect 20177 25857 20211 25891
rect 23489 25857 23523 25891
rect 23673 25857 23707 25891
rect 23765 25857 23799 25891
rect 23857 25857 23891 25891
rect 26157 25857 26191 25891
rect 26341 25857 26375 25891
rect 29745 25857 29779 25891
rect 31217 25857 31251 25891
rect 31401 25857 31435 25891
rect 31493 25857 31527 25891
rect 31585 25857 31619 25891
rect 32137 25857 32171 25891
rect 32321 25857 32355 25891
rect 32689 25857 32723 25891
rect 32965 25857 32999 25891
rect 33149 25857 33183 25891
rect 6561 25789 6595 25823
rect 13737 25789 13771 25823
rect 29469 25789 29503 25823
rect 32413 25789 32447 25823
rect 32505 25789 32539 25823
rect 7113 25721 7147 25755
rect 19717 25721 19751 25755
rect 13001 25653 13035 25687
rect 14565 25653 14599 25687
rect 15761 25653 15795 25687
rect 18981 25653 19015 25687
rect 19901 25653 19935 25687
rect 24133 25653 24167 25687
rect 26249 25653 26283 25687
rect 17693 25449 17727 25483
rect 17969 25449 18003 25483
rect 18705 25449 18739 25483
rect 20821 25449 20855 25483
rect 25421 25449 25455 25483
rect 30573 25449 30607 25483
rect 31033 25449 31067 25483
rect 33057 25449 33091 25483
rect 36737 25449 36771 25483
rect 37197 25449 37231 25483
rect 7941 25381 7975 25415
rect 9689 25381 9723 25415
rect 15669 25381 15703 25415
rect 17233 25381 17267 25415
rect 18337 25381 18371 25415
rect 1409 25313 1443 25347
rect 3157 25313 3191 25347
rect 4353 25313 4387 25347
rect 7297 25313 7331 25347
rect 8677 25313 8711 25347
rect 9045 25313 9079 25347
rect 10425 25313 10459 25347
rect 10609 25313 10643 25347
rect 12909 25313 12943 25347
rect 17601 25313 17635 25347
rect 19993 25313 20027 25347
rect 20269 25313 20303 25347
rect 20453 25313 20487 25347
rect 36921 25313 36955 25347
rect 4629 25245 4663 25279
rect 6653 25245 6687 25279
rect 6837 25245 6871 25279
rect 7113 25245 7147 25279
rect 7757 25245 7791 25279
rect 8401 25245 8435 25279
rect 11161 25245 11195 25279
rect 13093 25245 13127 25279
rect 13645 25245 13679 25279
rect 14289 25245 14323 25279
rect 14381 25245 14415 25279
rect 14657 25245 14691 25279
rect 15848 25245 15882 25279
rect 16037 25245 16071 25279
rect 16221 25245 16255 25279
rect 17417 25245 17451 25279
rect 17969 25245 18003 25279
rect 18061 25245 18095 25279
rect 18245 25245 18279 25279
rect 18521 25245 18555 25279
rect 18797 25245 18831 25279
rect 19901 25245 19935 25279
rect 20545 25245 20579 25279
rect 25053 25245 25087 25279
rect 25237 25245 25271 25279
rect 27261 25245 27295 25279
rect 27445 25245 27479 25279
rect 30481 25245 30515 25279
rect 30757 25245 30791 25279
rect 30849 25245 30883 25279
rect 31769 25245 31803 25279
rect 33333 25245 33367 25279
rect 33425 25245 33459 25279
rect 33517 25245 33551 25279
rect 33701 25245 33735 25279
rect 36277 25245 36311 25279
rect 36553 25245 36587 25279
rect 36829 25245 36863 25279
rect 37013 25245 37047 25279
rect 37105 25245 37139 25279
rect 37289 25245 37323 25279
rect 1685 25177 1719 25211
rect 4997 25177 5031 25211
rect 9229 25177 9263 25211
rect 10701 25177 10735 25211
rect 11437 25177 11471 25211
rect 14473 25177 14507 25211
rect 15945 25177 15979 25211
rect 17693 25177 17727 25211
rect 3801 25109 3835 25143
rect 6469 25109 6503 25143
rect 6929 25109 6963 25143
rect 8033 25109 8067 25143
rect 8493 25109 8527 25143
rect 9321 25109 9355 25143
rect 11069 25109 11103 25143
rect 14105 25109 14139 25143
rect 17785 25109 17819 25143
rect 27353 25109 27387 25143
rect 31861 25109 31895 25143
rect 36369 25109 36403 25143
rect 2513 24905 2547 24939
rect 2881 24905 2915 24939
rect 4077 24905 4111 24939
rect 11529 24905 11563 24939
rect 11897 24905 11931 24939
rect 19901 24905 19935 24939
rect 22201 24905 22235 24939
rect 27905 24905 27939 24939
rect 28549 24905 28583 24939
rect 34069 24905 34103 24939
rect 14105 24837 14139 24871
rect 16957 24837 16991 24871
rect 23857 24837 23891 24871
rect 28641 24837 28675 24871
rect 30573 24837 30607 24871
rect 2697 24769 2731 24803
rect 2973 24769 3007 24803
rect 4445 24769 4479 24803
rect 4721 24769 4755 24803
rect 5365 24769 5399 24803
rect 6837 24769 6871 24803
rect 7297 24769 7331 24803
rect 8033 24769 8067 24803
rect 11713 24769 11747 24803
rect 12081 24769 12115 24803
rect 13829 24769 13863 24803
rect 14013 24769 14047 24803
rect 14249 24769 14283 24803
rect 14749 24769 14783 24803
rect 14841 24769 14875 24803
rect 14933 24769 14967 24803
rect 15117 24769 15151 24803
rect 16865 24769 16899 24803
rect 17049 24769 17083 24803
rect 17233 24769 17267 24803
rect 18613 24769 18647 24803
rect 19533 24769 19567 24803
rect 22293 24769 22327 24803
rect 22845 24769 22879 24803
rect 23029 24769 23063 24803
rect 23121 24769 23155 24803
rect 23213 24769 23247 24803
rect 23673 24769 23707 24803
rect 23765 24769 23799 24803
rect 24041 24769 24075 24803
rect 24133 24769 24167 24803
rect 24317 24769 24351 24803
rect 24409 24769 24443 24803
rect 24506 24769 24540 24803
rect 24961 24769 24995 24803
rect 25881 24769 25915 24803
rect 26985 24769 27019 24803
rect 27169 24769 27203 24803
rect 27261 24769 27295 24803
rect 27445 24769 27479 24803
rect 27537 24769 27571 24803
rect 27629 24769 27663 24803
rect 29929 24769 29963 24803
rect 30205 24769 30239 24803
rect 30389 24769 30423 24803
rect 33241 24769 33275 24803
rect 33425 24769 33459 24803
rect 33609 24769 33643 24803
rect 34437 24769 34471 24803
rect 36369 24769 36403 24803
rect 36461 24769 36495 24803
rect 4353 24701 4387 24735
rect 4537 24701 4571 24735
rect 4905 24701 4939 24735
rect 5549 24701 5583 24735
rect 6653 24701 6687 24735
rect 7021 24701 7055 24735
rect 7481 24701 7515 24735
rect 8309 24701 8343 24735
rect 10057 24701 10091 24735
rect 12265 24701 12299 24735
rect 18705 24701 18739 24735
rect 18981 24701 19015 24735
rect 19441 24701 19475 24735
rect 22385 24701 22419 24735
rect 24702 24701 24736 24735
rect 26433 24701 26467 24735
rect 27905 24701 27939 24735
rect 28733 24701 28767 24735
rect 29745 24701 29779 24735
rect 34161 24701 34195 24735
rect 36553 24701 36587 24735
rect 36645 24701 36679 24735
rect 5181 24633 5215 24667
rect 28181 24633 28215 24667
rect 34345 24633 34379 24667
rect 4261 24565 4295 24599
rect 7113 24565 7147 24599
rect 14381 24565 14415 24599
rect 14565 24565 14599 24599
rect 16681 24565 16715 24599
rect 21833 24565 21867 24599
rect 23397 24565 23431 24599
rect 23489 24565 23523 24599
rect 27721 24565 27755 24599
rect 30113 24565 30147 24599
rect 33241 24565 33275 24599
rect 33701 24565 33735 24599
rect 34253 24565 34287 24599
rect 36829 24565 36863 24599
rect 6561 24361 6595 24395
rect 11897 24361 11931 24395
rect 25421 24361 25455 24395
rect 26801 24361 26835 24395
rect 27077 24361 27111 24395
rect 27721 24361 27755 24395
rect 28641 24361 28675 24395
rect 29101 24361 29135 24395
rect 31033 24361 31067 24395
rect 33149 24361 33183 24395
rect 34897 24361 34931 24395
rect 11989 24293 12023 24327
rect 15117 24293 15151 24327
rect 16037 24293 16071 24327
rect 21833 24293 21867 24327
rect 23673 24293 23707 24327
rect 35633 24293 35667 24327
rect 2973 24225 3007 24259
rect 4537 24225 4571 24259
rect 5549 24225 5583 24259
rect 13277 24225 13311 24259
rect 14473 24225 14507 24259
rect 22385 24225 22419 24259
rect 22585 24225 22619 24259
rect 27905 24225 27939 24259
rect 31769 24225 31803 24259
rect 35725 24225 35759 24259
rect 2697 24157 2731 24191
rect 3801 24157 3835 24191
rect 4721 24157 4755 24191
rect 5089 24157 5123 24191
rect 5733 24157 5767 24191
rect 5917 24157 5951 24191
rect 6745 24157 6779 24191
rect 6929 24157 6963 24191
rect 9229 24157 9263 24191
rect 9505 24157 9539 24191
rect 12357 24157 12391 24191
rect 13185 24157 13219 24191
rect 13461 24157 13495 24191
rect 13645 24157 13679 24191
rect 14105 24157 14139 24191
rect 15392 24157 15426 24191
rect 15485 24157 15519 24191
rect 15577 24157 15611 24191
rect 15761 24157 15795 24191
rect 16037 24157 16071 24191
rect 16405 24157 16439 24191
rect 16773 24157 16807 24191
rect 21281 24157 21315 24191
rect 21465 24157 21499 24191
rect 21654 24157 21688 24191
rect 22293 24157 22327 24191
rect 23121 24157 23155 24191
rect 23305 24157 23339 24191
rect 23397 24157 23431 24191
rect 23541 24157 23575 24191
rect 24501 24157 24535 24191
rect 24869 24157 24903 24191
rect 25053 24157 25087 24191
rect 25329 24157 25363 24191
rect 26065 24157 26099 24191
rect 26157 24157 26191 24191
rect 26341 24157 26375 24191
rect 27261 24157 27295 24191
rect 27353 24157 27387 24191
rect 27537 24157 27571 24191
rect 27629 24157 27663 24191
rect 27997 24157 28031 24191
rect 28089 24157 28123 24191
rect 28181 24157 28215 24191
rect 28365 24157 28399 24191
rect 28457 24157 28491 24191
rect 28733 24157 28767 24191
rect 28917 24157 28951 24191
rect 29009 24157 29043 24191
rect 29193 24157 29227 24191
rect 30481 24157 30515 24191
rect 30849 24157 30883 24191
rect 31953 24157 31987 24191
rect 32873 24167 32907 24201
rect 33701 24157 33735 24191
rect 33977 24157 34011 24191
rect 34713 24157 34747 24191
rect 34897 24157 34931 24191
rect 35203 24157 35237 24191
rect 36553 24157 36587 24191
rect 37197 24157 37231 24191
rect 9781 24089 9815 24123
rect 14289 24089 14323 24123
rect 21557 24089 21591 24123
rect 22845 24089 22879 24123
rect 23029 24089 23063 24123
rect 26525 24089 26559 24123
rect 26709 24089 26743 24123
rect 28641 24089 28675 24123
rect 30665 24089 30699 24123
rect 30757 24089 30791 24123
rect 33149 24089 33183 24123
rect 34529 24089 34563 24123
rect 2329 24021 2363 24055
rect 2789 24021 2823 24055
rect 4445 24021 4479 24055
rect 4997 24021 5031 24055
rect 9413 24021 9447 24055
rect 11253 24021 11287 24055
rect 22477 24021 22511 24055
rect 28825 24021 28859 24055
rect 32045 24021 32079 24055
rect 32413 24021 32447 24055
rect 32965 24021 32999 24055
rect 35081 24021 35115 24055
rect 35265 24021 35299 24055
rect 2789 23817 2823 23851
rect 13093 23817 13127 23851
rect 13461 23817 13495 23851
rect 16681 23817 16715 23851
rect 31033 23817 31067 23851
rect 34989 23817 35023 23851
rect 35817 23817 35851 23851
rect 36277 23817 36311 23851
rect 36737 23817 36771 23851
rect 2421 23749 2455 23783
rect 9413 23749 9447 23783
rect 13185 23749 13219 23783
rect 20913 23749 20947 23783
rect 23857 23749 23891 23783
rect 23949 23749 23983 23783
rect 25513 23749 25547 23783
rect 32873 23749 32907 23783
rect 36921 23749 36955 23783
rect 1961 23681 1995 23715
rect 2237 23681 2271 23715
rect 2513 23681 2547 23715
rect 2605 23681 2639 23715
rect 5457 23681 5491 23715
rect 6653 23681 6687 23715
rect 9321 23681 9355 23715
rect 11529 23681 11563 23715
rect 12909 23681 12943 23715
rect 13277 23681 13311 23715
rect 13737 23681 13771 23715
rect 14105 23681 14139 23715
rect 14473 23681 14507 23715
rect 17049 23681 17083 23715
rect 18429 23681 18463 23715
rect 18613 23681 18647 23715
rect 20637 23681 20671 23715
rect 20821 23681 20855 23715
rect 21005 23681 21039 23715
rect 23673 23681 23707 23715
rect 24046 23681 24080 23715
rect 25605 23681 25639 23715
rect 29561 23681 29595 23715
rect 30941 23681 30975 23715
rect 31125 23681 31159 23715
rect 32137 23681 32171 23715
rect 32285 23681 32319 23715
rect 32413 23681 32447 23715
rect 32505 23681 32539 23715
rect 32602 23681 32636 23715
rect 33149 23681 33183 23715
rect 33333 23681 33367 23715
rect 35265 23681 35299 23715
rect 35725 23681 35759 23715
rect 35909 23681 35943 23715
rect 36461 23681 36495 23715
rect 36553 23681 36587 23715
rect 36645 23681 36679 23715
rect 3525 23613 3559 23647
rect 5089 23613 5123 23647
rect 6929 23613 6963 23647
rect 11897 23613 11931 23647
rect 17141 23613 17175 23647
rect 17325 23613 17359 23647
rect 25421 23613 25455 23647
rect 29377 23613 29411 23647
rect 29745 23613 29779 23647
rect 35173 23613 35207 23647
rect 35633 23613 35667 23647
rect 36277 23613 36311 23647
rect 3663 23545 3697 23579
rect 8401 23545 8435 23579
rect 21189 23545 21223 23579
rect 36921 23545 36955 23579
rect 1777 23477 1811 23511
rect 2881 23477 2915 23511
rect 18521 23477 18555 23511
rect 24225 23477 24259 23511
rect 25973 23477 26007 23511
rect 32781 23477 32815 23511
rect 32965 23477 32999 23511
rect 33517 23477 33551 23511
rect 3157 23273 3191 23307
rect 3893 23273 3927 23307
rect 4261 23273 4295 23307
rect 7021 23273 7055 23307
rect 9597 23273 9631 23307
rect 9781 23273 9815 23307
rect 15853 23273 15887 23307
rect 16773 23273 16807 23307
rect 16957 23273 16991 23307
rect 19257 23273 19291 23307
rect 20177 23273 20211 23307
rect 22385 23273 22419 23307
rect 24961 23273 24995 23307
rect 27629 23273 27663 23307
rect 30297 23273 30331 23307
rect 36461 23273 36495 23307
rect 7297 23205 7331 23239
rect 13461 23205 13495 23239
rect 17693 23205 17727 23239
rect 24869 23205 24903 23239
rect 32229 23205 32263 23239
rect 1685 23137 1719 23171
rect 7941 23137 7975 23171
rect 12633 23137 12667 23171
rect 18337 23137 18371 23171
rect 19717 23137 19751 23171
rect 19901 23137 19935 23171
rect 22569 23137 22603 23171
rect 25053 23137 25087 23171
rect 27997 23137 28031 23171
rect 28089 23137 28123 23171
rect 29193 23137 29227 23171
rect 29929 23137 29963 23171
rect 31677 23137 31711 23171
rect 1409 23069 1443 23103
rect 3985 23069 4019 23103
rect 4353 23069 4387 23103
rect 7205 23069 7239 23103
rect 7665 23069 7699 23103
rect 10885 23069 10919 23103
rect 11069 23069 11103 23103
rect 11989 23069 12023 23103
rect 12081 23069 12115 23103
rect 12265 23069 12299 23103
rect 13553 23069 13587 23103
rect 13737 23069 13771 23103
rect 14565 23069 14599 23103
rect 14933 23069 14967 23103
rect 15117 23069 15151 23103
rect 15669 23069 15703 23103
rect 15853 23069 15887 23103
rect 16497 23069 16531 23103
rect 16681 23069 16715 23103
rect 17233 23069 17267 23103
rect 17325 23069 17359 23103
rect 17417 23069 17451 23103
rect 17601 23069 17635 23103
rect 18521 23069 18555 23103
rect 18705 23069 18739 23103
rect 20269 23069 20303 23103
rect 20453 23069 20487 23103
rect 21005 23069 21039 23103
rect 21189 23069 21223 23103
rect 21373 23069 21407 23103
rect 22937 23069 22971 23103
rect 24777 23069 24811 23103
rect 26525 23069 26559 23103
rect 26709 23069 26743 23103
rect 26893 23069 26927 23103
rect 27813 23069 27847 23103
rect 27905 23069 27939 23103
rect 28825 23069 28859 23103
rect 29009 23069 29043 23103
rect 30113 23069 30147 23103
rect 30297 23069 30331 23103
rect 36645 23069 36679 23103
rect 36921 23069 36955 23103
rect 37105 23069 37139 23103
rect 7757 23001 7791 23035
rect 9965 23001 9999 23035
rect 11529 23001 11563 23035
rect 12817 23001 12851 23035
rect 13001 23001 13035 23035
rect 16865 23001 16899 23035
rect 18061 23001 18095 23035
rect 20729 23001 20763 23035
rect 29653 23001 29687 23035
rect 31861 23001 31895 23035
rect 9781 22933 9815 22967
rect 10609 22933 10643 22967
rect 12449 22933 12483 22967
rect 16037 22933 16071 22967
rect 18153 22933 18187 22967
rect 18613 22933 18647 22967
rect 19625 22933 19659 22967
rect 22753 22933 22787 22967
rect 30481 22933 30515 22967
rect 31769 22933 31803 22967
rect 6837 22729 6871 22763
rect 9229 22729 9263 22763
rect 14565 22729 14599 22763
rect 15945 22729 15979 22763
rect 16773 22729 16807 22763
rect 17601 22729 17635 22763
rect 19901 22729 19935 22763
rect 23689 22729 23723 22763
rect 23857 22729 23891 22763
rect 25973 22729 26007 22763
rect 31125 22729 31159 22763
rect 31309 22729 31343 22763
rect 35081 22729 35115 22763
rect 35265 22729 35299 22763
rect 36185 22729 36219 22763
rect 36651 22729 36685 22763
rect 6929 22661 6963 22695
rect 9597 22661 9631 22695
rect 12265 22661 12299 22695
rect 15761 22661 15795 22695
rect 22753 22661 22787 22695
rect 23489 22661 23523 22695
rect 26985 22661 27019 22695
rect 27169 22661 27203 22695
rect 27353 22661 27387 22695
rect 28641 22661 28675 22695
rect 29995 22661 30029 22695
rect 30113 22661 30147 22695
rect 30205 22661 30239 22695
rect 31861 22661 31895 22695
rect 33793 22661 33827 22695
rect 35173 22661 35207 22695
rect 36553 22661 36587 22695
rect 36737 22661 36771 22695
rect 9321 22593 9355 22627
rect 9413 22593 9447 22627
rect 9781 22593 9815 22627
rect 9965 22593 9999 22627
rect 11529 22593 11563 22627
rect 11621 22593 11655 22627
rect 11805 22593 11839 22627
rect 13921 22593 13955 22627
rect 14105 22593 14139 22627
rect 14197 22593 14231 22627
rect 14289 22593 14323 22627
rect 16681 22593 16715 22627
rect 16865 22593 16899 22627
rect 17509 22593 17543 22627
rect 17693 22593 17727 22627
rect 18429 22593 18463 22627
rect 19717 22593 19751 22627
rect 19993 22593 20027 22627
rect 20729 22593 20763 22627
rect 22017 22593 22051 22627
rect 22201 22593 22235 22627
rect 22293 22593 22327 22627
rect 22419 22593 22453 22627
rect 23029 22593 23063 22627
rect 23121 22593 23155 22627
rect 23213 22593 23247 22627
rect 23397 22593 23431 22627
rect 24133 22593 24167 22627
rect 24869 22593 24903 22627
rect 25513 22593 25547 22627
rect 25697 22593 25731 22627
rect 25789 22593 25823 22627
rect 26157 22593 26191 22627
rect 26341 22593 26375 22627
rect 28273 22593 28307 22627
rect 28457 22593 28491 22627
rect 30297 22593 30331 22627
rect 30573 22593 30607 22627
rect 30665 22593 30699 22627
rect 30849 22593 30883 22627
rect 30941 22593 30975 22627
rect 31493 22593 31527 22627
rect 31585 22593 31619 22627
rect 32137 22593 32171 22627
rect 32230 22593 32264 22627
rect 32413 22593 32447 22627
rect 32505 22593 32539 22627
rect 32643 22593 32677 22627
rect 33701 22593 33735 22627
rect 33885 22593 33919 22627
rect 34161 22593 34195 22627
rect 34345 22593 34379 22627
rect 34529 22593 34563 22627
rect 34713 22593 34747 22627
rect 35397 22593 35431 22627
rect 35541 22593 35575 22627
rect 35633 22593 35667 22627
rect 35817 22593 35851 22627
rect 35909 22593 35943 22627
rect 36001 22593 36035 22627
rect 36829 22593 36863 22627
rect 37657 22593 37691 22627
rect 7021 22525 7055 22559
rect 15393 22525 15427 22559
rect 18337 22525 18371 22559
rect 21097 22525 21131 22559
rect 24593 22525 24627 22559
rect 25605 22525 25639 22559
rect 26525 22525 26559 22559
rect 29837 22525 29871 22559
rect 30481 22525 30515 22559
rect 31953 22525 31987 22559
rect 34437 22525 34471 22559
rect 34897 22525 34931 22559
rect 37565 22525 37599 22559
rect 9045 22457 9079 22491
rect 22661 22457 22695 22491
rect 6469 22389 6503 22423
rect 9781 22389 9815 22423
rect 15761 22389 15795 22423
rect 18153 22389 18187 22423
rect 19533 22389 19567 22423
rect 23673 22389 23707 22423
rect 32781 22389 32815 22423
rect 37381 22389 37415 22423
rect 10149 22185 10183 22219
rect 13461 22185 13495 22219
rect 17141 22185 17175 22219
rect 17509 22185 17543 22219
rect 18153 22185 18187 22219
rect 23673 22185 23707 22219
rect 32321 22185 32355 22219
rect 33517 22185 33551 22219
rect 35449 22185 35483 22219
rect 35909 22185 35943 22219
rect 9505 22117 9539 22151
rect 17693 22117 17727 22151
rect 25973 22117 26007 22151
rect 27353 22117 27387 22151
rect 30113 22117 30147 22151
rect 33885 22117 33919 22151
rect 3157 22049 3191 22083
rect 4353 22049 4387 22083
rect 14381 22049 14415 22083
rect 17601 22049 17635 22083
rect 18245 22049 18279 22083
rect 20545 22049 20579 22083
rect 23397 22049 23431 22083
rect 25145 22049 25179 22083
rect 26893 22049 26927 22083
rect 27721 22049 27755 22083
rect 28825 22049 28859 22083
rect 33333 22049 33367 22083
rect 33793 22049 33827 22083
rect 2881 21981 2915 22015
rect 3525 21981 3559 22015
rect 4169 21981 4203 22015
rect 4997 21981 5031 22015
rect 5733 21981 5767 22015
rect 8401 21981 8435 22015
rect 8585 21981 8619 22015
rect 8769 21981 8803 22015
rect 8953 21981 8987 22015
rect 9137 21981 9171 22015
rect 9229 21981 9263 22015
rect 9965 21981 9999 22015
rect 10241 21981 10275 22015
rect 12357 21981 12391 22015
rect 12817 21981 12851 22015
rect 13553 21981 13587 22015
rect 14289 21981 14323 22015
rect 15853 21981 15887 22015
rect 17417 21981 17451 22015
rect 17877 21981 17911 22015
rect 18153 21981 18187 22015
rect 18613 21981 18647 22015
rect 20637 21981 20671 22015
rect 22109 21981 22143 22015
rect 22293 21981 22327 22015
rect 22845 21981 22879 22015
rect 23029 21981 23063 22015
rect 24593 21981 24627 22015
rect 25329 21981 25363 22015
rect 25789 21981 25823 22015
rect 26525 21981 26559 22015
rect 26709 21981 26743 22015
rect 27537 21981 27571 22015
rect 27813 21981 27847 22015
rect 28089 21981 28123 22015
rect 28273 21981 28307 22015
rect 28733 21981 28767 22015
rect 29561 21981 29595 22015
rect 29929 21981 29963 22015
rect 32045 21981 32079 22015
rect 32137 21981 32171 22015
rect 32689 21981 32723 22015
rect 32873 21981 32907 22015
rect 33149 21981 33183 22015
rect 33425 21981 33459 22015
rect 33701 21981 33735 22015
rect 34805 21981 34839 22015
rect 34898 21981 34932 22015
rect 35173 21981 35207 22015
rect 35270 21981 35304 22015
rect 35541 21981 35575 22015
rect 2973 21913 3007 21947
rect 6009 21913 6043 21947
rect 7757 21913 7791 21947
rect 9505 21913 9539 21947
rect 11897 21913 11931 21947
rect 11989 21913 12023 21947
rect 12449 21913 12483 21947
rect 13737 21913 13771 21947
rect 15577 21913 15611 21947
rect 16037 21913 16071 21947
rect 23489 21913 23523 21947
rect 23689 21913 23723 21947
rect 29745 21913 29779 21947
rect 29837 21913 29871 21947
rect 31677 21913 31711 21947
rect 31769 21913 31803 21947
rect 35081 21913 35115 21947
rect 35725 21913 35759 21947
rect 2513 21845 2547 21879
rect 3341 21845 3375 21879
rect 3801 21845 3835 21879
rect 4261 21845 4295 21879
rect 4813 21845 4847 21879
rect 9137 21845 9171 21879
rect 9321 21845 9355 21879
rect 9689 21845 9723 21879
rect 12909 21845 12943 21879
rect 15669 21845 15703 21879
rect 17969 21845 18003 21879
rect 20729 21845 20763 21879
rect 21097 21845 21131 21879
rect 23857 21845 23891 21879
rect 5181 21641 5215 21675
rect 6377 21641 6411 21675
rect 9137 21641 9171 21675
rect 9505 21641 9539 21675
rect 15025 21641 15059 21675
rect 17325 21641 17359 21675
rect 17693 21641 17727 21675
rect 18245 21641 18279 21675
rect 24501 21641 24535 21675
rect 25805 21641 25839 21675
rect 25973 21641 26007 21675
rect 26617 21641 26651 21675
rect 27629 21641 27663 21675
rect 28917 21641 28951 21675
rect 30021 21641 30055 21675
rect 34989 21641 35023 21675
rect 36737 21641 36771 21675
rect 3065 21573 3099 21607
rect 4813 21573 4847 21607
rect 10977 21573 11011 21607
rect 13461 21573 13495 21607
rect 14657 21573 14691 21607
rect 14749 21573 14783 21607
rect 17877 21573 17911 21607
rect 18061 21573 18095 21607
rect 21281 21573 21315 21607
rect 25605 21573 25639 21607
rect 1777 21505 1811 21539
rect 2145 21505 2179 21539
rect 2789 21505 2823 21539
rect 5549 21505 5583 21539
rect 5641 21505 5675 21539
rect 6561 21505 6595 21539
rect 8585 21505 8619 21539
rect 8677 21505 8711 21539
rect 8861 21505 8895 21539
rect 8953 21505 8987 21539
rect 9689 21505 9723 21539
rect 9873 21505 9907 21539
rect 10701 21505 10735 21539
rect 10885 21505 10919 21539
rect 11069 21505 11103 21539
rect 11161 21505 11195 21539
rect 11345 21505 11379 21539
rect 11621 21505 11655 21539
rect 11989 21505 12023 21539
rect 13645 21505 13679 21539
rect 13829 21505 13863 21539
rect 13921 21505 13955 21539
rect 14013 21505 14047 21539
rect 14381 21505 14415 21539
rect 14474 21505 14508 21539
rect 14887 21505 14921 21539
rect 15761 21505 15795 21539
rect 16129 21505 16163 21539
rect 16865 21505 16899 21539
rect 17141 21505 17175 21539
rect 17233 21505 17267 21539
rect 17417 21505 17451 21539
rect 18153 21505 18187 21539
rect 18337 21505 18371 21539
rect 19441 21505 19475 21539
rect 19809 21505 19843 21539
rect 20269 21505 20303 21539
rect 20637 21505 20671 21539
rect 20821 21505 20855 21539
rect 20913 21505 20947 21539
rect 21006 21511 21040 21545
rect 22661 21505 22695 21539
rect 23213 21505 23247 21539
rect 23305 21505 23339 21539
rect 24317 21505 24351 21539
rect 26801 21505 26835 21539
rect 26985 21505 27019 21539
rect 27261 21505 27295 21539
rect 27813 21505 27847 21539
rect 27997 21505 28031 21539
rect 28733 21505 28767 21539
rect 29561 21505 29595 21539
rect 29653 21505 29687 21539
rect 29837 21505 29871 21539
rect 34989 21505 35023 21539
rect 35166 21505 35200 21539
rect 36921 21505 36955 21539
rect 37105 21505 37139 21539
rect 37657 21505 37691 21539
rect 5825 21437 5859 21471
rect 9781 21437 9815 21471
rect 9965 21437 9999 21471
rect 10425 21437 10459 21471
rect 14289 21437 14323 21471
rect 15485 21437 15519 21471
rect 17049 21437 17083 21471
rect 24133 21437 24167 21471
rect 26249 21437 26283 21471
rect 26341 21437 26375 21471
rect 28549 21437 28583 21471
rect 16129 21369 16163 21403
rect 20361 21369 20395 21403
rect 22753 21369 22787 21403
rect 1501 21301 1535 21335
rect 1961 21301 1995 21335
rect 10149 21301 10183 21335
rect 10609 21301 10643 21335
rect 11161 21301 11195 21335
rect 16681 21301 16715 21335
rect 25789 21301 25823 21335
rect 27077 21301 27111 21335
rect 27537 21301 27571 21335
rect 37841 21301 37875 21335
rect 1672 21097 1706 21131
rect 6101 21097 6135 21131
rect 13737 21097 13771 21131
rect 13921 21097 13955 21131
rect 19533 21097 19567 21131
rect 25421 21097 25455 21131
rect 30757 21097 30791 21131
rect 32873 21097 32907 21131
rect 34713 21097 34747 21131
rect 14105 21029 14139 21063
rect 20821 21029 20855 21063
rect 31033 21029 31067 21063
rect 31493 21029 31527 21063
rect 34437 21029 34471 21063
rect 36737 21029 36771 21063
rect 36921 21029 36955 21063
rect 1409 20961 1443 20995
rect 4353 20961 4387 20995
rect 25237 20961 25271 20995
rect 31217 20961 31251 20995
rect 33333 20961 33367 20995
rect 33977 20961 34011 20995
rect 36277 20961 36311 20995
rect 36829 20961 36863 20995
rect 8033 20893 8067 20927
rect 9965 20893 9999 20927
rect 10977 20893 11011 20927
rect 11161 20893 11195 20927
rect 11529 20893 11563 20927
rect 11621 20893 11655 20927
rect 11897 20893 11931 20927
rect 14243 20893 14277 20927
rect 14381 20893 14415 20927
rect 14473 20893 14507 20927
rect 14656 20893 14690 20927
rect 14749 20893 14783 20927
rect 16497 20893 16531 20927
rect 19441 20893 19475 20927
rect 19809 20893 19843 20927
rect 20453 20893 20487 20927
rect 21189 20893 21223 20927
rect 25697 20893 25731 20927
rect 27261 20893 27295 20927
rect 30113 20893 30147 20927
rect 30297 20893 30331 20927
rect 30481 20893 30515 20927
rect 30941 20893 30975 20927
rect 31125 20893 31159 20927
rect 31401 20893 31435 20927
rect 31769 20893 31803 20927
rect 33057 20893 33091 20927
rect 33149 20893 33183 20927
rect 33425 20893 33459 20927
rect 34069 20893 34103 20927
rect 34713 20893 34747 20927
rect 34897 20893 34931 20927
rect 36369 20893 36403 20927
rect 37059 20893 37093 20927
rect 37197 20893 37231 20927
rect 4629 20825 4663 20859
rect 6285 20825 6319 20859
rect 12357 20825 12391 20859
rect 13553 20825 13587 20859
rect 15761 20825 15795 20859
rect 21373 20825 21407 20859
rect 21557 20825 21591 20859
rect 24409 20825 24443 20859
rect 25421 20825 25455 20859
rect 31493 20825 31527 20859
rect 31677 20825 31711 20859
rect 3157 20757 3191 20791
rect 9873 20757 9907 20791
rect 13753 20757 13787 20791
rect 25605 20757 25639 20791
rect 27077 20757 27111 20791
rect 6745 20553 6779 20587
rect 9413 20553 9447 20587
rect 9781 20553 9815 20587
rect 17049 20553 17083 20587
rect 19441 20553 19475 20587
rect 22661 20553 22695 20587
rect 23949 20553 23983 20587
rect 24041 20553 24075 20587
rect 24409 20553 24443 20587
rect 24685 20553 24719 20587
rect 30205 20553 30239 20587
rect 31033 20553 31067 20587
rect 33885 20553 33919 20587
rect 34069 20553 34103 20587
rect 37105 20553 37139 20587
rect 7113 20485 7147 20519
rect 7205 20485 7239 20519
rect 8493 20485 8527 20519
rect 15485 20485 15519 20519
rect 25849 20485 25883 20519
rect 26065 20485 26099 20519
rect 31953 20485 31987 20519
rect 36737 20485 36771 20519
rect 36937 20485 36971 20519
rect 6653 20417 6687 20451
rect 8125 20417 8159 20451
rect 9045 20417 9079 20451
rect 9321 20417 9355 20451
rect 9597 20417 9631 20451
rect 10701 20417 10735 20451
rect 13093 20417 13127 20451
rect 13461 20417 13495 20451
rect 13921 20417 13955 20451
rect 15669 20417 15703 20451
rect 17141 20417 17175 20451
rect 17785 20417 17819 20451
rect 18521 20417 18555 20451
rect 18705 20417 18739 20451
rect 19441 20417 19475 20451
rect 19901 20417 19935 20451
rect 21005 20417 21039 20451
rect 22569 20417 22603 20451
rect 24593 20417 24627 20451
rect 24777 20417 24811 20451
rect 27169 20417 27203 20451
rect 27905 20417 27939 20451
rect 29009 20417 29043 20451
rect 29101 20417 29135 20451
rect 29377 20417 29411 20451
rect 29561 20417 29595 20451
rect 29745 20417 29779 20451
rect 30113 20417 30147 20451
rect 30389 20417 30423 20451
rect 30481 20417 30515 20451
rect 30573 20417 30607 20451
rect 31126 20417 31160 20451
rect 31566 20417 31600 20451
rect 31677 20417 31711 20451
rect 31769 20417 31803 20451
rect 33701 20417 33735 20451
rect 33977 20417 34011 20451
rect 34161 20417 34195 20451
rect 7297 20349 7331 20383
rect 10793 20349 10827 20383
rect 14197 20349 14231 20383
rect 16865 20349 16899 20383
rect 20729 20349 20763 20383
rect 20913 20349 20947 20383
rect 22845 20349 22879 20383
rect 23765 20349 23799 20383
rect 29929 20349 29963 20383
rect 31473 20349 31507 20383
rect 33425 20349 33459 20383
rect 8677 20281 8711 20315
rect 31953 20281 31987 20315
rect 33517 20281 33551 20315
rect 6469 20213 6503 20247
rect 8493 20213 8527 20247
rect 9137 20213 9171 20247
rect 10701 20213 10735 20247
rect 11069 20213 11103 20247
rect 15853 20213 15887 20247
rect 17509 20213 17543 20247
rect 17693 20213 17727 20247
rect 18613 20213 18647 20247
rect 21373 20213 21407 20247
rect 22201 20213 22235 20247
rect 25697 20213 25731 20247
rect 25881 20213 25915 20247
rect 27353 20213 27387 20247
rect 36921 20213 36955 20247
rect 7941 20009 7975 20043
rect 14565 20009 14599 20043
rect 30389 20009 30423 20043
rect 30573 20009 30607 20043
rect 30849 20009 30883 20043
rect 31493 20009 31527 20043
rect 33885 20009 33919 20043
rect 34805 20009 34839 20043
rect 36093 20009 36127 20043
rect 36553 20009 36587 20043
rect 36737 20009 36771 20043
rect 2605 19941 2639 19975
rect 17601 19941 17635 19975
rect 28089 19941 28123 19975
rect 30113 19941 30147 19975
rect 32045 19941 32079 19975
rect 33241 19941 33275 19975
rect 3249 19873 3283 19907
rect 3801 19873 3835 19907
rect 6193 19873 6227 19907
rect 6469 19873 6503 19907
rect 9505 19873 9539 19907
rect 12817 19873 12851 19907
rect 13369 19873 13403 19907
rect 16957 19873 16991 19907
rect 17141 19873 17175 19907
rect 19993 19873 20027 19907
rect 20453 19873 20487 19907
rect 21649 19873 21683 19907
rect 22109 19873 22143 19907
rect 24593 19873 24627 19907
rect 24685 19873 24719 19907
rect 31125 19873 31159 19907
rect 31217 19873 31251 19907
rect 35265 19873 35299 19907
rect 35541 19873 35575 19907
rect 2145 19805 2179 19839
rect 2973 19805 3007 19839
rect 9413 19805 9447 19839
rect 9781 19805 9815 19839
rect 9873 19805 9907 19839
rect 12173 19805 12207 19839
rect 12357 19805 12391 19839
rect 12449 19805 12483 19839
rect 12541 19805 12575 19839
rect 13093 19805 13127 19839
rect 13185 19805 13219 19839
rect 13553 19805 13587 19839
rect 14197 19805 14231 19839
rect 14933 19805 14967 19839
rect 15117 19805 15151 19839
rect 15669 19805 15703 19839
rect 16129 19805 16163 19839
rect 17877 19805 17911 19839
rect 19073 19805 19107 19839
rect 20177 19805 20211 19839
rect 20545 19805 20579 19839
rect 21557 19805 21591 19839
rect 21833 19805 21867 19839
rect 25237 19805 25271 19839
rect 27261 19805 27295 19839
rect 27721 19805 27755 19839
rect 27905 19805 27939 19839
rect 28273 19805 28307 19839
rect 28641 19805 28675 19839
rect 29561 19805 29595 19839
rect 29837 19805 29871 19839
rect 29929 19805 29963 19839
rect 30665 19805 30699 19839
rect 30849 19805 30883 19839
rect 31033 19805 31067 19839
rect 31309 19805 31343 19839
rect 31769 19805 31803 19839
rect 31861 19805 31895 19839
rect 33425 19805 33459 19839
rect 33701 19805 33735 19839
rect 33793 19805 33827 19839
rect 33977 19805 34011 19839
rect 35173 19805 35207 19839
rect 35449 19805 35483 19839
rect 35817 19805 35851 19839
rect 35909 19805 35943 19839
rect 36369 19805 36403 19839
rect 36645 19805 36679 19839
rect 36829 19805 36863 19839
rect 30435 19771 30469 19805
rect 4077 19737 4111 19771
rect 10149 19737 10183 19771
rect 10517 19737 10551 19771
rect 18245 19737 18279 19771
rect 19533 19737 19567 19771
rect 19717 19737 19751 19771
rect 19901 19737 19935 19771
rect 21189 19737 21223 19771
rect 22385 19737 22419 19771
rect 24777 19737 24811 19771
rect 25513 19737 25547 19771
rect 29745 19737 29779 19771
rect 30205 19737 30239 19771
rect 32045 19737 32079 19771
rect 36185 19737 36219 19771
rect 1961 19669 1995 19703
rect 3065 19669 3099 19703
rect 5549 19669 5583 19703
rect 10057 19669 10091 19703
rect 10333 19669 10367 19703
rect 10425 19669 10459 19703
rect 10609 19669 10643 19703
rect 14565 19669 14599 19703
rect 14749 19669 14783 19703
rect 15209 19669 15243 19703
rect 15485 19669 15519 19703
rect 17233 19669 17267 19703
rect 17693 19669 17727 19703
rect 22017 19669 22051 19703
rect 23857 19669 23891 19703
rect 25145 19669 25179 19703
rect 33609 19669 33643 19703
rect 4077 19465 4111 19499
rect 4353 19465 4387 19499
rect 4813 19465 4847 19499
rect 6745 19465 6779 19499
rect 12659 19465 12693 19499
rect 18797 19465 18831 19499
rect 22017 19465 22051 19499
rect 22477 19465 22511 19499
rect 25053 19465 25087 19499
rect 25421 19465 25455 19499
rect 26985 19465 27019 19499
rect 30573 19465 30607 19499
rect 31493 19465 31527 19499
rect 35081 19465 35115 19499
rect 35449 19465 35483 19499
rect 1685 19397 1719 19431
rect 4721 19397 4755 19431
rect 10241 19397 10275 19431
rect 12449 19397 12483 19431
rect 13645 19397 13679 19431
rect 15945 19397 15979 19431
rect 27153 19397 27187 19431
rect 27353 19397 27387 19431
rect 34161 19397 34195 19431
rect 34989 19397 35023 19431
rect 1409 19329 1443 19363
rect 4261 19329 4295 19363
rect 6837 19329 6871 19363
rect 9689 19329 9723 19363
rect 10057 19329 10091 19363
rect 10333 19329 10367 19363
rect 11713 19329 11747 19363
rect 12081 19329 12115 19363
rect 12909 19329 12943 19363
rect 13093 19329 13127 19363
rect 14749 19329 14783 19363
rect 15301 19329 15335 19363
rect 15393 19329 15427 19363
rect 15577 19329 15611 19363
rect 17049 19329 17083 19363
rect 22385 19329 22419 19363
rect 24869 19329 24903 19363
rect 25513 19329 25547 19363
rect 26157 19329 26191 19363
rect 28365 19329 28399 19363
rect 30481 19329 30515 19363
rect 31401 19329 31435 19363
rect 31677 19329 31711 19363
rect 33793 19329 33827 19363
rect 33977 19329 34011 19363
rect 34437 19329 34471 19363
rect 34621 19329 34655 19363
rect 35449 19329 35483 19363
rect 35633 19329 35667 19363
rect 37933 19329 37967 19363
rect 3157 19261 3191 19295
rect 4905 19261 4939 19295
rect 6929 19261 6963 19295
rect 9505 19261 9539 19295
rect 9965 19261 9999 19295
rect 11621 19261 11655 19295
rect 17325 19261 17359 19295
rect 22661 19261 22695 19295
rect 26433 19261 26467 19295
rect 28549 19261 28583 19295
rect 31861 19261 31895 19295
rect 34805 19261 34839 19295
rect 12265 19193 12299 19227
rect 12817 19193 12851 19227
rect 6377 19125 6411 19159
rect 9873 19125 9907 19159
rect 10057 19125 10091 19159
rect 11989 19125 12023 19159
rect 12633 19125 12667 19159
rect 13093 19125 13127 19159
rect 13921 19125 13955 19159
rect 14657 19125 14691 19159
rect 25973 19125 26007 19159
rect 26341 19125 26375 19159
rect 27169 19125 27203 19159
rect 37749 19125 37783 19159
rect 9597 18921 9631 18955
rect 12725 18921 12759 18955
rect 13737 18921 13771 18955
rect 24409 18921 24443 18955
rect 33885 18921 33919 18955
rect 34253 18921 34287 18955
rect 34437 18921 34471 18955
rect 37565 18921 37599 18955
rect 8217 18853 8251 18887
rect 33793 18853 33827 18887
rect 1685 18785 1719 18819
rect 4261 18785 4295 18819
rect 4445 18785 4479 18819
rect 8493 18785 8527 18819
rect 12909 18785 12943 18819
rect 14841 18785 14875 18819
rect 18705 18785 18739 18819
rect 21925 18785 21959 18819
rect 23029 18785 23063 18819
rect 1409 18717 1443 18751
rect 2513 18717 2547 18751
rect 4169 18717 4203 18751
rect 5825 18717 5859 18751
rect 8401 18717 8435 18751
rect 9321 18717 9355 18751
rect 9505 18717 9539 18751
rect 9781 18717 9815 18751
rect 10057 18717 10091 18751
rect 10156 18717 10190 18751
rect 10303 18717 10337 18751
rect 12173 18717 12207 18751
rect 12541 18717 12575 18751
rect 12817 18717 12851 18751
rect 13093 18717 13127 18751
rect 13185 18717 13219 18751
rect 14381 18717 14415 18751
rect 14565 18717 14599 18751
rect 14933 18717 14967 18751
rect 15301 18717 15335 18751
rect 15761 18717 15795 18751
rect 16313 18717 16347 18751
rect 18613 18717 18647 18751
rect 18889 18717 18923 18751
rect 19441 18717 19475 18751
rect 19533 18717 19567 18751
rect 19717 18717 19751 18751
rect 21557 18717 21591 18751
rect 22109 18717 22143 18751
rect 22385 18717 22419 18751
rect 22477 18717 22511 18751
rect 24685 18717 24719 18751
rect 24777 18717 24811 18751
rect 24869 18717 24903 18751
rect 25053 18717 25087 18751
rect 28733 18717 28767 18751
rect 29009 18717 29043 18751
rect 29377 18717 29411 18751
rect 32413 18717 32447 18751
rect 32597 18717 32631 18751
rect 33149 18717 33183 18751
rect 33333 18717 33367 18751
rect 33425 18717 33459 18751
rect 33517 18717 33551 18751
rect 34069 18717 34103 18751
rect 34253 18717 34287 18751
rect 34345 18717 34379 18751
rect 34529 18717 34563 18751
rect 37381 18717 37415 18751
rect 7849 18649 7883 18683
rect 13553 18649 13587 18683
rect 13753 18649 13787 18683
rect 17141 18649 17175 18683
rect 19993 18649 20027 18683
rect 32505 18649 32539 18683
rect 2329 18581 2363 18615
rect 3801 18581 3835 18615
rect 5641 18581 5675 18615
rect 8309 18581 8343 18615
rect 9505 18581 9539 18615
rect 9965 18581 9999 18615
rect 10517 18581 10551 18615
rect 12357 18581 12391 18615
rect 13369 18581 13403 18615
rect 13921 18581 13955 18615
rect 19073 18581 19107 18615
rect 21465 18581 21499 18615
rect 28641 18581 28675 18615
rect 28917 18581 28951 18615
rect 29285 18581 29319 18615
rect 4077 18377 4111 18411
rect 5457 18377 5491 18411
rect 14657 18377 14691 18411
rect 19717 18377 19751 18411
rect 22201 18377 22235 18411
rect 25421 18377 25455 18411
rect 26065 18377 26099 18411
rect 33793 18377 33827 18411
rect 1869 18309 1903 18343
rect 18613 18309 18647 18343
rect 19349 18309 19383 18343
rect 19441 18309 19475 18343
rect 20545 18309 20579 18343
rect 1593 18241 1627 18275
rect 3617 18241 3651 18275
rect 7849 18241 7883 18275
rect 8401 18241 8435 18275
rect 10241 18241 10275 18275
rect 10425 18241 10459 18275
rect 14289 18241 14323 18275
rect 14473 18241 14507 18275
rect 16313 18241 16347 18275
rect 16865 18241 16899 18275
rect 17233 18241 17267 18275
rect 19165 18241 19199 18275
rect 19533 18241 19567 18275
rect 21281 18241 21315 18275
rect 21833 18241 21867 18275
rect 22017 18241 22051 18275
rect 23029 18241 23063 18275
rect 25329 18241 25363 18275
rect 26985 18241 27019 18275
rect 28733 18241 28767 18275
rect 30665 18241 30699 18275
rect 32229 18241 32263 18275
rect 32321 18241 32355 18275
rect 33333 18241 33367 18275
rect 33609 18241 33643 18275
rect 4169 18173 4203 18207
rect 4353 18173 4387 18207
rect 5549 18173 5583 18207
rect 5641 18173 5675 18207
rect 15853 18173 15887 18207
rect 16221 18173 16255 18207
rect 16957 18173 16991 18207
rect 17141 18173 17175 18207
rect 17877 18173 17911 18207
rect 21189 18173 21223 18207
rect 29009 18173 29043 18207
rect 31033 18173 31067 18207
rect 33701 18173 33735 18207
rect 24317 18105 24351 18139
rect 25697 18105 25731 18139
rect 25789 18105 25823 18139
rect 33425 18105 33459 18139
rect 3709 18037 3743 18071
rect 5089 18037 5123 18071
rect 10241 18037 10275 18071
rect 14289 18037 14323 18071
rect 16497 18037 16531 18071
rect 18889 18037 18923 18071
rect 21465 18037 21499 18071
rect 25605 18037 25639 18071
rect 27169 18037 27203 18071
rect 30481 18037 30515 18071
rect 32505 18037 32539 18071
rect 10885 17833 10919 17867
rect 17601 17833 17635 17867
rect 19073 17833 19107 17867
rect 21741 17833 21775 17867
rect 28733 17833 28767 17867
rect 29193 17833 29227 17867
rect 30941 17833 30975 17867
rect 12633 17765 12667 17799
rect 21649 17765 21683 17799
rect 26617 17765 26651 17799
rect 5089 17697 5123 17731
rect 16681 17697 16715 17731
rect 20361 17697 20395 17731
rect 20637 17697 20671 17731
rect 24409 17697 24443 17731
rect 25145 17697 25179 17731
rect 25237 17697 25271 17731
rect 27077 17697 27111 17731
rect 29745 17697 29779 17731
rect 30389 17697 30423 17731
rect 4813 17629 4847 17663
rect 7113 17629 7147 17663
rect 7205 17629 7239 17663
rect 10241 17629 10275 17663
rect 10425 17629 10459 17663
rect 10517 17629 10551 17663
rect 10609 17629 10643 17663
rect 12173 17629 12207 17663
rect 12265 17629 12299 17663
rect 12449 17629 12483 17663
rect 14749 17629 14783 17663
rect 14933 17629 14967 17663
rect 15393 17629 15427 17663
rect 15485 17629 15519 17663
rect 16313 17629 16347 17663
rect 16405 17629 16439 17663
rect 16773 17629 16807 17663
rect 17233 17629 17267 17663
rect 17877 17629 17911 17663
rect 17969 17629 18003 17663
rect 18061 17629 18095 17663
rect 18245 17629 18279 17663
rect 18797 17629 18831 17663
rect 18889 17629 18923 17663
rect 19257 17629 19291 17663
rect 19625 17629 19659 17663
rect 19993 17629 20027 17663
rect 20821 17629 20855 17663
rect 21097 17629 21131 17663
rect 21925 17629 21959 17663
rect 22443 17629 22477 17663
rect 22569 17629 22603 17663
rect 22661 17629 22695 17663
rect 22846 17607 22880 17641
rect 23121 17629 23155 17663
rect 23489 17629 23523 17663
rect 24501 17629 24535 17663
rect 25329 17629 25363 17663
rect 25605 17629 25639 17663
rect 25697 17629 25731 17663
rect 26525 17629 26559 17663
rect 26801 17629 26835 17663
rect 28917 17629 28951 17663
rect 29009 17629 29043 17663
rect 29285 17629 29319 17663
rect 30573 17629 30607 17663
rect 30757 17629 30791 17663
rect 5365 17561 5399 17595
rect 8033 17561 8067 17595
rect 16037 17561 16071 17595
rect 18337 17561 18371 17595
rect 21465 17561 21499 17595
rect 22201 17561 22235 17595
rect 22937 17561 22971 17595
rect 24777 17561 24811 17595
rect 24863 17561 24897 17595
rect 4629 17493 4663 17527
rect 17141 17493 17175 17527
rect 24685 17493 24719 17527
rect 25513 17493 25547 17527
rect 25973 17493 26007 17527
rect 28549 17493 28583 17527
rect 11897 17289 11931 17323
rect 12541 17289 12575 17323
rect 13185 17289 13219 17323
rect 15577 17289 15611 17323
rect 19165 17289 19199 17323
rect 20821 17289 20855 17323
rect 21189 17289 21223 17323
rect 24685 17289 24719 17323
rect 25329 17289 25363 17323
rect 26985 17289 27019 17323
rect 27445 17289 27479 17323
rect 30573 17289 30607 17323
rect 4353 17221 4387 17255
rect 7205 17221 7239 17255
rect 12081 17221 12115 17255
rect 12265 17221 12299 17255
rect 12449 17221 12483 17255
rect 14013 17221 14047 17255
rect 30113 17221 30147 17255
rect 35173 17221 35207 17255
rect 3157 17153 3191 17187
rect 4077 17153 4111 17187
rect 6377 17153 6411 17187
rect 7941 17153 7975 17187
rect 8769 17153 8803 17187
rect 8861 17153 8895 17187
rect 9229 17153 9263 17187
rect 9689 17153 9723 17187
rect 10241 17153 10275 17187
rect 10333 17153 10367 17187
rect 10793 17153 10827 17187
rect 10977 17153 11011 17187
rect 11989 17153 12023 17187
rect 13737 17153 13771 17187
rect 13921 17153 13955 17187
rect 14110 17153 14144 17187
rect 15579 17153 15613 17187
rect 16681 17153 16715 17187
rect 16774 17153 16808 17187
rect 16957 17153 16991 17187
rect 17049 17153 17083 17187
rect 17146 17153 17180 17187
rect 18889 17153 18923 17187
rect 18981 17153 19015 17187
rect 20453 17153 20487 17187
rect 21281 17153 21315 17187
rect 22477 17153 22511 17187
rect 22845 17153 22879 17187
rect 24133 17153 24167 17187
rect 24225 17153 24259 17187
rect 24317 17153 24351 17187
rect 24961 17153 24995 17187
rect 25421 17153 25455 17187
rect 27353 17153 27387 17187
rect 30205 17153 30239 17187
rect 30665 17153 30699 17187
rect 33425 17153 33459 17187
rect 33701 17153 33735 17187
rect 34345 17153 34379 17187
rect 5825 17085 5859 17119
rect 10609 17085 10643 17119
rect 10701 17085 10735 17119
rect 11529 17085 11563 17119
rect 12725 17085 12759 17119
rect 12817 17085 12851 17119
rect 15117 17085 15151 17119
rect 18705 17085 18739 17119
rect 18797 17085 18831 17119
rect 20545 17085 20579 17119
rect 20913 17085 20947 17119
rect 21097 17085 21131 17119
rect 22293 17085 22327 17119
rect 22753 17085 22787 17119
rect 23489 17085 23523 17119
rect 23857 17085 23891 17119
rect 25145 17085 25179 17119
rect 27537 17085 27571 17119
rect 29929 17085 29963 17119
rect 33977 17085 34011 17119
rect 9413 17017 9447 17051
rect 11713 17017 11747 17051
rect 21005 17017 21039 17051
rect 24593 17017 24627 17051
rect 25053 17017 25087 17051
rect 2973 16949 3007 16983
rect 10057 16949 10091 16983
rect 10793 16949 10827 16983
rect 14289 16949 14323 16983
rect 15209 16949 15243 16983
rect 15761 16949 15795 16983
rect 17325 16949 17359 16983
rect 20453 16949 20487 16983
rect 23949 16949 23983 16983
rect 30849 16949 30883 16983
rect 33241 16949 33275 16983
rect 12357 16745 12391 16779
rect 17141 16745 17175 16779
rect 26985 16745 27019 16779
rect 30928 16745 30962 16779
rect 32413 16745 32447 16779
rect 17325 16677 17359 16711
rect 22569 16677 22603 16711
rect 1869 16609 1903 16643
rect 2145 16609 2179 16643
rect 4905 16609 4939 16643
rect 6929 16609 6963 16643
rect 7297 16609 7331 16643
rect 8217 16609 8251 16643
rect 8309 16609 8343 16643
rect 14289 16609 14323 16643
rect 18153 16609 18187 16643
rect 21833 16609 21867 16643
rect 32965 16609 32999 16643
rect 6837 16541 6871 16575
rect 7849 16541 7883 16575
rect 8953 16541 8987 16575
rect 9137 16541 9171 16575
rect 9505 16541 9539 16575
rect 9653 16541 9687 16575
rect 9873 16541 9907 16575
rect 10011 16541 10045 16575
rect 10604 16541 10638 16575
rect 10701 16541 10735 16575
rect 10976 16541 11010 16575
rect 11069 16541 11103 16575
rect 12265 16541 12299 16575
rect 12449 16541 12483 16575
rect 13553 16541 13587 16575
rect 14381 16541 14415 16575
rect 14752 16541 14786 16575
rect 17417 16541 17451 16575
rect 17693 16541 17727 16575
rect 18705 16541 18739 16575
rect 22108 16541 22142 16575
rect 22201 16541 22235 16575
rect 22293 16541 22327 16575
rect 22477 16541 22511 16575
rect 22844 16541 22878 16575
rect 22937 16541 22971 16575
rect 23029 16541 23063 16575
rect 23213 16541 23247 16575
rect 25973 16541 26007 16575
rect 26341 16541 26375 16575
rect 30389 16541 30423 16575
rect 30481 16541 30515 16575
rect 30665 16541 30699 16575
rect 32689 16541 32723 16575
rect 4169 16473 4203 16507
rect 7757 16473 7791 16507
rect 9781 16473 9815 16507
rect 10793 16473 10827 16507
rect 13737 16473 13771 16507
rect 16957 16473 16991 16507
rect 17173 16473 17207 16507
rect 17785 16473 17819 16507
rect 18429 16473 18463 16507
rect 26157 16473 26191 16507
rect 26249 16473 26283 16507
rect 26617 16473 26651 16507
rect 26801 16473 26835 16507
rect 3617 16405 3651 16439
rect 6377 16405 6411 16439
rect 6745 16405 6779 16439
rect 9137 16405 9171 16439
rect 10149 16405 10183 16439
rect 10425 16405 10459 16439
rect 13921 16405 13955 16439
rect 14749 16405 14783 16439
rect 14933 16405 14967 16439
rect 17601 16405 17635 16439
rect 26525 16405 26559 16439
rect 34437 16405 34471 16439
rect 1961 16201 1995 16235
rect 7849 16201 7883 16235
rect 8585 16201 8619 16235
rect 10241 16201 10275 16235
rect 19717 16201 19751 16235
rect 22569 16201 22603 16235
rect 25237 16201 25271 16235
rect 26433 16201 26467 16235
rect 32873 16201 32907 16235
rect 33241 16201 33275 16235
rect 33609 16201 33643 16235
rect 1409 16133 1443 16167
rect 1777 16133 1811 16167
rect 9689 16133 9723 16167
rect 9781 16133 9815 16167
rect 30113 16133 30147 16167
rect 30205 16133 30239 16167
rect 31033 16133 31067 16167
rect 33701 16133 33735 16167
rect 2145 16065 2179 16099
rect 3893 16065 3927 16099
rect 5457 16065 5491 16099
rect 7205 16065 7239 16099
rect 7297 16065 7331 16099
rect 7665 16065 7699 16099
rect 8401 16065 8435 16099
rect 9572 16065 9606 16099
rect 9909 16065 9943 16099
rect 10057 16065 10091 16099
rect 10149 16065 10183 16099
rect 10425 16065 10459 16099
rect 10609 16065 10643 16099
rect 12357 16065 12391 16099
rect 12541 16065 12575 16099
rect 12725 16065 12759 16099
rect 12817 16065 12851 16099
rect 13185 16065 13219 16099
rect 13369 16065 13403 16099
rect 14381 16065 14415 16099
rect 14933 16065 14967 16099
rect 15761 16065 15795 16099
rect 16037 16065 16071 16099
rect 16497 16065 16531 16099
rect 17233 16065 17267 16099
rect 17509 16065 17543 16099
rect 18061 16065 18095 16099
rect 18797 16065 18831 16099
rect 19655 16065 19689 16099
rect 20448 16065 20482 16099
rect 20545 16065 20579 16099
rect 20637 16065 20671 16099
rect 20820 16065 20854 16099
rect 20913 16065 20947 16099
rect 22109 16065 22143 16099
rect 22201 16065 22235 16099
rect 22385 16065 22419 16099
rect 24041 16065 24075 16099
rect 24189 16065 24223 16099
rect 24317 16065 24351 16099
rect 24409 16065 24443 16099
rect 24506 16065 24540 16099
rect 24777 16065 24811 16099
rect 24869 16065 24903 16099
rect 25053 16065 25087 16099
rect 25789 16065 25823 16099
rect 25937 16065 25971 16099
rect 26065 16065 26099 16099
rect 26157 16065 26191 16099
rect 26254 16065 26288 16099
rect 27905 16065 27939 16099
rect 28641 16065 28675 16099
rect 29101 16065 29135 16099
rect 29561 16065 29595 16099
rect 29837 16065 29871 16099
rect 29985 16065 30019 16099
rect 30343 16065 30377 16099
rect 30849 16065 30883 16099
rect 32965 16065 32999 16099
rect 7941 15997 7975 16031
rect 8309 15997 8343 16031
rect 13829 15997 13863 16031
rect 14197 15997 14231 16031
rect 14749 15997 14783 16031
rect 18521 15997 18555 16031
rect 20177 15997 20211 16031
rect 27997 15997 28031 16031
rect 30573 15997 30607 16031
rect 33885 15997 33919 16031
rect 12449 15929 12483 15963
rect 14657 15929 14691 15963
rect 15853 15929 15887 15963
rect 18153 15929 18187 15963
rect 19533 15929 19567 15963
rect 20085 15929 20119 15963
rect 20269 15929 20303 15963
rect 29561 15929 29595 15963
rect 4077 15861 4111 15895
rect 5273 15861 5307 15895
rect 7665 15861 7699 15895
rect 9413 15861 9447 15895
rect 15209 15861 15243 15895
rect 24685 15861 24719 15895
rect 27905 15861 27939 15895
rect 28273 15861 28307 15895
rect 30481 15861 30515 15895
rect 30665 15861 30699 15895
rect 9781 15657 9815 15691
rect 11253 15657 11287 15691
rect 12357 15657 12391 15691
rect 12817 15657 12851 15691
rect 12909 15657 12943 15691
rect 21557 15657 21591 15691
rect 22293 15657 22327 15691
rect 22477 15657 22511 15691
rect 26157 15657 26191 15691
rect 26893 15657 26927 15691
rect 29101 15657 29135 15691
rect 30113 15657 30147 15691
rect 13093 15589 13127 15623
rect 16221 15589 16255 15623
rect 18061 15589 18095 15623
rect 19809 15589 19843 15623
rect 20453 15589 20487 15623
rect 28457 15589 28491 15623
rect 28825 15589 28859 15623
rect 4997 15521 5031 15555
rect 6745 15521 6779 15555
rect 9873 15521 9907 15555
rect 12909 15521 12943 15555
rect 14197 15521 14231 15555
rect 17233 15521 17267 15555
rect 18521 15521 18555 15555
rect 22569 15521 22603 15555
rect 25421 15521 25455 15555
rect 27169 15521 27203 15555
rect 4445 15453 4479 15487
rect 4537 15453 4571 15487
rect 4721 15453 4755 15487
rect 7481 15453 7515 15487
rect 7941 15453 7975 15487
rect 10057 15453 10091 15487
rect 11437 15453 11471 15487
rect 11529 15453 11563 15487
rect 11713 15453 11747 15487
rect 11897 15453 11931 15487
rect 11989 15453 12023 15487
rect 12081 15453 12115 15487
rect 12725 15453 12759 15487
rect 14289 15453 14323 15487
rect 14657 15453 14691 15487
rect 15393 15453 15427 15487
rect 15761 15453 15795 15487
rect 16037 15453 16071 15487
rect 16497 15453 16531 15487
rect 17509 15453 17543 15487
rect 18061 15453 18095 15487
rect 18245 15453 18279 15487
rect 18889 15453 18923 15487
rect 19257 15453 19291 15487
rect 19441 15453 19475 15487
rect 19533 15453 19567 15487
rect 19625 15453 19659 15487
rect 19901 15453 19935 15487
rect 20177 15453 20211 15487
rect 20269 15453 20303 15487
rect 20913 15453 20947 15487
rect 21006 15453 21040 15487
rect 21281 15453 21315 15487
rect 21419 15453 21453 15487
rect 22661 15453 22695 15487
rect 24869 15453 24903 15487
rect 25513 15453 25547 15487
rect 25606 15453 25640 15487
rect 25881 15453 25915 15487
rect 26019 15453 26053 15487
rect 26249 15453 26283 15487
rect 26433 15453 26467 15487
rect 26525 15453 26559 15487
rect 26617 15453 26651 15487
rect 27537 15453 27571 15487
rect 27721 15453 27755 15487
rect 27813 15453 27847 15487
rect 27906 15453 27940 15487
rect 28181 15453 28215 15487
rect 28278 15453 28312 15487
rect 28641 15453 28675 15487
rect 28733 15453 28767 15487
rect 28917 15453 28951 15487
rect 29561 15453 29595 15487
rect 29837 15453 29871 15487
rect 29929 15453 29963 15487
rect 30573 15453 30607 15487
rect 30849 15453 30883 15487
rect 33609 15453 33643 15487
rect 9781 15385 9815 15419
rect 15117 15385 15151 15419
rect 16405 15385 16439 15419
rect 16957 15385 16991 15419
rect 20085 15385 20119 15419
rect 20729 15385 20763 15419
rect 21189 15385 21223 15419
rect 25053 15385 25087 15419
rect 25789 15385 25823 15419
rect 27445 15385 27479 15419
rect 28089 15385 28123 15419
rect 29745 15385 29779 15419
rect 31125 15385 31159 15419
rect 7389 15317 7423 15351
rect 7757 15317 7791 15351
rect 10241 15317 10275 15351
rect 18981 15317 19015 15351
rect 20637 15317 20671 15351
rect 25145 15317 25179 15351
rect 25237 15317 25271 15351
rect 27353 15317 27387 15351
rect 30757 15317 30791 15351
rect 32597 15317 32631 15351
rect 33517 15317 33551 15351
rect 1777 15113 1811 15147
rect 9137 15113 9171 15147
rect 9505 15113 9539 15147
rect 11989 15113 12023 15147
rect 15025 15113 15059 15147
rect 20269 15113 20303 15147
rect 25421 15113 25455 15147
rect 26525 15113 26559 15147
rect 28641 15113 28675 15147
rect 30757 15113 30791 15147
rect 31033 15113 31067 15147
rect 33241 15113 33275 15147
rect 7481 15045 7515 15079
rect 15393 15045 15427 15079
rect 17417 15045 17451 15079
rect 18705 15045 18739 15079
rect 18797 15045 18831 15079
rect 19901 15045 19935 15079
rect 20821 15045 20855 15079
rect 20913 15045 20947 15079
rect 24501 15045 24535 15079
rect 25053 15045 25087 15079
rect 25145 15045 25179 15079
rect 28273 15045 28307 15079
rect 29101 15045 29135 15079
rect 33609 15045 33643 15079
rect 1961 14977 1995 15011
rect 10241 14977 10275 15011
rect 12173 14977 12207 15011
rect 12265 14977 12299 15011
rect 12449 14977 12483 15011
rect 12541 14977 12575 15011
rect 14749 14977 14783 15011
rect 14933 14977 14967 15011
rect 15209 14977 15243 15011
rect 15485 14977 15519 15011
rect 17141 14977 17175 15011
rect 17234 14977 17268 15011
rect 17509 14977 17543 15011
rect 17647 14977 17681 15011
rect 17877 14977 17911 15011
rect 17969 14977 18003 15011
rect 18153 14977 18187 15011
rect 18429 14977 18463 15011
rect 18521 14977 18555 15011
rect 18889 14977 18923 15011
rect 19625 14977 19659 15011
rect 19783 14977 19817 15011
rect 19993 14977 20027 15011
rect 20085 14977 20119 15011
rect 20545 14977 20579 15011
rect 20637 14977 20671 15011
rect 21005 14977 21039 15011
rect 22017 14977 22051 15011
rect 23397 14977 23431 15011
rect 24225 14977 24259 15011
rect 24409 14977 24443 15011
rect 24593 14977 24627 15011
rect 24869 14977 24903 15011
rect 25237 14977 25271 15011
rect 25963 14977 25997 15011
rect 26065 14977 26099 15011
rect 26249 14977 26283 15011
rect 26341 14977 26375 15011
rect 28089 14977 28123 15011
rect 28365 14977 28399 15011
rect 28457 14977 28491 15011
rect 28733 14977 28767 15011
rect 28917 14977 28951 15011
rect 30389 14977 30423 15011
rect 31125 14977 31159 15011
rect 33057 14977 33091 15011
rect 7205 14909 7239 14943
rect 8953 14909 8987 14943
rect 9597 14909 9631 14943
rect 9689 14909 9723 14943
rect 10425 14909 10459 14943
rect 15945 14909 15979 14943
rect 18981 14909 19015 14943
rect 21833 14909 21867 14943
rect 30113 14909 30147 14943
rect 30297 14909 30331 14943
rect 33333 14909 33367 14943
rect 17785 14841 17819 14875
rect 18337 14841 18371 14875
rect 20545 14841 20579 14875
rect 22201 14773 22235 14807
rect 23213 14773 23247 14807
rect 24777 14773 24811 14807
rect 35081 14773 35115 14807
rect 4169 14569 4203 14603
rect 12541 14569 12575 14603
rect 18153 14569 18187 14603
rect 21741 14569 21775 14603
rect 24225 14569 24259 14603
rect 32873 14569 32907 14603
rect 33241 14569 33275 14603
rect 37841 14569 37875 14603
rect 10057 14501 10091 14535
rect 6377 14433 6411 14467
rect 7021 14433 7055 14467
rect 7205 14433 7239 14467
rect 8033 14433 8067 14467
rect 8217 14433 8251 14467
rect 20177 14433 20211 14467
rect 22753 14433 22787 14467
rect 33793 14433 33827 14467
rect 4353 14365 4387 14399
rect 4537 14365 4571 14399
rect 4629 14365 4663 14399
rect 6929 14365 6963 14399
rect 9873 14365 9907 14399
rect 10517 14365 10551 14399
rect 11161 14365 11195 14399
rect 11989 14365 12023 14399
rect 12265 14365 12299 14399
rect 12357 14365 12391 14399
rect 15025 14365 15059 14399
rect 17785 14365 17819 14399
rect 17877 14365 17911 14399
rect 17969 14365 18003 14399
rect 20049 14359 20083 14393
rect 20269 14365 20303 14399
rect 21005 14365 21039 14399
rect 21373 14365 21407 14399
rect 21925 14365 21959 14399
rect 22017 14365 22051 14399
rect 22477 14365 22511 14399
rect 27721 14365 27755 14399
rect 28273 14365 28307 14399
rect 30849 14365 30883 14399
rect 30941 14365 30975 14399
rect 31125 14365 31159 14399
rect 35357 14365 35391 14399
rect 37657 14365 37691 14399
rect 4905 14297 4939 14331
rect 7941 14297 7975 14331
rect 12173 14297 12207 14331
rect 17601 14297 17635 14331
rect 20177 14297 20211 14331
rect 20453 14297 20487 14331
rect 21189 14297 21223 14331
rect 21281 14297 21315 14331
rect 21741 14297 21775 14331
rect 31401 14297 31435 14331
rect 6561 14229 6595 14263
rect 7573 14229 7607 14263
rect 14933 14229 14967 14263
rect 21557 14229 21591 14263
rect 22201 14229 22235 14263
rect 27813 14229 27847 14263
rect 33609 14229 33643 14263
rect 33701 14229 33735 14263
rect 35449 14229 35483 14263
rect 4813 14025 4847 14059
rect 5181 14025 5215 14059
rect 11897 14025 11931 14059
rect 13921 14025 13955 14059
rect 14289 14025 14323 14059
rect 19441 14025 19475 14059
rect 21833 14025 21867 14059
rect 22661 14025 22695 14059
rect 23397 14025 23431 14059
rect 23765 14025 23799 14059
rect 31401 14025 31435 14059
rect 32137 14025 32171 14059
rect 32505 14025 32539 14059
rect 32597 14025 32631 14059
rect 1777 13957 1811 13991
rect 11161 13957 11195 13991
rect 14381 13957 14415 13991
rect 17509 13957 17543 13991
rect 19165 13957 19199 13991
rect 21465 13957 21499 13991
rect 22201 13957 22235 13991
rect 23857 13957 23891 13991
rect 29929 13957 29963 13991
rect 4905 13889 4939 13923
rect 5365 13889 5399 13923
rect 7481 13889 7515 13923
rect 9873 13889 9907 13923
rect 10057 13889 10091 13923
rect 10149 13889 10183 13923
rect 10333 13889 10367 13923
rect 10885 13889 10919 13923
rect 12173 13889 12207 13923
rect 12265 13889 12299 13923
rect 12357 13889 12391 13923
rect 12541 13889 12575 13923
rect 13737 13889 13771 13923
rect 14749 13889 14783 13923
rect 17784 13889 17818 13923
rect 17877 13889 17911 13923
rect 17969 13889 18003 13923
rect 18153 13889 18187 13923
rect 18889 13889 18923 13923
rect 19073 13889 19107 13923
rect 19257 13889 19291 13923
rect 21097 13889 21131 13923
rect 21281 13889 21315 13923
rect 22017 13889 22051 13923
rect 22109 13889 22143 13923
rect 22385 13889 22419 13923
rect 22753 13889 22787 13923
rect 27537 13889 27571 13923
rect 29699 13889 29733 13923
rect 29837 13889 29871 13923
rect 30113 13889 30147 13923
rect 31585 13889 31619 13923
rect 35357 13889 35391 13923
rect 1501 13821 1535 13855
rect 10701 13821 10735 13855
rect 14473 13821 14507 13855
rect 23949 13821 23983 13855
rect 27629 13821 27663 13855
rect 32689 13821 32723 13855
rect 33609 13821 33643 13855
rect 10609 13753 10643 13787
rect 7297 13685 7331 13719
rect 10057 13685 10091 13719
rect 13553 13685 13587 13719
rect 15012 13685 15046 13719
rect 16497 13685 16531 13719
rect 27537 13685 27571 13719
rect 27905 13685 27939 13719
rect 29561 13685 29595 13719
rect 35093 13685 35127 13719
rect 8493 13481 8527 13515
rect 9873 13481 9907 13515
rect 12817 13481 12851 13515
rect 15209 13481 15243 13515
rect 17969 13481 18003 13515
rect 26249 13481 26283 13515
rect 27261 13481 27295 13515
rect 31125 13481 31159 13515
rect 33241 13481 33275 13515
rect 10517 13413 10551 13447
rect 12633 13413 12667 13447
rect 15577 13413 15611 13447
rect 17877 13413 17911 13447
rect 26893 13413 26927 13447
rect 27997 13413 28031 13447
rect 28365 13413 28399 13447
rect 30297 13413 30331 13447
rect 33333 13413 33367 13447
rect 5457 13345 5491 13379
rect 7021 13345 7055 13379
rect 11345 13345 11379 13379
rect 16129 13345 16163 13379
rect 20085 13345 20119 13379
rect 20177 13345 20211 13379
rect 28273 13345 28307 13379
rect 30205 13345 30239 13379
rect 33793 13345 33827 13379
rect 33885 13345 33919 13379
rect 3985 13277 4019 13311
rect 5273 13277 5307 13311
rect 6469 13277 6503 13311
rect 6561 13277 6595 13311
rect 6745 13277 6779 13311
rect 9597 13277 9631 13311
rect 9781 13277 9815 13311
rect 10057 13277 10091 13311
rect 10241 13277 10275 13311
rect 10701 13277 10735 13311
rect 10885 13277 10919 13311
rect 11253 13277 11287 13311
rect 11897 13277 11931 13311
rect 11989 13277 12023 13311
rect 12633 13277 12667 13311
rect 13001 13277 13035 13311
rect 13093 13277 13127 13311
rect 13277 13277 13311 13311
rect 13369 13277 13403 13311
rect 13645 13277 13679 13311
rect 15393 13277 15427 13311
rect 15945 13277 15979 13311
rect 17233 13277 17267 13311
rect 17326 13277 17360 13311
rect 17509 13277 17543 13311
rect 17698 13277 17732 13311
rect 18153 13277 18187 13311
rect 18429 13277 18463 13311
rect 20637 13277 20671 13311
rect 24685 13277 24719 13311
rect 24961 13277 24995 13311
rect 25053 13277 25087 13311
rect 25605 13277 25639 13311
rect 25698 13277 25732 13311
rect 25973 13277 26007 13311
rect 26070 13277 26104 13311
rect 26341 13277 26375 13311
rect 26709 13277 26743 13311
rect 26985 13277 27019 13311
rect 27169 13277 27203 13311
rect 27813 13277 27847 13311
rect 27905 13277 27939 13311
rect 28089 13277 28123 13311
rect 28549 13277 28583 13311
rect 28641 13277 28675 13311
rect 28917 13277 28951 13311
rect 29929 13277 29963 13311
rect 30297 13277 30331 13311
rect 30665 13277 30699 13311
rect 31309 13277 31343 13311
rect 31401 13277 31435 13311
rect 31493 13277 31527 13311
rect 31585 13277 31619 13311
rect 31769 13277 31803 13311
rect 32229 13277 32263 13311
rect 33057 13277 33091 13311
rect 5365 13209 5399 13243
rect 10609 13209 10643 13243
rect 13553 13209 13587 13243
rect 16037 13209 16071 13243
rect 17601 13209 17635 13243
rect 19993 13209 20027 13243
rect 24869 13209 24903 13243
rect 25881 13209 25915 13243
rect 26525 13209 26559 13243
rect 26617 13209 26651 13243
rect 28733 13209 28767 13243
rect 3893 13141 3927 13175
rect 4905 13141 4939 13175
rect 18337 13141 18371 13175
rect 19625 13141 19659 13175
rect 20545 13141 20579 13175
rect 25237 13141 25271 13175
rect 31953 13141 31987 13175
rect 32321 13141 32355 13175
rect 33701 13141 33735 13175
rect 9781 12937 9815 12971
rect 12725 12937 12759 12971
rect 14749 12937 14783 12971
rect 19533 12937 19567 12971
rect 21373 12937 21407 12971
rect 27905 12937 27939 12971
rect 28365 12937 28399 12971
rect 29929 12937 29963 12971
rect 31953 12937 31987 12971
rect 5549 12869 5583 12903
rect 9137 12869 9171 12903
rect 12357 12869 12391 12903
rect 13277 12869 13311 12903
rect 19901 12869 19935 12903
rect 24869 12869 24903 12903
rect 26525 12869 26559 12903
rect 27997 12869 28031 12903
rect 3525 12801 3559 12835
rect 8493 12801 8527 12835
rect 8677 12801 8711 12835
rect 8861 12801 8895 12835
rect 8953 12801 8987 12835
rect 9045 12801 9079 12835
rect 9229 12801 9263 12835
rect 9505 12801 9539 12835
rect 9873 12801 9907 12835
rect 10149 12801 10183 12835
rect 10333 12801 10367 12835
rect 10793 12801 10827 12835
rect 12173 12801 12207 12835
rect 12449 12801 12483 12835
rect 12541 12801 12575 12835
rect 13001 12801 13035 12835
rect 19349 12801 19383 12835
rect 22293 12801 22327 12835
rect 24593 12801 24627 12835
rect 24686 12801 24720 12835
rect 24961 12801 24995 12835
rect 25058 12801 25092 12835
rect 25329 12801 25363 12835
rect 25605 12801 25639 12835
rect 26295 12801 26329 12835
rect 26433 12801 26467 12835
rect 26653 12801 26687 12835
rect 26801 12801 26835 12835
rect 27261 12801 27295 12835
rect 27354 12801 27388 12835
rect 27537 12801 27571 12835
rect 27629 12801 27663 12835
rect 27767 12801 27801 12835
rect 28181 12801 28215 12835
rect 29377 12801 29411 12835
rect 29469 12801 29503 12835
rect 29580 12801 29614 12835
rect 29745 12801 29779 12835
rect 31585 12801 31619 12835
rect 32137 12801 32171 12835
rect 3801 12733 3835 12767
rect 9321 12733 9355 12767
rect 10977 12733 11011 12767
rect 19625 12733 19659 12767
rect 25513 12733 25547 12767
rect 25697 12733 25731 12767
rect 25789 12733 25823 12767
rect 25973 12733 26007 12767
rect 31309 12733 31343 12767
rect 31493 12733 31527 12767
rect 32413 12733 32447 12767
rect 8585 12665 8619 12699
rect 25237 12665 25271 12699
rect 26157 12665 26191 12699
rect 23581 12597 23615 12631
rect 33885 12597 33919 12631
rect 4169 12393 4203 12427
rect 16589 12393 16623 12427
rect 16865 12393 16899 12427
rect 22109 12393 22143 12427
rect 27077 12393 27111 12427
rect 31769 12393 31803 12427
rect 18061 12325 18095 12359
rect 23581 12325 23615 12359
rect 24961 12325 24995 12359
rect 25053 12325 25087 12359
rect 25605 12325 25639 12359
rect 27629 12325 27663 12359
rect 15853 12257 15887 12291
rect 33425 12257 33459 12291
rect 33517 12257 33551 12291
rect 4353 12189 4387 12223
rect 4905 12189 4939 12223
rect 4997 12189 5031 12223
rect 5181 12189 5215 12223
rect 9873 12189 9907 12223
rect 10149 12189 10183 12223
rect 10793 12189 10827 12223
rect 10885 12189 10919 12223
rect 11253 12189 11287 12223
rect 11345 12189 11379 12223
rect 12541 12189 12575 12223
rect 15209 12189 15243 12223
rect 15393 12189 15427 12223
rect 15485 12189 15519 12223
rect 15577 12189 15611 12223
rect 15945 12189 15979 12223
rect 16037 12189 16071 12223
rect 16313 12189 16347 12223
rect 16405 12189 16439 12223
rect 16957 12189 16991 12223
rect 17049 12189 17083 12223
rect 18336 12189 18370 12223
rect 18429 12189 18463 12223
rect 18521 12189 18555 12223
rect 18705 12189 18739 12223
rect 22385 12189 22419 12223
rect 22569 12189 22603 12223
rect 23673 12189 23707 12223
rect 24409 12189 24443 12223
rect 24685 12189 24719 12223
rect 24777 12189 24811 12223
rect 27353 12189 27387 12223
rect 27445 12189 27479 12223
rect 29745 12189 29779 12223
rect 29837 12189 29871 12223
rect 30021 12189 30055 12223
rect 34069 12189 34103 12223
rect 34345 12189 34379 12223
rect 5457 12121 5491 12155
rect 7205 12121 7239 12155
rect 16221 12121 16255 12155
rect 21925 12121 21959 12155
rect 24593 12121 24627 12155
rect 25421 12121 25455 12155
rect 27261 12121 27295 12155
rect 30297 12121 30331 12155
rect 33609 12121 33643 12155
rect 12449 12053 12483 12087
rect 16681 12053 16715 12087
rect 22109 12053 22143 12087
rect 25237 12053 25271 12087
rect 25329 12053 25363 12087
rect 33977 12053 34011 12087
rect 34161 12053 34195 12087
rect 34529 12053 34563 12087
rect 1961 11849 1995 11883
rect 5641 11849 5675 11883
rect 6837 11849 6871 11883
rect 9873 11849 9907 11883
rect 11253 11849 11287 11883
rect 14013 11849 14047 11883
rect 18613 11849 18647 11883
rect 22477 11849 22511 11883
rect 24409 11849 24443 11883
rect 24961 11849 24995 11883
rect 30113 11849 30147 11883
rect 1777 11781 1811 11815
rect 6745 11781 6779 11815
rect 9229 11781 9263 11815
rect 16129 11781 16163 11815
rect 16865 11781 16899 11815
rect 18153 11781 18187 11815
rect 18245 11781 18279 11815
rect 20821 11781 20855 11815
rect 21005 11781 21039 11815
rect 23673 11781 23707 11815
rect 23857 11781 23891 11815
rect 24225 11781 24259 11815
rect 24777 11781 24811 11815
rect 30757 11781 30791 11815
rect 34805 11781 34839 11815
rect 1409 11713 1443 11747
rect 2145 11713 2179 11747
rect 5825 11713 5859 11747
rect 7389 11713 7423 11747
rect 9045 11713 9079 11747
rect 9413 11713 9447 11747
rect 9689 11713 9723 11747
rect 10149 11713 10183 11747
rect 10793 11713 10827 11747
rect 11161 11713 11195 11747
rect 11529 11713 11563 11747
rect 12265 11713 12299 11747
rect 14289 11713 14323 11747
rect 15393 11713 15427 11747
rect 15485 11713 15519 11747
rect 15577 11713 15611 11747
rect 15853 11713 15887 11747
rect 17049 11713 17083 11747
rect 17877 11713 17911 11747
rect 18025 11713 18059 11747
rect 18342 11713 18376 11747
rect 18797 11713 18831 11747
rect 18981 11713 19015 11747
rect 19073 11713 19107 11747
rect 22845 11713 22879 11747
rect 23397 11713 23431 11747
rect 25237 11713 25271 11747
rect 29561 11713 29595 11747
rect 29745 11713 29779 11747
rect 29837 11713 29871 11747
rect 29929 11713 29963 11747
rect 31309 11713 31343 11747
rect 35081 11713 35115 11747
rect 37657 11713 37691 11747
rect 6929 11645 6963 11679
rect 8861 11645 8895 11679
rect 9965 11645 9999 11679
rect 10517 11645 10551 11679
rect 12541 11645 12575 11679
rect 14473 11645 14507 11679
rect 33333 11645 33367 11679
rect 6377 11577 6411 11611
rect 15761 11577 15795 11611
rect 37841 11577 37875 11611
rect 7205 11509 7239 11543
rect 11713 11509 11747 11543
rect 15209 11509 15243 11543
rect 16681 11509 16715 11543
rect 18521 11509 18555 11543
rect 21097 11509 21131 11543
rect 23857 11509 23891 11543
rect 24041 11509 24075 11543
rect 24409 11509 24443 11543
rect 24593 11509 24627 11543
rect 24961 11509 24995 11543
rect 4721 11305 4755 11339
rect 12817 11305 12851 11339
rect 14841 11305 14875 11339
rect 16773 11305 16807 11339
rect 17969 11305 18003 11339
rect 18889 11305 18923 11339
rect 26801 11305 26835 11339
rect 28365 11305 28399 11339
rect 29561 11305 29595 11339
rect 13185 11237 13219 11271
rect 15945 11237 15979 11271
rect 16957 11237 16991 11271
rect 20085 11237 20119 11271
rect 21741 11237 21775 11271
rect 23765 11237 23799 11271
rect 25329 11237 25363 11271
rect 28273 11237 28307 11271
rect 28733 11237 28767 11271
rect 7021 11169 7055 11203
rect 10885 11169 10919 11203
rect 13737 11169 13771 11203
rect 16221 11169 16255 11203
rect 16681 11169 16715 11203
rect 18337 11169 18371 11203
rect 18429 11169 18463 11203
rect 20729 11169 20763 11203
rect 26157 11169 26191 11203
rect 26341 11169 26375 11203
rect 28457 11169 28491 11203
rect 29929 11169 29963 11203
rect 30205 11169 30239 11203
rect 30389 11169 30423 11203
rect 4905 11101 4939 11135
rect 5089 11101 5123 11135
rect 6469 11101 6503 11135
rect 6561 11101 6595 11135
rect 6745 11101 6779 11135
rect 10149 11101 10183 11135
rect 10701 11101 10735 11135
rect 11897 11101 11931 11135
rect 11989 11101 12023 11135
rect 12173 11101 12207 11135
rect 12265 11101 12299 11135
rect 13001 11101 13035 11135
rect 13553 11101 13587 11135
rect 14197 11101 14231 11135
rect 14290 11101 14324 11135
rect 14703 11101 14737 11135
rect 15301 11101 15335 11135
rect 15394 11101 15428 11135
rect 15577 11101 15611 11135
rect 15669 11101 15703 11135
rect 15766 11101 15800 11135
rect 16037 11101 16071 11135
rect 16589 11101 16623 11135
rect 17325 11101 17359 11135
rect 17418 11101 17452 11135
rect 17790 11101 17824 11135
rect 18613 11101 18647 11135
rect 18705 11101 18739 11135
rect 19441 11101 19475 11135
rect 19809 11101 19843 11135
rect 20453 11101 20487 11135
rect 21005 11101 21039 11135
rect 21373 11101 21407 11135
rect 22201 11101 22235 11135
rect 22569 11101 22603 11135
rect 23109 11111 23143 11145
rect 23305 11101 23339 11135
rect 23397 11101 23431 11135
rect 23490 11079 23524 11113
rect 24777 11101 24811 11135
rect 24961 11101 24995 11135
rect 25145 11101 25179 11135
rect 25513 11101 25547 11135
rect 25697 11101 25731 11135
rect 25789 11101 25823 11135
rect 25881 11101 25915 11135
rect 25973 11101 26007 11135
rect 26249 11101 26283 11135
rect 26525 11101 26559 11135
rect 26617 11101 26651 11135
rect 27813 11101 27847 11135
rect 28089 11101 28123 11135
rect 28365 11101 28399 11135
rect 29745 11101 29779 11135
rect 29837 11101 29871 11135
rect 30021 11101 30055 11135
rect 30481 11101 30515 11135
rect 30573 11101 30607 11135
rect 30665 11101 30699 11135
rect 13645 11033 13679 11067
rect 14473 11033 14507 11067
rect 14565 11033 14599 11067
rect 17601 11033 17635 11067
rect 17693 11033 17727 11067
rect 19533 11033 19567 11067
rect 19625 11033 19659 11067
rect 25053 11033 25087 11067
rect 8493 10965 8527 10999
rect 11713 10965 11747 10999
rect 19257 10965 19291 10999
rect 27905 10965 27939 10999
rect 5273 10761 5307 10795
rect 7573 10761 7607 10795
rect 8033 10761 8067 10795
rect 8953 10761 8987 10795
rect 12265 10761 12299 10795
rect 14381 10761 14415 10795
rect 15669 10761 15703 10795
rect 16313 10761 16347 10795
rect 17601 10761 17635 10795
rect 18337 10761 18371 10795
rect 20913 10761 20947 10795
rect 22017 10761 22051 10795
rect 23305 10761 23339 10795
rect 26249 10761 26283 10795
rect 27721 10761 27755 10795
rect 29837 10761 29871 10795
rect 32137 10761 32171 10795
rect 33885 10761 33919 10795
rect 12541 10693 12575 10727
rect 15393 10693 15427 10727
rect 17233 10693 17267 10727
rect 21833 10693 21867 10727
rect 25881 10693 25915 10727
rect 27445 10693 27479 10727
rect 28825 10693 28859 10727
rect 29469 10693 29503 10727
rect 33517 10693 33551 10727
rect 5089 10625 5123 10659
rect 5641 10625 5675 10659
rect 5733 10625 5767 10659
rect 7941 10625 7975 10659
rect 9321 10625 9355 10659
rect 9965 10625 9999 10659
rect 11529 10625 11563 10659
rect 11713 10625 11747 10659
rect 11805 10625 11839 10659
rect 11897 10625 11931 10659
rect 12449 10625 12483 10659
rect 12633 10625 12667 10659
rect 12817 10625 12851 10659
rect 13921 10625 13955 10659
rect 14197 10625 14231 10659
rect 15117 10625 15151 10659
rect 15301 10625 15335 10659
rect 15531 10625 15565 10659
rect 15761 10625 15795 10659
rect 15945 10625 15979 10659
rect 16037 10625 16071 10659
rect 16129 10625 16163 10659
rect 17049 10625 17083 10659
rect 17325 10625 17359 10659
rect 17417 10625 17451 10659
rect 17693 10625 17727 10659
rect 17877 10625 17911 10659
rect 17969 10625 18003 10659
rect 18061 10625 18095 10659
rect 18521 10625 18555 10659
rect 18981 10625 19015 10659
rect 19073 10625 19107 10659
rect 21097 10625 21131 10659
rect 21281 10625 21315 10659
rect 21373 10625 21407 10659
rect 22293 10625 22327 10659
rect 22753 10625 22787 10659
rect 22845 10625 22879 10659
rect 23029 10625 23063 10659
rect 23121 10625 23155 10659
rect 23397 10625 23431 10659
rect 25605 10625 25639 10659
rect 25698 10625 25732 10659
rect 25973 10625 26007 10659
rect 26111 10625 26145 10659
rect 27261 10625 27295 10659
rect 28319 10625 28353 10659
rect 28457 10625 28491 10659
rect 28687 10625 28721 10659
rect 28917 10625 28951 10659
rect 29101 10625 29135 10659
rect 29285 10625 29319 10659
rect 29561 10625 29595 10659
rect 29653 10625 29687 10659
rect 31401 10625 31435 10659
rect 32505 10625 32539 10659
rect 33977 10625 34011 10659
rect 5917 10557 5951 10591
rect 8125 10557 8159 10591
rect 9413 10557 9447 10591
rect 9505 10557 9539 10591
rect 9873 10557 9907 10591
rect 18705 10557 18739 10591
rect 18797 10557 18831 10591
rect 20821 10557 20855 10591
rect 25145 10557 25179 10591
rect 28089 10557 28123 10591
rect 32597 10557 32631 10591
rect 32689 10557 32723 10591
rect 33241 10557 33275 10591
rect 33425 10557 33459 10591
rect 18245 10489 18279 10523
rect 18613 10489 18647 10523
rect 27997 10489 28031 10523
rect 4905 10421 4939 10455
rect 12173 10421 12207 10455
rect 14013 10421 14047 10455
rect 22017 10421 22051 10455
rect 27629 10421 27663 10455
rect 28181 10421 28215 10455
rect 28549 10421 28583 10455
rect 31217 10421 31251 10455
rect 34161 10421 34195 10455
rect 4616 10217 4650 10251
rect 10701 10217 10735 10251
rect 15393 10217 15427 10251
rect 15945 10217 15979 10251
rect 20637 10217 20671 10251
rect 22109 10217 22143 10251
rect 23581 10217 23615 10251
rect 25605 10217 25639 10251
rect 28457 10217 28491 10251
rect 28825 10217 28859 10251
rect 29009 10217 29043 10251
rect 32781 10217 32815 10251
rect 17509 10149 17543 10183
rect 6377 10081 6411 10115
rect 7757 10081 7791 10115
rect 7941 10081 7975 10115
rect 31309 10081 31343 10115
rect 4077 10013 4111 10047
rect 4169 10013 4203 10047
rect 4353 10013 4387 10047
rect 6653 10013 6687 10047
rect 7021 10013 7055 10047
rect 8309 10013 8343 10047
rect 8769 10013 8803 10047
rect 8953 10013 8987 10047
rect 12909 10013 12943 10047
rect 15209 10013 15243 10047
rect 15301 10013 15335 10047
rect 17417 10013 17451 10047
rect 17785 10013 17819 10047
rect 17877 10013 17911 10047
rect 18061 10013 18095 10047
rect 19993 10013 20027 10047
rect 20086 10013 20120 10047
rect 20361 10013 20395 10047
rect 20458 10013 20492 10047
rect 22293 10013 22327 10047
rect 22569 10013 22603 10047
rect 23765 10013 23799 10047
rect 23857 10013 23891 10047
rect 24133 10013 24167 10047
rect 24961 10013 24995 10047
rect 25054 10013 25088 10047
rect 25467 10013 25501 10047
rect 26065 10013 26099 10047
rect 27905 10013 27939 10047
rect 28089 10013 28123 10047
rect 28273 10013 28307 10047
rect 30757 10013 30791 10047
rect 30849 10013 30883 10047
rect 31033 10013 31067 10047
rect 33425 10013 33459 10047
rect 8677 9945 8711 9979
rect 9229 9945 9263 9979
rect 17693 9945 17727 9979
rect 20269 9945 20303 9979
rect 23949 9945 23983 9979
rect 25237 9945 25271 9979
rect 25329 9945 25363 9979
rect 28181 9945 28215 9979
rect 28641 9945 28675 9979
rect 6561 9877 6595 9911
rect 6837 9877 6871 9911
rect 7297 9877 7331 9911
rect 7665 9877 7699 9911
rect 8493 9877 8527 9911
rect 12817 9877 12851 9911
rect 15577 9877 15611 9911
rect 22477 9877 22511 9911
rect 27537 9877 27571 9911
rect 28841 9877 28875 9911
rect 33517 9877 33551 9911
rect 8125 9673 8159 9707
rect 16497 9673 16531 9707
rect 17785 9673 17819 9707
rect 18429 9673 18463 9707
rect 33333 9673 33367 9707
rect 6653 9605 6687 9639
rect 13921 9605 13955 9639
rect 17049 9605 17083 9639
rect 23949 9605 23983 9639
rect 24685 9605 24719 9639
rect 24869 9605 24903 9639
rect 25053 9605 25087 9639
rect 27353 9605 27387 9639
rect 29837 9605 29871 9639
rect 34805 9605 34839 9639
rect 6377 9537 6411 9571
rect 9597 9537 9631 9571
rect 11989 9537 12023 9571
rect 15853 9537 15887 9571
rect 15945 9537 15979 9571
rect 16129 9537 16163 9571
rect 16221 9537 16255 9571
rect 16313 9537 16347 9571
rect 17233 9537 17267 9571
rect 17325 9537 17359 9571
rect 17417 9537 17451 9571
rect 17693 9537 17727 9571
rect 17969 9537 18003 9571
rect 19349 9537 19383 9571
rect 22109 9537 22143 9571
rect 22753 9537 22787 9571
rect 23673 9537 23707 9571
rect 23857 9537 23891 9571
rect 24041 9537 24075 9571
rect 24501 9537 24535 9571
rect 24777 9537 24811 9571
rect 25876 9537 25910 9571
rect 25973 9537 26007 9571
rect 26065 9537 26099 9571
rect 26248 9537 26282 9571
rect 26341 9537 26375 9571
rect 27169 9537 27203 9571
rect 27261 9537 27295 9571
rect 27537 9537 27571 9571
rect 29653 9537 29687 9571
rect 29929 9537 29963 9571
rect 30021 9537 30055 9571
rect 32781 9537 32815 9571
rect 9873 9469 9907 9503
rect 22201 9469 22235 9503
rect 22569 9469 22603 9503
rect 30849 9469 30883 9503
rect 31493 9469 31527 9503
rect 32873 9469 32907 9503
rect 32965 9469 32999 9503
rect 35081 9469 35115 9503
rect 13737 9401 13771 9435
rect 17601 9401 17635 9435
rect 18061 9401 18095 9435
rect 22937 9401 22971 9435
rect 25697 9401 25731 9435
rect 26985 9401 27019 9435
rect 11345 9333 11379 9367
rect 12252 9333 12286 9367
rect 15209 9333 15243 9367
rect 18153 9333 18187 9367
rect 20637 9333 20671 9367
rect 22201 9333 22235 9367
rect 22477 9333 22511 9367
rect 24225 9333 24259 9367
rect 30205 9333 30239 9367
rect 32413 9333 32447 9367
rect 10517 9129 10551 9163
rect 11437 9129 11471 9163
rect 13093 9129 13127 9163
rect 16221 9129 16255 9163
rect 21005 9129 21039 9163
rect 22477 9129 22511 9163
rect 28825 9129 28859 9163
rect 29009 9129 29043 9163
rect 30113 9129 30147 9163
rect 31953 9129 31987 9163
rect 34437 9129 34471 9163
rect 14473 9061 14507 9095
rect 18521 9061 18555 9095
rect 19625 9061 19659 9095
rect 22109 9061 22143 9095
rect 12081 8993 12115 9027
rect 15117 8993 15151 9027
rect 22569 8993 22603 9027
rect 24409 8993 24443 9027
rect 26065 8993 26099 9027
rect 26249 8993 26283 9027
rect 30481 8993 30515 9027
rect 4629 8925 4663 8959
rect 10701 8925 10735 8959
rect 10793 8925 10827 8959
rect 10977 8925 11011 8959
rect 11069 8925 11103 8959
rect 11161 8925 11195 8959
rect 11989 8925 12023 8959
rect 13277 8925 13311 8959
rect 13553 8925 13587 8959
rect 13645 8925 13679 8959
rect 13737 8925 13771 8959
rect 13921 8925 13955 8959
rect 14933 8925 14967 8959
rect 15577 8925 15611 8959
rect 15761 8925 15795 8959
rect 15853 8925 15887 8959
rect 15945 8925 15979 8959
rect 17877 8925 17911 8959
rect 18061 8925 18095 8959
rect 18153 8925 18187 8959
rect 18279 8935 18313 8969
rect 19881 8925 19915 8959
rect 19990 8925 20024 8959
rect 20090 8925 20124 8959
rect 20269 8925 20303 8959
rect 20361 8925 20395 8959
rect 20545 8925 20579 8959
rect 20637 8925 20671 8959
rect 20729 8925 20763 8959
rect 21097 8925 21131 8959
rect 21557 8925 21591 8959
rect 21925 8925 21959 8959
rect 22753 8925 22787 8959
rect 24685 8925 24719 8959
rect 24961 8925 24995 8959
rect 25513 8925 25547 8959
rect 25789 8925 25823 8959
rect 25973 8925 26007 8959
rect 27813 8925 27847 8959
rect 27997 8925 28031 8959
rect 29561 8925 29595 8959
rect 29653 8925 29687 8959
rect 29837 8925 29871 8959
rect 29929 8925 29963 8959
rect 30205 8925 30239 8959
rect 32413 8925 32447 8959
rect 32689 8925 32723 8959
rect 14841 8857 14875 8891
rect 21281 8857 21315 8891
rect 21465 8857 21499 8891
rect 21741 8857 21775 8891
rect 21833 8857 21867 8891
rect 22477 8857 22511 8891
rect 27905 8857 27939 8891
rect 28457 8857 28491 8891
rect 28834 8857 28868 8891
rect 32965 8857 32999 8891
rect 4537 8789 4571 8823
rect 11529 8789 11563 8823
rect 11897 8789 11931 8823
rect 13369 8789 13403 8823
rect 22937 8789 22971 8823
rect 26249 8789 26283 8823
rect 32597 8789 32631 8823
rect 17693 8585 17727 8619
rect 18061 8585 18095 8619
rect 20545 8585 20579 8619
rect 20913 8585 20947 8619
rect 22385 8585 22419 8619
rect 22569 8585 22603 8619
rect 23213 8585 23247 8619
rect 28365 8585 28399 8619
rect 30389 8585 30423 8619
rect 32873 8585 32907 8619
rect 6193 8517 6227 8551
rect 14749 8517 14783 8551
rect 20085 8517 20119 8551
rect 20177 8517 20211 8551
rect 21281 8517 21315 8551
rect 22017 8517 22051 8551
rect 23489 8517 23523 8551
rect 26801 8517 26835 8551
rect 27879 8517 27913 8551
rect 28733 8517 28767 8551
rect 28917 8517 28951 8551
rect 4169 8449 4203 8483
rect 7849 8449 7883 8483
rect 9597 8449 9631 8483
rect 15025 8449 15059 8483
rect 15117 8449 15151 8483
rect 15209 8449 15243 8483
rect 17877 8449 17911 8483
rect 18153 8449 18187 8483
rect 19809 8449 19843 8483
rect 19902 8449 19936 8483
rect 20274 8449 20308 8483
rect 20729 8449 20763 8483
rect 21005 8449 21039 8483
rect 21097 8449 21131 8483
rect 21373 8449 21407 8483
rect 21465 8449 21499 8483
rect 21833 8449 21867 8483
rect 22109 8449 22143 8483
rect 22201 8449 22235 8483
rect 22753 8449 22787 8483
rect 22845 8449 22879 8483
rect 23029 8449 23063 8483
rect 23121 8449 23155 8483
rect 23351 8449 23385 8483
rect 23581 8449 23615 8483
rect 23764 8449 23798 8483
rect 23857 8449 23891 8483
rect 25237 8449 25271 8483
rect 25421 8449 25455 8483
rect 25697 8449 25731 8483
rect 25973 8449 26007 8483
rect 26166 8449 26200 8483
rect 26985 8449 27019 8483
rect 27169 8449 27203 8483
rect 27721 8449 27755 8483
rect 27997 8449 28031 8483
rect 28089 8449 28123 8483
rect 28181 8449 28215 8483
rect 28513 8449 28547 8483
rect 28641 8449 28675 8483
rect 30481 8449 30515 8483
rect 32965 8449 32999 8483
rect 4445 8381 4479 8415
rect 28825 8381 28859 8415
rect 13461 8313 13495 8347
rect 14841 8313 14875 8347
rect 20453 8313 20487 8347
rect 21649 8313 21683 8347
rect 26985 8313 27019 8347
rect 15393 8245 15427 8279
rect 4905 8041 4939 8075
rect 11529 8041 11563 8075
rect 14105 8041 14139 8075
rect 15669 8041 15703 8075
rect 16405 8041 16439 8075
rect 16773 8041 16807 8075
rect 17969 8041 18003 8075
rect 18705 8041 18739 8075
rect 20361 8041 20395 8075
rect 22937 8041 22971 8075
rect 23121 8041 23155 8075
rect 24777 8041 24811 8075
rect 27905 8041 27939 8075
rect 29561 8041 29595 8075
rect 30573 8041 30607 8075
rect 5365 7973 5399 8007
rect 20453 7973 20487 8007
rect 6009 7905 6043 7939
rect 8769 7905 8803 7939
rect 10425 7905 10459 7939
rect 12449 7905 12483 7939
rect 18245 7905 18279 7939
rect 30573 7905 30607 7939
rect 5089 7837 5123 7871
rect 5733 7837 5767 7871
rect 6745 7837 6779 7871
rect 6837 7837 6871 7871
rect 7021 7837 7055 7871
rect 9413 7837 9447 7871
rect 9689 7837 9723 7871
rect 11713 7837 11747 7871
rect 11805 7837 11839 7871
rect 11989 7837 12023 7871
rect 12081 7837 12115 7871
rect 12173 7837 12207 7871
rect 14749 7837 14783 7871
rect 15117 7837 15151 7871
rect 15485 7837 15519 7871
rect 15761 7837 15795 7871
rect 15945 7837 15979 7871
rect 16129 7837 16163 7871
rect 16405 7837 16439 7871
rect 16497 7837 16531 7871
rect 17325 7837 17359 7871
rect 17418 7837 17452 7871
rect 17693 7837 17727 7871
rect 17831 7837 17865 7871
rect 18153 7837 18187 7871
rect 18429 7837 18463 7871
rect 18521 7837 18555 7871
rect 19809 7837 19843 7871
rect 19901 7837 19935 7871
rect 20085 7837 20119 7871
rect 20177 7837 20211 7871
rect 20637 7837 20671 7871
rect 20821 7837 20855 7871
rect 21005 7837 21039 7871
rect 24961 7837 24995 7871
rect 25237 7837 25271 7871
rect 27813 7837 27847 7871
rect 27997 7837 28031 7871
rect 29745 7837 29779 7871
rect 29837 7837 29871 7871
rect 30021 7837 30055 7871
rect 30113 7837 30147 7871
rect 30205 7837 30239 7871
rect 30389 7837 30423 7871
rect 30481 7837 30515 7871
rect 32413 7837 32447 7871
rect 7297 7769 7331 7803
rect 10149 7769 10183 7803
rect 15301 7769 15335 7803
rect 15393 7769 15427 7803
rect 16037 7769 16071 7803
rect 17601 7769 17635 7803
rect 20729 7769 20763 7803
rect 22753 7769 22787 7803
rect 22969 7769 23003 7803
rect 5825 7701 5859 7735
rect 9321 7701 9355 7735
rect 9505 7701 9539 7735
rect 9781 7701 9815 7735
rect 10241 7701 10275 7735
rect 13921 7701 13955 7735
rect 16313 7701 16347 7735
rect 25145 7701 25179 7735
rect 32321 7701 32355 7735
rect 6377 7497 6411 7531
rect 6837 7497 6871 7531
rect 7665 7497 7699 7531
rect 8401 7497 8435 7531
rect 12357 7497 12391 7531
rect 16037 7497 16071 7531
rect 18337 7497 18371 7531
rect 20177 7497 20211 7531
rect 22385 7497 22419 7531
rect 23305 7497 23339 7531
rect 25329 7497 25363 7531
rect 26249 7497 26283 7531
rect 29377 7497 29411 7531
rect 30389 7497 30423 7531
rect 31585 7497 31619 7531
rect 6745 7429 6779 7463
rect 9413 7429 9447 7463
rect 11805 7429 11839 7463
rect 13001 7429 13035 7463
rect 14749 7429 14783 7463
rect 18061 7429 18095 7463
rect 23397 7429 23431 7463
rect 29009 7429 29043 7463
rect 6101 7361 6135 7395
rect 7849 7361 7883 7395
rect 8493 7361 8527 7395
rect 9137 7361 9171 7395
rect 11621 7361 11655 7395
rect 11897 7361 11931 7395
rect 11989 7361 12023 7395
rect 12449 7361 12483 7395
rect 15393 7361 15427 7395
rect 15486 7361 15520 7395
rect 15669 7361 15703 7395
rect 15761 7361 15795 7395
rect 15899 7361 15933 7395
rect 16313 7361 16347 7395
rect 16497 7361 16531 7395
rect 17049 7361 17083 7395
rect 17233 7361 17267 7395
rect 17325 7361 17359 7395
rect 17417 7361 17451 7395
rect 17693 7361 17727 7395
rect 17786 7361 17820 7395
rect 17969 7361 18003 7395
rect 18158 7361 18192 7395
rect 18449 7361 18483 7395
rect 18613 7361 18647 7395
rect 18705 7361 18739 7395
rect 18797 7361 18831 7395
rect 20637 7361 20671 7395
rect 21281 7361 21315 7395
rect 21833 7361 21867 7395
rect 22017 7361 22051 7395
rect 22109 7361 22143 7395
rect 22201 7361 22235 7395
rect 22753 7361 22787 7395
rect 22937 7361 22971 7395
rect 23029 7361 23063 7395
rect 23121 7361 23155 7395
rect 25508 7361 25542 7395
rect 25605 7361 25639 7395
rect 25697 7361 25731 7395
rect 25880 7361 25914 7395
rect 25973 7361 26007 7395
rect 26065 7361 26099 7395
rect 26341 7361 26375 7395
rect 28825 7361 28859 7395
rect 29101 7361 29135 7395
rect 29193 7361 29227 7395
rect 29745 7361 29779 7395
rect 29838 7361 29872 7395
rect 30021 7361 30055 7395
rect 30113 7361 30147 7395
rect 30210 7361 30244 7395
rect 32137 7361 32171 7395
rect 6929 7293 6963 7327
rect 8585 7293 8619 7327
rect 10885 7293 10919 7327
rect 31401 7293 31435 7327
rect 31493 7293 31527 7327
rect 32413 7293 32447 7327
rect 8033 7225 8067 7259
rect 12173 7225 12207 7259
rect 16129 7225 16163 7259
rect 26065 7225 26099 7259
rect 5917 7157 5951 7191
rect 17601 7157 17635 7191
rect 18981 7157 19015 7191
rect 24685 7157 24719 7191
rect 31953 7157 31987 7191
rect 33885 7157 33919 7191
rect 5720 6953 5754 6987
rect 7205 6953 7239 6987
rect 18153 6953 18187 6987
rect 25881 6953 25915 6987
rect 29745 6953 29779 6987
rect 31769 6953 31803 6987
rect 18429 6885 18463 6919
rect 14105 6817 14139 6851
rect 18521 6817 18555 6851
rect 20269 6817 20303 6851
rect 28273 6817 28307 6851
rect 28549 6817 28583 6851
rect 5181 6749 5215 6783
rect 5273 6749 5307 6783
rect 5457 6749 5491 6783
rect 11897 6749 11931 6783
rect 14197 6749 14231 6783
rect 14381 6749 14415 6783
rect 14565 6749 14599 6783
rect 14657 6749 14691 6783
rect 14750 6749 14784 6783
rect 15122 6749 15156 6783
rect 16865 6749 16899 6783
rect 17141 6749 17175 6783
rect 17233 6749 17267 6783
rect 18337 6749 18371 6783
rect 18613 6749 18647 6783
rect 18797 6749 18831 6783
rect 20085 6749 20119 6783
rect 21557 6749 21591 6783
rect 21650 6749 21684 6783
rect 21833 6749 21867 6783
rect 21925 6749 21959 6783
rect 22063 6749 22097 6783
rect 22293 6749 22327 6783
rect 22386 6749 22420 6783
rect 22799 6749 22833 6783
rect 23208 6749 23242 6783
rect 23580 6749 23614 6783
rect 23673 6749 23707 6783
rect 24961 6749 24995 6783
rect 25053 6749 25087 6783
rect 25329 6749 25363 6783
rect 25697 6749 25731 6783
rect 26019 6749 26053 6783
rect 26157 6749 26191 6783
rect 26249 6749 26283 6783
rect 26432 6749 26466 6783
rect 26525 6749 26559 6783
rect 27261 6749 27295 6783
rect 27629 6749 27663 6783
rect 27813 6749 27847 6783
rect 27905 6749 27939 6783
rect 27997 6749 28031 6783
rect 28365 6749 28399 6783
rect 28641 6749 28675 6783
rect 28733 6749 28767 6783
rect 28825 6749 28859 6783
rect 29009 6749 29043 6783
rect 31585 6749 31619 6783
rect 14933 6681 14967 6715
rect 15025 6681 15059 6715
rect 17049 6681 17083 6715
rect 22569 6681 22603 6715
rect 22661 6681 22695 6715
rect 23305 6681 23339 6715
rect 23397 6681 23431 6715
rect 24777 6681 24811 6715
rect 25421 6681 25455 6715
rect 25513 6681 25547 6715
rect 26985 6681 27019 6715
rect 27537 6681 27571 6715
rect 29929 6681 29963 6715
rect 11805 6613 11839 6647
rect 15301 6613 15335 6647
rect 17417 6613 17451 6647
rect 22201 6613 22235 6647
rect 22937 6613 22971 6647
rect 23029 6613 23063 6647
rect 25053 6613 25087 6647
rect 25145 6613 25179 6647
rect 27169 6613 27203 6647
rect 27353 6613 27387 6647
rect 29561 6613 29595 6647
rect 29719 6613 29753 6647
rect 13369 6409 13403 6443
rect 13829 6409 13863 6443
rect 17049 6409 17083 6443
rect 17233 6409 17267 6443
rect 17601 6409 17635 6443
rect 18245 6409 18279 6443
rect 20177 6409 20211 6443
rect 21281 6409 21315 6443
rect 21649 6409 21683 6443
rect 23489 6409 23523 6443
rect 24409 6409 24443 6443
rect 24501 6409 24535 6443
rect 24869 6409 24903 6443
rect 25513 6409 25547 6443
rect 28089 6409 28123 6443
rect 13921 6341 13955 6375
rect 21465 6341 21499 6375
rect 26065 6341 26099 6375
rect 27721 6341 27755 6375
rect 8953 6273 8987 6307
rect 10517 6273 10551 6307
rect 11621 6273 11655 6307
rect 15025 6273 15059 6307
rect 17141 6273 17175 6307
rect 17509 6273 17543 6307
rect 17785 6273 17819 6307
rect 17969 6273 18003 6307
rect 19993 6273 20027 6307
rect 21373 6273 21407 6307
rect 21925 6273 21959 6307
rect 22109 6273 22143 6307
rect 22201 6273 22235 6307
rect 22293 6273 22327 6307
rect 22385 6273 22419 6307
rect 23213 6273 23247 6307
rect 23305 6273 23339 6307
rect 24593 6273 24627 6307
rect 25145 6273 25179 6307
rect 25605 6273 25639 6307
rect 25881 6273 25915 6307
rect 25973 6273 26007 6307
rect 26249 6273 26283 6307
rect 27813 6273 27847 6307
rect 27905 6273 27939 6307
rect 30205 6273 30239 6307
rect 11897 6205 11931 6239
rect 14013 6205 14047 6239
rect 19809 6205 19843 6239
rect 22937 6205 22971 6239
rect 24225 6205 24259 6239
rect 25329 6205 25363 6239
rect 16865 6137 16899 6171
rect 17417 6137 17451 6171
rect 17877 6137 17911 6171
rect 21097 6137 21131 6171
rect 24777 6137 24811 6171
rect 27537 6137 27571 6171
rect 8861 6069 8895 6103
rect 10425 6069 10459 6103
rect 13461 6069 13495 6103
rect 14933 6069 14967 6103
rect 22569 6069 22603 6103
rect 23029 6069 23063 6103
rect 25237 6069 25271 6103
rect 25697 6069 25731 6103
rect 30021 6069 30055 6103
rect 12357 5865 12391 5899
rect 24777 5865 24811 5899
rect 9321 5797 9355 5831
rect 25329 5797 25363 5831
rect 5549 5729 5583 5763
rect 6561 5729 6595 5763
rect 6745 5729 6779 5763
rect 8769 5729 8803 5763
rect 9781 5729 9815 5763
rect 9965 5729 9999 5763
rect 10241 5729 10275 5763
rect 12265 5729 12299 5763
rect 14749 5729 14783 5763
rect 15577 5729 15611 5763
rect 29929 5729 29963 5763
rect 5365 5661 5399 5695
rect 6653 5661 6687 5695
rect 9229 5661 9263 5695
rect 12541 5661 12575 5695
rect 13093 5661 13127 5695
rect 14473 5661 14507 5695
rect 15301 5661 15335 5695
rect 17233 5661 17267 5695
rect 17509 5661 17543 5695
rect 17601 5661 17635 5695
rect 19441 5661 19475 5695
rect 19533 5661 19567 5695
rect 24961 5661 24995 5695
rect 29653 5661 29687 5695
rect 31493 5661 31527 5695
rect 7021 5593 7055 5627
rect 9689 5593 9723 5627
rect 10517 5593 10551 5627
rect 25145 5593 25179 5627
rect 31769 5593 31803 5627
rect 5181 5525 5215 5559
rect 9045 5525 9079 5559
rect 13001 5525 13035 5559
rect 14105 5525 14139 5559
rect 14565 5525 14599 5559
rect 14933 5525 14967 5559
rect 15393 5525 15427 5559
rect 17417 5525 17451 5559
rect 17785 5525 17819 5559
rect 19257 5525 19291 5559
rect 19625 5525 19659 5559
rect 25053 5525 25087 5559
rect 31401 5525 31435 5559
rect 33241 5525 33275 5559
rect 5549 5321 5583 5355
rect 27445 5321 27479 5355
rect 29837 5321 29871 5355
rect 30021 5321 30055 5355
rect 30389 5321 30423 5355
rect 31677 5321 31711 5355
rect 32505 5321 32539 5355
rect 8033 5253 8067 5287
rect 8953 5253 8987 5287
rect 10701 5253 10735 5287
rect 11989 5253 12023 5287
rect 22385 5253 22419 5287
rect 1961 5185 1995 5219
rect 5365 5185 5399 5219
rect 7481 5185 7515 5219
rect 10977 5185 11011 5219
rect 11897 5185 11931 5219
rect 18981 5185 19015 5219
rect 22293 5185 22327 5219
rect 23857 5185 23891 5219
rect 26985 5185 27019 5219
rect 27261 5185 27295 5219
rect 27721 5185 27755 5219
rect 28089 5185 28123 5219
rect 29929 5185 29963 5219
rect 30481 5185 30515 5219
rect 31309 5185 31343 5219
rect 31769 5185 31803 5219
rect 8125 5117 8159 5151
rect 8217 5117 8251 5151
rect 8677 5117 8711 5151
rect 12081 5117 12115 5151
rect 12817 5117 12851 5151
rect 13093 5117 13127 5151
rect 14565 5117 14599 5151
rect 14749 5117 14783 5151
rect 15025 5117 15059 5151
rect 16497 5117 16531 5151
rect 19257 5117 19291 5151
rect 22569 5117 22603 5151
rect 23673 5117 23707 5151
rect 23765 5117 23799 5151
rect 30573 5117 30607 5151
rect 32597 5117 32631 5151
rect 32689 5117 32723 5151
rect 7297 5049 7331 5083
rect 7665 5049 7699 5083
rect 10793 5049 10827 5083
rect 11529 5049 11563 5083
rect 31493 5049 31527 5083
rect 32137 5049 32171 5083
rect 1777 4981 1811 5015
rect 20729 4981 20763 5015
rect 21925 4981 21959 5015
rect 24225 4981 24259 5015
rect 27169 4981 27203 5015
rect 27629 4981 27663 5015
rect 27997 4981 28031 5015
rect 1593 4777 1627 4811
rect 22845 4777 22879 4811
rect 26157 4777 26191 4811
rect 27169 4777 27203 4811
rect 13369 4709 13403 4743
rect 15025 4709 15059 4743
rect 23949 4709 23983 4743
rect 29193 4709 29227 4743
rect 19901 4641 19935 4675
rect 20913 4641 20947 4675
rect 21097 4641 21131 4675
rect 23489 4641 23523 4675
rect 24133 4641 24167 4675
rect 24409 4641 24443 4675
rect 24685 4641 24719 4675
rect 26525 4641 26559 4675
rect 8953 4573 8987 4607
rect 13553 4573 13587 4607
rect 15209 4573 15243 4607
rect 16957 4573 16991 4607
rect 19809 4573 19843 4607
rect 21005 4573 21039 4607
rect 23305 4573 23339 4607
rect 23765 4573 23799 4607
rect 24225 4573 24259 4607
rect 26709 4573 26743 4607
rect 27445 4573 27479 4607
rect 1501 4505 1535 4539
rect 21373 4505 21407 4539
rect 27721 4505 27755 4539
rect 9137 4437 9171 4471
rect 16865 4437 16899 4471
rect 19349 4437 19383 4471
rect 19717 4437 19751 4471
rect 22937 4437 22971 4471
rect 23397 4437 23431 4471
rect 26801 4437 26835 4471
rect 21833 4233 21867 4267
rect 26985 4233 27019 4267
rect 29561 4233 29595 4267
rect 27353 4165 27387 4199
rect 12265 4097 12299 4131
rect 12541 4097 12575 4131
rect 16313 4097 16347 4131
rect 22017 4097 22051 4131
rect 27445 4097 27479 4131
rect 16681 4029 16715 4063
rect 16957 4029 16991 4063
rect 27537 4029 27571 4063
rect 27813 4029 27847 4063
rect 28089 4029 28123 4063
rect 16497 3961 16531 3995
rect 12173 3893 12207 3927
rect 12357 3893 12391 3927
rect 18429 3893 18463 3927
rect 7113 3689 7147 3723
rect 17141 3689 17175 3723
rect 37657 3689 37691 3723
rect 15209 3621 15243 3655
rect 17969 3621 18003 3655
rect 18245 3621 18279 3655
rect 20453 3621 20487 3655
rect 11897 3553 11931 3587
rect 12173 3553 12207 3587
rect 14473 3553 14507 3587
rect 15853 3553 15887 3587
rect 17693 3553 17727 3587
rect 18797 3553 18831 3587
rect 19809 3553 19843 3587
rect 24593 3553 24627 3587
rect 24777 3553 24811 3587
rect 25329 3553 25363 3587
rect 26065 3553 26099 3587
rect 26249 3553 26283 3587
rect 6929 3485 6963 3519
rect 9045 3485 9079 3519
rect 9137 3485 9171 3519
rect 9321 3485 9355 3519
rect 11621 3485 11655 3519
rect 11713 3485 11747 3519
rect 14289 3485 14323 3519
rect 14657 3485 14691 3519
rect 15117 3485 15151 3519
rect 16865 3485 16899 3519
rect 18153 3485 18187 3519
rect 18613 3485 18647 3519
rect 19993 3485 20027 3519
rect 20729 3485 20763 3519
rect 21005 3485 21039 3519
rect 22109 3485 22143 3519
rect 22385 3485 22419 3519
rect 23949 3485 23983 3519
rect 25513 3485 25547 3519
rect 27261 3485 27295 3519
rect 28181 3485 28215 3519
rect 28365 3485 28399 3519
rect 37473 3485 37507 3519
rect 9597 3417 9631 3451
rect 11345 3417 11379 3451
rect 13921 3417 13955 3451
rect 11437 3349 11471 3383
rect 14105 3349 14139 3383
rect 14749 3349 14783 3383
rect 14933 3349 14967 3383
rect 15577 3349 15611 3383
rect 15669 3349 15703 3383
rect 16957 3349 16991 3383
rect 17509 3349 17543 3383
rect 17601 3349 17635 3383
rect 18705 3349 18739 3383
rect 20085 3349 20119 3383
rect 20545 3349 20579 3383
rect 20913 3349 20947 3383
rect 22017 3349 22051 3383
rect 22201 3349 22235 3383
rect 24041 3349 24075 3383
rect 24869 3349 24903 3383
rect 25237 3349 25271 3383
rect 25697 3349 25731 3383
rect 26341 3349 26375 3383
rect 26709 3349 26743 3383
rect 27169 3349 27203 3383
rect 28549 3349 28583 3383
rect 23581 3145 23615 3179
rect 31861 3145 31895 3179
rect 1777 3077 1811 3111
rect 12725 3077 12759 3111
rect 14473 3077 14507 3111
rect 14841 3077 14875 3111
rect 17601 3077 17635 3111
rect 20085 3077 20119 3111
rect 22109 3077 22143 3111
rect 25881 3077 25915 3111
rect 37565 3077 37599 3111
rect 2145 3009 2179 3043
rect 7021 3009 7055 3043
rect 10057 3009 10091 3043
rect 10793 3009 10827 3043
rect 10885 3009 10919 3043
rect 11529 3009 11563 3043
rect 11621 3009 11655 3043
rect 11805 3009 11839 3043
rect 12173 3009 12207 3043
rect 12265 3009 12299 3043
rect 14565 3009 14599 3043
rect 17325 3009 17359 3043
rect 19553 3009 19587 3043
rect 19809 3009 19843 3043
rect 21833 3009 21867 3043
rect 23857 3009 23891 3043
rect 25973 3009 26007 3043
rect 26433 3009 26467 3043
rect 26985 3009 27019 3043
rect 30849 3009 30883 3043
rect 31033 3009 31067 3043
rect 31217 3009 31251 3043
rect 31677 3009 31711 3043
rect 36921 3009 36955 3043
rect 10977 2941 11011 2975
rect 11989 2941 12023 2975
rect 19073 2941 19107 2975
rect 19349 2941 19383 2975
rect 24133 2941 24167 2975
rect 27261 2941 27295 2975
rect 9873 2873 9907 2907
rect 10425 2873 10459 2907
rect 12633 2873 12667 2907
rect 21557 2873 21591 2907
rect 26617 2873 26651 2907
rect 1501 2805 1535 2839
rect 1961 2805 1995 2839
rect 6837 2805 6871 2839
rect 11713 2805 11747 2839
rect 16313 2805 16347 2839
rect 19717 2805 19751 2839
rect 26157 2805 26191 2839
rect 28733 2805 28767 2839
rect 37105 2805 37139 2839
rect 37841 2805 37875 2839
rect 13231 2601 13265 2635
rect 25145 2601 25179 2635
rect 12633 2465 12667 2499
rect 14381 2465 14415 2499
rect 16129 2465 16163 2499
rect 31217 2465 31251 2499
rect 1777 2397 1811 2431
rect 2421 2397 2455 2431
rect 4353 2397 4387 2431
rect 6929 2397 6963 2431
rect 10885 2397 10919 2431
rect 12081 2397 12115 2431
rect 12265 2397 12299 2431
rect 12449 2397 12483 2431
rect 12541 2397 12575 2431
rect 13001 2397 13035 2431
rect 15117 2397 15151 2431
rect 16313 2397 16347 2431
rect 16497 2397 16531 2431
rect 16865 2397 16899 2431
rect 19809 2397 19843 2431
rect 24685 2397 24719 2431
rect 25329 2397 25363 2431
rect 27077 2397 27111 2431
rect 31033 2397 31067 2431
rect 35541 2397 35575 2431
rect 37381 2397 37415 2431
rect 1409 2329 1443 2363
rect 2053 2329 2087 2363
rect 3985 2329 4019 2363
rect 6561 2329 6595 2363
rect 11621 2329 11655 2363
rect 15577 2329 15611 2363
rect 15945 2329 15979 2363
rect 20177 2329 20211 2363
rect 11069 2261 11103 2295
rect 11713 2261 11747 2295
rect 16681 2261 16715 2295
rect 19993 2261 20027 2295
rect 20269 2261 20303 2295
rect 24961 2261 24995 2295
rect 27169 2261 27203 2295
rect 35725 2261 35759 2295
rect 37657 2261 37691 2295
<< metal1 >>
rect 1104 39194 38272 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 35594 39194
rect 35646 39142 35658 39194
rect 35710 39142 35722 39194
rect 35774 39142 35786 39194
rect 35838 39142 35850 39194
rect 35902 39142 38272 39194
rect 1104 39120 38272 39142
rect 658 39040 664 39092
rect 716 39080 722 39092
rect 1489 39083 1547 39089
rect 1489 39080 1501 39083
rect 716 39052 1501 39080
rect 716 39040 722 39052
rect 1489 39049 1501 39052
rect 1535 39049 1547 39083
rect 1489 39043 1547 39049
rect 2133 39083 2191 39089
rect 2133 39049 2145 39083
rect 2179 39049 2191 39083
rect 2133 39043 2191 39049
rect 1118 38972 1124 39024
rect 1176 39012 1182 39024
rect 2148 39012 2176 39043
rect 5258 39040 5264 39092
rect 5316 39080 5322 39092
rect 5353 39083 5411 39089
rect 5353 39080 5365 39083
rect 5316 39052 5365 39080
rect 5316 39040 5322 39052
rect 5353 39049 5365 39052
rect 5399 39049 5411 39083
rect 5353 39043 5411 39049
rect 9766 39040 9772 39092
rect 9824 39080 9830 39092
rect 9861 39083 9919 39089
rect 9861 39080 9873 39083
rect 9824 39052 9873 39080
rect 9824 39040 9830 39052
rect 9861 39049 9873 39052
rect 9907 39049 9919 39083
rect 9861 39043 9919 39049
rect 14182 39040 14188 39092
rect 14240 39080 14246 39092
rect 14553 39083 14611 39089
rect 14553 39080 14565 39083
rect 14240 39052 14565 39080
rect 14240 39040 14246 39052
rect 14553 39049 14565 39052
rect 14599 39049 14611 39083
rect 14553 39043 14611 39049
rect 17586 39040 17592 39092
rect 17644 39040 17650 39092
rect 23198 39040 23204 39092
rect 23256 39080 23262 39092
rect 23477 39083 23535 39089
rect 23477 39080 23489 39083
rect 23256 39052 23489 39080
rect 23256 39040 23262 39052
rect 23477 39049 23489 39052
rect 23523 39049 23535 39083
rect 23477 39043 23535 39049
rect 25130 39040 25136 39092
rect 25188 39080 25194 39092
rect 25409 39083 25467 39089
rect 25409 39080 25421 39083
rect 25188 39052 25421 39080
rect 25188 39040 25194 39052
rect 25409 39049 25421 39052
rect 25455 39049 25467 39083
rect 25409 39043 25467 39049
rect 27338 39040 27344 39092
rect 27396 39040 27402 39092
rect 31846 39040 31852 39092
rect 31904 39080 31910 39092
rect 32309 39083 32367 39089
rect 32309 39080 32321 39083
rect 31904 39052 32321 39080
rect 31904 39040 31910 39052
rect 32309 39049 32321 39052
rect 32355 39049 32367 39083
rect 32309 39043 32367 39049
rect 34146 39040 34152 39092
rect 34204 39080 34210 39092
rect 34885 39083 34943 39089
rect 34885 39080 34897 39083
rect 34204 39052 34897 39080
rect 34204 39040 34210 39052
rect 34885 39049 34897 39052
rect 34931 39049 34943 39083
rect 34885 39043 34943 39049
rect 36354 39040 36360 39092
rect 36412 39040 36418 39092
rect 1176 38984 2176 39012
rect 1176 38972 1182 38984
rect 20714 38972 20720 39024
rect 20772 39012 20778 39024
rect 20901 39015 20959 39021
rect 20901 39012 20913 39015
rect 20772 38984 20913 39012
rect 20772 38972 20778 38984
rect 20901 38981 20913 38984
rect 20947 38981 20959 39015
rect 20901 38975 20959 38981
rect 23934 38972 23940 39024
rect 23992 39012 23998 39024
rect 23992 38984 36308 39012
rect 23992 38972 23998 38984
rect 1762 38904 1768 38956
rect 1820 38904 1826 38956
rect 2038 38904 2044 38956
rect 2096 38904 2102 38956
rect 5629 38947 5687 38953
rect 5629 38913 5641 38947
rect 5675 38944 5687 38947
rect 9674 38944 9680 38956
rect 5675 38916 9680 38944
rect 5675 38913 5687 38916
rect 5629 38907 5687 38913
rect 9674 38904 9680 38916
rect 9732 38904 9738 38956
rect 10134 38904 10140 38956
rect 10192 38904 10198 38956
rect 14734 38904 14740 38956
rect 14792 38904 14798 38956
rect 17770 38904 17776 38956
rect 17828 38904 17834 38956
rect 23382 38904 23388 38956
rect 23440 38904 23446 38956
rect 25222 38904 25228 38956
rect 25280 38904 25286 38956
rect 27246 38904 27252 38956
rect 27304 38904 27310 38956
rect 32217 38947 32275 38953
rect 32217 38944 32229 38947
rect 31726 38916 32229 38944
rect 14826 38836 14832 38888
rect 14884 38876 14890 38888
rect 31726 38876 31754 38916
rect 32217 38913 32229 38916
rect 32263 38913 32275 38947
rect 32217 38907 32275 38913
rect 33594 38904 33600 38956
rect 33652 38944 33658 38956
rect 34793 38947 34851 38953
rect 34793 38944 34805 38947
rect 33652 38916 34805 38944
rect 33652 38904 33658 38916
rect 34793 38913 34805 38916
rect 34839 38913 34851 38947
rect 34793 38907 34851 38913
rect 36173 38947 36231 38953
rect 36173 38913 36185 38947
rect 36219 38913 36231 38947
rect 36280 38944 36308 38984
rect 37182 38972 37188 39024
rect 37240 39012 37246 39024
rect 37829 39015 37887 39021
rect 37829 39012 37841 39015
rect 37240 38984 37841 39012
rect 37240 38972 37246 38984
rect 37829 38981 37841 38984
rect 37875 38981 37887 39015
rect 37829 38975 37887 38981
rect 37645 38947 37703 38953
rect 37645 38944 37657 38947
rect 36280 38916 37657 38944
rect 36173 38907 36231 38913
rect 37645 38913 37657 38916
rect 37691 38913 37703 38947
rect 37645 38907 37703 38913
rect 14884 38848 31754 38876
rect 14884 38836 14890 38848
rect 13906 38768 13912 38820
rect 13964 38808 13970 38820
rect 20717 38811 20775 38817
rect 20717 38808 20729 38811
rect 13964 38780 20729 38808
rect 13964 38768 13970 38780
rect 20717 38777 20729 38780
rect 20763 38777 20775 38811
rect 36188 38808 36216 38907
rect 20717 38771 20775 38777
rect 22066 38780 36216 38808
rect 14642 38700 14648 38752
rect 14700 38740 14706 38752
rect 22066 38740 22094 38780
rect 14700 38712 22094 38740
rect 14700 38700 14706 38712
rect 1104 38650 38272 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 38272 38650
rect 1104 38576 38272 38598
rect 1949 38539 2007 38545
rect 1949 38505 1961 38539
rect 1995 38536 2007 38539
rect 2038 38536 2044 38548
rect 1995 38508 2044 38536
rect 1995 38505 2007 38508
rect 1949 38499 2007 38505
rect 2038 38496 2044 38508
rect 2096 38496 2102 38548
rect 9674 38496 9680 38548
rect 9732 38536 9738 38548
rect 11425 38539 11483 38545
rect 11425 38536 11437 38539
rect 9732 38508 11437 38536
rect 9732 38496 9738 38508
rect 11425 38505 11437 38508
rect 11471 38505 11483 38539
rect 11425 38499 11483 38505
rect 19426 38496 19432 38548
rect 19484 38536 19490 38548
rect 21082 38536 21088 38548
rect 19484 38508 21088 38536
rect 19484 38496 19490 38508
rect 21082 38496 21088 38508
rect 21140 38536 21146 38548
rect 21140 38508 23244 38536
rect 21140 38496 21146 38508
rect 23216 38480 23244 38508
rect 21560 38440 21864 38468
rect 17313 38403 17371 38409
rect 17313 38400 17325 38403
rect 15028 38372 17325 38400
rect 1765 38335 1823 38341
rect 1765 38301 1777 38335
rect 1811 38332 1823 38335
rect 1811 38304 2774 38332
rect 1811 38301 1823 38304
rect 1765 38295 1823 38301
rect 2746 38196 2774 38304
rect 11606 38292 11612 38344
rect 11664 38292 11670 38344
rect 14182 38292 14188 38344
rect 14240 38332 14246 38344
rect 15028 38341 15056 38372
rect 17313 38369 17325 38372
rect 17359 38400 17371 38403
rect 17954 38400 17960 38412
rect 17359 38372 17960 38400
rect 17359 38369 17371 38372
rect 17313 38363 17371 38369
rect 17954 38360 17960 38372
rect 18012 38400 18018 38412
rect 19705 38403 19763 38409
rect 19705 38400 19717 38403
rect 18012 38372 19717 38400
rect 18012 38360 18018 38372
rect 19705 38369 19717 38372
rect 19751 38400 19763 38403
rect 21560 38400 21588 38440
rect 21836 38409 21864 38440
rect 23198 38428 23204 38480
rect 23256 38468 23262 38480
rect 23474 38468 23480 38480
rect 23256 38440 23480 38468
rect 23256 38428 23262 38440
rect 23474 38428 23480 38440
rect 23532 38428 23538 38480
rect 24213 38471 24271 38477
rect 24213 38437 24225 38471
rect 24259 38468 24271 38471
rect 24259 38440 24532 38468
rect 24259 38437 24271 38440
rect 24213 38431 24271 38437
rect 19751 38372 21588 38400
rect 21821 38403 21879 38409
rect 19751 38369 19763 38372
rect 19705 38363 19763 38369
rect 21821 38369 21833 38403
rect 21867 38400 21879 38403
rect 24397 38403 24455 38409
rect 24397 38400 24409 38403
rect 21867 38372 24409 38400
rect 21867 38369 21879 38372
rect 21821 38363 21879 38369
rect 24397 38369 24409 38372
rect 24443 38369 24455 38403
rect 24504 38400 24532 38440
rect 24673 38403 24731 38409
rect 24673 38400 24685 38403
rect 24504 38372 24685 38400
rect 24397 38363 24455 38369
rect 24673 38369 24685 38372
rect 24719 38369 24731 38403
rect 24673 38363 24731 38369
rect 15013 38335 15071 38341
rect 15013 38332 15025 38335
rect 14240 38304 15025 38332
rect 14240 38292 14246 38304
rect 15013 38301 15025 38304
rect 15059 38301 15071 38335
rect 15013 38295 15071 38301
rect 21082 38292 21088 38344
rect 21140 38292 21146 38344
rect 23198 38292 23204 38344
rect 23256 38292 23262 38344
rect 24026 38292 24032 38344
rect 24084 38292 24090 38344
rect 15286 38224 15292 38276
rect 15344 38224 15350 38276
rect 15838 38224 15844 38276
rect 15896 38224 15902 38276
rect 17586 38224 17592 38276
rect 17644 38224 17650 38276
rect 19426 38264 19432 38276
rect 18814 38236 19432 38264
rect 19426 38224 19432 38236
rect 19484 38224 19490 38276
rect 19978 38224 19984 38276
rect 20036 38224 20042 38276
rect 22094 38224 22100 38276
rect 22152 38224 22158 38276
rect 23474 38224 23480 38276
rect 23532 38264 23538 38276
rect 24118 38264 24124 38276
rect 23532 38236 24124 38264
rect 23532 38224 23538 38236
rect 24118 38224 24124 38236
rect 24176 38264 24182 38276
rect 24176 38236 25162 38264
rect 24176 38224 24182 38236
rect 10318 38196 10324 38208
rect 2746 38168 10324 38196
rect 10318 38156 10324 38168
rect 10376 38156 10382 38208
rect 16758 38156 16764 38208
rect 16816 38156 16822 38208
rect 19058 38156 19064 38208
rect 19116 38156 19122 38208
rect 20714 38156 20720 38208
rect 20772 38196 20778 38208
rect 21450 38196 21456 38208
rect 20772 38168 21456 38196
rect 20772 38156 20778 38168
rect 21450 38156 21456 38168
rect 21508 38156 21514 38208
rect 22922 38156 22928 38208
rect 22980 38196 22986 38208
rect 23569 38199 23627 38205
rect 23569 38196 23581 38199
rect 22980 38168 23581 38196
rect 22980 38156 22986 38168
rect 23569 38165 23581 38168
rect 23615 38165 23627 38199
rect 23569 38159 23627 38165
rect 25038 38156 25044 38208
rect 25096 38196 25102 38208
rect 26050 38196 26056 38208
rect 25096 38168 26056 38196
rect 25096 38156 25102 38168
rect 26050 38156 26056 38168
rect 26108 38196 26114 38208
rect 26145 38199 26203 38205
rect 26145 38196 26157 38199
rect 26108 38168 26157 38196
rect 26108 38156 26114 38168
rect 26145 38165 26157 38168
rect 26191 38165 26203 38199
rect 26145 38159 26203 38165
rect 1104 38106 38272 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 35594 38106
rect 35646 38054 35658 38106
rect 35710 38054 35722 38106
rect 35774 38054 35786 38106
rect 35838 38054 35850 38106
rect 35902 38054 38272 38106
rect 1104 38032 38272 38054
rect 10134 37952 10140 38004
rect 10192 37992 10198 38004
rect 10229 37995 10287 38001
rect 10229 37992 10241 37995
rect 10192 37964 10241 37992
rect 10192 37952 10198 37964
rect 10229 37961 10241 37964
rect 10275 37961 10287 37995
rect 10229 37955 10287 37961
rect 10318 37952 10324 38004
rect 10376 37992 10382 38004
rect 12805 37995 12863 38001
rect 12805 37992 12817 37995
rect 10376 37964 12817 37992
rect 10376 37952 10382 37964
rect 12805 37961 12817 37964
rect 12851 37961 12863 37995
rect 12805 37955 12863 37961
rect 15286 37952 15292 38004
rect 15344 37992 15350 38004
rect 15565 37995 15623 38001
rect 15565 37992 15577 37995
rect 15344 37964 15577 37992
rect 15344 37952 15350 37964
rect 15565 37961 15577 37964
rect 15611 37961 15623 37995
rect 16390 37992 16396 38004
rect 15565 37955 15623 37961
rect 15672 37964 16396 37992
rect 13998 37884 14004 37936
rect 14056 37924 14062 37936
rect 15672 37924 15700 37964
rect 16390 37952 16396 37964
rect 16448 37952 16454 38004
rect 16669 37995 16727 38001
rect 16669 37961 16681 37995
rect 16715 37961 16727 37995
rect 16669 37955 16727 37961
rect 16684 37924 16712 37955
rect 16758 37952 16764 38004
rect 16816 37992 16822 38004
rect 17037 37995 17095 38001
rect 17037 37992 17049 37995
rect 16816 37964 17049 37992
rect 16816 37952 16822 37964
rect 17037 37961 17049 37964
rect 17083 37961 17095 37995
rect 17037 37955 17095 37961
rect 17589 37995 17647 38001
rect 17589 37961 17601 37995
rect 17635 37992 17647 37995
rect 17770 37992 17776 38004
rect 17635 37964 17776 37992
rect 17635 37961 17647 37964
rect 17589 37955 17647 37961
rect 17770 37952 17776 37964
rect 17828 37952 17834 38004
rect 17957 37995 18015 38001
rect 17957 37961 17969 37995
rect 18003 37992 18015 37995
rect 19058 37992 19064 38004
rect 18003 37964 19064 37992
rect 18003 37961 18015 37964
rect 17957 37955 18015 37961
rect 14056 37896 15700 37924
rect 15764 37896 16712 37924
rect 14056 37884 14062 37896
rect 1765 37859 1823 37865
rect 1765 37825 1777 37859
rect 1811 37856 1823 37859
rect 10413 37859 10471 37865
rect 1811 37828 2774 37856
rect 1811 37825 1823 37828
rect 1765 37819 1823 37825
rect 2746 37788 2774 37828
rect 10413 37825 10425 37859
rect 10459 37856 10471 37859
rect 12066 37856 12072 37868
rect 10459 37828 12072 37856
rect 10459 37825 10471 37828
rect 10413 37819 10471 37825
rect 12066 37816 12072 37828
rect 12124 37816 12130 37868
rect 12986 37816 12992 37868
rect 13044 37816 13050 37868
rect 15764 37865 15792 37896
rect 17678 37884 17684 37936
rect 17736 37924 17742 37936
rect 17972 37924 18000 37955
rect 19058 37952 19064 37964
rect 19116 37952 19122 38004
rect 19978 37952 19984 38004
rect 20036 37992 20042 38004
rect 20073 37995 20131 38001
rect 20073 37992 20085 37995
rect 20036 37964 20085 37992
rect 20036 37952 20042 37964
rect 20073 37961 20085 37964
rect 20119 37961 20131 37995
rect 20073 37955 20131 37961
rect 20714 37952 20720 38004
rect 20772 37952 20778 38004
rect 22094 37952 22100 38004
rect 22152 37992 22158 38004
rect 22281 37995 22339 38001
rect 22281 37992 22293 37995
rect 22152 37964 22293 37992
rect 22152 37952 22158 37964
rect 22281 37961 22293 37964
rect 22327 37961 22339 37995
rect 22281 37955 22339 37961
rect 22557 37995 22615 38001
rect 22557 37961 22569 37995
rect 22603 37961 22615 37995
rect 22557 37955 22615 37961
rect 17736 37896 18000 37924
rect 19812 37896 20852 37924
rect 17736 37884 17742 37896
rect 15749 37859 15807 37865
rect 13096 37828 15700 37856
rect 13096 37788 13124 37828
rect 2746 37760 13124 37788
rect 13173 37791 13231 37797
rect 13173 37757 13185 37791
rect 13219 37788 13231 37791
rect 13998 37788 14004 37800
rect 13219 37760 14004 37788
rect 13219 37757 13231 37760
rect 13173 37751 13231 37757
rect 13998 37748 14004 37760
rect 14056 37748 14062 37800
rect 15672 37788 15700 37828
rect 15749 37825 15761 37859
rect 15795 37825 15807 37859
rect 15749 37819 15807 37825
rect 16114 37816 16120 37868
rect 16172 37816 16178 37868
rect 16206 37816 16212 37868
rect 16264 37816 16270 37868
rect 16298 37816 16304 37868
rect 16356 37816 16362 37868
rect 16390 37816 16396 37868
rect 16448 37856 16454 37868
rect 16485 37859 16543 37865
rect 16485 37856 16497 37859
rect 16448 37828 16497 37856
rect 16448 37816 16454 37828
rect 16485 37825 16497 37828
rect 16531 37825 16543 37859
rect 16485 37819 16543 37825
rect 17328 37828 18184 37856
rect 17328 37800 17356 37828
rect 15672 37760 17080 37788
rect 17052 37720 17080 37760
rect 17126 37748 17132 37800
rect 17184 37748 17190 37800
rect 17310 37748 17316 37800
rect 17368 37748 17374 37800
rect 18046 37748 18052 37800
rect 18104 37748 18110 37800
rect 18156 37797 18184 37828
rect 19812 37800 19840 37896
rect 20257 37859 20315 37865
rect 20257 37825 20269 37859
rect 20303 37856 20315 37859
rect 20824 37856 20852 37896
rect 22465 37859 22523 37865
rect 20303 37828 20392 37856
rect 20824 37828 20944 37856
rect 20303 37825 20315 37828
rect 20257 37819 20315 37825
rect 18141 37791 18199 37797
rect 18141 37757 18153 37791
rect 18187 37788 18199 37791
rect 19794 37788 19800 37800
rect 18187 37760 19800 37788
rect 18187 37757 18199 37760
rect 18141 37751 18199 37757
rect 19794 37748 19800 37760
rect 19852 37748 19858 37800
rect 19978 37720 19984 37732
rect 2746 37692 15884 37720
rect 17052 37692 19984 37720
rect 934 37612 940 37664
rect 992 37652 998 37664
rect 1489 37655 1547 37661
rect 1489 37652 1501 37655
rect 992 37624 1501 37652
rect 992 37612 998 37624
rect 1489 37621 1501 37624
rect 1535 37621 1547 37655
rect 1489 37615 1547 37621
rect 1762 37612 1768 37664
rect 1820 37652 1826 37664
rect 2746 37652 2774 37692
rect 15856 37661 15884 37692
rect 19978 37680 19984 37692
rect 20036 37680 20042 37732
rect 20364 37729 20392 37828
rect 20806 37748 20812 37800
rect 20864 37748 20870 37800
rect 20916 37797 20944 37828
rect 22465 37825 22477 37859
rect 22511 37856 22523 37859
rect 22572 37856 22600 37955
rect 22922 37952 22928 38004
rect 22980 37952 22986 38004
rect 24026 37952 24032 38004
rect 24084 37992 24090 38004
rect 24397 37995 24455 38001
rect 24397 37992 24409 37995
rect 24084 37964 24409 37992
rect 24084 37952 24090 37964
rect 24397 37961 24409 37964
rect 24443 37961 24455 37995
rect 24397 37955 24455 37961
rect 24765 37995 24823 38001
rect 24765 37961 24777 37995
rect 24811 37992 24823 37995
rect 25038 37992 25044 38004
rect 24811 37964 25044 37992
rect 24811 37961 24823 37964
rect 24765 37955 24823 37961
rect 25038 37952 25044 37964
rect 25096 37952 25102 38004
rect 25222 37952 25228 38004
rect 25280 37952 25286 38004
rect 26605 37995 26663 38001
rect 26605 37961 26617 37995
rect 26651 37992 26663 37995
rect 27246 37992 27252 38004
rect 26651 37964 27252 37992
rect 26651 37961 26663 37964
rect 26605 37955 26663 37961
rect 27246 37952 27252 37964
rect 27304 37952 27310 38004
rect 25608 37896 26280 37924
rect 25608 37868 25636 37896
rect 22511 37828 22600 37856
rect 25501 37859 25559 37865
rect 22511 37825 22523 37828
rect 22465 37819 22523 37825
rect 25501 37825 25513 37859
rect 25547 37825 25559 37859
rect 25501 37819 25559 37825
rect 20901 37791 20959 37797
rect 20901 37757 20913 37791
rect 20947 37788 20959 37791
rect 20947 37760 22094 37788
rect 20947 37757 20959 37760
rect 20901 37751 20959 37757
rect 20349 37723 20407 37729
rect 20349 37689 20361 37723
rect 20395 37689 20407 37723
rect 22066 37720 22094 37760
rect 23014 37748 23020 37800
rect 23072 37748 23078 37800
rect 23201 37791 23259 37797
rect 23201 37757 23213 37791
rect 23247 37788 23259 37791
rect 23750 37788 23756 37800
rect 23247 37760 23756 37788
rect 23247 37757 23259 37760
rect 23201 37751 23259 37757
rect 23216 37720 23244 37751
rect 23750 37748 23756 37760
rect 23808 37748 23814 37800
rect 24854 37748 24860 37800
rect 24912 37748 24918 37800
rect 24949 37791 25007 37797
rect 24949 37757 24961 37791
rect 24995 37757 25007 37791
rect 25516 37788 25544 37819
rect 25590 37816 25596 37868
rect 25648 37816 25654 37868
rect 25682 37816 25688 37868
rect 25740 37816 25746 37868
rect 25869 37859 25927 37865
rect 25869 37825 25881 37859
rect 25915 37856 25927 37859
rect 25961 37859 26019 37865
rect 25961 37856 25973 37859
rect 25915 37828 25973 37856
rect 25915 37825 25927 37828
rect 25869 37819 25927 37825
rect 25961 37825 25973 37828
rect 26007 37825 26019 37859
rect 25961 37819 26019 37825
rect 25774 37788 25780 37800
rect 25516 37760 25780 37788
rect 24949 37751 25007 37757
rect 22066 37692 23244 37720
rect 23768 37720 23796 37748
rect 24964 37720 24992 37751
rect 25774 37748 25780 37760
rect 25832 37748 25838 37800
rect 23768 37692 24992 37720
rect 20349 37683 20407 37689
rect 1820 37624 2774 37652
rect 15841 37655 15899 37661
rect 1820 37612 1826 37624
rect 15841 37621 15853 37655
rect 15887 37621 15899 37655
rect 15841 37615 15899 37621
rect 24946 37612 24952 37664
rect 25004 37652 25010 37664
rect 25884 37652 25912 37819
rect 26142 37816 26148 37868
rect 26200 37816 26206 37868
rect 26252 37865 26280 37896
rect 26237 37859 26295 37865
rect 26237 37825 26249 37859
rect 26283 37825 26295 37859
rect 26237 37819 26295 37825
rect 26329 37859 26387 37865
rect 26329 37825 26341 37859
rect 26375 37856 26387 37859
rect 27246 37856 27252 37868
rect 26375 37828 27252 37856
rect 26375 37825 26387 37828
rect 26329 37819 26387 37825
rect 27246 37816 27252 37828
rect 27304 37816 27310 37868
rect 37642 37816 37648 37868
rect 37700 37816 37706 37868
rect 25004 37624 25912 37652
rect 25004 37612 25010 37624
rect 37826 37612 37832 37664
rect 37884 37612 37890 37664
rect 1104 37562 38272 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38272 37562
rect 1104 37488 38272 37510
rect 11606 37408 11612 37460
rect 11664 37408 11670 37460
rect 12066 37408 12072 37460
rect 12124 37408 12130 37460
rect 16114 37408 16120 37460
rect 16172 37408 16178 37460
rect 16298 37408 16304 37460
rect 16356 37448 16362 37460
rect 16393 37451 16451 37457
rect 16393 37448 16405 37451
rect 16356 37420 16405 37448
rect 16356 37408 16362 37420
rect 16393 37417 16405 37420
rect 16439 37417 16451 37451
rect 16393 37411 16451 37417
rect 19978 37408 19984 37460
rect 20036 37408 20042 37460
rect 20346 37408 20352 37460
rect 20404 37448 20410 37460
rect 21082 37448 21088 37460
rect 20404 37420 21088 37448
rect 20404 37408 20410 37420
rect 21082 37408 21088 37420
rect 21140 37448 21146 37460
rect 22830 37448 22836 37460
rect 21140 37420 22836 37448
rect 21140 37408 21146 37420
rect 22830 37408 22836 37420
rect 22888 37408 22894 37460
rect 25409 37451 25467 37457
rect 25409 37417 25421 37451
rect 25455 37448 25467 37451
rect 25682 37448 25688 37460
rect 25455 37420 25688 37448
rect 25455 37417 25467 37420
rect 25409 37411 25467 37417
rect 25682 37408 25688 37420
rect 25740 37408 25746 37460
rect 25869 37451 25927 37457
rect 25869 37417 25881 37451
rect 25915 37448 25927 37451
rect 26142 37448 26148 37460
rect 25915 37420 26148 37448
rect 25915 37417 25927 37420
rect 25869 37411 25927 37417
rect 26142 37408 26148 37420
rect 26200 37408 26206 37460
rect 16132 37380 16160 37408
rect 24670 37380 24676 37392
rect 16132 37352 24676 37380
rect 24670 37340 24676 37352
rect 24728 37340 24734 37392
rect 2590 37272 2596 37324
rect 2648 37312 2654 37324
rect 8478 37312 8484 37324
rect 2648 37284 8484 37312
rect 2648 37272 2654 37284
rect 8478 37272 8484 37284
rect 8536 37272 8542 37324
rect 11974 37272 11980 37324
rect 12032 37272 12038 37324
rect 14458 37272 14464 37324
rect 14516 37312 14522 37324
rect 16114 37312 16120 37324
rect 14516 37284 16120 37312
rect 14516 37272 14522 37284
rect 16114 37272 16120 37284
rect 16172 37272 16178 37324
rect 20162 37312 20168 37324
rect 19306 37284 20168 37312
rect 11793 37247 11851 37253
rect 11793 37244 11805 37247
rect 11624 37216 11805 37244
rect 11624 37120 11652 37216
rect 11793 37213 11805 37216
rect 11839 37244 11851 37247
rect 12253 37247 12311 37253
rect 12253 37244 12265 37247
rect 11839 37216 12265 37244
rect 11839 37213 11851 37216
rect 11793 37207 11851 37213
rect 12253 37213 12265 37216
rect 12299 37213 12311 37247
rect 12253 37207 12311 37213
rect 12434 37204 12440 37256
rect 12492 37204 12498 37256
rect 12710 37204 12716 37256
rect 12768 37204 12774 37256
rect 16209 37247 16267 37253
rect 16209 37213 16221 37247
rect 16255 37244 16267 37247
rect 16298 37244 16304 37256
rect 16255 37216 16304 37244
rect 16255 37213 16267 37216
rect 16209 37207 16267 37213
rect 16298 37204 16304 37216
rect 16356 37244 16362 37256
rect 16758 37244 16764 37256
rect 16356 37216 16764 37244
rect 16356 37204 16362 37216
rect 16758 37204 16764 37216
rect 16816 37204 16822 37256
rect 19306 37244 19334 37284
rect 20162 37272 20168 37284
rect 20220 37272 20226 37324
rect 21542 37272 21548 37324
rect 21600 37312 21606 37324
rect 21600 37284 25728 37312
rect 21600 37272 21606 37284
rect 19260 37216 19334 37244
rect 13538 37136 13544 37188
rect 13596 37176 13602 37188
rect 16025 37179 16083 37185
rect 16025 37176 16037 37179
rect 13596 37148 16037 37176
rect 13596 37136 13602 37148
rect 16025 37145 16037 37148
rect 16071 37176 16083 37179
rect 19260 37176 19288 37216
rect 19886 37204 19892 37256
rect 19944 37244 19950 37256
rect 20257 37247 20315 37253
rect 20257 37244 20269 37247
rect 19944 37216 20269 37244
rect 19944 37204 19950 37216
rect 20257 37213 20269 37216
rect 20303 37213 20315 37247
rect 20257 37207 20315 37213
rect 20349 37247 20407 37253
rect 20349 37213 20361 37247
rect 20395 37213 20407 37247
rect 20349 37207 20407 37213
rect 20441 37247 20499 37253
rect 20441 37213 20453 37247
rect 20487 37213 20499 37247
rect 20441 37207 20499 37213
rect 16071 37148 19288 37176
rect 16071 37145 16083 37148
rect 16025 37139 16083 37145
rect 19334 37136 19340 37188
rect 19392 37176 19398 37188
rect 20364 37176 20392 37207
rect 19392 37148 20392 37176
rect 20456 37176 20484 37207
rect 20530 37204 20536 37256
rect 20588 37244 20594 37256
rect 20625 37247 20683 37253
rect 20625 37244 20637 37247
rect 20588 37216 20637 37244
rect 20588 37204 20594 37216
rect 20625 37213 20637 37216
rect 20671 37213 20683 37247
rect 20625 37207 20683 37213
rect 20901 37247 20959 37253
rect 20901 37213 20913 37247
rect 20947 37244 20959 37247
rect 20990 37244 20996 37256
rect 20947 37216 20996 37244
rect 20947 37213 20959 37216
rect 20901 37207 20959 37213
rect 20990 37204 20996 37216
rect 21048 37244 21054 37256
rect 22922 37244 22928 37256
rect 21048 37216 22928 37244
rect 21048 37204 21054 37216
rect 22922 37204 22928 37216
rect 22980 37204 22986 37256
rect 25501 37247 25559 37253
rect 25501 37244 25513 37247
rect 25056 37216 25513 37244
rect 20717 37179 20775 37185
rect 20717 37176 20729 37179
rect 20456 37148 20729 37176
rect 19392 37136 19398 37148
rect 20717 37145 20729 37148
rect 20763 37145 20775 37179
rect 20717 37139 20775 37145
rect 21082 37136 21088 37188
rect 21140 37136 21146 37188
rect 22830 37136 22836 37188
rect 22888 37176 22894 37188
rect 25056 37185 25084 37216
rect 25501 37213 25513 37216
rect 25547 37213 25559 37247
rect 25501 37207 25559 37213
rect 25041 37179 25099 37185
rect 25041 37176 25053 37179
rect 22888 37148 25053 37176
rect 22888 37136 22894 37148
rect 25041 37145 25053 37148
rect 25087 37145 25099 37179
rect 25041 37139 25099 37145
rect 25130 37136 25136 37188
rect 25188 37176 25194 37188
rect 25700 37185 25728 37284
rect 25225 37179 25283 37185
rect 25225 37176 25237 37179
rect 25188 37148 25237 37176
rect 25188 37136 25194 37148
rect 25225 37145 25237 37148
rect 25271 37145 25283 37179
rect 25225 37139 25283 37145
rect 25685 37179 25743 37185
rect 25685 37145 25697 37179
rect 25731 37145 25743 37179
rect 25685 37139 25743 37145
rect 11606 37068 11612 37120
rect 11664 37068 11670 37120
rect 12894 37068 12900 37120
rect 12952 37068 12958 37120
rect 19058 37068 19064 37120
rect 19116 37108 19122 37120
rect 21542 37108 21548 37120
rect 19116 37080 21548 37108
rect 19116 37068 19122 37080
rect 21542 37068 21548 37080
rect 21600 37068 21606 37120
rect 1104 37018 38272 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 38272 37018
rect 1104 36944 38272 36966
rect 12710 36864 12716 36916
rect 12768 36864 12774 36916
rect 12894 36864 12900 36916
rect 12952 36904 12958 36916
rect 20717 36907 20775 36913
rect 12952 36876 13124 36904
rect 12952 36864 12958 36876
rect 12986 36836 12992 36848
rect 12084 36808 12992 36836
rect 10686 36660 10692 36712
rect 10744 36700 10750 36712
rect 12084 36709 12112 36808
rect 12986 36796 12992 36808
rect 13044 36796 13050 36848
rect 13096 36845 13124 36876
rect 20717 36873 20729 36907
rect 20763 36904 20775 36907
rect 20806 36904 20812 36916
rect 20763 36876 20812 36904
rect 20763 36873 20775 36876
rect 20717 36867 20775 36873
rect 20806 36864 20812 36876
rect 20864 36864 20870 36916
rect 21266 36864 21272 36916
rect 21324 36904 21330 36916
rect 21726 36904 21732 36916
rect 21324 36876 21732 36904
rect 21324 36864 21330 36876
rect 21726 36864 21732 36876
rect 21784 36904 21790 36916
rect 21784 36876 22968 36904
rect 21784 36864 21790 36876
rect 13081 36839 13139 36845
rect 13081 36805 13093 36839
rect 13127 36805 13139 36839
rect 13081 36799 13139 36805
rect 19426 36796 19432 36848
rect 19484 36796 19490 36848
rect 21450 36796 21456 36848
rect 21508 36836 21514 36848
rect 21910 36836 21916 36848
rect 21508 36808 21916 36836
rect 21508 36796 21514 36808
rect 21910 36796 21916 36808
rect 21968 36836 21974 36848
rect 22157 36839 22215 36845
rect 22157 36836 22169 36839
rect 21968 36808 22169 36836
rect 21968 36796 21974 36808
rect 22157 36805 22169 36808
rect 22203 36805 22215 36839
rect 22157 36799 22215 36805
rect 22373 36839 22431 36845
rect 22373 36805 22385 36839
rect 22419 36836 22431 36839
rect 22940 36836 22968 36876
rect 23014 36864 23020 36916
rect 23072 36904 23078 36916
rect 23293 36907 23351 36913
rect 23293 36904 23305 36907
rect 23072 36876 23305 36904
rect 23072 36864 23078 36876
rect 23293 36873 23305 36876
rect 23339 36873 23351 36907
rect 23293 36867 23351 36873
rect 33594 36864 33600 36916
rect 33652 36864 33658 36916
rect 37553 36907 37611 36913
rect 37553 36873 37565 36907
rect 37599 36904 37611 36907
rect 37642 36904 37648 36916
rect 37599 36876 37648 36904
rect 37599 36873 37611 36876
rect 37553 36867 37611 36873
rect 37642 36864 37648 36876
rect 37700 36864 37706 36916
rect 22419 36808 22784 36836
rect 22940 36808 23796 36836
rect 22419 36805 22431 36808
rect 22373 36799 22431 36805
rect 12342 36728 12348 36780
rect 12400 36728 12406 36780
rect 14090 36728 14096 36780
rect 14148 36768 14154 36780
rect 15838 36768 15844 36780
rect 14148 36740 15844 36768
rect 14148 36728 14154 36740
rect 15838 36728 15844 36740
rect 15896 36728 15902 36780
rect 17954 36728 17960 36780
rect 18012 36768 18018 36780
rect 18141 36771 18199 36777
rect 18141 36768 18153 36771
rect 18012 36740 18153 36768
rect 18012 36728 18018 36740
rect 18141 36737 18153 36740
rect 18187 36737 18199 36771
rect 18141 36731 18199 36737
rect 21085 36771 21143 36777
rect 21085 36737 21097 36771
rect 21131 36768 21143 36771
rect 21358 36768 21364 36780
rect 21131 36740 21364 36768
rect 21131 36737 21143 36740
rect 21085 36731 21143 36737
rect 21358 36728 21364 36740
rect 21416 36728 21422 36780
rect 22756 36777 22784 36808
rect 22741 36771 22799 36777
rect 22741 36737 22753 36771
rect 22787 36768 22799 36771
rect 22922 36768 22928 36780
rect 22787 36740 22928 36768
rect 22787 36737 22799 36740
rect 22741 36731 22799 36737
rect 22922 36728 22928 36740
rect 22980 36728 22986 36780
rect 23658 36728 23664 36780
rect 23716 36728 23722 36780
rect 23768 36768 23796 36808
rect 23768 36740 23888 36768
rect 12069 36703 12127 36709
rect 12069 36700 12081 36703
rect 10744 36672 12081 36700
rect 10744 36660 10750 36672
rect 12069 36669 12081 36672
rect 12115 36669 12127 36703
rect 12069 36663 12127 36669
rect 12253 36703 12311 36709
rect 12253 36669 12265 36703
rect 12299 36700 12311 36703
rect 12710 36700 12716 36712
rect 12299 36672 12716 36700
rect 12299 36669 12311 36672
rect 12253 36663 12311 36669
rect 12710 36660 12716 36672
rect 12768 36660 12774 36712
rect 12805 36703 12863 36709
rect 12805 36669 12817 36703
rect 12851 36700 12863 36703
rect 12851 36672 14228 36700
rect 12851 36669 12863 36672
rect 12805 36663 12863 36669
rect 14200 36576 14228 36672
rect 18414 36660 18420 36712
rect 18472 36660 18478 36712
rect 21174 36660 21180 36712
rect 21232 36660 21238 36712
rect 21266 36660 21272 36712
rect 21324 36660 21330 36712
rect 23860 36709 23888 36740
rect 25130 36728 25136 36780
rect 25188 36728 25194 36780
rect 25317 36771 25375 36777
rect 25317 36737 25329 36771
rect 25363 36768 25375 36771
rect 25363 36740 26004 36768
rect 25363 36737 25375 36740
rect 25317 36731 25375 36737
rect 22649 36703 22707 36709
rect 22649 36669 22661 36703
rect 22695 36669 22707 36703
rect 22649 36663 22707 36669
rect 23109 36703 23167 36709
rect 23109 36669 23121 36703
rect 23155 36700 23167 36703
rect 23753 36703 23811 36709
rect 23753 36700 23765 36703
rect 23155 36672 23765 36700
rect 23155 36669 23167 36672
rect 23109 36663 23167 36669
rect 23753 36669 23765 36672
rect 23799 36669 23811 36703
rect 23753 36663 23811 36669
rect 23845 36703 23903 36709
rect 23845 36669 23857 36703
rect 23891 36700 23903 36703
rect 25406 36700 25412 36712
rect 23891 36672 25412 36700
rect 23891 36669 23903 36672
rect 23845 36663 23903 36669
rect 22664 36632 22692 36663
rect 25406 36660 25412 36672
rect 25464 36660 25470 36712
rect 21284 36604 22692 36632
rect 21284 36576 21312 36604
rect 14182 36524 14188 36576
rect 14240 36524 14246 36576
rect 14550 36524 14556 36576
rect 14608 36524 14614 36576
rect 19889 36567 19947 36573
rect 19889 36533 19901 36567
rect 19935 36564 19947 36567
rect 21266 36564 21272 36576
rect 19935 36536 21272 36564
rect 19935 36533 19947 36536
rect 19889 36527 19947 36533
rect 21266 36524 21272 36536
rect 21324 36524 21330 36576
rect 22002 36524 22008 36576
rect 22060 36524 22066 36576
rect 22204 36573 22232 36604
rect 25976 36576 26004 36740
rect 28442 36728 28448 36780
rect 28500 36768 28506 36780
rect 33413 36771 33471 36777
rect 33413 36768 33425 36771
rect 28500 36740 33425 36768
rect 28500 36728 28506 36740
rect 33413 36737 33425 36740
rect 33459 36737 33471 36771
rect 33413 36731 33471 36737
rect 37366 36728 37372 36780
rect 37424 36728 37430 36780
rect 22189 36567 22247 36573
rect 22189 36533 22201 36567
rect 22235 36564 22247 36567
rect 22235 36536 22269 36564
rect 22235 36533 22247 36536
rect 22189 36527 22247 36533
rect 25314 36524 25320 36576
rect 25372 36524 25378 36576
rect 25958 36524 25964 36576
rect 26016 36524 26022 36576
rect 1104 36474 38272 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38272 36474
rect 1104 36400 38272 36422
rect 14090 36360 14096 36372
rect 10888 36332 14096 36360
rect 9858 36184 9864 36236
rect 9916 36224 9922 36236
rect 10888 36224 10916 36332
rect 14090 36320 14096 36332
rect 14148 36320 14154 36372
rect 14826 36320 14832 36372
rect 14884 36320 14890 36372
rect 16761 36363 16819 36369
rect 16761 36329 16773 36363
rect 16807 36360 16819 36363
rect 17126 36360 17132 36372
rect 16807 36332 17132 36360
rect 16807 36329 16819 36332
rect 16761 36323 16819 36329
rect 17126 36320 17132 36332
rect 17184 36320 17190 36372
rect 18414 36320 18420 36372
rect 18472 36360 18478 36372
rect 18509 36363 18567 36369
rect 18509 36360 18521 36363
rect 18472 36332 18521 36360
rect 18472 36320 18478 36332
rect 18509 36329 18521 36332
rect 18555 36329 18567 36363
rect 18509 36323 18567 36329
rect 21174 36320 21180 36372
rect 21232 36360 21238 36372
rect 21729 36363 21787 36369
rect 21729 36360 21741 36363
rect 21232 36332 21741 36360
rect 21232 36320 21238 36332
rect 21729 36329 21741 36332
rect 21775 36329 21787 36363
rect 21729 36323 21787 36329
rect 24854 36320 24860 36372
rect 24912 36320 24918 36372
rect 25314 36320 25320 36372
rect 25372 36320 25378 36372
rect 25958 36320 25964 36372
rect 26016 36320 26022 36372
rect 28442 36320 28448 36372
rect 28500 36320 28506 36372
rect 28997 36363 29055 36369
rect 28997 36329 29009 36363
rect 29043 36360 29055 36363
rect 37366 36360 37372 36372
rect 29043 36332 37372 36360
rect 29043 36329 29055 36332
rect 28997 36323 29055 36329
rect 37366 36320 37372 36332
rect 37424 36320 37430 36372
rect 12986 36252 12992 36304
rect 13044 36292 13050 36304
rect 17310 36292 17316 36304
rect 13044 36264 17316 36292
rect 13044 36252 13050 36264
rect 9916 36196 10916 36224
rect 9916 36184 9922 36196
rect 8294 36116 8300 36168
rect 8352 36156 8358 36168
rect 9214 36156 9220 36168
rect 8352 36128 9220 36156
rect 8352 36116 8358 36128
rect 9214 36116 9220 36128
rect 9272 36156 9278 36168
rect 9493 36159 9551 36165
rect 9493 36156 9505 36159
rect 9272 36128 9505 36156
rect 9272 36116 9278 36128
rect 9493 36125 9505 36128
rect 9539 36125 9551 36159
rect 10888 36142 10916 36196
rect 13909 36227 13967 36233
rect 13909 36193 13921 36227
rect 13955 36224 13967 36227
rect 13955 36196 14412 36224
rect 13955 36193 13967 36196
rect 13909 36187 13967 36193
rect 9493 36119 9551 36125
rect 11624 36128 13860 36156
rect 11624 36100 11652 36128
rect 9766 36048 9772 36100
rect 9824 36048 9830 36100
rect 11606 36048 11612 36100
rect 11664 36048 11670 36100
rect 13538 36048 13544 36100
rect 13596 36048 13602 36100
rect 13725 36091 13783 36097
rect 13725 36057 13737 36091
rect 13771 36057 13783 36091
rect 13832 36088 13860 36128
rect 14090 36116 14096 36168
rect 14148 36156 14154 36168
rect 14384 36165 14412 36196
rect 15378 36184 15384 36236
rect 15436 36184 15442 36236
rect 15488 36233 15516 36264
rect 17310 36252 17316 36264
rect 17368 36252 17374 36304
rect 19245 36295 19303 36301
rect 19245 36261 19257 36295
rect 19291 36261 19303 36295
rect 19245 36255 19303 36261
rect 15473 36227 15531 36233
rect 15473 36193 15485 36227
rect 15519 36193 15531 36227
rect 15473 36187 15531 36193
rect 16393 36227 16451 36233
rect 16393 36193 16405 36227
rect 16439 36224 16451 36227
rect 16574 36224 16580 36236
rect 16439 36196 16580 36224
rect 16439 36193 16451 36196
rect 16393 36187 16451 36193
rect 16574 36184 16580 36196
rect 16632 36184 16638 36236
rect 16669 36227 16727 36233
rect 16669 36193 16681 36227
rect 16715 36224 16727 36227
rect 17221 36227 17279 36233
rect 17221 36224 17233 36227
rect 16715 36196 17233 36224
rect 16715 36193 16727 36196
rect 16669 36187 16727 36193
rect 17221 36193 17233 36196
rect 17267 36193 17279 36227
rect 17221 36187 17279 36193
rect 17405 36227 17463 36233
rect 17405 36193 17417 36227
rect 17451 36224 17463 36227
rect 18782 36224 18788 36236
rect 17451 36196 18788 36224
rect 17451 36193 17463 36196
rect 17405 36187 17463 36193
rect 14185 36159 14243 36165
rect 14185 36156 14197 36159
rect 14148 36128 14197 36156
rect 14148 36116 14154 36128
rect 14185 36125 14197 36128
rect 14231 36125 14243 36159
rect 14185 36119 14243 36125
rect 14369 36159 14427 36165
rect 14369 36125 14381 36159
rect 14415 36125 14427 36159
rect 14369 36119 14427 36125
rect 14458 36116 14464 36168
rect 14516 36116 14522 36168
rect 14553 36159 14611 36165
rect 14553 36125 14565 36159
rect 14599 36156 14611 36159
rect 15194 36156 15200 36168
rect 14599 36128 15200 36156
rect 14599 36125 14611 36128
rect 14553 36119 14611 36125
rect 15194 36116 15200 36128
rect 15252 36116 15258 36168
rect 15289 36159 15347 36165
rect 15289 36125 15301 36159
rect 15335 36156 15347 36159
rect 15746 36156 15752 36168
rect 15335 36128 15752 36156
rect 15335 36125 15347 36128
rect 15289 36119 15347 36125
rect 15746 36116 15752 36128
rect 15804 36116 15810 36168
rect 16298 36116 16304 36168
rect 16356 36116 16362 36168
rect 16758 36116 16764 36168
rect 16816 36156 16822 36168
rect 17420 36156 17448 36187
rect 18782 36184 18788 36196
rect 18840 36184 18846 36236
rect 16816 36128 17448 36156
rect 18693 36159 18751 36165
rect 16816 36116 16822 36128
rect 18693 36125 18705 36159
rect 18739 36156 18751 36159
rect 19260 36156 19288 36255
rect 21266 36252 21272 36304
rect 21324 36252 21330 36304
rect 21453 36295 21511 36301
rect 21453 36261 21465 36295
rect 21499 36261 21511 36295
rect 21453 36255 21511 36261
rect 19794 36184 19800 36236
rect 19852 36184 19858 36236
rect 18739 36128 19288 36156
rect 18739 36125 18751 36128
rect 18693 36119 18751 36125
rect 19610 36116 19616 36168
rect 19668 36156 19674 36168
rect 21177 36159 21235 36165
rect 21177 36156 21189 36159
rect 19668 36128 21189 36156
rect 19668 36116 19674 36128
rect 21177 36125 21189 36128
rect 21223 36156 21235 36159
rect 21284 36156 21312 36252
rect 21223 36128 21312 36156
rect 21468 36156 21496 36255
rect 21910 36224 21916 36236
rect 21652 36196 21916 36224
rect 21545 36159 21603 36165
rect 21545 36156 21557 36159
rect 21468 36128 21557 36156
rect 21223 36125 21235 36128
rect 21177 36119 21235 36125
rect 21545 36125 21557 36128
rect 21591 36125 21603 36159
rect 21545 36119 21603 36125
rect 13832 36060 15167 36088
rect 13725 36051 13783 36057
rect 11238 35980 11244 36032
rect 11296 35980 11302 36032
rect 12618 35980 12624 36032
rect 12676 36020 12682 36032
rect 13740 36020 13768 36051
rect 12676 35992 13768 36020
rect 12676 35980 12682 35992
rect 14918 35980 14924 36032
rect 14976 35980 14982 36032
rect 15139 36020 15167 36060
rect 15304 36060 19840 36088
rect 15304 36020 15332 36060
rect 15139 35992 15332 36020
rect 17126 35980 17132 36032
rect 17184 35980 17190 36032
rect 19702 35980 19708 36032
rect 19760 35980 19766 36032
rect 19812 36020 19840 36060
rect 20990 36048 20996 36100
rect 21048 36088 21054 36100
rect 21269 36091 21327 36097
rect 21269 36088 21281 36091
rect 21048 36060 21281 36088
rect 21048 36048 21054 36060
rect 21269 36057 21281 36060
rect 21315 36057 21327 36091
rect 21269 36051 21327 36057
rect 21453 36091 21511 36097
rect 21453 36057 21465 36091
rect 21499 36088 21511 36091
rect 21652 36088 21680 36196
rect 21910 36184 21916 36196
rect 21968 36224 21974 36236
rect 25332 36233 25360 36320
rect 25317 36227 25375 36233
rect 21968 36196 22968 36224
rect 21968 36184 21974 36196
rect 21729 36159 21787 36165
rect 21729 36125 21741 36159
rect 21775 36156 21787 36159
rect 22094 36156 22100 36168
rect 21775 36128 22100 36156
rect 21775 36125 21787 36128
rect 21729 36119 21787 36125
rect 22094 36116 22100 36128
rect 22152 36116 22158 36168
rect 22940 36165 22968 36196
rect 25317 36193 25329 36227
rect 25363 36193 25375 36227
rect 25317 36187 25375 36193
rect 25406 36184 25412 36236
rect 25464 36184 25470 36236
rect 25884 36196 28856 36224
rect 22925 36159 22983 36165
rect 22925 36125 22937 36159
rect 22971 36125 22983 36159
rect 22925 36119 22983 36125
rect 25682 36116 25688 36168
rect 25740 36116 25746 36168
rect 21499 36060 21680 36088
rect 22741 36091 22799 36097
rect 21499 36057 21511 36060
rect 21453 36051 21511 36057
rect 22741 36057 22753 36091
rect 22787 36088 22799 36091
rect 22830 36088 22836 36100
rect 22787 36060 22836 36088
rect 22787 36057 22799 36060
rect 22741 36051 22799 36057
rect 22830 36048 22836 36060
rect 22888 36048 22894 36100
rect 25884 36088 25912 36196
rect 25961 36159 26019 36165
rect 25961 36125 25973 36159
rect 26007 36156 26019 36159
rect 26050 36156 26056 36168
rect 26007 36128 26056 36156
rect 26007 36125 26019 36128
rect 25961 36119 26019 36125
rect 26050 36116 26056 36128
rect 26108 36116 26114 36168
rect 27798 36116 27804 36168
rect 27856 36156 27862 36168
rect 28276 36165 28304 36196
rect 28077 36159 28135 36165
rect 28077 36156 28089 36159
rect 27856 36128 28089 36156
rect 27856 36116 27862 36128
rect 28077 36125 28089 36128
rect 28123 36125 28135 36159
rect 28077 36119 28135 36125
rect 28261 36159 28319 36165
rect 28261 36125 28273 36159
rect 28307 36125 28319 36159
rect 28261 36119 28319 36125
rect 28626 36116 28632 36168
rect 28684 36116 28690 36168
rect 28828 36165 28856 36196
rect 28813 36159 28871 36165
rect 28813 36125 28825 36159
rect 28859 36125 28871 36159
rect 28813 36119 28871 36125
rect 23032 36060 25912 36088
rect 23032 36020 23060 36060
rect 19812 35992 23060 36020
rect 23106 35980 23112 36032
rect 23164 35980 23170 36032
rect 25222 35980 25228 36032
rect 25280 35980 25286 36032
rect 25777 36023 25835 36029
rect 25777 35989 25789 36023
rect 25823 36020 25835 36023
rect 25866 36020 25872 36032
rect 25823 35992 25872 36020
rect 25823 35989 25835 35992
rect 25777 35983 25835 35989
rect 25866 35980 25872 35992
rect 25924 35980 25930 36032
rect 1104 35930 38272 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 38272 35930
rect 1104 35856 38272 35878
rect 9766 35776 9772 35828
rect 9824 35816 9830 35828
rect 10045 35819 10103 35825
rect 10045 35816 10057 35819
rect 9824 35788 10057 35816
rect 9824 35776 9830 35788
rect 10045 35785 10057 35788
rect 10091 35785 10103 35819
rect 10045 35779 10103 35785
rect 10597 35819 10655 35825
rect 10597 35785 10609 35819
rect 10643 35785 10655 35819
rect 10597 35779 10655 35785
rect 10965 35819 11023 35825
rect 10965 35785 10977 35819
rect 11011 35816 11023 35819
rect 11238 35816 11244 35828
rect 11011 35788 11244 35816
rect 11011 35785 11023 35788
rect 10965 35779 11023 35785
rect 9858 35748 9864 35760
rect 9706 35720 9864 35748
rect 9858 35708 9864 35720
rect 9916 35708 9922 35760
rect 8202 35640 8208 35692
rect 8260 35640 8266 35692
rect 10229 35683 10287 35689
rect 10229 35649 10241 35683
rect 10275 35680 10287 35683
rect 10612 35680 10640 35779
rect 11238 35776 11244 35788
rect 11296 35776 11302 35828
rect 12618 35816 12624 35828
rect 11348 35788 12624 35816
rect 11348 35680 11376 35788
rect 12618 35776 12624 35788
rect 12676 35776 12682 35828
rect 12710 35776 12716 35828
rect 12768 35816 12774 35828
rect 13354 35816 13360 35828
rect 12768 35788 13360 35816
rect 12768 35776 12774 35788
rect 13354 35776 13360 35788
rect 13412 35776 13418 35828
rect 16574 35816 16580 35828
rect 16316 35788 16580 35816
rect 12897 35751 12955 35757
rect 12897 35748 12909 35751
rect 11992 35720 12909 35748
rect 11992 35689 12020 35720
rect 12897 35717 12909 35720
rect 12943 35748 12955 35751
rect 13446 35748 13452 35760
rect 12943 35720 13452 35748
rect 12943 35717 12955 35720
rect 12897 35711 12955 35717
rect 10275 35652 10640 35680
rect 10704 35652 11376 35680
rect 11977 35683 12035 35689
rect 10275 35649 10287 35652
rect 10229 35643 10287 35649
rect 8481 35615 8539 35621
rect 8481 35581 8493 35615
rect 8527 35612 8539 35615
rect 8938 35612 8944 35624
rect 8527 35584 8944 35612
rect 8527 35581 8539 35584
rect 8481 35575 8539 35581
rect 8938 35572 8944 35584
rect 8996 35572 9002 35624
rect 9950 35572 9956 35624
rect 10008 35612 10014 35624
rect 10704 35612 10732 35652
rect 11977 35649 11989 35683
rect 12023 35649 12035 35683
rect 11977 35643 12035 35649
rect 12253 35683 12311 35689
rect 12253 35649 12265 35683
rect 12299 35680 12311 35683
rect 12299 35652 12333 35680
rect 12299 35649 12311 35652
rect 12253 35643 12311 35649
rect 10008 35584 10732 35612
rect 10008 35572 10014 35584
rect 11054 35572 11060 35624
rect 11112 35572 11118 35624
rect 11149 35615 11207 35621
rect 11149 35581 11161 35615
rect 11195 35581 11207 35615
rect 11149 35575 11207 35581
rect 11164 35544 11192 35575
rect 11238 35572 11244 35624
rect 11296 35612 11302 35624
rect 12268 35612 12296 35643
rect 12434 35640 12440 35692
rect 12492 35680 12498 35692
rect 12713 35683 12771 35689
rect 12713 35680 12725 35683
rect 12492 35652 12725 35680
rect 12492 35640 12498 35652
rect 12713 35649 12725 35652
rect 12759 35680 12771 35683
rect 13081 35683 13139 35689
rect 12759 35652 13032 35680
rect 12759 35649 12771 35652
rect 12713 35643 12771 35649
rect 13004 35624 13032 35652
rect 13081 35649 13093 35683
rect 13127 35649 13139 35683
rect 13081 35643 13139 35649
rect 13275 35683 13333 35689
rect 13275 35649 13287 35683
rect 13321 35680 13333 35683
rect 13372 35680 13400 35720
rect 13446 35708 13452 35720
rect 13504 35708 13510 35760
rect 15838 35748 15844 35760
rect 15686 35720 15844 35748
rect 15838 35708 15844 35720
rect 15896 35708 15902 35760
rect 16316 35757 16344 35788
rect 16574 35776 16580 35788
rect 16632 35816 16638 35828
rect 17313 35819 17371 35825
rect 17313 35816 17325 35819
rect 16632 35788 17325 35816
rect 16632 35776 16638 35788
rect 17313 35785 17325 35788
rect 17359 35785 17371 35819
rect 17313 35779 17371 35785
rect 16285 35751 16344 35757
rect 16285 35717 16297 35751
rect 16331 35720 16344 35751
rect 16331 35717 16343 35720
rect 16285 35711 16343 35717
rect 16390 35708 16396 35760
rect 16448 35748 16454 35760
rect 16485 35751 16543 35757
rect 16485 35748 16497 35751
rect 16448 35720 16497 35748
rect 16448 35708 16454 35720
rect 16485 35717 16497 35720
rect 16531 35748 16543 35751
rect 17328 35748 17356 35779
rect 18046 35776 18052 35828
rect 18104 35816 18110 35828
rect 18141 35819 18199 35825
rect 18141 35816 18153 35819
rect 18104 35788 18153 35816
rect 18104 35776 18110 35788
rect 18141 35785 18153 35788
rect 18187 35785 18199 35819
rect 18141 35779 18199 35785
rect 19610 35776 19616 35828
rect 19668 35776 19674 35828
rect 25130 35816 25136 35828
rect 19812 35788 25136 35816
rect 16531 35720 16988 35748
rect 17328 35720 17908 35748
rect 16531 35717 16543 35720
rect 16485 35711 16543 35717
rect 16960 35689 16988 35720
rect 17880 35689 17908 35720
rect 13321 35652 13400 35680
rect 16945 35683 17003 35689
rect 13321 35649 13333 35652
rect 13275 35643 13333 35649
rect 16945 35649 16957 35683
rect 16991 35649 17003 35683
rect 16945 35643 17003 35649
rect 17037 35683 17095 35689
rect 17037 35649 17049 35683
rect 17083 35680 17095 35683
rect 17497 35683 17555 35689
rect 17083 35652 17448 35680
rect 17083 35649 17095 35652
rect 17037 35643 17095 35649
rect 12526 35612 12532 35624
rect 11296 35584 12532 35612
rect 11296 35572 11302 35584
rect 12526 35572 12532 35584
rect 12584 35572 12590 35624
rect 12986 35572 12992 35624
rect 13044 35572 13050 35624
rect 13096 35612 13124 35643
rect 13096 35584 13676 35612
rect 10704 35516 11192 35544
rect 10704 35488 10732 35516
rect 11790 35504 11796 35556
rect 11848 35544 11854 35556
rect 12069 35547 12127 35553
rect 12069 35544 12081 35547
rect 11848 35516 12081 35544
rect 11848 35504 11854 35516
rect 12069 35513 12081 35516
rect 12115 35513 12127 35547
rect 12069 35507 12127 35513
rect 10686 35436 10692 35488
rect 10744 35436 10750 35488
rect 11882 35436 11888 35488
rect 11940 35436 11946 35488
rect 12342 35436 12348 35488
rect 12400 35476 12406 35488
rect 13096 35476 13124 35584
rect 13648 35556 13676 35584
rect 14182 35572 14188 35624
rect 14240 35572 14246 35624
rect 14458 35572 14464 35624
rect 14516 35572 14522 35624
rect 16850 35572 16856 35624
rect 16908 35572 16914 35624
rect 17129 35615 17187 35621
rect 17129 35612 17141 35615
rect 16960 35584 17141 35612
rect 13630 35504 13636 35556
rect 13688 35504 13694 35556
rect 16960 35544 16988 35584
rect 17129 35581 17141 35584
rect 17175 35581 17187 35615
rect 17420 35612 17448 35652
rect 17497 35649 17509 35683
rect 17543 35680 17555 35683
rect 17865 35683 17923 35689
rect 17543 35652 17816 35680
rect 17543 35649 17555 35652
rect 17497 35643 17555 35649
rect 17678 35612 17684 35624
rect 17420 35584 17684 35612
rect 17129 35575 17187 35581
rect 17678 35572 17684 35584
rect 17736 35572 17742 35624
rect 17788 35612 17816 35652
rect 17865 35649 17877 35683
rect 17911 35649 17923 35683
rect 17865 35643 17923 35649
rect 18046 35640 18052 35692
rect 18104 35640 18110 35692
rect 18509 35683 18567 35689
rect 18509 35649 18521 35683
rect 18555 35680 18567 35683
rect 18874 35680 18880 35692
rect 18555 35652 18880 35680
rect 18555 35649 18567 35652
rect 18509 35643 18567 35649
rect 18874 35640 18880 35652
rect 18932 35640 18938 35692
rect 19628 35680 19656 35776
rect 19705 35683 19763 35689
rect 19705 35680 19717 35683
rect 19628 35652 19717 35680
rect 19705 35649 19717 35652
rect 19751 35649 19763 35683
rect 19705 35643 19763 35649
rect 17957 35615 18015 35621
rect 17788 35584 17908 35612
rect 17880 35556 17908 35584
rect 17957 35581 17969 35615
rect 18003 35612 18015 35615
rect 18601 35615 18659 35621
rect 18601 35612 18613 35615
rect 18003 35584 18613 35612
rect 18003 35581 18015 35584
rect 17957 35575 18015 35581
rect 18601 35581 18613 35584
rect 18647 35581 18659 35615
rect 18601 35575 18659 35581
rect 18782 35572 18788 35624
rect 18840 35572 18846 35624
rect 15948 35516 16988 35544
rect 12400 35448 13124 35476
rect 12400 35436 12406 35448
rect 13170 35436 13176 35488
rect 13228 35436 13234 35488
rect 15746 35436 15752 35488
rect 15804 35476 15810 35488
rect 15948 35485 15976 35516
rect 15933 35479 15991 35485
rect 15933 35476 15945 35479
rect 15804 35448 15945 35476
rect 15804 35436 15810 35448
rect 15933 35445 15945 35448
rect 15979 35445 15991 35479
rect 15933 35439 15991 35445
rect 16114 35436 16120 35488
rect 16172 35436 16178 35488
rect 16316 35485 16344 35516
rect 17862 35504 17868 35556
rect 17920 35544 17926 35556
rect 19812 35544 19840 35788
rect 25130 35776 25136 35788
rect 25188 35816 25194 35828
rect 25593 35819 25651 35825
rect 25593 35816 25605 35819
rect 25188 35788 25605 35816
rect 25188 35776 25194 35788
rect 25593 35785 25605 35788
rect 25639 35785 25651 35819
rect 25593 35779 25651 35785
rect 22094 35708 22100 35760
rect 22152 35708 22158 35760
rect 25682 35748 25688 35760
rect 25056 35720 25688 35748
rect 22112 35680 22140 35708
rect 22649 35683 22707 35689
rect 22649 35680 22661 35683
rect 22112 35652 22661 35680
rect 22649 35649 22661 35652
rect 22695 35680 22707 35683
rect 22738 35680 22744 35692
rect 22695 35652 22744 35680
rect 22695 35649 22707 35652
rect 22649 35643 22707 35649
rect 22738 35640 22744 35652
rect 22796 35640 22802 35692
rect 22462 35572 22468 35624
rect 22520 35572 22526 35624
rect 25056 35621 25084 35720
rect 25682 35708 25688 35720
rect 25740 35757 25746 35760
rect 25740 35751 25803 35757
rect 25740 35717 25757 35751
rect 25791 35717 25803 35751
rect 25740 35711 25803 35717
rect 25740 35708 25746 35711
rect 25866 35708 25872 35760
rect 25924 35748 25930 35760
rect 25961 35751 26019 35757
rect 25961 35748 25973 35751
rect 25924 35720 25973 35748
rect 25924 35708 25930 35720
rect 25961 35717 25973 35720
rect 26007 35717 26019 35751
rect 25961 35711 26019 35717
rect 25130 35640 25136 35692
rect 25188 35680 25194 35692
rect 25884 35680 25912 35708
rect 25188 35652 25912 35680
rect 25188 35640 25194 35652
rect 37642 35640 37648 35692
rect 37700 35640 37706 35692
rect 25041 35615 25099 35621
rect 25041 35612 25053 35615
rect 22848 35584 25053 35612
rect 17920 35516 19840 35544
rect 17920 35504 17926 35516
rect 16301 35479 16359 35485
rect 16301 35445 16313 35479
rect 16347 35445 16359 35479
rect 16301 35439 16359 35445
rect 16482 35436 16488 35488
rect 16540 35476 16546 35488
rect 16669 35479 16727 35485
rect 16669 35476 16681 35479
rect 16540 35448 16681 35476
rect 16540 35436 16546 35448
rect 16669 35445 16681 35448
rect 16715 35445 16727 35479
rect 16669 35439 16727 35445
rect 17678 35436 17684 35488
rect 17736 35476 17742 35488
rect 18138 35476 18144 35488
rect 17736 35448 18144 35476
rect 17736 35436 17742 35448
rect 18138 35436 18144 35448
rect 18196 35436 18202 35488
rect 19610 35436 19616 35488
rect 19668 35436 19674 35488
rect 22646 35436 22652 35488
rect 22704 35476 22710 35488
rect 22848 35485 22876 35584
rect 25041 35581 25053 35584
rect 25087 35581 25099 35615
rect 25041 35575 25099 35581
rect 22833 35479 22891 35485
rect 22833 35476 22845 35479
rect 22704 35448 22845 35476
rect 22704 35436 22710 35448
rect 22833 35445 22845 35448
rect 22879 35445 22891 35479
rect 22833 35439 22891 35445
rect 25498 35436 25504 35488
rect 25556 35436 25562 35488
rect 25777 35479 25835 35485
rect 25777 35445 25789 35479
rect 25823 35476 25835 35479
rect 26050 35476 26056 35488
rect 25823 35448 26056 35476
rect 25823 35445 25835 35448
rect 25777 35439 25835 35445
rect 26050 35436 26056 35448
rect 26108 35436 26114 35488
rect 37826 35436 37832 35488
rect 37884 35436 37890 35488
rect 1104 35386 38272 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38272 35386
rect 1104 35312 38272 35334
rect 8938 35232 8944 35284
rect 8996 35232 9002 35284
rect 9950 35232 9956 35284
rect 10008 35232 10014 35284
rect 11054 35232 11060 35284
rect 11112 35272 11118 35284
rect 11333 35275 11391 35281
rect 11333 35272 11345 35275
rect 11112 35244 11345 35272
rect 11112 35232 11118 35244
rect 11333 35241 11345 35244
rect 11379 35241 11391 35275
rect 11333 35235 11391 35241
rect 11790 35232 11796 35284
rect 11848 35232 11854 35284
rect 11882 35232 11888 35284
rect 11940 35232 11946 35284
rect 12434 35232 12440 35284
rect 12492 35232 12498 35284
rect 12618 35232 12624 35284
rect 12676 35232 12682 35284
rect 13354 35232 13360 35284
rect 13412 35232 13418 35284
rect 14458 35232 14464 35284
rect 14516 35272 14522 35284
rect 14645 35275 14703 35281
rect 14645 35272 14657 35275
rect 14516 35244 14657 35272
rect 14516 35232 14522 35244
rect 14645 35241 14657 35244
rect 14691 35241 14703 35275
rect 14645 35235 14703 35241
rect 15378 35232 15384 35284
rect 15436 35272 15442 35284
rect 16393 35275 16451 35281
rect 16393 35272 16405 35275
rect 15436 35244 16405 35272
rect 15436 35232 15442 35244
rect 16393 35241 16405 35244
rect 16439 35241 16451 35275
rect 16393 35235 16451 35241
rect 16850 35232 16856 35284
rect 16908 35272 16914 35284
rect 17862 35272 17868 35284
rect 16908 35244 17868 35272
rect 16908 35232 16914 35244
rect 17862 35232 17868 35244
rect 17920 35232 17926 35284
rect 17957 35275 18015 35281
rect 17957 35241 17969 35275
rect 18003 35272 18015 35275
rect 18046 35272 18052 35284
rect 18003 35244 18052 35272
rect 18003 35241 18015 35244
rect 17957 35235 18015 35241
rect 18046 35232 18052 35244
rect 18104 35232 18110 35284
rect 19702 35232 19708 35284
rect 19760 35272 19766 35284
rect 19981 35275 20039 35281
rect 19981 35272 19993 35275
rect 19760 35244 19993 35272
rect 19760 35232 19766 35244
rect 19981 35241 19993 35244
rect 20027 35241 20039 35275
rect 19981 35235 20039 35241
rect 20717 35275 20775 35281
rect 20717 35241 20729 35275
rect 20763 35272 20775 35275
rect 23382 35272 23388 35284
rect 20763 35244 23388 35272
rect 20763 35241 20775 35244
rect 20717 35235 20775 35241
rect 23382 35232 23388 35244
rect 23440 35232 23446 35284
rect 25498 35232 25504 35284
rect 25556 35232 25562 35284
rect 37553 35275 37611 35281
rect 37553 35241 37565 35275
rect 37599 35272 37611 35275
rect 37642 35272 37648 35284
rect 37599 35244 37648 35272
rect 37599 35241 37611 35244
rect 37553 35235 37611 35241
rect 37642 35232 37648 35244
rect 37700 35232 37706 35284
rect 9968 35204 9996 35232
rect 9784 35176 9996 35204
rect 9784 35077 9812 35176
rect 10045 35139 10103 35145
rect 10045 35105 10057 35139
rect 10091 35136 10103 35139
rect 10686 35136 10692 35148
rect 10091 35108 10692 35136
rect 10091 35105 10103 35108
rect 10045 35099 10103 35105
rect 10686 35096 10692 35108
rect 10744 35096 10750 35148
rect 11808 35136 11836 35232
rect 11532 35108 11836 35136
rect 11532 35077 11560 35108
rect 9125 35071 9183 35077
rect 9125 35037 9137 35071
rect 9171 35068 9183 35071
rect 9769 35071 9827 35077
rect 9171 35040 9444 35068
rect 9171 35037 9183 35040
rect 9125 35031 9183 35037
rect 934 34960 940 35012
rect 992 35000 998 35012
rect 1489 35003 1547 35009
rect 1489 35000 1501 35003
rect 992 34972 1501 35000
rect 992 34960 998 34972
rect 1489 34969 1501 34972
rect 1535 34969 1547 35003
rect 1489 34963 1547 34969
rect 1673 35003 1731 35009
rect 1673 34969 1685 35003
rect 1719 35000 1731 35003
rect 5994 35000 6000 35012
rect 1719 34972 6000 35000
rect 1719 34969 1731 34972
rect 1673 34963 1731 34969
rect 5994 34960 6000 34972
rect 6052 34960 6058 35012
rect 9416 34941 9444 35040
rect 9769 35037 9781 35071
rect 9815 35037 9827 35071
rect 9769 35031 9827 35037
rect 11517 35071 11575 35077
rect 11517 35037 11529 35071
rect 11563 35037 11575 35071
rect 11517 35031 11575 35037
rect 11609 35071 11667 35077
rect 11609 35037 11621 35071
rect 11655 35068 11667 35071
rect 11900 35068 11928 35232
rect 12253 35139 12311 35145
rect 12253 35105 12265 35139
rect 12299 35136 12311 35139
rect 12452 35136 12480 35232
rect 12299 35108 12480 35136
rect 12529 35139 12587 35145
rect 12299 35105 12311 35108
rect 12253 35099 12311 35105
rect 12529 35105 12541 35139
rect 12575 35136 12587 35139
rect 12636 35136 12664 35232
rect 16758 35204 16764 35216
rect 13004 35176 16764 35204
rect 12894 35136 12900 35148
rect 12575 35108 12900 35136
rect 12575 35105 12587 35108
rect 12529 35099 12587 35105
rect 12894 35096 12900 35108
rect 12952 35096 12958 35148
rect 13004 35080 13032 35176
rect 16758 35164 16764 35176
rect 16816 35164 16822 35216
rect 18782 35164 18788 35216
rect 18840 35204 18846 35216
rect 18840 35176 21772 35204
rect 18840 35164 18846 35176
rect 13262 35136 13268 35148
rect 13096 35108 13268 35136
rect 11655 35040 11928 35068
rect 11655 35037 11667 35040
rect 11609 35031 11667 35037
rect 11974 35028 11980 35080
rect 12032 35028 12038 35080
rect 12342 35028 12348 35080
rect 12400 35028 12406 35080
rect 12434 35028 12440 35080
rect 12492 35028 12498 35080
rect 12713 35071 12771 35077
rect 12713 35037 12725 35071
rect 12759 35037 12771 35071
rect 12713 35031 12771 35037
rect 11698 34960 11704 35012
rect 11756 34960 11762 35012
rect 11839 35003 11897 35009
rect 11839 34969 11851 35003
rect 11885 35000 11897 35003
rect 11885 34972 12480 35000
rect 11885 34969 11897 34972
rect 11839 34963 11897 34969
rect 9401 34935 9459 34941
rect 9401 34901 9413 34935
rect 9447 34901 9459 34935
rect 9401 34895 9459 34901
rect 9858 34892 9864 34944
rect 9916 34892 9922 34944
rect 11606 34892 11612 34944
rect 11664 34932 11670 34944
rect 12069 34935 12127 34941
rect 12069 34932 12081 34935
rect 11664 34904 12081 34932
rect 11664 34892 11670 34904
rect 12069 34901 12081 34904
rect 12115 34901 12127 34935
rect 12452 34932 12480 34972
rect 12526 34960 12532 35012
rect 12584 35000 12590 35012
rect 12728 35000 12756 35031
rect 12986 35028 12992 35080
rect 13044 35028 13050 35080
rect 13096 35077 13124 35108
rect 13262 35096 13268 35108
rect 13320 35096 13326 35148
rect 15838 35096 15844 35148
rect 15896 35136 15902 35148
rect 16117 35139 16175 35145
rect 16117 35136 16129 35139
rect 15896 35108 16129 35136
rect 15896 35096 15902 35108
rect 16117 35105 16129 35108
rect 16163 35105 16175 35139
rect 19334 35136 19340 35148
rect 16117 35099 16175 35105
rect 16224 35108 18092 35136
rect 13081 35071 13139 35077
rect 13081 35037 13093 35071
rect 13127 35037 13139 35071
rect 13081 35031 13139 35037
rect 13173 35071 13231 35077
rect 13173 35037 13185 35071
rect 13219 35068 13231 35071
rect 13219 35040 13400 35068
rect 13219 35037 13231 35040
rect 13173 35031 13231 35037
rect 12584 34972 12756 35000
rect 12871 35003 12929 35009
rect 12584 34960 12590 34972
rect 12871 34969 12883 35003
rect 12917 34969 12929 35003
rect 13372 35000 13400 35040
rect 13446 35028 13452 35080
rect 13504 35028 13510 35080
rect 13817 35071 13875 35077
rect 13817 35068 13829 35071
rect 13556 35040 13829 35068
rect 13556 35000 13584 35040
rect 13817 35037 13829 35040
rect 13863 35037 13875 35071
rect 13817 35031 13875 35037
rect 14829 35071 14887 35077
rect 14829 35037 14841 35071
rect 14875 35068 14887 35071
rect 14918 35068 14924 35080
rect 14875 35040 14924 35068
rect 14875 35037 14887 35040
rect 14829 35031 14887 35037
rect 14918 35028 14924 35040
rect 14976 35028 14982 35080
rect 16224 35068 16252 35108
rect 15028 35040 16252 35068
rect 13372 34972 13584 35000
rect 12871 34963 12929 34969
rect 12710 34932 12716 34944
rect 12452 34904 12716 34932
rect 12069 34895 12127 34901
rect 12710 34892 12716 34904
rect 12768 34932 12774 34944
rect 12886 34932 12914 34963
rect 13630 34960 13636 35012
rect 13688 35000 13694 35012
rect 14550 35000 14556 35012
rect 13688 34972 14556 35000
rect 13688 34960 13694 34972
rect 14550 34960 14556 34972
rect 14608 35000 14614 35012
rect 15028 35000 15056 35040
rect 16574 35028 16580 35080
rect 16632 35028 16638 35080
rect 16758 35028 16764 35080
rect 16816 35028 16822 35080
rect 17037 35071 17095 35077
rect 17037 35037 17049 35071
rect 17083 35037 17095 35071
rect 17037 35031 17095 35037
rect 14608 34972 15056 35000
rect 14608 34960 14614 34972
rect 15286 34960 15292 35012
rect 15344 35000 15350 35012
rect 15381 35003 15439 35009
rect 15381 35000 15393 35003
rect 15344 34972 15393 35000
rect 15344 34960 15350 34972
rect 15381 34969 15393 34972
rect 15427 34969 15439 35003
rect 15381 34963 15439 34969
rect 16666 34960 16672 35012
rect 16724 34960 16730 35012
rect 16850 34960 16856 35012
rect 16908 35009 16914 35012
rect 16908 35003 16937 35009
rect 16925 34969 16937 35003
rect 17052 35000 17080 35031
rect 17862 35028 17868 35080
rect 17920 35068 17926 35080
rect 17957 35071 18015 35077
rect 17957 35068 17969 35071
rect 17920 35040 17969 35068
rect 17920 35028 17926 35040
rect 17957 35037 17969 35040
rect 18003 35037 18015 35071
rect 17957 35031 18015 35037
rect 18064 35000 18092 35108
rect 18892 35108 19340 35136
rect 18138 35028 18144 35080
rect 18196 35028 18202 35080
rect 18230 35028 18236 35080
rect 18288 35068 18294 35080
rect 18892 35077 18920 35108
rect 19334 35096 19340 35108
rect 19392 35096 19398 35148
rect 19444 35145 19472 35176
rect 21744 35148 21772 35176
rect 22462 35164 22468 35216
rect 22520 35204 22526 35216
rect 22520 35176 22968 35204
rect 22520 35164 22526 35176
rect 19429 35139 19487 35145
rect 19429 35105 19441 35139
rect 19475 35105 19487 35139
rect 19429 35099 19487 35105
rect 19521 35139 19579 35145
rect 19521 35105 19533 35139
rect 19567 35136 19579 35139
rect 19610 35136 19616 35148
rect 19567 35108 19616 35136
rect 19567 35105 19579 35108
rect 19521 35099 19579 35105
rect 18877 35071 18935 35077
rect 18877 35068 18889 35071
rect 18288 35040 18889 35068
rect 18288 35028 18294 35040
rect 18877 35037 18889 35040
rect 18923 35037 18935 35071
rect 18877 35031 18935 35037
rect 19061 35071 19119 35077
rect 19061 35037 19073 35071
rect 19107 35068 19119 35071
rect 19536 35068 19564 35099
rect 19610 35096 19616 35108
rect 19668 35096 19674 35148
rect 20530 35136 20536 35148
rect 20088 35108 20536 35136
rect 20088 35077 20116 35108
rect 20530 35096 20536 35108
rect 20588 35096 20594 35148
rect 21726 35096 21732 35148
rect 21784 35096 21790 35148
rect 22833 35139 22891 35145
rect 22833 35136 22845 35139
rect 22480 35108 22845 35136
rect 19107 35040 19564 35068
rect 20073 35071 20131 35077
rect 19107 35037 19119 35040
rect 19061 35031 19119 35037
rect 20073 35037 20085 35071
rect 20119 35037 20131 35071
rect 20073 35031 20131 35037
rect 20254 35028 20260 35080
rect 20312 35028 20318 35080
rect 20346 35028 20352 35080
rect 20404 35028 20410 35080
rect 20441 35071 20499 35077
rect 20441 35037 20453 35071
rect 20487 35037 20499 35071
rect 20441 35031 20499 35037
rect 20456 35000 20484 35031
rect 21174 35028 21180 35080
rect 21232 35028 21238 35080
rect 22480 35077 22508 35108
rect 22833 35105 22845 35108
rect 22879 35105 22891 35139
rect 22833 35099 22891 35105
rect 22465 35071 22523 35077
rect 22465 35037 22477 35071
rect 22511 35037 22523 35071
rect 22465 35031 22523 35037
rect 22646 35028 22652 35080
rect 22704 35028 22710 35080
rect 22738 35028 22744 35080
rect 22796 35028 22802 35080
rect 22940 35077 22968 35176
rect 23750 35096 23756 35148
rect 23808 35136 23814 35148
rect 24949 35139 25007 35145
rect 24949 35136 24961 35139
rect 23808 35108 24961 35136
rect 23808 35096 23814 35108
rect 24949 35105 24961 35108
rect 24995 35105 25007 35139
rect 24949 35099 25007 35105
rect 25406 35096 25412 35148
rect 25464 35096 25470 35148
rect 25516 35136 25544 35232
rect 25685 35139 25743 35145
rect 25685 35136 25697 35139
rect 25516 35108 25697 35136
rect 25685 35105 25697 35108
rect 25731 35105 25743 35139
rect 25685 35099 25743 35105
rect 25777 35139 25835 35145
rect 25777 35105 25789 35139
rect 25823 35105 25835 35139
rect 25777 35099 25835 35105
rect 22925 35071 22983 35077
rect 22925 35037 22937 35071
rect 22971 35037 22983 35071
rect 22925 35031 22983 35037
rect 24765 35071 24823 35077
rect 24765 35037 24777 35071
rect 24811 35068 24823 35071
rect 25130 35068 25136 35080
rect 24811 35040 25136 35068
rect 24811 35037 24823 35040
rect 24765 35031 24823 35037
rect 25130 35028 25136 35040
rect 25188 35028 25194 35080
rect 25424 35068 25452 35096
rect 25792 35068 25820 35099
rect 25424 35040 25820 35068
rect 37366 35028 37372 35080
rect 37424 35028 37430 35080
rect 17052 34972 17908 35000
rect 18064 34972 20484 35000
rect 21913 35003 21971 35009
rect 16908 34963 16937 34969
rect 16908 34960 16914 34963
rect 17880 34944 17908 34972
rect 21913 34969 21925 35003
rect 21959 35000 21971 35003
rect 22557 35003 22615 35009
rect 22557 35000 22569 35003
rect 21959 34972 22569 35000
rect 21959 34969 21971 34972
rect 21913 34963 21971 34969
rect 22557 34969 22569 34972
rect 22603 34969 22615 35003
rect 22557 34963 22615 34969
rect 12768 34904 12914 34932
rect 12768 34892 12774 34904
rect 17862 34892 17868 34944
rect 17920 34892 17926 34944
rect 19058 34892 19064 34944
rect 19116 34892 19122 34944
rect 19613 34935 19671 34941
rect 19613 34901 19625 34935
rect 19659 34932 19671 34935
rect 20162 34932 20168 34944
rect 19659 34904 20168 34932
rect 19659 34901 19671 34904
rect 19613 34895 19671 34901
rect 20162 34892 20168 34904
rect 20220 34892 20226 34944
rect 20990 34892 20996 34944
rect 21048 34892 21054 34944
rect 21266 34892 21272 34944
rect 21324 34932 21330 34944
rect 22005 34935 22063 34941
rect 22005 34932 22017 34935
rect 21324 34904 22017 34932
rect 21324 34892 21330 34904
rect 22005 34901 22017 34904
rect 22051 34901 22063 34935
rect 22005 34895 22063 34901
rect 22370 34892 22376 34944
rect 22428 34892 22434 34944
rect 24394 34892 24400 34944
rect 24452 34892 24458 34944
rect 24857 34935 24915 34941
rect 24857 34901 24869 34935
rect 24903 34932 24915 34935
rect 25225 34935 25283 34941
rect 25225 34932 25237 34935
rect 24903 34904 25237 34932
rect 24903 34901 24915 34904
rect 24857 34895 24915 34901
rect 25225 34901 25237 34904
rect 25271 34901 25283 34935
rect 25225 34895 25283 34901
rect 25590 34892 25596 34944
rect 25648 34892 25654 34944
rect 1104 34842 38272 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 38272 34842
rect 1104 34768 38272 34790
rect 9858 34688 9864 34740
rect 9916 34728 9922 34740
rect 11517 34731 11575 34737
rect 11517 34728 11529 34731
rect 9916 34700 11529 34728
rect 9916 34688 9922 34700
rect 11517 34697 11529 34700
rect 11563 34697 11575 34731
rect 11517 34691 11575 34697
rect 11698 34688 11704 34740
rect 11756 34728 11762 34740
rect 12973 34731 13031 34737
rect 11756 34700 12480 34728
rect 11756 34688 11762 34700
rect 11900 34669 11928 34700
rect 11241 34663 11299 34669
rect 11241 34629 11253 34663
rect 11287 34660 11299 34663
rect 11793 34663 11851 34669
rect 11793 34660 11805 34663
rect 11287 34632 11805 34660
rect 11287 34629 11299 34632
rect 11241 34623 11299 34629
rect 11793 34629 11805 34632
rect 11839 34629 11851 34663
rect 11793 34623 11851 34629
rect 11885 34663 11943 34669
rect 11885 34629 11897 34663
rect 11931 34629 11943 34663
rect 12342 34660 12348 34672
rect 11885 34623 11943 34629
rect 12176 34632 12348 34660
rect 11333 34595 11391 34601
rect 11333 34561 11345 34595
rect 11379 34561 11391 34595
rect 11333 34555 11391 34561
rect 11348 34388 11376 34555
rect 11606 34552 11612 34604
rect 11664 34592 11670 34604
rect 12176 34601 12204 34632
rect 12342 34620 12348 34632
rect 12400 34620 12406 34672
rect 12452 34669 12480 34700
rect 12973 34697 12985 34731
rect 13019 34728 13031 34731
rect 13446 34728 13452 34740
rect 13019 34700 13452 34728
rect 13019 34697 13031 34700
rect 12973 34691 13031 34697
rect 13446 34688 13452 34700
rect 13504 34688 13510 34740
rect 14366 34688 14372 34740
rect 14424 34688 14430 34740
rect 16209 34731 16267 34737
rect 16209 34697 16221 34731
rect 16255 34728 16267 34731
rect 16666 34728 16672 34740
rect 16255 34700 16672 34728
rect 16255 34697 16267 34700
rect 16209 34691 16267 34697
rect 16666 34688 16672 34700
rect 16724 34688 16730 34740
rect 20073 34731 20131 34737
rect 20073 34697 20085 34731
rect 20119 34728 20131 34731
rect 20254 34728 20260 34740
rect 20119 34700 20260 34728
rect 20119 34697 20131 34700
rect 20073 34691 20131 34697
rect 20254 34688 20260 34700
rect 20312 34688 20318 34740
rect 20346 34688 20352 34740
rect 20404 34688 20410 34740
rect 21174 34688 21180 34740
rect 21232 34728 21238 34740
rect 21821 34731 21879 34737
rect 21821 34728 21833 34731
rect 21232 34700 21833 34728
rect 21232 34688 21238 34700
rect 21821 34697 21833 34700
rect 21867 34697 21879 34731
rect 21821 34691 21879 34697
rect 22281 34731 22339 34737
rect 22281 34697 22293 34731
rect 22327 34728 22339 34731
rect 22370 34728 22376 34740
rect 22327 34700 22376 34728
rect 22327 34697 22339 34700
rect 22281 34691 22339 34697
rect 22370 34688 22376 34700
rect 22428 34688 22434 34740
rect 22462 34688 22468 34740
rect 22520 34688 22526 34740
rect 25041 34731 25099 34737
rect 25041 34697 25053 34731
rect 25087 34728 25099 34731
rect 25130 34728 25136 34740
rect 25087 34700 25136 34728
rect 25087 34697 25099 34700
rect 25041 34691 25099 34697
rect 25130 34688 25136 34700
rect 25188 34688 25194 34740
rect 26602 34688 26608 34740
rect 26660 34728 26666 34740
rect 27522 34728 27528 34740
rect 26660 34700 27528 34728
rect 26660 34688 26666 34700
rect 27522 34688 27528 34700
rect 27580 34728 27586 34740
rect 29733 34731 29791 34737
rect 29733 34728 29745 34731
rect 27580 34700 29745 34728
rect 27580 34688 27586 34700
rect 29733 34697 29745 34700
rect 29779 34728 29791 34731
rect 29779 34700 29960 34728
rect 29779 34697 29791 34700
rect 29733 34691 29791 34697
rect 12437 34663 12495 34669
rect 12437 34629 12449 34663
rect 12483 34660 12495 34663
rect 13173 34663 13231 34669
rect 12483 34632 13032 34660
rect 12483 34629 12495 34632
rect 12437 34623 12495 34629
rect 13004 34604 13032 34632
rect 13173 34629 13185 34663
rect 13219 34660 13231 34663
rect 13630 34660 13636 34672
rect 13219 34632 13636 34660
rect 13219 34629 13231 34632
rect 13173 34623 13231 34629
rect 13630 34620 13636 34632
rect 13688 34620 13694 34672
rect 14384 34660 14412 34688
rect 18230 34660 18236 34672
rect 14384 34632 18236 34660
rect 18230 34620 18236 34632
rect 18288 34620 18294 34672
rect 20364 34660 20392 34688
rect 19904 34632 20392 34660
rect 22189 34663 22247 34669
rect 11701 34595 11759 34601
rect 11701 34592 11713 34595
rect 11664 34564 11713 34592
rect 11664 34552 11670 34564
rect 11701 34561 11713 34564
rect 11747 34561 11759 34595
rect 11701 34555 11759 34561
rect 12023 34595 12081 34601
rect 12023 34561 12035 34595
rect 12069 34561 12081 34595
rect 12023 34555 12081 34561
rect 12161 34595 12219 34601
rect 12161 34561 12173 34595
rect 12207 34561 12219 34595
rect 12161 34555 12219 34561
rect 12038 34468 12066 34555
rect 12250 34552 12256 34604
rect 12308 34592 12314 34604
rect 12713 34595 12771 34601
rect 12713 34592 12725 34595
rect 12308 34564 12725 34592
rect 12308 34552 12314 34564
rect 12713 34561 12725 34564
rect 12759 34561 12771 34595
rect 12713 34555 12771 34561
rect 12986 34552 12992 34604
rect 13044 34552 13050 34604
rect 15286 34552 15292 34604
rect 15344 34552 15350 34604
rect 16114 34552 16120 34604
rect 16172 34552 16178 34604
rect 19904 34601 19932 34632
rect 22189 34629 22201 34663
rect 22235 34660 22247 34663
rect 22480 34660 22508 34688
rect 22235 34632 22508 34660
rect 22235 34629 22247 34632
rect 22189 34623 22247 34629
rect 24118 34620 24124 34672
rect 24176 34620 24182 34672
rect 29549 34663 29607 34669
rect 29549 34629 29561 34663
rect 29595 34660 29607 34663
rect 29595 34632 29776 34660
rect 29595 34629 29607 34632
rect 29549 34623 29607 34629
rect 19889 34595 19947 34601
rect 19889 34561 19901 34595
rect 19935 34561 19947 34595
rect 19889 34555 19947 34561
rect 19978 34552 19984 34604
rect 20036 34592 20042 34604
rect 20073 34595 20131 34601
rect 20073 34592 20085 34595
rect 20036 34564 20085 34592
rect 20036 34552 20042 34564
rect 20073 34561 20085 34564
rect 20119 34561 20131 34595
rect 20073 34555 20131 34561
rect 29362 34552 29368 34604
rect 29420 34552 29426 34604
rect 29641 34595 29699 34601
rect 29641 34592 29653 34595
rect 29564 34564 29653 34592
rect 15304 34524 15332 34552
rect 19426 34524 19432 34536
rect 15304 34496 19432 34524
rect 19426 34484 19432 34496
rect 19484 34524 19490 34536
rect 21450 34524 21456 34536
rect 19484 34496 21456 34524
rect 19484 34484 19490 34496
rect 21450 34484 21456 34496
rect 21508 34484 21514 34536
rect 22465 34527 22523 34533
rect 22465 34493 22477 34527
rect 22511 34493 22523 34527
rect 22465 34487 22523 34493
rect 11974 34416 11980 34468
rect 12032 34456 12066 34468
rect 12710 34456 12716 34468
rect 12032 34428 12716 34456
rect 12032 34416 12038 34428
rect 12710 34416 12716 34428
rect 12768 34456 12774 34468
rect 16850 34456 16856 34468
rect 12768 34428 16856 34456
rect 12768 34416 12774 34428
rect 16850 34416 16856 34428
rect 16908 34416 16914 34468
rect 12618 34388 12624 34400
rect 11348 34360 12624 34388
rect 12618 34348 12624 34360
rect 12676 34388 12682 34400
rect 12805 34391 12863 34397
rect 12805 34388 12817 34391
rect 12676 34360 12817 34388
rect 12676 34348 12682 34360
rect 12805 34357 12817 34360
rect 12851 34357 12863 34391
rect 12805 34351 12863 34357
rect 12894 34348 12900 34400
rect 12952 34388 12958 34400
rect 12989 34391 13047 34397
rect 12989 34388 13001 34391
rect 12952 34360 13001 34388
rect 12952 34348 12958 34360
rect 12989 34357 13001 34360
rect 13035 34357 13047 34391
rect 12989 34351 13047 34357
rect 15194 34348 15200 34400
rect 15252 34388 15258 34400
rect 18230 34388 18236 34400
rect 15252 34360 18236 34388
rect 15252 34348 15258 34360
rect 18230 34348 18236 34360
rect 18288 34348 18294 34400
rect 22480 34388 22508 34487
rect 23290 34484 23296 34536
rect 23348 34484 23354 34536
rect 23566 34484 23572 34536
rect 23624 34484 23630 34536
rect 28902 34484 28908 34536
rect 28960 34524 28966 34536
rect 29181 34527 29239 34533
rect 29181 34524 29193 34527
rect 28960 34496 29193 34524
rect 28960 34484 28966 34496
rect 29181 34493 29193 34496
rect 29227 34524 29239 34527
rect 29227 34496 29408 34524
rect 29227 34493 29239 34496
rect 29181 34487 29239 34493
rect 29380 34456 29408 34496
rect 29564 34456 29592 34564
rect 29641 34561 29653 34564
rect 29687 34561 29699 34595
rect 29641 34555 29699 34561
rect 29748 34524 29776 34632
rect 29822 34552 29828 34604
rect 29880 34552 29886 34604
rect 29932 34601 29960 34700
rect 29917 34595 29975 34601
rect 29917 34561 29929 34595
rect 29963 34561 29975 34595
rect 29917 34555 29975 34561
rect 30101 34595 30159 34601
rect 30101 34561 30113 34595
rect 30147 34561 30159 34595
rect 30101 34555 30159 34561
rect 30116 34524 30144 34555
rect 29748 34496 30144 34524
rect 29380 34428 29592 34456
rect 23750 34388 23756 34400
rect 22480 34360 23756 34388
rect 23750 34348 23756 34360
rect 23808 34348 23814 34400
rect 30098 34348 30104 34400
rect 30156 34348 30162 34400
rect 1104 34298 38272 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38272 34298
rect 1104 34224 38272 34246
rect 14734 34144 14740 34196
rect 14792 34144 14798 34196
rect 17862 34144 17868 34196
rect 17920 34144 17926 34196
rect 22462 34144 22468 34196
rect 22520 34144 22526 34196
rect 23566 34144 23572 34196
rect 23624 34184 23630 34196
rect 23753 34187 23811 34193
rect 23753 34184 23765 34187
rect 23624 34156 23765 34184
rect 23624 34144 23630 34156
rect 23753 34153 23765 34156
rect 23799 34153 23811 34187
rect 23753 34147 23811 34153
rect 26786 34144 26792 34196
rect 26844 34184 26850 34196
rect 26881 34187 26939 34193
rect 26881 34184 26893 34187
rect 26844 34156 26893 34184
rect 26844 34144 26850 34156
rect 26881 34153 26893 34156
rect 26927 34184 26939 34187
rect 26927 34156 27476 34184
rect 26927 34153 26939 34156
rect 26881 34147 26939 34153
rect 6914 34076 6920 34128
rect 6972 34116 6978 34128
rect 17880 34116 17908 34144
rect 6972 34088 17908 34116
rect 6972 34076 6978 34088
rect 23014 34076 23020 34128
rect 23072 34116 23078 34128
rect 26513 34119 26571 34125
rect 23072 34088 25452 34116
rect 23072 34076 23078 34088
rect 12434 34008 12440 34060
rect 12492 34048 12498 34060
rect 12986 34048 12992 34060
rect 12492 34020 12992 34048
rect 12492 34008 12498 34020
rect 12986 34008 12992 34020
rect 13044 34008 13050 34060
rect 14182 34008 14188 34060
rect 14240 34048 14246 34060
rect 20717 34051 20775 34057
rect 20717 34048 20729 34051
rect 14240 34020 20729 34048
rect 14240 34008 14246 34020
rect 20717 34017 20729 34020
rect 20763 34048 20775 34051
rect 23290 34048 23296 34060
rect 20763 34020 23296 34048
rect 20763 34017 20775 34020
rect 20717 34011 20775 34017
rect 23290 34008 23296 34020
rect 23348 34008 23354 34060
rect 4062 33940 4068 33992
rect 4120 33980 4126 33992
rect 5169 33983 5227 33989
rect 5169 33980 5181 33983
rect 4120 33952 5181 33980
rect 4120 33940 4126 33952
rect 5169 33949 5181 33952
rect 5215 33949 5227 33983
rect 5169 33943 5227 33949
rect 14090 33940 14096 33992
rect 14148 33940 14154 33992
rect 14277 33983 14335 33989
rect 14277 33949 14289 33983
rect 14323 33949 14335 33983
rect 14277 33943 14335 33949
rect 5445 33915 5503 33921
rect 5445 33881 5457 33915
rect 5491 33912 5503 33915
rect 5718 33912 5724 33924
rect 5491 33884 5724 33912
rect 5491 33881 5503 33884
rect 5445 33875 5503 33881
rect 5718 33872 5724 33884
rect 5776 33872 5782 33924
rect 5828 33884 5934 33912
rect 5350 33804 5356 33856
rect 5408 33844 5414 33856
rect 5828 33844 5856 33884
rect 12894 33872 12900 33924
rect 12952 33912 12958 33924
rect 14292 33912 14320 33943
rect 14366 33940 14372 33992
rect 14424 33940 14430 33992
rect 14461 33983 14519 33989
rect 14461 33949 14473 33983
rect 14507 33949 14519 33983
rect 14461 33943 14519 33949
rect 12952 33884 14320 33912
rect 14476 33912 14504 33943
rect 15378 33940 15384 33992
rect 15436 33940 15442 33992
rect 15470 33940 15476 33992
rect 15528 33980 15534 33992
rect 15565 33983 15623 33989
rect 15565 33980 15577 33983
rect 15528 33952 15577 33980
rect 15528 33940 15534 33952
rect 15565 33949 15577 33952
rect 15611 33949 15623 33983
rect 17773 33983 17831 33989
rect 17773 33980 17785 33983
rect 15565 33943 15623 33949
rect 17420 33952 17785 33980
rect 15102 33912 15108 33924
rect 14476 33884 15108 33912
rect 12952 33872 12958 33884
rect 15102 33872 15108 33884
rect 15160 33912 15166 33924
rect 15654 33912 15660 33924
rect 15160 33884 15660 33912
rect 15160 33872 15166 33884
rect 15654 33872 15660 33884
rect 15712 33872 15718 33924
rect 15749 33915 15807 33921
rect 15749 33881 15761 33915
rect 15795 33912 15807 33915
rect 15930 33912 15936 33924
rect 15795 33884 15936 33912
rect 15795 33881 15807 33884
rect 15749 33875 15807 33881
rect 15930 33872 15936 33884
rect 15988 33872 15994 33924
rect 17420 33856 17448 33952
rect 17773 33949 17785 33952
rect 17819 33949 17831 33983
rect 17773 33943 17831 33949
rect 17957 33983 18015 33989
rect 17957 33949 17969 33983
rect 18003 33980 18015 33983
rect 18138 33980 18144 33992
rect 18003 33952 18144 33980
rect 18003 33949 18015 33952
rect 17957 33943 18015 33949
rect 18138 33940 18144 33952
rect 18196 33940 18202 33992
rect 22462 33940 22468 33992
rect 22520 33980 22526 33992
rect 23109 33983 23167 33989
rect 23109 33980 23121 33983
rect 22520 33952 23121 33980
rect 22520 33940 22526 33952
rect 23109 33949 23121 33952
rect 23155 33949 23167 33983
rect 23109 33943 23167 33949
rect 23937 33983 23995 33989
rect 23937 33949 23949 33983
rect 23983 33980 23995 33983
rect 24394 33980 24400 33992
rect 23983 33952 24400 33980
rect 23983 33949 23995 33952
rect 23937 33943 23995 33949
rect 24394 33940 24400 33952
rect 24452 33940 24458 33992
rect 25130 33940 25136 33992
rect 25188 33980 25194 33992
rect 25424 33989 25452 34088
rect 26513 34085 26525 34119
rect 26559 34116 26571 34119
rect 27338 34116 27344 34128
rect 26559 34088 27344 34116
rect 26559 34085 26571 34088
rect 26513 34079 26571 34085
rect 27338 34076 27344 34088
rect 27396 34076 27402 34128
rect 27448 34116 27476 34156
rect 27522 34144 27528 34196
rect 27580 34144 27586 34196
rect 27448 34088 30604 34116
rect 26329 34051 26387 34057
rect 26329 34017 26341 34051
rect 26375 34048 26387 34051
rect 26418 34048 26424 34060
rect 26375 34020 26424 34048
rect 26375 34017 26387 34020
rect 26329 34011 26387 34017
rect 26418 34008 26424 34020
rect 26476 34048 26482 34060
rect 26476 34020 26740 34048
rect 26476 34008 26482 34020
rect 25225 33983 25283 33989
rect 25225 33980 25237 33983
rect 25188 33952 25237 33980
rect 25188 33940 25194 33952
rect 25225 33949 25237 33952
rect 25271 33949 25283 33983
rect 25225 33943 25283 33949
rect 25409 33983 25467 33989
rect 25409 33949 25421 33983
rect 25455 33949 25467 33983
rect 25409 33943 25467 33949
rect 26602 33940 26608 33992
rect 26660 33940 26666 33992
rect 26712 33980 26740 34020
rect 30098 34008 30104 34060
rect 30156 34048 30162 34060
rect 30576 34057 30604 34088
rect 30193 34051 30251 34057
rect 30193 34048 30205 34051
rect 30156 34020 30205 34048
rect 30156 34008 30162 34020
rect 30193 34017 30205 34020
rect 30239 34017 30251 34051
rect 30193 34011 30251 34017
rect 30561 34051 30619 34057
rect 30561 34017 30573 34051
rect 30607 34048 30619 34051
rect 31386 34048 31392 34060
rect 30607 34020 31392 34048
rect 30607 34017 30619 34020
rect 30561 34011 30619 34017
rect 27341 33983 27399 33989
rect 26712 33976 27200 33980
rect 27341 33976 27353 33983
rect 26712 33952 27353 33976
rect 27172 33949 27353 33952
rect 27387 33949 27399 33983
rect 27172 33948 27399 33949
rect 27341 33943 27399 33948
rect 27522 33940 27528 33992
rect 27580 33980 27586 33992
rect 29730 33980 29736 33992
rect 27580 33952 29736 33980
rect 27580 33940 27586 33952
rect 29730 33940 29736 33952
rect 29788 33980 29794 33992
rect 29825 33983 29883 33989
rect 29825 33980 29837 33983
rect 29788 33952 29837 33980
rect 29788 33940 29794 33952
rect 29825 33949 29837 33952
rect 29871 33949 29883 33983
rect 29825 33943 29883 33949
rect 30009 33983 30067 33989
rect 30009 33949 30021 33983
rect 30055 33949 30067 33983
rect 30208 33980 30236 34011
rect 31386 34008 31392 34020
rect 31444 34008 31450 34060
rect 30285 33983 30343 33989
rect 30285 33980 30297 33983
rect 30208 33952 30297 33980
rect 30009 33943 30067 33949
rect 30285 33949 30297 33952
rect 30331 33949 30343 33983
rect 30285 33943 30343 33949
rect 30377 33983 30435 33989
rect 30377 33949 30389 33983
rect 30423 33980 30435 33983
rect 31754 33980 31760 33992
rect 30423 33952 31760 33980
rect 30423 33949 30435 33952
rect 30377 33943 30435 33949
rect 20990 33872 20996 33924
rect 21048 33872 21054 33924
rect 21450 33872 21456 33924
rect 21508 33872 21514 33924
rect 22925 33915 22983 33921
rect 22925 33881 22937 33915
rect 22971 33912 22983 33915
rect 23014 33912 23020 33924
rect 22971 33884 23020 33912
rect 22971 33881 22983 33884
rect 22925 33875 22983 33881
rect 23014 33872 23020 33884
rect 23072 33872 23078 33924
rect 26697 33915 26755 33921
rect 23124 33884 24164 33912
rect 5408 33816 5856 33844
rect 5408 33804 5414 33816
rect 17402 33804 17408 33856
rect 17460 33804 17466 33856
rect 17770 33804 17776 33856
rect 17828 33804 17834 33856
rect 17862 33804 17868 33856
rect 17920 33844 17926 33856
rect 23124 33844 23152 33884
rect 24136 33856 24164 33884
rect 26697 33881 26709 33915
rect 26743 33912 26755 33915
rect 29086 33912 29092 33924
rect 26743 33884 27200 33912
rect 26743 33881 26755 33884
rect 26697 33875 26755 33881
rect 17920 33816 23152 33844
rect 17920 33804 17926 33816
rect 23290 33804 23296 33856
rect 23348 33804 23354 33856
rect 24118 33804 24124 33856
rect 24176 33804 24182 33856
rect 25038 33804 25044 33856
rect 25096 33804 25102 33856
rect 26326 33804 26332 33856
rect 26384 33844 26390 33856
rect 26897 33847 26955 33853
rect 26897 33844 26909 33847
rect 26384 33816 26909 33844
rect 26384 33804 26390 33816
rect 26897 33813 26909 33816
rect 26943 33813 26955 33847
rect 26897 33807 26955 33813
rect 27062 33804 27068 33856
rect 27120 33804 27126 33856
rect 27172 33853 27200 33884
rect 27264 33884 29092 33912
rect 27264 33856 27292 33884
rect 29086 33872 29092 33884
rect 29144 33872 29150 33924
rect 30024 33912 30052 33943
rect 30392 33912 30420 33943
rect 31754 33940 31760 33952
rect 31812 33940 31818 33992
rect 30024 33884 30420 33912
rect 27157 33847 27215 33853
rect 27157 33813 27169 33847
rect 27203 33813 27215 33847
rect 27157 33807 27215 33813
rect 27246 33804 27252 33856
rect 27304 33804 27310 33856
rect 27890 33804 27896 33856
rect 27948 33844 27954 33856
rect 30466 33844 30472 33856
rect 27948 33816 30472 33844
rect 27948 33804 27954 33816
rect 30466 33804 30472 33816
rect 30524 33804 30530 33856
rect 30558 33804 30564 33856
rect 30616 33804 30622 33856
rect 1104 33754 38272 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 38272 33754
rect 1104 33680 38272 33702
rect 5718 33600 5724 33652
rect 5776 33640 5782 33652
rect 5905 33643 5963 33649
rect 5905 33640 5917 33643
rect 5776 33612 5917 33640
rect 5776 33600 5782 33612
rect 5905 33609 5917 33612
rect 5951 33609 5963 33643
rect 5905 33603 5963 33609
rect 6917 33643 6975 33649
rect 6917 33609 6929 33643
rect 6963 33609 6975 33643
rect 6917 33603 6975 33609
rect 4341 33575 4399 33581
rect 4341 33541 4353 33575
rect 4387 33572 4399 33575
rect 4614 33572 4620 33584
rect 4387 33544 4620 33572
rect 4387 33541 4399 33544
rect 4341 33535 4399 33541
rect 4614 33532 4620 33544
rect 4672 33532 4678 33584
rect 5350 33532 5356 33584
rect 5408 33532 5414 33584
rect 6932 33572 6960 33603
rect 8294 33600 8300 33652
rect 8352 33640 8358 33652
rect 8757 33643 8815 33649
rect 8757 33640 8769 33643
rect 8352 33612 8769 33640
rect 8352 33600 8358 33612
rect 8757 33609 8769 33612
rect 8803 33640 8815 33643
rect 11790 33640 11796 33652
rect 8803 33612 11796 33640
rect 8803 33609 8815 33612
rect 8757 33603 8815 33609
rect 11790 33600 11796 33612
rect 11848 33600 11854 33652
rect 12250 33640 12256 33652
rect 11900 33612 12256 33640
rect 7285 33575 7343 33581
rect 7285 33572 7297 33575
rect 6932 33544 7297 33572
rect 7285 33541 7297 33544
rect 7331 33541 7343 33575
rect 7285 33535 7343 33541
rect 9493 33575 9551 33581
rect 9493 33541 9505 33575
rect 9539 33572 9551 33575
rect 9766 33572 9772 33584
rect 9539 33544 9772 33572
rect 9539 33541 9551 33544
rect 9493 33535 9551 33541
rect 9766 33532 9772 33544
rect 9824 33532 9830 33584
rect 9950 33532 9956 33584
rect 10008 33532 10014 33584
rect 11900 33516 11928 33612
rect 12250 33600 12256 33612
rect 12308 33600 12314 33652
rect 12894 33600 12900 33652
rect 12952 33600 12958 33652
rect 14182 33600 14188 33652
rect 14240 33640 14246 33652
rect 14277 33643 14335 33649
rect 14277 33640 14289 33643
rect 14240 33612 14289 33640
rect 14240 33600 14246 33612
rect 14277 33609 14289 33612
rect 14323 33609 14335 33643
rect 14277 33603 14335 33609
rect 15013 33643 15071 33649
rect 15013 33609 15025 33643
rect 15059 33640 15071 33643
rect 15378 33640 15384 33652
rect 15059 33612 15384 33640
rect 15059 33609 15071 33612
rect 15013 33603 15071 33609
rect 11974 33532 11980 33584
rect 12032 33581 12038 33584
rect 12032 33575 12061 33581
rect 12049 33541 12061 33575
rect 12032 33535 12061 33541
rect 12529 33575 12587 33581
rect 12529 33541 12541 33575
rect 12575 33572 12587 33575
rect 13538 33572 13544 33584
rect 12575 33544 13544 33572
rect 12575 33541 12587 33544
rect 12529 33535 12587 33541
rect 12032 33532 12038 33535
rect 13188 33516 13216 33544
rect 13538 33532 13544 33544
rect 13596 33532 13602 33584
rect 6086 33464 6092 33516
rect 6144 33464 6150 33516
rect 6730 33464 6736 33516
rect 6788 33464 6794 33516
rect 8938 33504 8944 33516
rect 8418 33476 8944 33504
rect 8938 33464 8944 33476
rect 8996 33504 9002 33516
rect 8996 33476 9168 33504
rect 8996 33464 9002 33476
rect 4062 33396 4068 33448
rect 4120 33396 4126 33448
rect 7006 33396 7012 33448
rect 7064 33396 7070 33448
rect 9140 33368 9168 33476
rect 11698 33464 11704 33516
rect 11756 33464 11762 33516
rect 11790 33464 11796 33516
rect 11848 33464 11854 33516
rect 11882 33464 11888 33516
rect 11940 33464 11946 33516
rect 12710 33464 12716 33516
rect 12768 33464 12774 33516
rect 12989 33507 13047 33513
rect 12989 33473 13001 33507
rect 13035 33473 13047 33507
rect 12989 33467 13047 33473
rect 9214 33396 9220 33448
rect 9272 33396 9278 33448
rect 9950 33436 9956 33448
rect 9324 33408 9956 33436
rect 9324 33368 9352 33408
rect 9950 33396 9956 33408
rect 10008 33396 10014 33448
rect 11606 33396 11612 33448
rect 11664 33436 11670 33448
rect 12161 33439 12219 33445
rect 12161 33436 12173 33439
rect 11664 33408 12173 33436
rect 11664 33396 11670 33408
rect 12161 33405 12173 33408
rect 12207 33405 12219 33439
rect 12161 33399 12219 33405
rect 12434 33396 12440 33448
rect 12492 33436 12498 33448
rect 13004 33436 13032 33467
rect 13170 33464 13176 33516
rect 13228 33464 13234 33516
rect 14826 33464 14832 33516
rect 14884 33464 14890 33516
rect 15010 33464 15016 33516
rect 15068 33464 15074 33516
rect 15120 33513 15148 33612
rect 15378 33600 15384 33612
rect 15436 33600 15442 33652
rect 15654 33600 15660 33652
rect 15712 33600 15718 33652
rect 17126 33600 17132 33652
rect 17184 33640 17190 33652
rect 21634 33640 21640 33652
rect 17184 33612 21640 33640
rect 17184 33600 17190 33612
rect 21634 33600 21640 33612
rect 21692 33600 21698 33652
rect 24670 33600 24676 33652
rect 24728 33600 24734 33652
rect 26329 33643 26387 33649
rect 26329 33609 26341 33643
rect 26375 33640 26387 33643
rect 26418 33640 26424 33652
rect 26375 33612 26424 33640
rect 26375 33609 26387 33612
rect 26329 33603 26387 33609
rect 26418 33600 26424 33612
rect 26476 33600 26482 33652
rect 27062 33600 27068 33652
rect 27120 33600 27126 33652
rect 28261 33643 28319 33649
rect 28261 33609 28273 33643
rect 28307 33609 28319 33643
rect 28261 33603 28319 33609
rect 28467 33612 28948 33640
rect 15473 33575 15531 33581
rect 15473 33541 15485 33575
rect 15519 33572 15531 33575
rect 24688 33572 24716 33600
rect 15519 33544 16160 33572
rect 15519 33541 15531 33544
rect 15473 33535 15531 33541
rect 15105 33507 15163 33513
rect 15105 33473 15117 33507
rect 15151 33473 15163 33507
rect 15105 33467 15163 33473
rect 15289 33507 15347 33513
rect 15289 33473 15301 33507
rect 15335 33473 15347 33507
rect 15289 33467 15347 33473
rect 15381 33507 15439 33513
rect 15381 33473 15393 33507
rect 15427 33473 15439 33507
rect 15381 33467 15439 33473
rect 15565 33507 15623 33513
rect 15565 33473 15577 33507
rect 15611 33504 15623 33507
rect 15930 33504 15936 33516
rect 15611 33476 15936 33504
rect 15611 33473 15623 33476
rect 15565 33467 15623 33473
rect 12492 33408 13032 33436
rect 12492 33396 12498 33408
rect 15304 33368 15332 33467
rect 15396 33436 15424 33467
rect 15930 33464 15936 33476
rect 15988 33464 15994 33516
rect 16022 33464 16028 33516
rect 16080 33464 16086 33516
rect 16132 33513 16160 33544
rect 18340 33544 18828 33572
rect 18340 33516 18368 33544
rect 16117 33507 16175 33513
rect 16117 33473 16129 33507
rect 16163 33473 16175 33507
rect 16117 33467 16175 33473
rect 16301 33507 16359 33513
rect 16301 33473 16313 33507
rect 16347 33504 16359 33507
rect 17678 33504 17684 33516
rect 16347 33476 17684 33504
rect 16347 33473 16359 33476
rect 16301 33467 16359 33473
rect 17678 33464 17684 33476
rect 17736 33464 17742 33516
rect 18141 33507 18199 33513
rect 18141 33473 18153 33507
rect 18187 33504 18199 33507
rect 18322 33504 18328 33516
rect 18187 33476 18328 33504
rect 18187 33473 18199 33476
rect 18141 33467 18199 33473
rect 18322 33464 18328 33476
rect 18380 33464 18386 33516
rect 18800 33513 18828 33544
rect 19812 33544 20116 33572
rect 24688 33544 27016 33572
rect 18509 33507 18567 33513
rect 18509 33473 18521 33507
rect 18555 33473 18567 33507
rect 18509 33467 18567 33473
rect 18693 33507 18751 33513
rect 18693 33473 18705 33507
rect 18739 33473 18751 33507
rect 18693 33467 18751 33473
rect 18785 33507 18843 33513
rect 18785 33473 18797 33507
rect 18831 33473 18843 33507
rect 18785 33467 18843 33473
rect 16040 33436 16068 33464
rect 15396 33408 16068 33436
rect 17402 33396 17408 33448
rect 17460 33396 17466 33448
rect 18046 33396 18052 33448
rect 18104 33436 18110 33448
rect 18524 33436 18552 33467
rect 18104 33408 18552 33436
rect 18708 33436 18736 33467
rect 19334 33464 19340 33516
rect 19392 33464 19398 33516
rect 19610 33464 19616 33516
rect 19668 33504 19674 33516
rect 19812 33513 19840 33544
rect 20088 33516 20116 33544
rect 19797 33507 19855 33513
rect 19797 33504 19809 33507
rect 19668 33476 19809 33504
rect 19668 33464 19674 33476
rect 19797 33473 19809 33476
rect 19843 33473 19855 33507
rect 19797 33467 19855 33473
rect 19981 33507 20039 33513
rect 19981 33473 19993 33507
rect 20027 33473 20039 33507
rect 19981 33467 20039 33473
rect 18877 33439 18935 33445
rect 18877 33436 18889 33439
rect 18708 33408 18889 33436
rect 18104 33396 18110 33408
rect 18877 33405 18889 33408
rect 18923 33405 18935 33439
rect 19352 33436 19380 33464
rect 19996 33436 20024 33467
rect 20070 33464 20076 33516
rect 20128 33464 20134 33516
rect 25866 33464 25872 33516
rect 25924 33464 25930 33516
rect 26053 33507 26111 33513
rect 26053 33473 26065 33507
rect 26099 33473 26111 33507
rect 26053 33467 26111 33473
rect 26145 33507 26203 33513
rect 26145 33473 26157 33507
rect 26191 33504 26203 33507
rect 26326 33504 26332 33516
rect 26191 33476 26332 33504
rect 26191 33473 26203 33476
rect 26145 33467 26203 33473
rect 19352 33408 20024 33436
rect 26068 33436 26096 33467
rect 26326 33464 26332 33476
rect 26384 33464 26390 33516
rect 26510 33464 26516 33516
rect 26568 33464 26574 33516
rect 26988 33513 27016 33544
rect 26973 33507 27031 33513
rect 26973 33473 26985 33507
rect 27019 33473 27031 33507
rect 27080 33504 27108 33600
rect 27709 33575 27767 33581
rect 27709 33572 27721 33575
rect 27356 33544 27721 33572
rect 27356 33513 27384 33544
rect 27709 33541 27721 33544
rect 27755 33541 27767 33575
rect 28276 33572 28304 33603
rect 28467 33572 28495 33612
rect 28276 33544 28495 33572
rect 28558 33544 28764 33572
rect 27709 33535 27767 33541
rect 27249 33507 27307 33513
rect 27249 33504 27261 33507
rect 27080 33476 27261 33504
rect 26973 33467 27031 33473
rect 27249 33473 27261 33476
rect 27295 33473 27307 33507
rect 27249 33467 27307 33473
rect 27341 33507 27399 33513
rect 27341 33473 27353 33507
rect 27387 33473 27399 33507
rect 27341 33467 27399 33473
rect 27522 33464 27528 33516
rect 27580 33504 27586 33516
rect 27580 33476 28028 33504
rect 27580 33464 27586 33476
rect 26602 33436 26608 33448
rect 26068 33408 26608 33436
rect 18877 33399 18935 33405
rect 26602 33396 26608 33408
rect 26660 33436 26666 33448
rect 26697 33439 26755 33445
rect 26697 33436 26709 33439
rect 26660 33408 26709 33436
rect 26660 33396 26666 33408
rect 26697 33405 26709 33408
rect 26743 33405 26755 33439
rect 26697 33399 26755 33405
rect 27890 33396 27896 33448
rect 27948 33396 27954 33448
rect 28000 33436 28028 33476
rect 28166 33464 28172 33516
rect 28224 33504 28230 33516
rect 28445 33507 28503 33513
rect 28445 33504 28457 33507
rect 28224 33476 28457 33504
rect 28224 33464 28230 33476
rect 28445 33473 28457 33476
rect 28491 33504 28503 33507
rect 28558 33504 28586 33544
rect 28736 33513 28764 33544
rect 28920 33513 28948 33612
rect 29086 33600 29092 33652
rect 29144 33600 29150 33652
rect 29730 33600 29736 33652
rect 29788 33600 29794 33652
rect 30558 33600 30564 33652
rect 30616 33600 30622 33652
rect 31754 33600 31760 33652
rect 31812 33600 31818 33652
rect 28491 33476 28586 33504
rect 28629 33507 28687 33513
rect 28491 33473 28503 33476
rect 28445 33467 28503 33473
rect 28629 33473 28641 33507
rect 28675 33473 28687 33507
rect 28629 33467 28687 33473
rect 28721 33507 28779 33513
rect 28721 33473 28733 33507
rect 28767 33473 28779 33507
rect 28905 33507 28963 33513
rect 28905 33504 28917 33507
rect 28863 33476 28917 33504
rect 28721 33467 28779 33473
rect 28905 33473 28917 33476
rect 28951 33504 28963 33507
rect 29178 33504 29184 33516
rect 28951 33476 29184 33504
rect 28951 33473 28963 33476
rect 28905 33467 28963 33473
rect 28537 33439 28595 33445
rect 28537 33436 28549 33439
rect 28000 33408 28549 33436
rect 28537 33405 28549 33408
rect 28583 33405 28595 33439
rect 28644 33436 28672 33467
rect 29178 33464 29184 33476
rect 29236 33464 29242 33516
rect 29270 33464 29276 33516
rect 29328 33464 29334 33516
rect 29748 33504 29776 33600
rect 29825 33507 29883 33513
rect 29825 33504 29837 33507
rect 29748 33476 29837 33504
rect 29825 33473 29837 33476
rect 29871 33473 29883 33507
rect 29825 33467 29883 33473
rect 29917 33507 29975 33513
rect 29917 33473 29929 33507
rect 29963 33504 29975 33507
rect 30576 33504 30604 33600
rect 29963 33476 30604 33504
rect 31113 33507 31171 33513
rect 29963 33473 29975 33476
rect 29917 33467 29975 33473
rect 31113 33473 31125 33507
rect 31159 33473 31171 33507
rect 31113 33467 31171 33473
rect 31389 33507 31447 33513
rect 31389 33473 31401 33507
rect 31435 33473 31447 33507
rect 31389 33467 31447 33473
rect 30193 33439 30251 33445
rect 30193 33436 30205 33439
rect 28644 33408 30205 33436
rect 28537 33399 28595 33405
rect 30193 33405 30205 33408
rect 30239 33405 30251 33439
rect 30193 33399 30251 33405
rect 9140 33340 9352 33368
rect 10888 33340 12388 33368
rect 15304 33340 15424 33368
rect 5810 33260 5816 33312
rect 5868 33300 5874 33312
rect 10888 33300 10916 33340
rect 12360 33312 12388 33340
rect 15396 33312 15424 33340
rect 20806 33328 20812 33380
rect 20864 33368 20870 33380
rect 27246 33368 27252 33380
rect 20864 33340 25912 33368
rect 20864 33328 20870 33340
rect 5868 33272 10916 33300
rect 5868 33260 5874 33272
rect 10962 33260 10968 33312
rect 11020 33260 11026 33312
rect 11514 33260 11520 33312
rect 11572 33260 11578 33312
rect 12342 33260 12348 33312
rect 12400 33260 12406 33312
rect 15194 33260 15200 33312
rect 15252 33260 15258 33312
rect 15378 33260 15384 33312
rect 15436 33260 15442 33312
rect 18506 33260 18512 33312
rect 18564 33260 18570 33312
rect 19794 33260 19800 33312
rect 19852 33260 19858 33312
rect 25682 33260 25688 33312
rect 25740 33260 25746 33312
rect 25884 33300 25912 33340
rect 26528 33340 27252 33368
rect 26528 33300 26556 33340
rect 27246 33328 27252 33340
rect 27304 33328 27310 33380
rect 27430 33328 27436 33380
rect 27488 33328 27494 33380
rect 28074 33328 28080 33380
rect 28132 33368 28138 33380
rect 28905 33371 28963 33377
rect 28905 33368 28917 33371
rect 28132 33340 28917 33368
rect 28132 33328 28138 33340
rect 28905 33337 28917 33340
rect 28951 33337 28963 33371
rect 30098 33368 30104 33380
rect 28905 33331 28963 33337
rect 29564 33340 30104 33368
rect 25884 33272 26556 33300
rect 27985 33303 28043 33309
rect 27985 33269 27997 33303
rect 28031 33300 28043 33303
rect 29564 33300 29592 33340
rect 30098 33328 30104 33340
rect 30156 33328 30162 33380
rect 28031 33272 29592 33300
rect 28031 33269 28043 33272
rect 27985 33263 28043 33269
rect 29638 33260 29644 33312
rect 29696 33260 29702 33312
rect 30208 33300 30236 33399
rect 30282 33396 30288 33448
rect 30340 33396 30346 33448
rect 30466 33396 30472 33448
rect 30524 33436 30530 33448
rect 31128 33436 31156 33467
rect 31202 33436 31208 33448
rect 30524 33408 31208 33436
rect 30524 33396 30530 33408
rect 31202 33396 31208 33408
rect 31260 33396 31266 33448
rect 31404 33436 31432 33467
rect 31478 33464 31484 33516
rect 31536 33464 31542 33516
rect 31632 33507 31690 33513
rect 31632 33473 31644 33507
rect 31678 33504 31690 33507
rect 31678 33476 31754 33504
rect 31678 33473 31690 33476
rect 31632 33467 31690 33473
rect 31726 33436 31754 33476
rect 31846 33464 31852 33516
rect 31904 33504 31910 33516
rect 32306 33504 32312 33516
rect 31904 33476 32312 33504
rect 31904 33464 31910 33476
rect 32306 33464 32312 33476
rect 32364 33504 32370 33516
rect 32585 33507 32643 33513
rect 32585 33504 32597 33507
rect 32364 33476 32597 33504
rect 32364 33464 32370 33476
rect 32585 33473 32597 33476
rect 32631 33473 32643 33507
rect 32585 33467 32643 33473
rect 32030 33436 32036 33448
rect 31404 33408 31524 33436
rect 31726 33408 32036 33436
rect 31496 33380 31524 33408
rect 32030 33396 32036 33408
rect 32088 33436 32094 33448
rect 32493 33439 32551 33445
rect 32493 33436 32505 33439
rect 32088 33408 32505 33436
rect 32088 33396 32094 33408
rect 32493 33405 32505 33408
rect 32539 33405 32551 33439
rect 32493 33399 32551 33405
rect 31113 33371 31171 33377
rect 31113 33337 31125 33371
rect 31159 33368 31171 33371
rect 31386 33368 31392 33380
rect 31159 33340 31392 33368
rect 31159 33337 31171 33340
rect 31113 33331 31171 33337
rect 31386 33328 31392 33340
rect 31444 33328 31450 33380
rect 31478 33328 31484 33380
rect 31536 33328 31542 33380
rect 31941 33371 31999 33377
rect 31941 33337 31953 33371
rect 31987 33368 31999 33371
rect 33134 33368 33140 33380
rect 31987 33340 33140 33368
rect 31987 33337 31999 33340
rect 31941 33331 31999 33337
rect 33134 33328 33140 33340
rect 33192 33368 33198 33380
rect 34146 33368 34152 33380
rect 33192 33340 34152 33368
rect 33192 33328 33198 33340
rect 34146 33328 34152 33340
rect 34204 33328 34210 33380
rect 31754 33300 31760 33312
rect 30208 33272 31760 33300
rect 31754 33260 31760 33272
rect 31812 33260 31818 33312
rect 32861 33303 32919 33309
rect 32861 33269 32873 33303
rect 32907 33300 32919 33303
rect 34054 33300 34060 33312
rect 32907 33272 34060 33300
rect 32907 33269 32919 33272
rect 32861 33263 32919 33269
rect 34054 33260 34060 33272
rect 34112 33260 34118 33312
rect 1104 33210 38272 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38272 33210
rect 1104 33136 38272 33158
rect 4433 33099 4491 33105
rect 4433 33065 4445 33099
rect 4479 33096 4491 33099
rect 4614 33096 4620 33108
rect 4479 33068 4620 33096
rect 4479 33065 4491 33068
rect 4433 33059 4491 33065
rect 4614 33056 4620 33068
rect 4672 33056 4678 33108
rect 5813 33099 5871 33105
rect 5813 33065 5825 33099
rect 5859 33096 5871 33099
rect 6086 33096 6092 33108
rect 5859 33068 6092 33096
rect 5859 33065 5871 33068
rect 5813 33059 5871 33065
rect 6086 33056 6092 33068
rect 6144 33056 6150 33108
rect 6730 33056 6736 33108
rect 6788 33096 6794 33108
rect 6825 33099 6883 33105
rect 6825 33096 6837 33099
rect 6788 33068 6837 33096
rect 6788 33056 6794 33068
rect 6825 33065 6837 33068
rect 6871 33065 6883 33099
rect 6825 33059 6883 33065
rect 9766 33056 9772 33108
rect 9824 33056 9830 33108
rect 11698 33056 11704 33108
rect 11756 33056 11762 33108
rect 11790 33056 11796 33108
rect 11848 33056 11854 33108
rect 14369 33099 14427 33105
rect 14369 33065 14381 33099
rect 14415 33096 14427 33099
rect 14415 33068 15056 33096
rect 14415 33065 14427 33068
rect 14369 33059 14427 33065
rect 8389 33031 8447 33037
rect 8389 32997 8401 33031
rect 8435 32997 8447 33031
rect 11716 33028 11744 33056
rect 15028 33040 15056 33068
rect 16022 33056 16028 33108
rect 16080 33056 16086 33108
rect 17494 33096 17500 33108
rect 16132 33068 17500 33096
rect 12253 33031 12311 33037
rect 12253 33028 12265 33031
rect 11716 33000 12265 33028
rect 8389 32991 8447 32997
rect 12253 32997 12265 33000
rect 12299 32997 12311 33031
rect 12253 32991 12311 32997
rect 13725 33031 13783 33037
rect 13725 32997 13737 33031
rect 13771 33028 13783 33031
rect 13771 33000 14136 33028
rect 13771 32997 13783 33000
rect 13725 32991 13783 32997
rect 5261 32963 5319 32969
rect 5261 32929 5273 32963
rect 5307 32960 5319 32963
rect 6457 32963 6515 32969
rect 6457 32960 6469 32963
rect 5307 32932 6469 32960
rect 5307 32929 5319 32932
rect 5261 32923 5319 32929
rect 6457 32929 6469 32932
rect 6503 32960 6515 32963
rect 7466 32960 7472 32972
rect 6503 32932 7472 32960
rect 6503 32929 6515 32932
rect 6457 32923 6515 32929
rect 7466 32920 7472 32932
rect 7524 32960 7530 32972
rect 7745 32963 7803 32969
rect 7745 32960 7757 32963
rect 7524 32932 7757 32960
rect 7524 32920 7530 32932
rect 7745 32929 7757 32932
rect 7791 32929 7803 32963
rect 7745 32923 7803 32929
rect 4617 32895 4675 32901
rect 4617 32861 4629 32895
rect 4663 32892 4675 32895
rect 5077 32895 5135 32901
rect 4663 32864 4752 32892
rect 4663 32861 4675 32864
rect 4617 32855 4675 32861
rect 4724 32765 4752 32864
rect 5077 32861 5089 32895
rect 5123 32892 5135 32895
rect 5350 32892 5356 32904
rect 5123 32864 5356 32892
rect 5123 32861 5135 32864
rect 5077 32855 5135 32861
rect 5350 32852 5356 32864
rect 5408 32852 5414 32904
rect 5810 32852 5816 32904
rect 5868 32852 5874 32904
rect 6273 32895 6331 32901
rect 6273 32861 6285 32895
rect 6319 32892 6331 32895
rect 6914 32892 6920 32904
rect 6319 32864 6920 32892
rect 6319 32861 6331 32864
rect 6273 32855 6331 32861
rect 6914 32852 6920 32864
rect 6972 32852 6978 32904
rect 7098 32852 7104 32904
rect 7156 32892 7162 32904
rect 8021 32895 8079 32901
rect 8021 32892 8033 32895
rect 7156 32864 8033 32892
rect 7156 32852 7162 32864
rect 8021 32861 8033 32864
rect 8067 32861 8079 32895
rect 8294 32892 8300 32904
rect 8021 32855 8079 32861
rect 8128 32864 8300 32892
rect 5169 32827 5227 32833
rect 5169 32793 5181 32827
rect 5215 32824 5227 32827
rect 5828 32824 5856 32852
rect 5215 32796 5856 32824
rect 5215 32793 5227 32796
rect 5169 32787 5227 32793
rect 7926 32784 7932 32836
rect 7984 32784 7990 32836
rect 4709 32759 4767 32765
rect 4709 32725 4721 32759
rect 4755 32725 4767 32759
rect 4709 32719 4767 32725
rect 5718 32716 5724 32768
rect 5776 32756 5782 32768
rect 6181 32759 6239 32765
rect 6181 32756 6193 32759
rect 5776 32728 6193 32756
rect 5776 32716 5782 32728
rect 6181 32725 6193 32728
rect 6227 32725 6239 32759
rect 6181 32719 6239 32725
rect 6730 32716 6736 32768
rect 6788 32756 6794 32768
rect 7193 32759 7251 32765
rect 7193 32756 7205 32759
rect 6788 32728 7205 32756
rect 6788 32716 6794 32728
rect 7193 32725 7205 32728
rect 7239 32725 7251 32759
rect 7193 32719 7251 32725
rect 7285 32759 7343 32765
rect 7285 32725 7297 32759
rect 7331 32756 7343 32759
rect 8128 32756 8156 32864
rect 8294 32852 8300 32864
rect 8352 32852 8358 32904
rect 8404 32892 8432 32991
rect 10686 32920 10692 32972
rect 10744 32960 10750 32972
rect 10965 32963 11023 32969
rect 10965 32960 10977 32963
rect 10744 32932 10977 32960
rect 10744 32920 10750 32932
rect 10965 32929 10977 32932
rect 11011 32929 11023 32963
rect 10965 32923 11023 32929
rect 11514 32920 11520 32972
rect 11572 32920 11578 32972
rect 11606 32920 11612 32972
rect 11664 32960 11670 32972
rect 14108 32960 14136 33000
rect 14826 32988 14832 33040
rect 14884 32988 14890 33040
rect 15010 32988 15016 33040
rect 15068 33028 15074 33040
rect 16132 33028 16160 33068
rect 17494 33056 17500 33068
rect 17552 33056 17558 33108
rect 18138 33056 18144 33108
rect 18196 33096 18202 33108
rect 18325 33099 18383 33105
rect 18325 33096 18337 33099
rect 18196 33068 18337 33096
rect 18196 33056 18202 33068
rect 18325 33065 18337 33068
rect 18371 33065 18383 33099
rect 18325 33059 18383 33065
rect 19058 33056 19064 33108
rect 19116 33096 19122 33108
rect 19702 33096 19708 33108
rect 19116 33068 19708 33096
rect 19116 33056 19122 33068
rect 19702 33056 19708 33068
rect 19760 33056 19766 33108
rect 19978 33056 19984 33108
rect 20036 33056 20042 33108
rect 20070 33056 20076 33108
rect 20128 33056 20134 33108
rect 21726 33056 21732 33108
rect 21784 33096 21790 33108
rect 23842 33096 23848 33108
rect 21784 33068 23848 33096
rect 21784 33056 21790 33068
rect 23842 33056 23848 33068
rect 23900 33056 23906 33108
rect 26510 33056 26516 33108
rect 26568 33056 26574 33108
rect 26602 33056 26608 33108
rect 26660 33096 26666 33108
rect 26697 33099 26755 33105
rect 26697 33096 26709 33099
rect 26660 33068 26709 33096
rect 26660 33056 26666 33068
rect 26697 33065 26709 33068
rect 26743 33065 26755 33099
rect 26697 33059 26755 33065
rect 29178 33056 29184 33108
rect 29236 33056 29242 33108
rect 29270 33056 29276 33108
rect 29328 33096 29334 33108
rect 29549 33099 29607 33105
rect 29549 33096 29561 33099
rect 29328 33068 29561 33096
rect 29328 33056 29334 33068
rect 29549 33065 29561 33068
rect 29595 33065 29607 33099
rect 29549 33059 29607 33065
rect 30006 33056 30012 33108
rect 30064 33056 30070 33108
rect 33042 33096 33048 33108
rect 31404 33068 33048 33096
rect 17221 33031 17279 33037
rect 17221 33028 17233 33031
rect 15068 33000 16160 33028
rect 17052 33000 17233 33028
rect 15068 32988 15074 33000
rect 14844 32960 14872 32988
rect 11664 32932 13492 32960
rect 11664 32920 11670 32932
rect 8665 32895 8723 32901
rect 8665 32892 8677 32895
rect 8404 32864 8677 32892
rect 8665 32861 8677 32864
rect 8711 32861 8723 32895
rect 8665 32855 8723 32861
rect 9953 32895 10011 32901
rect 9953 32861 9965 32895
rect 9999 32892 10011 32895
rect 9999 32864 10456 32892
rect 9999 32861 10011 32864
rect 9953 32855 10011 32861
rect 7331 32728 8156 32756
rect 7331 32725 7343 32728
rect 7285 32719 7343 32725
rect 8202 32716 8208 32768
rect 8260 32756 8266 32768
rect 10428 32765 10456 32864
rect 8481 32759 8539 32765
rect 8481 32756 8493 32759
rect 8260 32728 8493 32756
rect 8260 32716 8266 32728
rect 8481 32725 8493 32728
rect 8527 32725 8539 32759
rect 8481 32719 8539 32725
rect 10413 32759 10471 32765
rect 10413 32725 10425 32759
rect 10459 32725 10471 32759
rect 10704 32756 10732 32920
rect 10781 32895 10839 32901
rect 10781 32861 10793 32895
rect 10827 32861 10839 32895
rect 10781 32855 10839 32861
rect 10873 32895 10931 32901
rect 10873 32861 10885 32895
rect 10919 32892 10931 32895
rect 11532 32892 11560 32920
rect 10919 32864 11560 32892
rect 10919 32861 10931 32864
rect 10873 32855 10931 32861
rect 10796 32824 10824 32855
rect 11698 32852 11704 32904
rect 11756 32852 11762 32904
rect 11885 32895 11943 32901
rect 11885 32861 11897 32895
rect 11931 32892 11943 32895
rect 12437 32895 12495 32901
rect 12437 32892 12449 32895
rect 11931 32864 12449 32892
rect 11931 32861 11943 32864
rect 11885 32855 11943 32861
rect 10796 32796 10916 32824
rect 10778 32756 10784 32768
rect 10704 32728 10784 32756
rect 10413 32719 10471 32725
rect 10778 32716 10784 32728
rect 10836 32716 10842 32768
rect 10888 32756 10916 32796
rect 11992 32768 12020 32864
rect 12437 32861 12449 32864
rect 12483 32892 12495 32895
rect 12710 32892 12716 32904
rect 12483 32864 12716 32892
rect 12483 32861 12495 32864
rect 12437 32855 12495 32861
rect 12710 32852 12716 32864
rect 12768 32852 12774 32904
rect 13464 32901 13492 32932
rect 14108 32932 14964 32960
rect 13173 32895 13231 32901
rect 13173 32861 13185 32895
rect 13219 32861 13231 32895
rect 13173 32855 13231 32861
rect 13449 32895 13507 32901
rect 13449 32861 13461 32895
rect 13495 32861 13507 32895
rect 13449 32855 13507 32861
rect 12250 32784 12256 32836
rect 12308 32824 12314 32836
rect 12618 32824 12624 32836
rect 12308 32796 12624 32824
rect 12308 32784 12314 32796
rect 12618 32784 12624 32796
rect 12676 32784 12682 32836
rect 10962 32756 10968 32768
rect 10888 32728 10968 32756
rect 10962 32716 10968 32728
rect 11020 32756 11026 32768
rect 11974 32756 11980 32768
rect 11020 32728 11980 32756
rect 11020 32716 11026 32728
rect 11974 32716 11980 32728
rect 12032 32716 12038 32768
rect 13188 32756 13216 32855
rect 13538 32852 13544 32904
rect 13596 32852 13602 32904
rect 14108 32901 14136 32932
rect 14936 32901 14964 32932
rect 15120 32901 15148 33000
rect 17052 32972 17080 33000
rect 17221 32997 17233 33000
rect 17267 32997 17279 33031
rect 17221 32991 17279 32997
rect 17512 33000 19012 33028
rect 15212 32932 15792 32960
rect 15212 32904 15240 32932
rect 14093 32895 14151 32901
rect 14093 32861 14105 32895
rect 14139 32861 14151 32895
rect 14093 32855 14151 32861
rect 14829 32895 14887 32901
rect 14829 32861 14841 32895
rect 14875 32861 14887 32895
rect 14829 32855 14887 32861
rect 14921 32895 14979 32901
rect 14921 32861 14933 32895
rect 14967 32861 14979 32895
rect 14921 32855 14979 32861
rect 15105 32895 15163 32901
rect 15105 32861 15117 32895
rect 15151 32861 15163 32895
rect 15105 32855 15163 32861
rect 13262 32784 13268 32836
rect 13320 32824 13326 32836
rect 13357 32827 13415 32833
rect 13357 32824 13369 32827
rect 13320 32796 13369 32824
rect 13320 32784 13326 32796
rect 13357 32793 13369 32796
rect 13403 32793 13415 32827
rect 14737 32827 14795 32833
rect 14737 32824 14749 32827
rect 13357 32787 13415 32793
rect 14476 32796 14749 32824
rect 14476 32768 14504 32796
rect 14737 32793 14749 32796
rect 14783 32793 14795 32827
rect 14844 32824 14872 32855
rect 15194 32852 15200 32904
rect 15252 32852 15258 32904
rect 15470 32852 15476 32904
rect 15528 32852 15534 32904
rect 15764 32901 15792 32932
rect 16298 32920 16304 32972
rect 16356 32960 16362 32972
rect 16577 32963 16635 32969
rect 16577 32960 16589 32963
rect 16356 32932 16589 32960
rect 16356 32920 16362 32932
rect 16577 32929 16589 32932
rect 16623 32929 16635 32963
rect 16577 32923 16635 32929
rect 17034 32920 17040 32972
rect 17092 32920 17098 32972
rect 15749 32895 15807 32901
rect 15749 32861 15761 32895
rect 15795 32861 15807 32895
rect 15749 32855 15807 32861
rect 16393 32895 16451 32901
rect 16393 32861 16405 32895
rect 16439 32892 16451 32895
rect 17052 32892 17080 32920
rect 17512 32901 17540 33000
rect 18138 32960 18144 32972
rect 17880 32932 18144 32960
rect 16439 32864 17080 32892
rect 17497 32895 17555 32901
rect 16439 32861 16451 32864
rect 16393 32855 16451 32861
rect 17497 32861 17509 32895
rect 17543 32861 17555 32895
rect 17497 32855 17555 32861
rect 17589 32895 17647 32901
rect 17589 32861 17601 32895
rect 17635 32892 17647 32895
rect 17678 32892 17684 32904
rect 17635 32864 17684 32892
rect 17635 32861 17647 32864
rect 17589 32855 17647 32861
rect 15013 32827 15071 32833
rect 15013 32824 15025 32827
rect 14844 32796 15025 32824
rect 14737 32787 14795 32793
rect 15013 32793 15025 32796
rect 15059 32793 15071 32827
rect 15013 32787 15071 32793
rect 14366 32756 14372 32768
rect 13188 32728 14372 32756
rect 14366 32716 14372 32728
rect 14424 32716 14430 32768
rect 14458 32716 14464 32768
rect 14516 32716 14522 32768
rect 14550 32716 14556 32768
rect 14608 32716 14614 32768
rect 14752 32756 14780 32787
rect 15488 32756 15516 32852
rect 15565 32827 15623 32833
rect 15565 32793 15577 32827
rect 15611 32824 15623 32827
rect 16408 32824 16436 32855
rect 17678 32852 17684 32864
rect 17736 32852 17742 32904
rect 17770 32852 17776 32904
rect 17828 32852 17834 32904
rect 17880 32901 17908 32932
rect 18138 32920 18144 32932
rect 18196 32920 18202 32972
rect 18230 32920 18236 32972
rect 18288 32920 18294 32972
rect 18877 32963 18935 32969
rect 18877 32960 18889 32963
rect 18616 32932 18889 32960
rect 17865 32895 17923 32901
rect 17865 32861 17877 32895
rect 17911 32861 17923 32895
rect 17865 32855 17923 32861
rect 17954 32852 17960 32904
rect 18012 32892 18018 32904
rect 18506 32892 18512 32904
rect 18012 32864 18057 32892
rect 18156 32864 18512 32892
rect 18012 32852 18018 32864
rect 15611 32796 16436 32824
rect 17221 32827 17279 32833
rect 15611 32793 15623 32796
rect 15565 32787 15623 32793
rect 17221 32793 17233 32827
rect 17267 32824 17279 32827
rect 18156 32824 18184 32864
rect 18506 32852 18512 32864
rect 18564 32852 18570 32904
rect 17267 32796 18184 32824
rect 17267 32793 17279 32796
rect 17221 32787 17279 32793
rect 14752 32728 15516 32756
rect 15930 32716 15936 32768
rect 15988 32716 15994 32768
rect 16022 32716 16028 32768
rect 16080 32756 16086 32768
rect 16298 32756 16304 32768
rect 16080 32728 16304 32756
rect 16080 32716 16086 32728
rect 16298 32716 16304 32728
rect 16356 32716 16362 32768
rect 16482 32716 16488 32768
rect 16540 32716 16546 32768
rect 17402 32716 17408 32768
rect 17460 32756 17466 32768
rect 17862 32756 17868 32768
rect 17460 32728 17868 32756
rect 17460 32716 17466 32728
rect 17862 32716 17868 32728
rect 17920 32716 17926 32768
rect 17954 32716 17960 32768
rect 18012 32756 18018 32768
rect 18616 32756 18644 32932
rect 18877 32929 18889 32932
rect 18923 32929 18935 32963
rect 18877 32923 18935 32929
rect 18782 32852 18788 32904
rect 18840 32852 18846 32904
rect 18693 32827 18751 32833
rect 18693 32793 18705 32827
rect 18739 32824 18751 32827
rect 18984 32824 19012 33000
rect 19426 32988 19432 33040
rect 19484 33028 19490 33040
rect 19996 33028 20024 33056
rect 22738 33028 22744 33040
rect 19484 33000 20024 33028
rect 20640 33000 22744 33028
rect 19484 32988 19490 33000
rect 20640 32969 20668 33000
rect 22738 32988 22744 33000
rect 22796 32988 22802 33040
rect 26786 33028 26792 33040
rect 25516 33000 26792 33028
rect 20625 32963 20683 32969
rect 20625 32960 20637 32963
rect 20180 32932 20637 32960
rect 19334 32852 19340 32904
rect 19392 32852 19398 32904
rect 19610 32852 19616 32904
rect 19668 32852 19674 32904
rect 19705 32895 19763 32901
rect 19705 32861 19717 32895
rect 19751 32861 19763 32895
rect 19705 32855 19763 32861
rect 19242 32824 19248 32836
rect 18739 32796 19248 32824
rect 18739 32793 18751 32796
rect 18693 32787 18751 32793
rect 19242 32784 19248 32796
rect 19300 32784 19306 32836
rect 19352 32824 19380 32852
rect 19720 32824 19748 32855
rect 19794 32852 19800 32904
rect 19852 32892 19858 32904
rect 19889 32895 19947 32901
rect 19889 32892 19901 32895
rect 19852 32864 19901 32892
rect 19852 32852 19858 32864
rect 19889 32861 19901 32864
rect 19935 32861 19947 32895
rect 19889 32855 19947 32861
rect 19978 32852 19984 32904
rect 20036 32852 20042 32904
rect 19352 32796 19748 32824
rect 20180 32756 20208 32932
rect 20625 32929 20637 32932
rect 20671 32929 20683 32963
rect 20625 32923 20683 32929
rect 21174 32920 21180 32972
rect 21232 32960 21238 32972
rect 21232 32932 22200 32960
rect 21232 32920 21238 32932
rect 22172 32911 22200 32932
rect 22172 32905 22239 32911
rect 21726 32852 21732 32904
rect 21784 32852 21790 32904
rect 22002 32852 22008 32904
rect 22060 32901 22066 32904
rect 22060 32895 22109 32901
rect 22060 32861 22063 32895
rect 22097 32861 22109 32895
rect 22172 32871 22193 32905
rect 22227 32892 22239 32905
rect 23014 32892 23020 32904
rect 22227 32871 23020 32892
rect 22172 32864 23020 32871
rect 22060 32855 22109 32861
rect 22060 32852 22066 32855
rect 23014 32852 23020 32864
rect 23072 32852 23078 32904
rect 25516 32901 25544 33000
rect 26786 32988 26792 33000
rect 26844 32988 26850 33040
rect 28077 33031 28135 33037
rect 28077 32997 28089 33031
rect 28123 33028 28135 33031
rect 28166 33028 28172 33040
rect 28123 33000 28172 33028
rect 28123 32997 28135 33000
rect 28077 32991 28135 32997
rect 28166 32988 28172 33000
rect 28224 32988 28230 33040
rect 26160 32932 26832 32960
rect 25501 32895 25559 32901
rect 25501 32861 25513 32895
rect 25547 32861 25559 32895
rect 25501 32855 25559 32861
rect 25682 32852 25688 32904
rect 25740 32852 25746 32904
rect 26160 32901 26188 32932
rect 26804 32901 26832 32932
rect 27614 32920 27620 32972
rect 27672 32920 27678 32972
rect 29196 32960 29224 33056
rect 29730 32988 29736 33040
rect 29788 33028 29794 33040
rect 31404 33037 31432 33068
rect 33042 33056 33048 33068
rect 33100 33056 33106 33108
rect 33137 33099 33195 33105
rect 33137 33065 33149 33099
rect 33183 33096 33195 33099
rect 33318 33096 33324 33108
rect 33183 33068 33324 33096
rect 33183 33065 33195 33068
rect 33137 33059 33195 33065
rect 33318 33056 33324 33068
rect 33376 33056 33382 33108
rect 34072 33068 35388 33096
rect 31389 33031 31447 33037
rect 31389 33028 31401 33031
rect 29788 33000 31401 33028
rect 29788 32988 29794 33000
rect 31389 32997 31401 33000
rect 31435 32997 31447 33031
rect 31846 33028 31852 33040
rect 31389 32991 31447 32997
rect 31496 33000 31852 33028
rect 29273 32963 29331 32969
rect 29273 32960 29285 32963
rect 29196 32932 29285 32960
rect 29273 32929 29285 32932
rect 29319 32929 29331 32963
rect 29273 32923 29331 32929
rect 29638 32920 29644 32972
rect 29696 32960 29702 32972
rect 29825 32963 29883 32969
rect 29825 32960 29837 32963
rect 29696 32932 29837 32960
rect 29696 32920 29702 32932
rect 29825 32929 29837 32932
rect 29871 32929 29883 32963
rect 31496 32960 31524 33000
rect 31846 32988 31852 33000
rect 31904 33028 31910 33040
rect 32585 33031 32643 33037
rect 31904 33000 32260 33028
rect 31904 32988 31910 33000
rect 29825 32923 29883 32929
rect 30024 32932 30604 32960
rect 26145 32895 26203 32901
rect 26145 32861 26157 32895
rect 26191 32861 26203 32895
rect 26605 32895 26663 32901
rect 26605 32892 26617 32895
rect 26145 32855 26203 32861
rect 26528 32864 26617 32892
rect 26528 32836 26556 32864
rect 26605 32861 26617 32864
rect 26651 32861 26663 32895
rect 26605 32855 26663 32861
rect 26789 32895 26847 32901
rect 26789 32861 26801 32895
rect 26835 32892 26847 32895
rect 27154 32892 27160 32904
rect 26835 32864 27160 32892
rect 26835 32861 26847 32864
rect 26789 32855 26847 32861
rect 27154 32852 27160 32864
rect 27212 32852 27218 32904
rect 27709 32895 27767 32901
rect 27709 32861 27721 32895
rect 27755 32861 27767 32895
rect 29181 32895 29239 32901
rect 29181 32892 29193 32895
rect 27709 32855 27767 32861
rect 28828 32864 29193 32892
rect 21818 32784 21824 32836
rect 21876 32784 21882 32836
rect 21913 32827 21971 32833
rect 21913 32793 21925 32827
rect 21959 32824 21971 32827
rect 22370 32824 22376 32836
rect 21959 32796 22376 32824
rect 21959 32793 21971 32796
rect 21913 32787 21971 32793
rect 22370 32784 22376 32796
rect 22428 32784 22434 32836
rect 26329 32827 26387 32833
rect 26329 32793 26341 32827
rect 26375 32824 26387 32827
rect 26510 32824 26516 32836
rect 26375 32796 26516 32824
rect 26375 32793 26387 32796
rect 26329 32787 26387 32793
rect 26510 32784 26516 32796
rect 26568 32824 26574 32836
rect 27724 32824 27752 32855
rect 26568 32796 27752 32824
rect 26568 32784 26574 32796
rect 28828 32768 28856 32864
rect 29181 32861 29193 32864
rect 29227 32861 29239 32895
rect 29181 32855 29239 32861
rect 29365 32895 29423 32901
rect 29365 32861 29377 32895
rect 29411 32892 29423 32895
rect 30024 32892 30052 32932
rect 29411 32864 30052 32892
rect 29411 32861 29423 32864
rect 29365 32855 29423 32861
rect 29196 32824 29224 32855
rect 30098 32852 30104 32904
rect 30156 32852 30162 32904
rect 30282 32824 30288 32836
rect 29196 32796 30288 32824
rect 30282 32784 30288 32796
rect 30340 32824 30346 32836
rect 30576 32833 30604 32932
rect 31404 32932 31524 32960
rect 31726 32932 32168 32960
rect 31202 32852 31208 32904
rect 31260 32892 31266 32904
rect 31404 32901 31432 32932
rect 31389 32895 31447 32901
rect 31389 32892 31401 32895
rect 31260 32864 31401 32892
rect 31260 32852 31266 32864
rect 31389 32861 31401 32864
rect 31435 32861 31447 32895
rect 31389 32855 31447 32861
rect 31570 32852 31576 32904
rect 31628 32892 31634 32904
rect 31726 32892 31754 32932
rect 31628 32864 31754 32892
rect 31628 32852 31634 32864
rect 31938 32852 31944 32904
rect 31996 32892 32002 32904
rect 32140 32901 32168 32932
rect 32232 32901 32260 33000
rect 32585 32997 32597 33031
rect 32631 33028 32643 33031
rect 34072 33028 34100 33068
rect 32631 33000 34100 33028
rect 32631 32997 32643 33000
rect 32585 32991 32643 32997
rect 34146 32988 34152 33040
rect 34204 32988 34210 33040
rect 35158 33028 35164 33040
rect 34900 33000 35164 33028
rect 34900 32969 34928 33000
rect 35158 32988 35164 33000
rect 35216 32988 35222 33040
rect 34701 32963 34759 32969
rect 34701 32960 34713 32963
rect 33428 32932 34713 32960
rect 32125 32895 32183 32901
rect 31996 32864 32076 32892
rect 31996 32852 32002 32864
rect 30377 32827 30435 32833
rect 30377 32824 30389 32827
rect 30340 32796 30389 32824
rect 30340 32784 30346 32796
rect 30377 32793 30389 32796
rect 30423 32793 30435 32827
rect 30377 32787 30435 32793
rect 30561 32827 30619 32833
rect 30561 32793 30573 32827
rect 30607 32824 30619 32827
rect 32048 32824 32076 32864
rect 32125 32861 32137 32895
rect 32171 32861 32183 32895
rect 32125 32855 32183 32861
rect 32217 32895 32275 32901
rect 32217 32861 32229 32895
rect 32263 32861 32275 32895
rect 33045 32895 33103 32901
rect 33045 32892 33057 32895
rect 32217 32855 32275 32861
rect 32324 32864 33057 32892
rect 32324 32824 32352 32864
rect 33045 32861 33057 32864
rect 33091 32861 33103 32895
rect 33045 32855 33103 32861
rect 33134 32852 33140 32904
rect 33192 32892 33198 32904
rect 33428 32901 33456 32932
rect 34701 32929 34713 32932
rect 34747 32929 34759 32963
rect 34885 32963 34943 32969
rect 34885 32960 34897 32963
rect 34701 32923 34759 32929
rect 34808 32932 34897 32960
rect 33321 32895 33379 32901
rect 33321 32892 33333 32895
rect 33192 32864 33333 32892
rect 33192 32852 33198 32864
rect 33321 32861 33333 32864
rect 33367 32861 33379 32895
rect 33321 32855 33379 32861
rect 33413 32895 33471 32901
rect 33413 32861 33425 32895
rect 33459 32861 33471 32895
rect 33413 32855 33471 32861
rect 34054 32852 34060 32904
rect 34112 32892 34118 32904
rect 34149 32895 34207 32901
rect 34149 32892 34161 32895
rect 34112 32864 34161 32892
rect 34112 32852 34118 32864
rect 34149 32861 34161 32864
rect 34195 32861 34207 32895
rect 34149 32855 34207 32861
rect 34425 32895 34483 32901
rect 34425 32861 34437 32895
rect 34471 32892 34483 32895
rect 34808 32892 34836 32932
rect 34885 32929 34897 32932
rect 34931 32929 34943 32963
rect 34885 32923 34943 32929
rect 34471 32864 34836 32892
rect 34471 32861 34483 32864
rect 34425 32855 34483 32861
rect 30607 32796 31984 32824
rect 32048 32796 32352 32824
rect 30607 32793 30619 32796
rect 30561 32787 30619 32793
rect 18012 32728 20208 32756
rect 18012 32716 18018 32728
rect 20438 32716 20444 32768
rect 20496 32716 20502 32768
rect 20533 32759 20591 32765
rect 20533 32725 20545 32759
rect 20579 32756 20591 32759
rect 20714 32756 20720 32768
rect 20579 32728 20720 32756
rect 20579 32725 20591 32728
rect 20533 32719 20591 32725
rect 20714 32716 20720 32728
rect 20772 32716 20778 32768
rect 21450 32716 21456 32768
rect 21508 32756 21514 32768
rect 21545 32759 21603 32765
rect 21545 32756 21557 32759
rect 21508 32728 21557 32756
rect 21508 32716 21514 32728
rect 21545 32725 21557 32728
rect 21591 32725 21603 32759
rect 21545 32719 21603 32725
rect 22278 32716 22284 32768
rect 22336 32716 22342 32768
rect 23474 32716 23480 32768
rect 23532 32756 23538 32768
rect 24210 32756 24216 32768
rect 23532 32728 24216 32756
rect 23532 32716 23538 32728
rect 24210 32716 24216 32728
rect 24268 32716 24274 32768
rect 24302 32716 24308 32768
rect 24360 32756 24366 32768
rect 25501 32759 25559 32765
rect 25501 32756 25513 32759
rect 24360 32728 25513 32756
rect 24360 32716 24366 32728
rect 25501 32725 25513 32728
rect 25547 32725 25559 32759
rect 25501 32719 25559 32725
rect 28810 32716 28816 32768
rect 28868 32716 28874 32768
rect 29546 32716 29552 32768
rect 29604 32756 29610 32768
rect 30193 32759 30251 32765
rect 30193 32756 30205 32759
rect 29604 32728 30205 32756
rect 29604 32716 29610 32728
rect 30193 32725 30205 32728
rect 30239 32725 30251 32759
rect 30193 32719 30251 32725
rect 31754 32716 31760 32768
rect 31812 32756 31818 32768
rect 31849 32759 31907 32765
rect 31849 32756 31861 32759
rect 31812 32728 31861 32756
rect 31812 32716 31818 32728
rect 31849 32725 31861 32728
rect 31895 32725 31907 32759
rect 31956 32756 31984 32796
rect 32398 32784 32404 32836
rect 32456 32784 32462 32836
rect 33686 32824 33692 32836
rect 32508 32796 33692 32824
rect 32508 32756 32536 32796
rect 33686 32784 33692 32796
rect 33744 32784 33750 32836
rect 34164 32824 34192 32855
rect 34974 32852 34980 32904
rect 35032 32852 35038 32904
rect 35069 32895 35127 32901
rect 35069 32861 35081 32895
rect 35115 32861 35127 32895
rect 35069 32855 35127 32861
rect 35161 32895 35219 32901
rect 35161 32861 35173 32895
rect 35207 32892 35219 32895
rect 35360 32892 35388 33068
rect 36630 32892 36636 32904
rect 35207 32864 36636 32892
rect 35207 32861 35219 32864
rect 35161 32855 35219 32861
rect 35084 32824 35112 32855
rect 36630 32852 36636 32864
rect 36688 32852 36694 32904
rect 37921 32895 37979 32901
rect 37921 32861 37933 32895
rect 37967 32892 37979 32895
rect 38286 32892 38292 32904
rect 37967 32864 38292 32892
rect 37967 32861 37979 32864
rect 37921 32855 37979 32861
rect 38286 32852 38292 32864
rect 38344 32852 38350 32904
rect 34164 32796 35112 32824
rect 31956 32728 32536 32756
rect 31849 32719 31907 32725
rect 33594 32716 33600 32768
rect 33652 32716 33658 32768
rect 34333 32759 34391 32765
rect 34333 32725 34345 32759
rect 34379 32756 34391 32759
rect 34974 32756 34980 32768
rect 34379 32728 34980 32756
rect 34379 32725 34391 32728
rect 34333 32719 34391 32725
rect 34974 32716 34980 32728
rect 35032 32756 35038 32768
rect 35986 32756 35992 32768
rect 35032 32728 35992 32756
rect 35032 32716 35038 32728
rect 35986 32716 35992 32728
rect 36044 32716 36050 32768
rect 37734 32716 37740 32768
rect 37792 32716 37798 32768
rect 1104 32666 38272 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 38272 32666
rect 1104 32592 38272 32614
rect 8202 32512 8208 32564
rect 8260 32512 8266 32564
rect 17310 32512 17316 32564
rect 17368 32552 17374 32564
rect 18230 32552 18236 32564
rect 17368 32524 18236 32552
rect 17368 32512 17374 32524
rect 18230 32512 18236 32524
rect 18288 32512 18294 32564
rect 18782 32512 18788 32564
rect 18840 32552 18846 32564
rect 18877 32555 18935 32561
rect 18877 32552 18889 32555
rect 18840 32524 18889 32552
rect 18840 32512 18846 32524
rect 18877 32521 18889 32524
rect 18923 32521 18935 32555
rect 18877 32515 18935 32521
rect 18966 32512 18972 32564
rect 19024 32552 19030 32564
rect 20346 32552 20352 32564
rect 19024 32524 20352 32552
rect 19024 32512 19030 32524
rect 20346 32512 20352 32524
rect 20404 32512 20410 32564
rect 20438 32512 20444 32564
rect 20496 32512 20502 32564
rect 21818 32512 21824 32564
rect 21876 32512 21882 32564
rect 22278 32512 22284 32564
rect 22336 32512 22342 32564
rect 22370 32512 22376 32564
rect 22428 32552 22434 32564
rect 22428 32524 24256 32552
rect 22428 32512 22434 32524
rect 7929 32487 7987 32493
rect 7929 32453 7941 32487
rect 7975 32484 7987 32487
rect 8220 32484 8248 32512
rect 7975 32456 8248 32484
rect 7975 32453 7987 32456
rect 7929 32447 7987 32453
rect 8938 32444 8944 32496
rect 8996 32444 9002 32496
rect 12342 32444 12348 32496
rect 12400 32484 12406 32496
rect 12529 32487 12587 32493
rect 12529 32484 12541 32487
rect 12400 32456 12541 32484
rect 12400 32444 12406 32456
rect 12529 32453 12541 32456
rect 12575 32453 12587 32487
rect 21545 32487 21603 32493
rect 21545 32484 21557 32487
rect 12529 32447 12587 32453
rect 19720 32456 21557 32484
rect 11330 32376 11336 32428
rect 11388 32416 11394 32428
rect 12253 32419 12311 32425
rect 12253 32416 12265 32419
rect 11388 32388 12265 32416
rect 11388 32376 11394 32388
rect 12253 32385 12265 32388
rect 12299 32385 12311 32419
rect 12253 32379 12311 32385
rect 12437 32419 12495 32425
rect 12437 32385 12449 32419
rect 12483 32385 12495 32419
rect 12437 32379 12495 32385
rect 12673 32419 12731 32425
rect 12673 32385 12685 32419
rect 12719 32416 12731 32419
rect 12802 32416 12808 32428
rect 12719 32388 12808 32416
rect 12719 32385 12731 32388
rect 12673 32379 12731 32385
rect 7650 32308 7656 32360
rect 7708 32308 7714 32360
rect 7926 32308 7932 32360
rect 7984 32348 7990 32360
rect 9401 32351 9459 32357
rect 9401 32348 9413 32351
rect 7984 32320 9413 32348
rect 7984 32308 7990 32320
rect 9401 32317 9413 32320
rect 9447 32348 9459 32351
rect 11606 32348 11612 32360
rect 9447 32320 11612 32348
rect 9447 32317 9459 32320
rect 9401 32311 9459 32317
rect 11606 32308 11612 32320
rect 11664 32308 11670 32360
rect 12452 32348 12480 32379
rect 12802 32376 12808 32388
rect 12860 32416 12866 32428
rect 13538 32416 13544 32428
rect 12860 32388 13544 32416
rect 12860 32376 12866 32388
rect 13538 32376 13544 32388
rect 13596 32376 13602 32428
rect 17862 32376 17868 32428
rect 17920 32416 17926 32428
rect 18141 32419 18199 32425
rect 18141 32416 18153 32419
rect 17920 32388 18153 32416
rect 17920 32376 17926 32388
rect 18141 32385 18153 32388
rect 18187 32385 18199 32419
rect 18141 32379 18199 32385
rect 18693 32419 18751 32425
rect 18693 32385 18705 32419
rect 18739 32385 18751 32419
rect 18693 32379 18751 32385
rect 13262 32348 13268 32360
rect 12452 32320 13268 32348
rect 12636 32224 12664 32320
rect 13262 32308 13268 32320
rect 13320 32308 13326 32360
rect 16022 32308 16028 32360
rect 16080 32348 16086 32360
rect 17954 32348 17960 32360
rect 16080 32320 17960 32348
rect 16080 32308 16086 32320
rect 17954 32308 17960 32320
rect 18012 32308 18018 32360
rect 18046 32308 18052 32360
rect 18104 32348 18110 32360
rect 18598 32348 18604 32360
rect 18104 32320 18604 32348
rect 18104 32308 18110 32320
rect 18598 32308 18604 32320
rect 18656 32308 18662 32360
rect 18708 32348 18736 32379
rect 18782 32376 18788 32428
rect 18840 32416 18846 32428
rect 19334 32416 19340 32428
rect 18840 32388 19340 32416
rect 18840 32376 18846 32388
rect 19334 32376 19340 32388
rect 19392 32376 19398 32428
rect 19058 32348 19064 32360
rect 18708 32320 19064 32348
rect 19058 32308 19064 32320
rect 19116 32308 19122 32360
rect 19150 32308 19156 32360
rect 19208 32308 19214 32360
rect 19242 32308 19248 32360
rect 19300 32348 19306 32360
rect 19613 32351 19671 32357
rect 19613 32348 19625 32351
rect 19300 32320 19625 32348
rect 19300 32308 19306 32320
rect 19613 32317 19625 32320
rect 19659 32317 19671 32351
rect 19720 32348 19748 32456
rect 19797 32419 19855 32425
rect 19797 32385 19809 32419
rect 19843 32416 19855 32419
rect 20349 32419 20407 32425
rect 20349 32416 20361 32419
rect 19843 32388 20361 32416
rect 19843 32385 19855 32388
rect 19797 32379 19855 32385
rect 20349 32385 20361 32388
rect 20395 32416 20407 32419
rect 20438 32416 20444 32428
rect 20395 32388 20444 32416
rect 20395 32385 20407 32388
rect 20349 32379 20407 32385
rect 20438 32376 20444 32388
rect 20496 32376 20502 32428
rect 20548 32425 20576 32456
rect 21545 32453 21557 32456
rect 21591 32484 21603 32487
rect 22296 32484 22324 32512
rect 21591 32456 21956 32484
rect 22296 32456 22600 32484
rect 21591 32453 21603 32456
rect 21545 32447 21603 32453
rect 20533 32419 20591 32425
rect 20533 32385 20545 32419
rect 20579 32385 20591 32419
rect 20533 32379 20591 32385
rect 20622 32376 20628 32428
rect 20680 32376 20686 32428
rect 21177 32419 21235 32425
rect 21177 32385 21189 32419
rect 21223 32385 21235 32419
rect 21177 32379 21235 32385
rect 21361 32419 21419 32425
rect 21361 32385 21373 32419
rect 21407 32414 21419 32419
rect 21450 32414 21456 32428
rect 21407 32386 21456 32414
rect 21407 32385 21419 32386
rect 21361 32379 21419 32385
rect 19889 32351 19947 32357
rect 19889 32348 19901 32351
rect 19720 32320 19901 32348
rect 19613 32311 19671 32317
rect 19889 32317 19901 32320
rect 19935 32317 19947 32351
rect 19889 32311 19947 32317
rect 19981 32351 20039 32357
rect 19981 32317 19993 32351
rect 20027 32317 20039 32351
rect 19981 32311 20039 32317
rect 14366 32240 14372 32292
rect 14424 32280 14430 32292
rect 19996 32280 20024 32311
rect 20070 32308 20076 32360
rect 20128 32308 20134 32360
rect 21192 32348 21220 32379
rect 21450 32376 21456 32386
rect 21508 32416 21514 32428
rect 21637 32419 21695 32425
rect 21508 32388 21553 32416
rect 21508 32376 21514 32388
rect 21637 32385 21649 32419
rect 21683 32416 21695 32419
rect 21928 32416 21956 32456
rect 22572 32425 22600 32456
rect 22646 32444 22652 32496
rect 22704 32444 22710 32496
rect 23661 32487 23719 32493
rect 23661 32484 23673 32487
rect 22756 32456 22968 32484
rect 22373 32419 22431 32425
rect 22373 32416 22385 32419
rect 21683 32414 21772 32416
rect 21683 32388 21864 32414
rect 21928 32388 22385 32416
rect 21683 32385 21695 32388
rect 21744 32386 21864 32388
rect 21637 32379 21695 32385
rect 21836 32348 21864 32386
rect 22373 32385 22385 32388
rect 22419 32385 22431 32419
rect 22373 32379 22431 32385
rect 22557 32419 22615 32425
rect 22557 32385 22569 32419
rect 22603 32385 22615 32419
rect 22557 32379 22615 32385
rect 22278 32348 22284 32360
rect 21192 32320 22284 32348
rect 22278 32308 22284 32320
rect 22336 32308 22342 32360
rect 20717 32283 20775 32289
rect 20717 32280 20729 32283
rect 14424 32252 18644 32280
rect 19996 32252 20729 32280
rect 14424 32240 14430 32252
rect 12618 32172 12624 32224
rect 12676 32172 12682 32224
rect 12805 32215 12863 32221
rect 12805 32181 12817 32215
rect 12851 32212 12863 32215
rect 18046 32212 18052 32224
rect 12851 32184 18052 32212
rect 12851 32181 12863 32184
rect 12805 32175 12863 32181
rect 18046 32172 18052 32184
rect 18104 32172 18110 32224
rect 18233 32215 18291 32221
rect 18233 32181 18245 32215
rect 18279 32212 18291 32215
rect 18506 32212 18512 32224
rect 18279 32184 18512 32212
rect 18279 32181 18291 32184
rect 18233 32175 18291 32181
rect 18506 32172 18512 32184
rect 18564 32172 18570 32224
rect 18616 32212 18644 32252
rect 20717 32249 20729 32252
rect 20763 32249 20775 32283
rect 20717 32243 20775 32249
rect 21174 32240 21180 32292
rect 21232 32280 21238 32292
rect 21361 32283 21419 32289
rect 21361 32280 21373 32283
rect 21232 32252 21373 32280
rect 21232 32240 21238 32252
rect 21361 32249 21373 32252
rect 21407 32249 21419 32283
rect 21361 32243 21419 32249
rect 21450 32240 21456 32292
rect 21508 32280 21514 32292
rect 21913 32283 21971 32289
rect 21913 32280 21925 32283
rect 21508 32252 21925 32280
rect 21508 32240 21514 32252
rect 21913 32249 21925 32252
rect 21959 32249 21971 32283
rect 22756 32280 22784 32456
rect 22940 32425 22968 32456
rect 23216 32456 23673 32484
rect 23216 32428 23244 32456
rect 23661 32453 23673 32456
rect 23707 32453 23719 32487
rect 23661 32447 23719 32453
rect 23842 32444 23848 32496
rect 23900 32484 23906 32496
rect 23900 32456 24072 32484
rect 23900 32444 23906 32456
rect 22833 32419 22891 32425
rect 22833 32385 22845 32419
rect 22879 32385 22891 32419
rect 22833 32379 22891 32385
rect 22925 32419 22983 32425
rect 22925 32385 22937 32419
rect 22971 32385 22983 32419
rect 22925 32379 22983 32385
rect 22848 32348 22876 32379
rect 23014 32376 23020 32428
rect 23072 32416 23078 32428
rect 23109 32419 23167 32425
rect 23109 32416 23121 32419
rect 23072 32388 23121 32416
rect 23072 32376 23078 32388
rect 23109 32385 23121 32388
rect 23155 32385 23167 32419
rect 23109 32379 23167 32385
rect 23198 32376 23204 32428
rect 23256 32376 23262 32428
rect 23566 32376 23572 32428
rect 23624 32376 23630 32428
rect 24044 32425 24072 32456
rect 24118 32444 24124 32496
rect 24176 32444 24182 32496
rect 24228 32493 24256 32524
rect 29546 32512 29552 32564
rect 29604 32552 29610 32564
rect 29841 32555 29899 32561
rect 29841 32552 29853 32555
rect 29604 32524 29853 32552
rect 29604 32512 29610 32524
rect 29841 32521 29853 32524
rect 29887 32521 29899 32555
rect 29841 32515 29899 32521
rect 30006 32512 30012 32564
rect 30064 32512 30070 32564
rect 30190 32512 30196 32564
rect 30248 32512 30254 32564
rect 31478 32512 31484 32564
rect 31536 32552 31542 32564
rect 31536 32524 32444 32552
rect 31536 32512 31542 32524
rect 24213 32487 24271 32493
rect 24213 32453 24225 32487
rect 24259 32453 24271 32487
rect 25041 32487 25099 32493
rect 25041 32484 25053 32487
rect 24213 32447 24271 32453
rect 24320 32456 25053 32484
rect 23753 32419 23811 32425
rect 23753 32385 23765 32419
rect 23799 32385 23811 32419
rect 23753 32379 23811 32385
rect 24029 32419 24087 32425
rect 24029 32385 24041 32419
rect 24075 32385 24087 32419
rect 24029 32379 24087 32385
rect 23382 32348 23388 32360
rect 22848 32320 23388 32348
rect 23382 32308 23388 32320
rect 23440 32308 23446 32360
rect 23768 32348 23796 32379
rect 24320 32348 24348 32456
rect 25041 32453 25053 32456
rect 25087 32453 25099 32487
rect 25041 32447 25099 32453
rect 29178 32444 29184 32496
rect 29236 32484 29242 32496
rect 29641 32487 29699 32493
rect 29641 32484 29653 32487
rect 29236 32456 29653 32484
rect 29236 32444 29242 32456
rect 29641 32453 29653 32456
rect 29687 32453 29699 32487
rect 30208 32484 30236 32512
rect 31570 32484 31576 32496
rect 30208 32456 31576 32484
rect 29641 32447 29699 32453
rect 31570 32444 31576 32456
rect 31628 32484 31634 32496
rect 32309 32487 32367 32493
rect 32309 32484 32321 32487
rect 31628 32456 32321 32484
rect 31628 32444 31634 32456
rect 32309 32453 32321 32456
rect 32355 32453 32367 32487
rect 32309 32447 32367 32453
rect 32416 32428 32444 32524
rect 33594 32484 33600 32496
rect 33244 32456 33600 32484
rect 24394 32376 24400 32428
rect 24452 32376 24458 32428
rect 24489 32419 24547 32425
rect 24489 32385 24501 32419
rect 24535 32385 24547 32419
rect 24489 32379 24547 32385
rect 23768 32320 24348 32348
rect 23750 32280 23756 32292
rect 22756 32252 23756 32280
rect 21913 32243 21971 32249
rect 23750 32240 23756 32252
rect 23808 32240 23814 32292
rect 24504 32280 24532 32379
rect 24578 32376 24584 32428
rect 24636 32416 24642 32428
rect 24673 32419 24731 32425
rect 24673 32416 24685 32419
rect 24636 32388 24685 32416
rect 24636 32376 24642 32388
rect 24673 32385 24685 32388
rect 24719 32416 24731 32419
rect 24949 32419 25007 32425
rect 24949 32416 24961 32419
rect 24719 32388 24961 32416
rect 24719 32385 24731 32388
rect 24673 32379 24731 32385
rect 24949 32385 24961 32388
rect 24995 32385 25007 32419
rect 24949 32379 25007 32385
rect 25130 32376 25136 32428
rect 25188 32416 25194 32428
rect 25188 32388 31754 32416
rect 25188 32376 25194 32388
rect 31726 32348 31754 32388
rect 32122 32376 32128 32428
rect 32180 32376 32186 32428
rect 32398 32376 32404 32428
rect 32456 32416 32462 32428
rect 32858 32416 32864 32428
rect 32456 32388 32864 32416
rect 32456 32376 32462 32388
rect 32858 32376 32864 32388
rect 32916 32376 32922 32428
rect 33244 32425 33272 32456
rect 33594 32444 33600 32456
rect 33652 32444 33658 32496
rect 33229 32419 33287 32425
rect 33229 32385 33241 32419
rect 33275 32385 33287 32419
rect 33229 32379 33287 32385
rect 33686 32376 33692 32428
rect 33744 32376 33750 32428
rect 33965 32419 34023 32425
rect 33965 32385 33977 32419
rect 34011 32416 34023 32419
rect 34425 32419 34483 32425
rect 34425 32416 34437 32419
rect 34011 32388 34437 32416
rect 34011 32385 34023 32388
rect 33965 32379 34023 32385
rect 34425 32385 34437 32388
rect 34471 32385 34483 32419
rect 34425 32379 34483 32385
rect 31726 32320 33364 32348
rect 24136 32252 24532 32280
rect 24596 32252 24992 32280
rect 24136 32224 24164 32252
rect 22002 32212 22008 32224
rect 18616 32184 22008 32212
rect 22002 32172 22008 32184
rect 22060 32172 22066 32224
rect 22462 32172 22468 32224
rect 22520 32172 22526 32224
rect 23014 32172 23020 32224
rect 23072 32212 23078 32224
rect 23474 32212 23480 32224
rect 23072 32184 23480 32212
rect 23072 32172 23078 32184
rect 23474 32172 23480 32184
rect 23532 32172 23538 32224
rect 23566 32172 23572 32224
rect 23624 32212 23630 32224
rect 23845 32215 23903 32221
rect 23845 32212 23857 32215
rect 23624 32184 23857 32212
rect 23624 32172 23630 32184
rect 23845 32181 23857 32184
rect 23891 32212 23903 32215
rect 24118 32212 24124 32224
rect 23891 32184 24124 32212
rect 23891 32181 23903 32184
rect 23845 32175 23903 32181
rect 24118 32172 24124 32184
rect 24176 32172 24182 32224
rect 24210 32172 24216 32224
rect 24268 32212 24274 32224
rect 24596 32212 24624 32252
rect 24268 32184 24624 32212
rect 24268 32172 24274 32184
rect 24854 32172 24860 32224
rect 24912 32172 24918 32224
rect 24964 32212 24992 32252
rect 26050 32240 26056 32292
rect 26108 32280 26114 32292
rect 32861 32283 32919 32289
rect 32861 32280 32873 32283
rect 26108 32252 32873 32280
rect 26108 32240 26114 32252
rect 32861 32249 32873 32252
rect 32907 32249 32919 32283
rect 33336 32280 33364 32320
rect 33410 32308 33416 32360
rect 33468 32308 33474 32360
rect 33704 32348 33732 32376
rect 34330 32348 34336 32360
rect 33704 32320 34336 32348
rect 34330 32308 34336 32320
rect 34388 32308 34394 32360
rect 34606 32308 34612 32360
rect 34664 32308 34670 32360
rect 34698 32308 34704 32360
rect 34756 32308 34762 32360
rect 35069 32351 35127 32357
rect 35069 32317 35081 32351
rect 35115 32348 35127 32351
rect 35342 32348 35348 32360
rect 35115 32320 35348 32348
rect 35115 32317 35127 32320
rect 35069 32311 35127 32317
rect 35342 32308 35348 32320
rect 35400 32308 35406 32360
rect 37734 32308 37740 32360
rect 37792 32308 37798 32360
rect 37752 32280 37780 32308
rect 33336 32252 37780 32280
rect 32861 32243 32919 32249
rect 27798 32212 27804 32224
rect 24964 32184 27804 32212
rect 27798 32172 27804 32184
rect 27856 32172 27862 32224
rect 29730 32172 29736 32224
rect 29788 32212 29794 32224
rect 29825 32215 29883 32221
rect 29825 32212 29837 32215
rect 29788 32184 29837 32212
rect 29788 32172 29794 32184
rect 29825 32181 29837 32184
rect 29871 32181 29883 32215
rect 29825 32175 29883 32181
rect 32493 32215 32551 32221
rect 32493 32181 32505 32215
rect 32539 32212 32551 32215
rect 33318 32212 33324 32224
rect 32539 32184 33324 32212
rect 32539 32181 32551 32184
rect 32493 32175 32551 32181
rect 33318 32172 33324 32184
rect 33376 32172 33382 32224
rect 1104 32122 38272 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38272 32122
rect 1104 32048 38272 32070
rect 3789 32011 3847 32017
rect 3789 31977 3801 32011
rect 3835 32008 3847 32011
rect 4798 32008 4804 32020
rect 3835 31980 4804 32008
rect 3835 31977 3847 31980
rect 3789 31971 3847 31977
rect 4798 31968 4804 31980
rect 4856 31968 4862 32020
rect 19058 31968 19064 32020
rect 19116 32008 19122 32020
rect 20714 32008 20720 32020
rect 19116 31980 20720 32008
rect 19116 31968 19122 31980
rect 20714 31968 20720 31980
rect 20772 32008 20778 32020
rect 21453 32011 21511 32017
rect 21453 32008 21465 32011
rect 20772 31980 21465 32008
rect 20772 31968 20778 31980
rect 21453 31977 21465 31980
rect 21499 31977 21511 32011
rect 21453 31971 21511 31977
rect 21818 31968 21824 32020
rect 21876 31968 21882 32020
rect 23014 32008 23020 32020
rect 22066 31980 23020 32008
rect 14550 31900 14556 31952
rect 14608 31900 14614 31952
rect 19076 31940 19104 31968
rect 18156 31912 19104 31940
rect 4062 31872 4068 31884
rect 3988 31844 4068 31872
rect 3326 31764 3332 31816
rect 3384 31804 3390 31816
rect 3988 31804 4016 31844
rect 4062 31832 4068 31844
rect 4120 31872 4126 31884
rect 5537 31875 5595 31881
rect 5537 31872 5549 31875
rect 4120 31844 5549 31872
rect 4120 31832 4126 31844
rect 5537 31841 5549 31844
rect 5583 31872 5595 31875
rect 6365 31875 6423 31881
rect 6365 31872 6377 31875
rect 5583 31844 6377 31872
rect 5583 31841 5595 31844
rect 5537 31835 5595 31841
rect 6365 31841 6377 31844
rect 6411 31872 6423 31875
rect 7006 31872 7012 31884
rect 6411 31844 7012 31872
rect 6411 31841 6423 31844
rect 6365 31835 6423 31841
rect 7006 31832 7012 31844
rect 7064 31872 7070 31884
rect 7650 31872 7656 31884
rect 7064 31844 7656 31872
rect 7064 31832 7070 31844
rect 7650 31832 7656 31844
rect 7708 31832 7714 31884
rect 8478 31832 8484 31884
rect 8536 31872 8542 31884
rect 12986 31872 12992 31884
rect 8536 31844 12992 31872
rect 8536 31832 8542 31844
rect 12986 31832 12992 31844
rect 13044 31832 13050 31884
rect 3384 31776 4016 31804
rect 3384 31764 3390 31776
rect 4154 31764 4160 31816
rect 4212 31764 4218 31816
rect 8662 31804 8668 31816
rect 7774 31790 8668 31804
rect 7760 31776 8668 31790
rect 4172 31668 4200 31764
rect 5258 31696 5264 31748
rect 5316 31696 5322 31748
rect 6638 31696 6644 31748
rect 6696 31696 6702 31748
rect 5442 31668 5448 31680
rect 4172 31640 5448 31668
rect 5442 31628 5448 31640
rect 5500 31668 5506 31680
rect 7760 31668 7788 31776
rect 8662 31764 8668 31776
rect 8720 31804 8726 31816
rect 9582 31804 9588 31816
rect 8720 31776 9588 31804
rect 8720 31764 8726 31776
rect 9582 31764 9588 31776
rect 9640 31764 9646 31816
rect 11514 31764 11520 31816
rect 11572 31804 11578 31816
rect 11609 31807 11667 31813
rect 11609 31804 11621 31807
rect 11572 31776 11621 31804
rect 11572 31764 11578 31776
rect 11609 31773 11621 31776
rect 11655 31773 11667 31807
rect 11609 31767 11667 31773
rect 11790 31764 11796 31816
rect 11848 31764 11854 31816
rect 11974 31764 11980 31816
rect 12032 31764 12038 31816
rect 12069 31807 12127 31813
rect 12069 31773 12081 31807
rect 12115 31804 12127 31807
rect 12250 31804 12256 31816
rect 12115 31776 12256 31804
rect 12115 31773 12127 31776
rect 12069 31767 12127 31773
rect 11698 31696 11704 31748
rect 11756 31736 11762 31748
rect 12084 31736 12112 31767
rect 12250 31764 12256 31776
rect 12308 31764 12314 31816
rect 12342 31764 12348 31816
rect 12400 31804 12406 31816
rect 12526 31804 12532 31816
rect 12400 31776 12532 31804
rect 12400 31764 12406 31776
rect 12526 31764 12532 31776
rect 12584 31764 12590 31816
rect 14568 31804 14596 31900
rect 14921 31875 14979 31881
rect 14921 31841 14933 31875
rect 14967 31872 14979 31875
rect 16482 31872 16488 31884
rect 14967 31844 15976 31872
rect 14967 31841 14979 31844
rect 14921 31835 14979 31841
rect 14826 31804 14832 31816
rect 14568 31776 14832 31804
rect 14826 31764 14832 31776
rect 14884 31764 14890 31816
rect 15948 31813 15976 31844
rect 16224 31844 16488 31872
rect 16224 31816 16252 31844
rect 16482 31832 16488 31844
rect 16540 31872 16546 31884
rect 18156 31881 18184 31912
rect 19886 31900 19892 31952
rect 19944 31940 19950 31952
rect 21726 31940 21732 31952
rect 19944 31912 21732 31940
rect 19944 31900 19950 31912
rect 21726 31900 21732 31912
rect 21784 31900 21790 31952
rect 17957 31875 18015 31881
rect 17957 31872 17969 31875
rect 16540 31844 17969 31872
rect 16540 31832 16546 31844
rect 17957 31841 17969 31844
rect 18003 31841 18015 31875
rect 17957 31835 18015 31841
rect 18141 31875 18199 31881
rect 18141 31841 18153 31875
rect 18187 31841 18199 31875
rect 18141 31835 18199 31841
rect 18325 31875 18383 31881
rect 18325 31841 18337 31875
rect 18371 31872 18383 31875
rect 18506 31872 18512 31884
rect 18371 31844 18512 31872
rect 18371 31841 18383 31844
rect 18325 31835 18383 31841
rect 18506 31832 18512 31844
rect 18564 31832 18570 31884
rect 15841 31807 15899 31813
rect 15841 31804 15853 31807
rect 15488 31776 15853 31804
rect 11756 31708 12112 31736
rect 11756 31696 11762 31708
rect 5500 31640 7788 31668
rect 5500 31628 5506 31640
rect 8110 31628 8116 31680
rect 8168 31668 8174 31680
rect 12360 31668 12388 31764
rect 15488 31680 15516 31776
rect 15841 31773 15853 31776
rect 15887 31773 15899 31807
rect 15841 31767 15899 31773
rect 15933 31807 15991 31813
rect 15933 31773 15945 31807
rect 15979 31773 15991 31807
rect 15933 31767 15991 31773
rect 16114 31764 16120 31816
rect 16172 31764 16178 31816
rect 16206 31764 16212 31816
rect 16264 31764 16270 31816
rect 18233 31807 18291 31813
rect 18233 31773 18245 31807
rect 18279 31804 18291 31807
rect 18417 31807 18475 31813
rect 18279 31776 18368 31804
rect 18279 31773 18291 31776
rect 18233 31767 18291 31773
rect 18340 31736 18368 31776
rect 18417 31773 18429 31807
rect 18463 31804 18475 31807
rect 19058 31804 19064 31816
rect 18463 31776 19064 31804
rect 18463 31773 18475 31776
rect 18417 31767 18475 31773
rect 19058 31764 19064 31776
rect 19116 31764 19122 31816
rect 21637 31807 21695 31813
rect 21637 31773 21649 31807
rect 21683 31804 21695 31807
rect 21836 31804 21864 31968
rect 22066 31884 22094 31980
rect 23014 31968 23020 31980
rect 23072 31968 23078 32020
rect 23198 31968 23204 32020
rect 23256 31968 23262 32020
rect 24397 32011 24455 32017
rect 24397 32008 24409 32011
rect 23400 31980 24409 32008
rect 22002 31832 22008 31884
rect 22060 31844 22094 31884
rect 22060 31832 22066 31844
rect 22738 31832 22744 31884
rect 22796 31832 22802 31884
rect 21683 31776 21864 31804
rect 21913 31807 21971 31813
rect 21683 31773 21695 31776
rect 21637 31767 21695 31773
rect 21913 31773 21925 31807
rect 21959 31804 21971 31807
rect 22649 31807 22707 31813
rect 22649 31804 22661 31807
rect 21959 31776 22661 31804
rect 21959 31773 21971 31776
rect 21913 31767 21971 31773
rect 22649 31773 22661 31776
rect 22695 31804 22707 31807
rect 23109 31807 23167 31813
rect 22695 31776 23060 31804
rect 22695 31773 22707 31776
rect 22649 31767 22707 31773
rect 18782 31736 18788 31748
rect 18340 31708 18788 31736
rect 18782 31696 18788 31708
rect 18840 31696 18846 31748
rect 21821 31739 21879 31745
rect 21821 31705 21833 31739
rect 21867 31736 21879 31739
rect 22462 31736 22468 31748
rect 21867 31708 22468 31736
rect 21867 31705 21879 31708
rect 21821 31699 21879 31705
rect 22462 31696 22468 31708
rect 22520 31696 22526 31748
rect 23032 31736 23060 31776
rect 23109 31773 23121 31807
rect 23155 31804 23167 31807
rect 23216 31804 23244 31968
rect 23400 31940 23428 31980
rect 24397 31977 24409 31980
rect 24443 31977 24455 32011
rect 24397 31971 24455 31977
rect 24854 31968 24860 32020
rect 24912 31968 24918 32020
rect 25777 32011 25835 32017
rect 25777 31977 25789 32011
rect 25823 32008 25835 32011
rect 27154 32008 27160 32020
rect 25823 31980 27160 32008
rect 25823 31977 25835 31980
rect 25777 31971 25835 31977
rect 27154 31968 27160 31980
rect 27212 31968 27218 32020
rect 32309 32011 32367 32017
rect 32309 32008 32321 32011
rect 32048 31980 32321 32008
rect 23750 31940 23756 31952
rect 23155 31776 23244 31804
rect 23308 31912 23428 31940
rect 23492 31912 23756 31940
rect 23155 31773 23167 31776
rect 23109 31767 23167 31773
rect 23308 31736 23336 31912
rect 23382 31764 23388 31816
rect 23440 31764 23446 31816
rect 23492 31804 23520 31912
rect 23750 31900 23756 31912
rect 23808 31900 23814 31952
rect 24872 31940 24900 31968
rect 24228 31912 24900 31940
rect 23676 31844 24164 31872
rect 23676 31813 23704 31844
rect 23569 31807 23627 31813
rect 23569 31804 23581 31807
rect 23492 31776 23581 31804
rect 23032 31708 23336 31736
rect 8168 31640 12388 31668
rect 8168 31628 8174 31640
rect 13814 31628 13820 31680
rect 13872 31668 13878 31680
rect 14090 31668 14096 31680
rect 13872 31640 14096 31668
rect 13872 31628 13878 31640
rect 14090 31628 14096 31640
rect 14148 31668 14154 31680
rect 15286 31668 15292 31680
rect 14148 31640 15292 31668
rect 14148 31628 14154 31640
rect 15286 31628 15292 31640
rect 15344 31628 15350 31680
rect 15470 31628 15476 31680
rect 15528 31628 15534 31680
rect 16390 31628 16396 31680
rect 16448 31628 16454 31680
rect 16574 31628 16580 31680
rect 16632 31668 16638 31680
rect 20162 31668 20168 31680
rect 16632 31640 20168 31668
rect 16632 31628 16638 31640
rect 20162 31628 20168 31640
rect 20220 31628 20226 31680
rect 22186 31628 22192 31680
rect 22244 31628 22250 31680
rect 22557 31671 22615 31677
rect 22557 31637 22569 31671
rect 22603 31668 22615 31671
rect 23207 31671 23265 31677
rect 23207 31668 23219 31671
rect 22603 31640 23219 31668
rect 22603 31637 22615 31640
rect 22557 31631 22615 31637
rect 23207 31637 23219 31640
rect 23253 31637 23265 31671
rect 23207 31631 23265 31637
rect 23293 31671 23351 31677
rect 23293 31637 23305 31671
rect 23339 31668 23351 31671
rect 23492 31668 23520 31776
rect 23569 31773 23581 31776
rect 23615 31773 23627 31807
rect 23569 31767 23627 31773
rect 23661 31807 23719 31813
rect 23661 31773 23673 31807
rect 23707 31773 23719 31807
rect 23661 31767 23719 31773
rect 23750 31764 23756 31816
rect 23808 31804 23814 31816
rect 23845 31807 23903 31813
rect 23845 31804 23857 31807
rect 23808 31776 23857 31804
rect 23808 31764 23814 31776
rect 23845 31773 23857 31776
rect 23891 31773 23903 31807
rect 23845 31767 23903 31773
rect 24029 31807 24087 31813
rect 24029 31773 24041 31807
rect 24075 31773 24087 31807
rect 24029 31767 24087 31773
rect 23339 31640 23520 31668
rect 24044 31668 24072 31767
rect 24136 31736 24164 31844
rect 24228 31813 24256 31912
rect 27798 31900 27804 31952
rect 27856 31900 27862 31952
rect 24578 31832 24584 31884
rect 24636 31872 24642 31884
rect 24688 31872 24900 31880
rect 27709 31875 27767 31881
rect 24636 31852 26280 31872
rect 24636 31844 24716 31852
rect 24872 31844 26280 31852
rect 24636 31832 24642 31844
rect 24213 31807 24271 31813
rect 24213 31773 24225 31807
rect 24259 31773 24271 31807
rect 24213 31767 24271 31773
rect 24673 31807 24731 31813
rect 24673 31773 24685 31807
rect 24719 31773 24731 31807
rect 24673 31767 24731 31773
rect 25685 31807 25743 31813
rect 25685 31773 25697 31807
rect 25731 31773 25743 31807
rect 25685 31767 25743 31773
rect 25869 31807 25927 31813
rect 25869 31773 25881 31807
rect 25915 31773 25927 31807
rect 26252 31804 26280 31844
rect 27709 31841 27721 31875
rect 27755 31872 27767 31875
rect 29730 31872 29736 31884
rect 27755 31844 29736 31872
rect 27755 31841 27767 31844
rect 27709 31835 27767 31841
rect 29730 31832 29736 31844
rect 29788 31832 29794 31884
rect 31570 31832 31576 31884
rect 31628 31832 31634 31884
rect 27890 31804 27896 31816
rect 26252 31776 27896 31804
rect 25869 31767 25927 31773
rect 24688 31736 24716 31767
rect 24136 31708 24716 31736
rect 25700 31680 25728 31767
rect 24394 31668 24400 31680
rect 24044 31640 24400 31668
rect 23339 31637 23351 31640
rect 23293 31631 23351 31637
rect 24394 31628 24400 31640
rect 24452 31668 24458 31680
rect 25041 31671 25099 31677
rect 25041 31668 25053 31671
rect 24452 31640 25053 31668
rect 24452 31628 24458 31640
rect 25041 31637 25053 31640
rect 25087 31637 25099 31671
rect 25041 31631 25099 31637
rect 25682 31628 25688 31680
rect 25740 31628 25746 31680
rect 25774 31628 25780 31680
rect 25832 31668 25838 31680
rect 25884 31668 25912 31767
rect 27890 31764 27896 31776
rect 27948 31764 27954 31816
rect 27985 31807 28043 31813
rect 27985 31773 27997 31807
rect 28031 31804 28043 31807
rect 28074 31804 28080 31816
rect 28031 31776 28080 31804
rect 28031 31773 28043 31776
rect 27985 31767 28043 31773
rect 28074 31764 28080 31776
rect 28132 31764 28138 31816
rect 31478 31764 31484 31816
rect 31536 31804 31542 31816
rect 32048 31804 32076 31980
rect 32309 31977 32321 31980
rect 32355 31977 32367 32011
rect 32309 31971 32367 31977
rect 34698 31968 34704 32020
rect 34756 31968 34762 32020
rect 32122 31900 32128 31952
rect 32180 31940 32186 31952
rect 34716 31940 34744 31968
rect 32180 31912 34744 31940
rect 32180 31900 32186 31912
rect 32140 31813 32168 31900
rect 32306 31832 32312 31884
rect 32364 31832 32370 31884
rect 31536 31776 32076 31804
rect 32125 31807 32183 31813
rect 31536 31764 31542 31776
rect 32125 31773 32137 31807
rect 32171 31773 32183 31807
rect 32125 31767 32183 31773
rect 32324 31804 32352 31832
rect 32401 31807 32459 31813
rect 32401 31804 32413 31807
rect 32324 31776 32413 31804
rect 30006 31696 30012 31748
rect 30064 31736 30070 31748
rect 32324 31736 32352 31776
rect 32401 31773 32413 31776
rect 32447 31773 32459 31807
rect 32401 31767 32459 31773
rect 33781 31807 33839 31813
rect 33781 31773 33793 31807
rect 33827 31804 33839 31807
rect 33888 31804 33916 31912
rect 34146 31832 34152 31884
rect 34204 31832 34210 31884
rect 34330 31832 34336 31884
rect 34388 31832 34394 31884
rect 33827 31776 33916 31804
rect 34057 31807 34115 31813
rect 33827 31773 33839 31776
rect 33781 31767 33839 31773
rect 34057 31773 34069 31807
rect 34103 31804 34115 31807
rect 34103 31776 34376 31804
rect 34103 31773 34115 31776
rect 34057 31767 34115 31773
rect 30064 31708 32352 31736
rect 30064 31696 30070 31708
rect 34348 31680 34376 31776
rect 25832 31640 25912 31668
rect 25832 31628 25838 31640
rect 26326 31628 26332 31680
rect 26384 31668 26390 31680
rect 34238 31668 34244 31680
rect 26384 31640 34244 31668
rect 26384 31628 26390 31640
rect 34238 31628 34244 31640
rect 34296 31628 34302 31680
rect 34330 31628 34336 31680
rect 34388 31628 34394 31680
rect 1104 31578 38272 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 38272 31578
rect 1104 31504 38272 31526
rect 4893 31467 4951 31473
rect 4893 31433 4905 31467
rect 4939 31464 4951 31467
rect 5258 31464 5264 31476
rect 4939 31436 5264 31464
rect 4939 31433 4951 31436
rect 4893 31427 4951 31433
rect 5258 31424 5264 31436
rect 5316 31424 5322 31476
rect 6549 31467 6607 31473
rect 6549 31433 6561 31467
rect 6595 31464 6607 31467
rect 6638 31464 6644 31476
rect 6595 31436 6644 31464
rect 6595 31433 6607 31436
rect 6549 31427 6607 31433
rect 6638 31424 6644 31436
rect 6696 31424 6702 31476
rect 7650 31424 7656 31476
rect 7708 31464 7714 31476
rect 8757 31467 8815 31473
rect 8757 31464 8769 31467
rect 7708 31436 8769 31464
rect 7708 31424 7714 31436
rect 8757 31433 8769 31436
rect 8803 31464 8815 31467
rect 9214 31464 9220 31476
rect 8803 31436 9220 31464
rect 8803 31433 8815 31436
rect 8757 31427 8815 31433
rect 9214 31424 9220 31436
rect 9272 31424 9278 31476
rect 12434 31464 12440 31476
rect 9692 31436 12440 31464
rect 2622 31368 4200 31396
rect 4172 31340 4200 31368
rect 6454 31356 6460 31408
rect 6512 31396 6518 31408
rect 7009 31399 7067 31405
rect 7009 31396 7021 31399
rect 6512 31368 7021 31396
rect 6512 31356 6518 31368
rect 7009 31365 7021 31368
rect 7055 31365 7067 31399
rect 7009 31359 7067 31365
rect 7466 31356 7472 31408
rect 7524 31396 7530 31408
rect 9692 31396 9720 31436
rect 12434 31424 12440 31436
rect 12492 31424 12498 31476
rect 12618 31464 12624 31476
rect 12544 31436 12624 31464
rect 7524 31368 9720 31396
rect 7524 31356 7530 31368
rect 9858 31356 9864 31408
rect 9916 31396 9922 31408
rect 11241 31399 11299 31405
rect 9916 31368 10074 31396
rect 9916 31356 9922 31368
rect 11241 31365 11253 31399
rect 11287 31396 11299 31399
rect 11793 31399 11851 31405
rect 11793 31396 11805 31399
rect 11287 31368 11805 31396
rect 11287 31365 11299 31368
rect 11241 31359 11299 31365
rect 11793 31365 11805 31368
rect 11839 31365 11851 31399
rect 11793 31359 11851 31365
rect 11882 31356 11888 31408
rect 11940 31356 11946 31408
rect 12158 31356 12164 31408
rect 12216 31396 12222 31408
rect 12216 31368 12388 31396
rect 12216 31356 12222 31368
rect 3326 31288 3332 31340
rect 3384 31288 3390 31340
rect 4154 31288 4160 31340
rect 4212 31328 4218 31340
rect 4982 31328 4988 31340
rect 4212 31300 4988 31328
rect 4212 31288 4218 31300
rect 4982 31288 4988 31300
rect 5040 31288 5046 31340
rect 6365 31331 6423 31337
rect 6365 31297 6377 31331
rect 6411 31328 6423 31331
rect 7101 31331 7159 31337
rect 6411 31300 6684 31328
rect 6411 31297 6423 31300
rect 6365 31291 6423 31297
rect 3050 31220 3056 31272
rect 3108 31220 3114 31272
rect 3418 31220 3424 31272
rect 3476 31220 3482 31272
rect 4341 31263 4399 31269
rect 4341 31229 4353 31263
rect 4387 31260 4399 31263
rect 4614 31260 4620 31272
rect 4387 31232 4620 31260
rect 4387 31229 4399 31232
rect 4341 31223 4399 31229
rect 4614 31220 4620 31232
rect 4672 31220 4678 31272
rect 5074 31220 5080 31272
rect 5132 31260 5138 31272
rect 5629 31263 5687 31269
rect 5629 31260 5641 31263
rect 5132 31232 5641 31260
rect 5132 31220 5138 31232
rect 5629 31229 5641 31232
rect 5675 31229 5687 31263
rect 5629 31223 5687 31229
rect 1581 31127 1639 31133
rect 1581 31093 1593 31127
rect 1627 31124 1639 31127
rect 3436 31124 3464 31220
rect 6656 31201 6684 31300
rect 7101 31297 7113 31331
rect 7147 31328 7159 31331
rect 8110 31328 8116 31340
rect 7147 31300 8116 31328
rect 7147 31297 7159 31300
rect 7101 31291 7159 31297
rect 8110 31288 8116 31300
rect 8168 31288 8174 31340
rect 9214 31288 9220 31340
rect 9272 31328 9278 31340
rect 9309 31331 9367 31337
rect 9309 31328 9321 31331
rect 9272 31300 9321 31328
rect 9272 31288 9278 31300
rect 9309 31297 9321 31300
rect 9355 31297 9367 31331
rect 9309 31291 9367 31297
rect 11146 31288 11152 31340
rect 11204 31288 11210 31340
rect 11514 31288 11520 31340
rect 11572 31328 11578 31340
rect 12066 31337 12072 31340
rect 11701 31331 11759 31337
rect 11701 31328 11713 31331
rect 11572 31300 11713 31328
rect 11572 31288 11578 31300
rect 11701 31297 11713 31300
rect 11747 31297 11759 31331
rect 11701 31291 11759 31297
rect 12023 31331 12072 31337
rect 12023 31297 12035 31331
rect 12069 31297 12072 31331
rect 12023 31291 12072 31297
rect 12038 31290 12072 31291
rect 12066 31288 12072 31290
rect 12124 31288 12130 31340
rect 12360 31337 12388 31368
rect 12544 31340 12572 31436
rect 12618 31424 12624 31436
rect 12676 31464 12682 31476
rect 13538 31464 13544 31476
rect 12676 31436 13544 31464
rect 12676 31424 12682 31436
rect 13538 31424 13544 31436
rect 13596 31424 13602 31476
rect 13633 31467 13691 31473
rect 13633 31433 13645 31467
rect 13679 31464 13691 31467
rect 14274 31464 14280 31476
rect 13679 31436 14280 31464
rect 13679 31433 13691 31436
rect 13633 31427 13691 31433
rect 14274 31424 14280 31436
rect 14332 31464 14338 31476
rect 15013 31467 15071 31473
rect 15013 31464 15025 31467
rect 14332 31436 15025 31464
rect 14332 31424 14338 31436
rect 15013 31433 15025 31436
rect 15059 31433 15071 31467
rect 15013 31427 15071 31433
rect 15562 31424 15568 31476
rect 15620 31424 15626 31476
rect 15749 31467 15807 31473
rect 15749 31433 15761 31467
rect 15795 31464 15807 31467
rect 16390 31464 16396 31476
rect 15795 31436 16396 31464
rect 15795 31433 15807 31436
rect 15749 31427 15807 31433
rect 13648 31368 14044 31396
rect 13648 31340 13676 31368
rect 12345 31331 12403 31337
rect 12345 31297 12357 31331
rect 12391 31297 12403 31331
rect 12345 31291 12403 31297
rect 12526 31288 12532 31340
rect 12584 31288 12590 31340
rect 12621 31331 12679 31337
rect 12621 31297 12633 31331
rect 12667 31297 12679 31331
rect 12621 31291 12679 31297
rect 12713 31331 12771 31337
rect 12713 31297 12725 31331
rect 12759 31328 12771 31331
rect 12802 31328 12808 31340
rect 12759 31300 12808 31328
rect 12759 31297 12771 31300
rect 12713 31291 12771 31297
rect 6914 31220 6920 31272
rect 6972 31260 6978 31272
rect 7193 31263 7251 31269
rect 7193 31260 7205 31263
rect 6972 31232 7205 31260
rect 6972 31220 6978 31232
rect 7193 31229 7205 31232
rect 7239 31260 7251 31263
rect 7374 31260 7380 31272
rect 7239 31232 7380 31260
rect 7239 31229 7251 31232
rect 7193 31223 7251 31229
rect 7374 31220 7380 31232
rect 7432 31220 7438 31272
rect 9582 31220 9588 31272
rect 9640 31220 9646 31272
rect 12161 31263 12219 31269
rect 12161 31260 12173 31263
rect 10704 31232 12173 31260
rect 6641 31195 6699 31201
rect 6641 31161 6653 31195
rect 6687 31161 6699 31195
rect 6641 31155 6699 31161
rect 1627 31096 3464 31124
rect 1627 31093 1639 31096
rect 1581 31087 1639 31093
rect 4062 31084 4068 31136
rect 4120 31084 4126 31136
rect 5077 31127 5135 31133
rect 5077 31093 5089 31127
rect 5123 31124 5135 31127
rect 5258 31124 5264 31136
rect 5123 31096 5264 31124
rect 5123 31093 5135 31096
rect 5077 31087 5135 31093
rect 5258 31084 5264 31096
rect 5316 31084 5322 31136
rect 9398 31084 9404 31136
rect 9456 31124 9462 31136
rect 10704 31124 10732 31232
rect 12161 31229 12173 31232
rect 12207 31260 12219 31263
rect 12636 31260 12664 31291
rect 12802 31288 12808 31300
rect 12860 31288 12866 31340
rect 13449 31331 13507 31337
rect 13449 31328 13461 31331
rect 12912 31300 13461 31328
rect 12207 31232 12664 31260
rect 12207 31229 12219 31232
rect 12161 31223 12219 31229
rect 12342 31152 12348 31204
rect 12400 31192 12406 31204
rect 12710 31192 12716 31204
rect 12400 31164 12716 31192
rect 12400 31152 12406 31164
rect 12710 31152 12716 31164
rect 12768 31152 12774 31204
rect 12912 31201 12940 31300
rect 13449 31297 13461 31300
rect 13495 31297 13507 31331
rect 13449 31291 13507 31297
rect 12897 31195 12955 31201
rect 12897 31161 12909 31195
rect 12943 31161 12955 31195
rect 12897 31155 12955 31161
rect 9456 31096 10732 31124
rect 9456 31084 9462 31096
rect 11054 31084 11060 31136
rect 11112 31084 11118 31136
rect 11514 31084 11520 31136
rect 11572 31084 11578 31136
rect 13464 31124 13492 31291
rect 13630 31288 13636 31340
rect 13688 31288 13694 31340
rect 13722 31288 13728 31340
rect 13780 31288 13786 31340
rect 13814 31288 13820 31340
rect 13872 31318 13878 31340
rect 14016 31337 14044 31368
rect 14090 31356 14096 31408
rect 14148 31356 14154 31408
rect 15381 31399 15439 31405
rect 15381 31396 15393 31399
rect 14476 31368 15393 31396
rect 13909 31331 13967 31337
rect 13909 31318 13921 31331
rect 13872 31297 13921 31318
rect 13955 31297 13967 31331
rect 13872 31291 13967 31297
rect 14001 31331 14059 31337
rect 14001 31297 14013 31331
rect 14047 31297 14059 31331
rect 14185 31331 14243 31337
rect 14185 31328 14197 31331
rect 14001 31291 14059 31297
rect 14108 31300 14197 31328
rect 13872 31290 13952 31291
rect 13872 31288 13878 31290
rect 13814 31152 13820 31204
rect 13872 31192 13878 31204
rect 13909 31195 13967 31201
rect 13909 31192 13921 31195
rect 13872 31164 13921 31192
rect 13872 31152 13878 31164
rect 13909 31161 13921 31164
rect 13955 31161 13967 31195
rect 13909 31155 13967 31161
rect 14108 31124 14136 31300
rect 14185 31297 14197 31300
rect 14231 31297 14243 31331
rect 14185 31291 14243 31297
rect 14324 31331 14382 31337
rect 14324 31297 14336 31331
rect 14370 31328 14382 31331
rect 14476 31328 14504 31368
rect 15381 31365 15393 31368
rect 15427 31365 15439 31399
rect 15580 31396 15608 31424
rect 15381 31359 15439 31365
rect 15488 31368 15608 31396
rect 14370 31300 14504 31328
rect 14370 31297 14382 31300
rect 14324 31291 14382 31297
rect 14550 31288 14556 31340
rect 14608 31288 14614 31340
rect 14662 31334 14720 31337
rect 14660 31331 14780 31334
rect 14660 31300 14674 31331
rect 14662 31297 14674 31300
rect 14708 31306 14780 31331
rect 14708 31297 14720 31306
rect 14662 31291 14720 31297
rect 14752 31260 14780 31306
rect 14826 31288 14832 31340
rect 14884 31328 14890 31340
rect 14921 31331 14979 31337
rect 14921 31328 14933 31331
rect 14884 31300 14933 31328
rect 14884 31288 14890 31300
rect 14921 31297 14933 31300
rect 14967 31297 14979 31331
rect 14921 31291 14979 31297
rect 15010 31288 15016 31340
rect 15068 31328 15074 31340
rect 15488 31337 15516 31368
rect 15200 31331 15258 31337
rect 15068 31300 15167 31328
rect 15068 31288 15074 31300
rect 15139 31269 15167 31300
rect 15200 31297 15212 31331
rect 15246 31297 15258 31331
rect 15200 31291 15258 31297
rect 15473 31331 15531 31337
rect 15473 31297 15485 31331
rect 15519 31297 15531 31331
rect 15473 31291 15531 31297
rect 15565 31331 15623 31337
rect 15565 31297 15577 31331
rect 15611 31297 15623 31331
rect 15565 31291 15623 31297
rect 15124 31263 15182 31269
rect 14752 31232 14964 31260
rect 14826 31152 14832 31204
rect 14884 31152 14890 31204
rect 14369 31127 14427 31133
rect 14369 31124 14381 31127
rect 13464 31096 14381 31124
rect 14369 31093 14381 31096
rect 14415 31093 14427 31127
rect 14936 31124 14964 31232
rect 15124 31229 15136 31263
rect 15170 31229 15182 31263
rect 15124 31223 15182 31229
rect 15215 31192 15243 31291
rect 15580 31260 15608 31291
rect 15838 31288 15844 31340
rect 15896 31328 15902 31340
rect 16224 31337 16252 31436
rect 16390 31424 16396 31436
rect 16448 31424 16454 31476
rect 17972 31436 18736 31464
rect 16117 31331 16175 31337
rect 16117 31328 16129 31331
rect 15896 31300 16129 31328
rect 15896 31288 15902 31300
rect 16117 31297 16129 31300
rect 16163 31297 16175 31331
rect 16117 31291 16175 31297
rect 16209 31331 16267 31337
rect 16209 31297 16221 31331
rect 16255 31297 16267 31331
rect 16209 31291 16267 31297
rect 16393 31331 16451 31337
rect 16393 31297 16405 31331
rect 16439 31328 16451 31331
rect 16574 31328 16580 31340
rect 16439 31300 16580 31328
rect 16439 31297 16451 31300
rect 16393 31291 16451 31297
rect 16574 31288 16580 31300
rect 16632 31288 16638 31340
rect 16666 31288 16672 31340
rect 16724 31328 16730 31340
rect 16761 31331 16819 31337
rect 16761 31328 16773 31331
rect 16724 31300 16773 31328
rect 16724 31288 16730 31300
rect 16761 31297 16773 31300
rect 16807 31297 16819 31331
rect 16761 31291 16819 31297
rect 17034 31288 17040 31340
rect 17092 31288 17098 31340
rect 17972 31337 18000 31436
rect 18138 31356 18144 31408
rect 18196 31356 18202 31408
rect 18598 31356 18604 31408
rect 18656 31356 18662 31408
rect 18708 31396 18736 31436
rect 19058 31424 19064 31476
rect 19116 31424 19122 31476
rect 19334 31424 19340 31476
rect 19392 31464 19398 31476
rect 19981 31467 20039 31473
rect 19981 31464 19993 31467
rect 19392 31436 19993 31464
rect 19392 31424 19398 31436
rect 19981 31433 19993 31436
rect 20027 31464 20039 31467
rect 20622 31464 20628 31476
rect 20027 31436 20628 31464
rect 20027 31433 20039 31436
rect 19981 31427 20039 31433
rect 20622 31424 20628 31436
rect 20680 31424 20686 31476
rect 21545 31467 21603 31473
rect 21545 31433 21557 31467
rect 21591 31464 21603 31467
rect 22462 31464 22468 31476
rect 21591 31436 22468 31464
rect 21591 31433 21603 31436
rect 21545 31427 21603 31433
rect 19153 31399 19211 31405
rect 19153 31396 19165 31399
rect 18708 31368 19165 31396
rect 19153 31365 19165 31368
rect 19199 31365 19211 31399
rect 19153 31359 19211 31365
rect 20162 31356 20168 31408
rect 20220 31396 20226 31408
rect 21361 31399 21419 31405
rect 21361 31396 21373 31399
rect 20220 31368 21373 31396
rect 20220 31356 20226 31368
rect 21361 31365 21373 31368
rect 21407 31365 21419 31399
rect 21361 31359 21419 31365
rect 21652 31368 21956 31396
rect 17957 31331 18015 31337
rect 17957 31297 17969 31331
rect 18003 31297 18015 31331
rect 17957 31291 18015 31297
rect 16298 31260 16304 31272
rect 15396 31232 16304 31260
rect 15286 31192 15292 31204
rect 15215 31164 15292 31192
rect 15286 31152 15292 31164
rect 15344 31152 15350 31204
rect 15194 31124 15200 31136
rect 14936 31096 15200 31124
rect 14369 31087 14427 31093
rect 15194 31084 15200 31096
rect 15252 31124 15258 31136
rect 15396 31124 15424 31232
rect 16298 31220 16304 31232
rect 16356 31260 16362 31272
rect 16945 31263 17003 31269
rect 16945 31260 16957 31263
rect 16356 31232 16957 31260
rect 16356 31220 16362 31232
rect 16945 31229 16957 31232
rect 16991 31229 17003 31263
rect 16945 31223 17003 31229
rect 15565 31195 15623 31201
rect 15565 31161 15577 31195
rect 15611 31192 15623 31195
rect 16574 31192 16580 31204
rect 15611 31164 16580 31192
rect 15611 31161 15623 31164
rect 15565 31155 15623 31161
rect 16574 31152 16580 31164
rect 16632 31152 16638 31204
rect 16853 31195 16911 31201
rect 16853 31161 16865 31195
rect 16899 31161 16911 31195
rect 16853 31155 16911 31161
rect 15252 31096 15424 31124
rect 15252 31084 15258 31096
rect 15930 31084 15936 31136
rect 15988 31084 15994 31136
rect 16022 31084 16028 31136
rect 16080 31124 16086 31136
rect 16868 31124 16896 31155
rect 17972 31136 18000 31291
rect 18230 31288 18236 31340
rect 18288 31288 18294 31340
rect 18325 31331 18383 31337
rect 18325 31297 18337 31331
rect 18371 31328 18383 31331
rect 18616 31328 18644 31356
rect 18693 31331 18751 31337
rect 18693 31328 18705 31331
rect 18371 31300 18705 31328
rect 18371 31297 18383 31300
rect 18325 31291 18383 31297
rect 18693 31297 18705 31300
rect 18739 31297 18751 31331
rect 18693 31291 18751 31297
rect 18877 31331 18935 31337
rect 18877 31297 18889 31331
rect 18923 31297 18935 31331
rect 18877 31291 18935 31297
rect 18248 31260 18276 31288
rect 18598 31260 18604 31272
rect 18248 31232 18604 31260
rect 18598 31220 18604 31232
rect 18656 31220 18662 31272
rect 18509 31195 18567 31201
rect 18509 31161 18521 31195
rect 18555 31192 18567 31195
rect 18892 31192 18920 31291
rect 19058 31288 19064 31340
rect 19116 31328 19122 31340
rect 21652 31337 21680 31368
rect 19337 31331 19395 31337
rect 19337 31328 19349 31331
rect 19116 31300 19349 31328
rect 19116 31288 19122 31300
rect 19337 31297 19349 31300
rect 19383 31297 19395 31331
rect 19337 31291 19395 31297
rect 19521 31331 19579 31337
rect 19521 31297 19533 31331
rect 19567 31328 19579 31331
rect 19797 31331 19855 31337
rect 19797 31328 19809 31331
rect 19567 31300 19809 31328
rect 19567 31297 19579 31300
rect 19521 31291 19579 31297
rect 19797 31297 19809 31300
rect 19843 31297 19855 31331
rect 19797 31291 19855 31297
rect 21637 31331 21695 31337
rect 21637 31297 21649 31331
rect 21683 31297 21695 31331
rect 21637 31291 21695 31297
rect 21821 31331 21879 31337
rect 21821 31297 21833 31331
rect 21867 31297 21879 31331
rect 21928 31328 21956 31368
rect 22186 31337 22192 31340
rect 22152 31331 22192 31337
rect 22152 31328 22164 31331
rect 21928 31300 22164 31328
rect 21821 31291 21879 31297
rect 22152 31297 22164 31300
rect 22152 31291 22192 31297
rect 19613 31263 19671 31269
rect 19613 31260 19625 31263
rect 19168 31232 19625 31260
rect 19168 31204 19196 31232
rect 19613 31229 19625 31232
rect 19659 31229 19671 31263
rect 19613 31223 19671 31229
rect 18555 31164 18920 31192
rect 18555 31161 18567 31164
rect 18509 31155 18567 31161
rect 19150 31152 19156 31204
rect 19208 31152 19214 31204
rect 21361 31195 21419 31201
rect 21361 31161 21373 31195
rect 21407 31192 21419 31195
rect 21836 31192 21864 31291
rect 22186 31288 22192 31291
rect 22244 31288 22250 31340
rect 22388 31337 22416 31436
rect 22462 31424 22468 31436
rect 22520 31424 22526 31476
rect 24305 31467 24363 31473
rect 24305 31433 24317 31467
rect 24351 31464 24363 31467
rect 24394 31464 24400 31476
rect 24351 31436 24400 31464
rect 24351 31433 24363 31436
rect 24305 31427 24363 31433
rect 24394 31424 24400 31436
rect 24452 31424 24458 31476
rect 26326 31424 26332 31476
rect 26384 31424 26390 31476
rect 27614 31424 27620 31476
rect 27672 31464 27678 31476
rect 27709 31467 27767 31473
rect 27709 31464 27721 31467
rect 27672 31436 27721 31464
rect 27672 31424 27678 31436
rect 27709 31433 27721 31436
rect 27755 31433 27767 31467
rect 27709 31427 27767 31433
rect 29089 31467 29147 31473
rect 29089 31433 29101 31467
rect 29135 31464 29147 31467
rect 30098 31464 30104 31476
rect 29135 31436 30104 31464
rect 29135 31433 29147 31436
rect 29089 31427 29147 31433
rect 30098 31424 30104 31436
rect 30156 31424 30162 31476
rect 31481 31467 31539 31473
rect 31481 31433 31493 31467
rect 31527 31464 31539 31467
rect 31527 31436 31754 31464
rect 31527 31433 31539 31436
rect 31481 31427 31539 31433
rect 25038 31356 25044 31408
rect 25096 31396 25102 31408
rect 25590 31396 25596 31408
rect 25096 31368 25596 31396
rect 25096 31356 25102 31368
rect 22373 31331 22431 31337
rect 22373 31297 22385 31331
rect 22419 31297 22431 31331
rect 22373 31291 22431 31297
rect 24118 31288 24124 31340
rect 24176 31288 24182 31340
rect 24305 31331 24363 31337
rect 24305 31297 24317 31331
rect 24351 31328 24363 31331
rect 24486 31328 24492 31340
rect 24351 31300 24492 31328
rect 24351 31297 24363 31300
rect 24305 31291 24363 31297
rect 24486 31288 24492 31300
rect 24544 31288 24550 31340
rect 24946 31288 24952 31340
rect 25004 31288 25010 31340
rect 25130 31288 25136 31340
rect 25188 31288 25194 31340
rect 25240 31337 25268 31368
rect 25590 31356 25596 31368
rect 25648 31356 25654 31408
rect 25225 31331 25283 31337
rect 25225 31297 25237 31331
rect 25271 31297 25283 31331
rect 25225 31291 25283 31297
rect 25317 31331 25375 31337
rect 25317 31297 25329 31331
rect 25363 31328 25375 31331
rect 26344 31328 26372 31424
rect 27341 31399 27399 31405
rect 27341 31365 27353 31399
rect 27387 31396 27399 31399
rect 31726 31396 31754 31436
rect 32306 31424 32312 31476
rect 32364 31464 32370 31476
rect 32861 31467 32919 31473
rect 32364 31436 32720 31464
rect 32364 31424 32370 31436
rect 27387 31368 28948 31396
rect 27387 31365 27399 31368
rect 27341 31359 27399 31365
rect 25363 31300 26372 31328
rect 25363 31297 25375 31300
rect 25317 31291 25375 31297
rect 21407 31164 21864 31192
rect 21407 31161 21419 31164
rect 21361 31155 21419 31161
rect 21910 31152 21916 31204
rect 21968 31152 21974 31204
rect 16080 31096 16896 31124
rect 16080 31084 16086 31096
rect 17218 31084 17224 31136
rect 17276 31084 17282 31136
rect 17954 31084 17960 31136
rect 18012 31084 18018 31136
rect 18598 31084 18604 31136
rect 18656 31124 18662 31136
rect 19168 31124 19196 31152
rect 18656 31096 19196 31124
rect 18656 31084 18662 31096
rect 21818 31084 21824 31136
rect 21876 31124 21882 31136
rect 25332 31124 25360 31291
rect 27154 31288 27160 31340
rect 27212 31288 27218 31340
rect 28000 31337 28028 31368
rect 28920 31340 28948 31368
rect 29840 31368 30236 31396
rect 31726 31368 32352 31396
rect 27985 31331 28043 31337
rect 27985 31297 27997 31331
rect 28031 31297 28043 31331
rect 27985 31291 28043 31297
rect 28350 31288 28356 31340
rect 28408 31288 28414 31340
rect 28534 31288 28540 31340
rect 28592 31288 28598 31340
rect 28902 31288 28908 31340
rect 28960 31288 28966 31340
rect 29840 31337 29868 31368
rect 30208 31340 30236 31368
rect 29825 31331 29883 31337
rect 29825 31297 29837 31331
rect 29871 31297 29883 31331
rect 29825 31291 29883 31297
rect 29914 31288 29920 31340
rect 29972 31288 29978 31340
rect 30006 31288 30012 31340
rect 30064 31328 30070 31340
rect 30101 31331 30159 31337
rect 30101 31328 30113 31331
rect 30064 31300 30113 31328
rect 30064 31288 30070 31300
rect 30101 31297 30113 31300
rect 30147 31297 30159 31331
rect 30101 31291 30159 31297
rect 30190 31288 30196 31340
rect 30248 31328 30254 31340
rect 30377 31331 30435 31337
rect 30377 31328 30389 31331
rect 30248 31300 30389 31328
rect 30248 31288 30254 31300
rect 30377 31297 30389 31300
rect 30423 31297 30435 31331
rect 30377 31291 30435 31297
rect 30653 31331 30711 31337
rect 30653 31297 30665 31331
rect 30699 31297 30711 31331
rect 30653 31291 30711 31297
rect 30837 31331 30895 31337
rect 30837 31297 30849 31331
rect 30883 31328 30895 31331
rect 31113 31331 31171 31337
rect 31113 31328 31125 31331
rect 30883 31300 31125 31328
rect 30883 31297 30895 31300
rect 30837 31291 30895 31297
rect 31113 31297 31125 31300
rect 31159 31328 31171 31331
rect 31478 31328 31484 31340
rect 31159 31300 31484 31328
rect 31159 31297 31171 31300
rect 31113 31291 31171 31297
rect 26970 31220 26976 31272
rect 27028 31220 27034 31272
rect 27246 31220 27252 31272
rect 27304 31260 27310 31272
rect 27709 31263 27767 31269
rect 27709 31260 27721 31263
rect 27304 31232 27721 31260
rect 27304 31220 27310 31232
rect 27709 31229 27721 31232
rect 27755 31229 27767 31263
rect 27709 31223 27767 31229
rect 28442 31220 28448 31272
rect 28500 31260 28506 31272
rect 28629 31263 28687 31269
rect 28629 31260 28641 31263
rect 28500 31232 28641 31260
rect 28500 31220 28506 31232
rect 28629 31229 28641 31232
rect 28675 31229 28687 31263
rect 28629 31223 28687 31229
rect 28721 31263 28779 31269
rect 28721 31229 28733 31263
rect 28767 31260 28779 31263
rect 30668 31260 30696 31291
rect 31478 31288 31484 31300
rect 31536 31288 31542 31340
rect 32324 31337 32352 31368
rect 32692 31337 32720 31436
rect 32861 31433 32873 31467
rect 32907 31464 32919 31467
rect 33410 31464 33416 31476
rect 32907 31436 33416 31464
rect 32907 31433 32919 31436
rect 32861 31427 32919 31433
rect 33410 31424 33416 31436
rect 33468 31424 33474 31476
rect 33965 31467 34023 31473
rect 33965 31433 33977 31467
rect 34011 31464 34023 31467
rect 34011 31436 34560 31464
rect 34011 31433 34023 31436
rect 33965 31427 34023 31433
rect 33042 31356 33048 31408
rect 33100 31396 33106 31408
rect 34057 31399 34115 31405
rect 33100 31368 33732 31396
rect 33100 31356 33106 31368
rect 32125 31331 32183 31337
rect 32125 31328 32137 31331
rect 31726 31300 32137 31328
rect 31018 31260 31024 31272
rect 28767 31232 30328 31260
rect 30668 31232 31024 31260
rect 28767 31229 28779 31232
rect 28721 31223 28779 31229
rect 27893 31195 27951 31201
rect 27893 31161 27905 31195
rect 27939 31192 27951 31195
rect 29086 31192 29092 31204
rect 27939 31164 29092 31192
rect 27939 31161 27951 31164
rect 27893 31155 27951 31161
rect 29086 31152 29092 31164
rect 29144 31152 29150 31204
rect 21876 31096 25360 31124
rect 25593 31127 25651 31133
rect 21876 31084 21882 31096
rect 25593 31093 25605 31127
rect 25639 31124 25651 31127
rect 28626 31124 28632 31136
rect 25639 31096 28632 31124
rect 25639 31093 25651 31096
rect 25593 31087 25651 31093
rect 28626 31084 28632 31096
rect 28684 31084 28690 31136
rect 28718 31084 28724 31136
rect 28776 31124 28782 31136
rect 30193 31127 30251 31133
rect 30193 31124 30205 31127
rect 28776 31096 30205 31124
rect 28776 31084 28782 31096
rect 30193 31093 30205 31096
rect 30239 31093 30251 31127
rect 30300 31124 30328 31232
rect 31018 31220 31024 31232
rect 31076 31220 31082 31272
rect 31294 31220 31300 31272
rect 31352 31260 31358 31272
rect 31726 31260 31754 31300
rect 32125 31297 32137 31300
rect 32171 31297 32183 31331
rect 32125 31291 32183 31297
rect 32309 31331 32367 31337
rect 32309 31297 32321 31331
rect 32355 31328 32367 31331
rect 32677 31331 32735 31337
rect 32355 31300 32628 31328
rect 32355 31297 32367 31300
rect 32309 31291 32367 31297
rect 31352 31232 31754 31260
rect 32401 31263 32459 31269
rect 31352 31220 31358 31232
rect 32401 31229 32413 31263
rect 32447 31229 32459 31263
rect 32401 31223 32459 31229
rect 30374 31152 30380 31204
rect 30432 31192 30438 31204
rect 32416 31192 32444 31223
rect 32490 31220 32496 31272
rect 32548 31220 32554 31272
rect 32600 31260 32628 31300
rect 32677 31297 32689 31331
rect 32723 31297 32735 31331
rect 32677 31291 32735 31297
rect 32858 31288 32864 31340
rect 32916 31328 32922 31340
rect 33229 31331 33287 31337
rect 33229 31328 33241 31331
rect 32916 31300 33241 31328
rect 32916 31288 32922 31300
rect 33229 31297 33241 31300
rect 33275 31297 33287 31331
rect 33229 31291 33287 31297
rect 33321 31331 33379 31337
rect 33321 31297 33333 31331
rect 33367 31297 33379 31331
rect 33321 31291 33379 31297
rect 33336 31260 33364 31291
rect 33410 31288 33416 31340
rect 33468 31288 33474 31340
rect 33594 31288 33600 31340
rect 33652 31288 33658 31340
rect 33704 31337 33732 31368
rect 34057 31365 34069 31399
rect 34103 31396 34115 31399
rect 34103 31368 34376 31396
rect 34103 31365 34115 31368
rect 34057 31359 34115 31365
rect 34348 31340 34376 31368
rect 33689 31331 33747 31337
rect 33689 31297 33701 31331
rect 33735 31297 33747 31331
rect 33689 31291 33747 31297
rect 32600 31232 33364 31260
rect 33704 31260 33732 31291
rect 34146 31288 34152 31340
rect 34204 31288 34210 31340
rect 34330 31288 34336 31340
rect 34388 31288 34394 31340
rect 34532 31337 34560 31436
rect 35434 31424 35440 31476
rect 35492 31424 35498 31476
rect 35897 31467 35955 31473
rect 35897 31433 35909 31467
rect 35943 31464 35955 31467
rect 35986 31464 35992 31476
rect 35943 31436 35992 31464
rect 35943 31433 35955 31436
rect 35897 31427 35955 31433
rect 35986 31424 35992 31436
rect 36044 31424 36050 31476
rect 35342 31396 35348 31408
rect 34716 31368 35348 31396
rect 34517 31331 34575 31337
rect 34517 31297 34529 31331
rect 34563 31297 34575 31331
rect 34517 31291 34575 31297
rect 34606 31288 34612 31340
rect 34664 31288 34670 31340
rect 34716 31260 34744 31368
rect 35342 31356 35348 31368
rect 35400 31356 35406 31408
rect 35452 31396 35480 31424
rect 36449 31399 36507 31405
rect 36449 31396 36461 31399
rect 35452 31368 36461 31396
rect 34790 31288 34796 31340
rect 34848 31288 34854 31340
rect 34885 31331 34943 31337
rect 34885 31297 34897 31331
rect 34931 31328 34943 31331
rect 34931 31300 35204 31328
rect 34931 31297 34943 31300
rect 34885 31291 34943 31297
rect 35176 31269 35204 31300
rect 35434 31288 35440 31340
rect 35492 31288 35498 31340
rect 35636 31337 35664 31368
rect 36449 31365 36461 31368
rect 36495 31365 36507 31399
rect 36449 31359 36507 31365
rect 35529 31331 35587 31337
rect 35529 31297 35541 31331
rect 35575 31297 35587 31331
rect 35529 31291 35587 31297
rect 35621 31331 35679 31337
rect 35621 31297 35633 31331
rect 35667 31297 35679 31331
rect 35621 31291 35679 31297
rect 33704 31232 34744 31260
rect 35161 31263 35219 31269
rect 35161 31229 35173 31263
rect 35207 31229 35219 31263
rect 35544 31260 35572 31291
rect 35710 31288 35716 31340
rect 35768 31328 35774 31340
rect 35805 31331 35863 31337
rect 35805 31328 35817 31331
rect 35768 31300 35817 31328
rect 35768 31288 35774 31300
rect 35805 31297 35817 31300
rect 35851 31297 35863 31331
rect 35805 31291 35863 31297
rect 36078 31288 36084 31340
rect 36136 31288 36142 31340
rect 36262 31288 36268 31340
rect 36320 31288 36326 31340
rect 36354 31288 36360 31340
rect 36412 31288 36418 31340
rect 36538 31288 36544 31340
rect 36596 31288 36602 31340
rect 36556 31260 36584 31288
rect 35544 31232 36584 31260
rect 35161 31223 35219 31229
rect 30432 31164 34008 31192
rect 30432 31152 30438 31164
rect 33980 31136 34008 31164
rect 34238 31152 34244 31204
rect 34296 31192 34302 31204
rect 34333 31195 34391 31201
rect 34333 31192 34345 31195
rect 34296 31164 34345 31192
rect 34296 31152 34302 31164
rect 34333 31161 34345 31164
rect 34379 31161 34391 31195
rect 34333 31155 34391 31161
rect 32490 31124 32496 31136
rect 30300 31096 32496 31124
rect 30193 31087 30251 31093
rect 32490 31084 32496 31096
rect 32548 31084 32554 31136
rect 32950 31084 32956 31136
rect 33008 31084 33014 31136
rect 33962 31084 33968 31136
rect 34020 31084 34026 31136
rect 1104 31034 38272 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38272 31034
rect 1104 30960 38272 30982
rect 3050 30880 3056 30932
rect 3108 30920 3114 30932
rect 3145 30923 3203 30929
rect 3145 30920 3157 30923
rect 3108 30892 3157 30920
rect 3108 30880 3114 30892
rect 3145 30889 3157 30892
rect 3191 30889 3203 30923
rect 4062 30920 4068 30932
rect 3145 30883 3203 30889
rect 3528 30892 4068 30920
rect 3326 30676 3332 30728
rect 3384 30676 3390 30728
rect 3528 30725 3556 30892
rect 4062 30880 4068 30892
rect 4120 30880 4126 30932
rect 4433 30923 4491 30929
rect 4433 30889 4445 30923
rect 4479 30920 4491 30923
rect 4614 30920 4620 30932
rect 4479 30892 4620 30920
rect 4479 30889 4491 30892
rect 4433 30883 4491 30889
rect 4614 30880 4620 30892
rect 4672 30880 4678 30932
rect 5074 30880 5080 30932
rect 5132 30880 5138 30932
rect 9582 30880 9588 30932
rect 9640 30920 9646 30932
rect 9769 30923 9827 30929
rect 9769 30920 9781 30923
rect 9640 30892 9781 30920
rect 9640 30880 9646 30892
rect 9769 30889 9781 30892
rect 9815 30889 9827 30923
rect 11514 30920 11520 30932
rect 9769 30883 9827 30889
rect 10796 30892 11520 30920
rect 4522 30852 4528 30864
rect 3620 30824 4528 30852
rect 3620 30725 3648 30824
rect 4522 30812 4528 30824
rect 4580 30812 4586 30864
rect 5092 30784 5120 30880
rect 8680 30824 9536 30852
rect 4172 30756 5120 30784
rect 6825 30787 6883 30793
rect 3970 30725 3976 30728
rect 3513 30719 3571 30725
rect 3513 30685 3525 30719
rect 3559 30685 3571 30719
rect 3513 30679 3571 30685
rect 3605 30719 3663 30725
rect 3605 30685 3617 30719
rect 3651 30685 3663 30719
rect 3605 30679 3663 30685
rect 3789 30719 3847 30725
rect 3789 30685 3801 30719
rect 3835 30685 3847 30719
rect 3789 30679 3847 30685
rect 3937 30719 3976 30725
rect 3937 30685 3949 30719
rect 3937 30679 3976 30685
rect 3804 30580 3832 30679
rect 3970 30676 3976 30679
rect 4028 30676 4034 30728
rect 4062 30608 4068 30660
rect 4120 30608 4126 30660
rect 4172 30657 4200 30756
rect 4338 30725 4344 30728
rect 4295 30719 4344 30725
rect 4295 30685 4307 30719
rect 4341 30685 4344 30719
rect 4295 30679 4344 30685
rect 4338 30676 4344 30679
rect 4396 30676 4402 30728
rect 4157 30651 4215 30657
rect 4157 30617 4169 30651
rect 4203 30617 4215 30651
rect 4632 30648 4660 30756
rect 6825 30753 6837 30787
rect 6871 30784 6883 30787
rect 7006 30784 7012 30796
rect 6871 30756 7012 30784
rect 6871 30753 6883 30756
rect 6825 30747 6883 30753
rect 7006 30744 7012 30756
rect 7064 30744 7070 30796
rect 7374 30744 7380 30796
rect 7432 30784 7438 30796
rect 8680 30784 8708 30824
rect 7432 30756 8708 30784
rect 8757 30787 8815 30793
rect 7432 30744 7438 30756
rect 8757 30753 8769 30787
rect 8803 30784 8815 30787
rect 9398 30784 9404 30796
rect 8803 30756 9404 30784
rect 8803 30753 8815 30756
rect 8757 30747 8815 30753
rect 9398 30744 9404 30756
rect 9456 30744 9462 30796
rect 9508 30793 9536 30824
rect 10796 30793 10824 30892
rect 11514 30880 11520 30892
rect 11572 30880 11578 30932
rect 11609 30923 11667 30929
rect 11609 30889 11621 30923
rect 11655 30920 11667 30923
rect 11790 30920 11796 30932
rect 11655 30892 11796 30920
rect 11655 30889 11667 30892
rect 11609 30883 11667 30889
rect 11146 30812 11152 30864
rect 11204 30852 11210 30864
rect 11425 30855 11483 30861
rect 11425 30852 11437 30855
rect 11204 30824 11437 30852
rect 11204 30812 11210 30824
rect 11425 30821 11437 30824
rect 11471 30821 11483 30855
rect 11624 30852 11652 30883
rect 11790 30880 11796 30892
rect 11848 30920 11854 30932
rect 11848 30892 13308 30920
rect 11848 30880 11854 30892
rect 11425 30815 11483 30821
rect 11532 30824 11652 30852
rect 9493 30787 9551 30793
rect 9493 30753 9505 30787
rect 9539 30753 9551 30787
rect 9493 30747 9551 30753
rect 10781 30787 10839 30793
rect 10781 30753 10793 30787
rect 10827 30753 10839 30787
rect 10781 30747 10839 30753
rect 10870 30744 10876 30796
rect 10928 30744 10934 30796
rect 11532 30784 11560 30824
rect 12526 30812 12532 30864
rect 12584 30812 12590 30864
rect 13170 30852 13176 30864
rect 13096 30824 13176 30852
rect 11072 30756 11560 30784
rect 11072 30728 11100 30756
rect 4798 30676 4804 30728
rect 4856 30716 4862 30728
rect 4893 30719 4951 30725
rect 4893 30716 4905 30719
rect 4856 30688 4905 30716
rect 4856 30676 4862 30688
rect 4893 30685 4905 30688
rect 4939 30685 4951 30719
rect 8662 30716 8668 30728
rect 8418 30688 8668 30716
rect 4893 30679 4951 30685
rect 8662 30676 8668 30688
rect 8720 30676 8726 30728
rect 9953 30719 10011 30725
rect 9953 30685 9965 30719
rect 9999 30716 10011 30719
rect 10689 30719 10747 30725
rect 9999 30688 10364 30716
rect 9999 30685 10011 30688
rect 9953 30679 10011 30685
rect 4706 30648 4712 30660
rect 4632 30620 4712 30648
rect 4157 30611 4215 30617
rect 4706 30608 4712 30620
rect 4764 30608 4770 30660
rect 4982 30608 4988 30660
rect 5040 30648 5046 30660
rect 5040 30620 5382 30648
rect 5040 30608 5046 30620
rect 6546 30608 6552 30660
rect 6604 30608 6610 30660
rect 7282 30608 7288 30660
rect 7340 30608 7346 30660
rect 4430 30580 4436 30592
rect 3804 30552 4436 30580
rect 4430 30540 4436 30552
rect 4488 30540 4494 30592
rect 8938 30540 8944 30592
rect 8996 30540 9002 30592
rect 9306 30540 9312 30592
rect 9364 30540 9370 30592
rect 10336 30589 10364 30688
rect 10689 30685 10701 30719
rect 10735 30716 10747 30719
rect 11054 30716 11060 30728
rect 10735 30688 11060 30716
rect 10735 30685 10747 30688
rect 10689 30679 10747 30685
rect 11054 30676 11060 30688
rect 11112 30676 11118 30728
rect 12437 30719 12495 30725
rect 12437 30685 12449 30719
rect 12483 30685 12495 30719
rect 12544 30716 12572 30812
rect 12621 30719 12679 30725
rect 12621 30716 12633 30719
rect 12544 30688 12633 30716
rect 12437 30679 12495 30685
rect 12621 30685 12633 30688
rect 12667 30685 12679 30719
rect 12621 30679 12679 30685
rect 11577 30651 11635 30657
rect 11577 30617 11589 30651
rect 11623 30648 11635 30651
rect 11698 30648 11704 30660
rect 11623 30620 11704 30648
rect 11623 30617 11635 30620
rect 11577 30611 11635 30617
rect 11698 30608 11704 30620
rect 11756 30608 11762 30660
rect 11793 30651 11851 30657
rect 11793 30617 11805 30651
rect 11839 30648 11851 30651
rect 11974 30648 11980 30660
rect 11839 30620 11980 30648
rect 11839 30617 11851 30620
rect 11793 30611 11851 30617
rect 11974 30608 11980 30620
rect 12032 30608 12038 30660
rect 12452 30648 12480 30679
rect 12710 30676 12716 30728
rect 12768 30676 12774 30728
rect 12802 30676 12808 30728
rect 12860 30676 12866 30728
rect 12526 30648 12532 30660
rect 12452 30620 12532 30648
rect 12526 30608 12532 30620
rect 12584 30608 12590 30660
rect 12820 30648 12848 30676
rect 13096 30657 13124 30824
rect 13170 30812 13176 30824
rect 13228 30812 13234 30864
rect 13280 30725 13308 30892
rect 13722 30880 13728 30932
rect 13780 30920 13786 30932
rect 14185 30923 14243 30929
rect 14185 30920 14197 30923
rect 13780 30892 14197 30920
rect 13780 30880 13786 30892
rect 14185 30889 14197 30892
rect 14231 30889 14243 30923
rect 14185 30883 14243 30889
rect 14274 30880 14280 30932
rect 14332 30880 14338 30932
rect 15930 30880 15936 30932
rect 15988 30880 15994 30932
rect 16206 30880 16212 30932
rect 16264 30920 16270 30932
rect 16264 30892 16896 30920
rect 16264 30880 16270 30892
rect 14292 30725 14320 30880
rect 15948 30852 15976 30880
rect 16868 30861 16896 30892
rect 18598 30880 18604 30932
rect 18656 30880 18662 30932
rect 19429 30923 19487 30929
rect 19429 30889 19441 30923
rect 19475 30920 19487 30923
rect 20070 30920 20076 30932
rect 19475 30892 20076 30920
rect 19475 30889 19487 30892
rect 19429 30883 19487 30889
rect 20070 30880 20076 30892
rect 20128 30880 20134 30932
rect 25593 30923 25651 30929
rect 25593 30889 25605 30923
rect 25639 30920 25651 30923
rect 26970 30920 26976 30932
rect 25639 30892 26976 30920
rect 25639 30889 25651 30892
rect 25593 30883 25651 30889
rect 26970 30880 26976 30892
rect 27028 30880 27034 30932
rect 32950 30880 32956 30932
rect 33008 30880 33014 30932
rect 34606 30880 34612 30932
rect 34664 30920 34670 30932
rect 34701 30923 34759 30929
rect 34701 30920 34713 30923
rect 34664 30892 34713 30920
rect 34664 30880 34670 30892
rect 34701 30889 34713 30892
rect 34747 30889 34759 30923
rect 34701 30883 34759 30889
rect 36173 30923 36231 30929
rect 36173 30889 36185 30923
rect 36219 30920 36231 30923
rect 36354 30920 36360 30932
rect 36219 30892 36360 30920
rect 36219 30889 36231 30892
rect 36173 30883 36231 30889
rect 36354 30880 36360 30892
rect 36412 30880 36418 30932
rect 16853 30855 16911 30861
rect 15948 30824 16804 30852
rect 15010 30744 15016 30796
rect 15068 30744 15074 30796
rect 15930 30744 15936 30796
rect 15988 30744 15994 30796
rect 16022 30744 16028 30796
rect 16080 30744 16086 30796
rect 16114 30744 16120 30796
rect 16172 30744 16178 30796
rect 16298 30744 16304 30796
rect 16356 30744 16362 30796
rect 13254 30719 13312 30725
rect 13254 30685 13266 30719
rect 13300 30685 13312 30719
rect 13254 30679 13312 30685
rect 14277 30719 14335 30725
rect 14277 30685 14289 30719
rect 14323 30685 14335 30719
rect 15028 30716 15056 30744
rect 16040 30716 16068 30744
rect 16209 30719 16267 30725
rect 16209 30716 16221 30719
rect 15028 30688 15976 30716
rect 16040 30688 16221 30716
rect 14277 30679 14335 30685
rect 12728 30620 12848 30648
rect 13081 30651 13139 30657
rect 12728 30592 12756 30620
rect 13081 30617 13093 30651
rect 13127 30617 13139 30651
rect 15948 30648 15976 30688
rect 16209 30685 16221 30688
rect 16255 30685 16267 30719
rect 16209 30679 16267 30685
rect 16393 30719 16451 30725
rect 16393 30685 16405 30719
rect 16439 30685 16451 30719
rect 16393 30679 16451 30685
rect 16408 30648 16436 30679
rect 16574 30676 16580 30728
rect 16632 30676 16638 30728
rect 16776 30725 16804 30824
rect 16853 30821 16865 30855
rect 16899 30821 16911 30855
rect 16853 30815 16911 30821
rect 17586 30812 17592 30864
rect 17644 30852 17650 30864
rect 25222 30852 25228 30864
rect 17644 30824 25228 30852
rect 17644 30812 17650 30824
rect 25222 30812 25228 30824
rect 25280 30812 25286 30864
rect 25682 30812 25688 30864
rect 25740 30852 25746 30864
rect 32493 30855 32551 30861
rect 25740 30824 27016 30852
rect 25740 30812 25746 30824
rect 19058 30784 19064 30796
rect 18248 30756 19064 30784
rect 18248 30728 18276 30756
rect 16761 30719 16819 30725
rect 16761 30685 16773 30719
rect 16807 30685 16819 30719
rect 16761 30679 16819 30685
rect 18230 30676 18236 30728
rect 18288 30676 18294 30728
rect 18708 30725 18736 30756
rect 19058 30744 19064 30756
rect 19116 30744 19122 30796
rect 20070 30744 20076 30796
rect 20128 30784 20134 30796
rect 22370 30784 22376 30796
rect 20128 30756 22376 30784
rect 20128 30744 20134 30756
rect 22370 30744 22376 30756
rect 22428 30744 22434 30796
rect 18509 30719 18567 30725
rect 18509 30685 18521 30719
rect 18555 30685 18567 30719
rect 18509 30679 18567 30685
rect 18693 30719 18751 30725
rect 18693 30685 18705 30719
rect 18739 30716 18751 30719
rect 18877 30719 18935 30725
rect 18877 30716 18889 30719
rect 18739 30688 18889 30716
rect 18739 30685 18751 30688
rect 18693 30679 18751 30685
rect 18877 30685 18889 30688
rect 18923 30685 18935 30719
rect 18877 30679 18935 30685
rect 18969 30719 19027 30725
rect 18969 30685 18981 30719
rect 19015 30716 19027 30719
rect 19245 30719 19303 30725
rect 19245 30716 19257 30719
rect 19015 30688 19257 30716
rect 19015 30685 19027 30688
rect 18969 30679 19027 30685
rect 19245 30685 19257 30688
rect 19291 30685 19303 30719
rect 19245 30679 19303 30685
rect 19429 30719 19487 30725
rect 19429 30685 19441 30719
rect 19475 30685 19487 30719
rect 19429 30679 19487 30685
rect 25225 30719 25283 30725
rect 25225 30685 25237 30719
rect 25271 30716 25283 30719
rect 25700 30716 25728 30812
rect 25271 30688 25728 30716
rect 26237 30719 26295 30725
rect 25271 30685 25283 30688
rect 25225 30679 25283 30685
rect 26237 30685 26249 30719
rect 26283 30685 26295 30719
rect 26237 30679 26295 30685
rect 26789 30719 26847 30725
rect 26789 30685 26801 30719
rect 26835 30716 26847 30719
rect 26988 30716 27016 30824
rect 32493 30821 32505 30855
rect 32539 30852 32551 30855
rect 32539 30824 32812 30852
rect 32539 30821 32551 30824
rect 32493 30815 32551 30821
rect 32784 30796 32812 30824
rect 28166 30784 28172 30796
rect 27908 30756 28172 30784
rect 26835 30688 27016 30716
rect 26835 30685 26847 30688
rect 26789 30679 26847 30685
rect 17954 30648 17960 30660
rect 13081 30611 13139 30617
rect 13372 30620 15148 30648
rect 15948 30620 16436 30648
rect 16592 30620 17960 30648
rect 10321 30583 10379 30589
rect 10321 30549 10333 30583
rect 10367 30549 10379 30583
rect 10321 30543 10379 30549
rect 12710 30540 12716 30592
rect 12768 30540 12774 30592
rect 12989 30583 13047 30589
rect 12989 30549 13001 30583
rect 13035 30580 13047 30583
rect 13372 30580 13400 30620
rect 13035 30552 13400 30580
rect 13035 30549 13047 30552
rect 12989 30543 13047 30549
rect 13446 30540 13452 30592
rect 13504 30540 13510 30592
rect 15120 30580 15148 30620
rect 16592 30580 16620 30620
rect 17954 30608 17960 30620
rect 18012 30648 18018 30660
rect 18524 30648 18552 30679
rect 19444 30648 19472 30679
rect 18012 30620 19472 30648
rect 25409 30651 25467 30657
rect 18012 30608 18018 30620
rect 25409 30617 25421 30651
rect 25455 30648 25467 30651
rect 25774 30648 25780 30660
rect 25455 30620 25780 30648
rect 25455 30617 25467 30620
rect 25409 30611 25467 30617
rect 25774 30608 25780 30620
rect 25832 30648 25838 30660
rect 26252 30648 26280 30679
rect 25832 30620 26280 30648
rect 25832 30608 25838 30620
rect 26694 30608 26700 30660
rect 26752 30648 26758 30660
rect 26804 30648 26832 30679
rect 27706 30676 27712 30728
rect 27764 30676 27770 30728
rect 27908 30725 27936 30756
rect 28166 30744 28172 30756
rect 28224 30784 28230 30796
rect 28718 30784 28724 30796
rect 28224 30756 28724 30784
rect 28224 30744 28230 30756
rect 28718 30744 28724 30756
rect 28776 30744 28782 30796
rect 29273 30787 29331 30793
rect 29273 30784 29285 30787
rect 28828 30756 29285 30784
rect 28828 30728 28856 30756
rect 29273 30753 29285 30756
rect 29319 30753 29331 30787
rect 30374 30784 30380 30796
rect 29273 30747 29331 30753
rect 29564 30756 30380 30784
rect 27893 30719 27951 30725
rect 27893 30685 27905 30719
rect 27939 30685 27951 30719
rect 27893 30679 27951 30685
rect 27985 30719 28043 30725
rect 27985 30685 27997 30719
rect 28031 30716 28043 30719
rect 28258 30716 28264 30728
rect 28031 30688 28264 30716
rect 28031 30685 28043 30688
rect 27985 30679 28043 30685
rect 26752 30620 26832 30648
rect 27617 30651 27675 30657
rect 26752 30608 26758 30620
rect 27617 30617 27629 30651
rect 27663 30648 27675 30651
rect 28000 30648 28028 30679
rect 28258 30676 28264 30688
rect 28316 30716 28322 30728
rect 28537 30719 28595 30725
rect 28537 30716 28549 30719
rect 28316 30688 28549 30716
rect 28316 30676 28322 30688
rect 28537 30685 28549 30688
rect 28583 30685 28595 30719
rect 28537 30679 28595 30685
rect 28810 30676 28816 30728
rect 28868 30676 28874 30728
rect 28905 30719 28963 30725
rect 28905 30685 28917 30719
rect 28951 30716 28963 30719
rect 29086 30716 29092 30728
rect 28951 30688 29092 30716
rect 28951 30685 28963 30688
rect 28905 30679 28963 30685
rect 29086 30676 29092 30688
rect 29144 30676 29150 30728
rect 27663 30620 28028 30648
rect 27663 30617 27675 30620
rect 27617 30611 27675 30617
rect 28442 30608 28448 30660
rect 28500 30648 28506 30660
rect 29564 30648 29592 30756
rect 30374 30744 30380 30756
rect 30432 30744 30438 30796
rect 32766 30744 32772 30796
rect 32824 30744 32830 30796
rect 31938 30716 31944 30728
rect 28500 30620 29592 30648
rect 30392 30688 31944 30716
rect 28500 30608 28506 30620
rect 15120 30552 16620 30580
rect 20162 30540 20168 30592
rect 20220 30580 20226 30592
rect 23566 30580 23572 30592
rect 20220 30552 23572 30580
rect 20220 30540 20226 30552
rect 23566 30540 23572 30552
rect 23624 30580 23630 30592
rect 30392 30580 30420 30688
rect 31938 30676 31944 30688
rect 31996 30716 32002 30728
rect 32217 30719 32275 30725
rect 32217 30716 32229 30719
rect 31996 30688 32229 30716
rect 31996 30676 32002 30688
rect 32217 30685 32229 30688
rect 32263 30685 32275 30719
rect 32217 30679 32275 30685
rect 32493 30719 32551 30725
rect 32493 30685 32505 30719
rect 32539 30716 32551 30719
rect 32968 30716 32996 30880
rect 34606 30744 34612 30796
rect 34664 30784 34670 30796
rect 35710 30784 35716 30796
rect 34664 30756 35716 30784
rect 34664 30744 34670 30756
rect 35710 30744 35716 30756
rect 35768 30744 35774 30796
rect 35986 30744 35992 30796
rect 36044 30744 36050 30796
rect 35069 30719 35127 30725
rect 35069 30716 35081 30719
rect 32539 30688 32996 30716
rect 34072 30688 35081 30716
rect 32539 30685 32551 30688
rect 32493 30679 32551 30685
rect 32232 30648 32260 30679
rect 34072 30660 34100 30688
rect 35069 30685 35081 30688
rect 35115 30685 35127 30719
rect 35069 30679 35127 30685
rect 35434 30676 35440 30728
rect 35492 30716 35498 30728
rect 35897 30719 35955 30725
rect 35897 30716 35909 30719
rect 35492 30688 35909 30716
rect 35492 30676 35498 30688
rect 35897 30685 35909 30688
rect 35943 30716 35955 30719
rect 36078 30716 36084 30728
rect 35943 30688 36084 30716
rect 35943 30685 35955 30688
rect 35897 30679 35955 30685
rect 36078 30676 36084 30688
rect 36136 30676 36142 30728
rect 33502 30648 33508 30660
rect 32232 30620 33508 30648
rect 33502 30608 33508 30620
rect 33560 30608 33566 30660
rect 34054 30608 34060 30660
rect 34112 30608 34118 30660
rect 34330 30608 34336 30660
rect 34388 30648 34394 30660
rect 34885 30651 34943 30657
rect 34885 30648 34897 30651
rect 34388 30620 34897 30648
rect 34388 30608 34394 30620
rect 34885 30617 34897 30620
rect 34931 30617 34943 30651
rect 34885 30611 34943 30617
rect 23624 30552 30420 30580
rect 23624 30540 23630 30552
rect 30926 30540 30932 30592
rect 30984 30580 30990 30592
rect 32309 30583 32367 30589
rect 32309 30580 32321 30583
rect 30984 30552 32321 30580
rect 30984 30540 30990 30552
rect 32309 30549 32321 30552
rect 32355 30549 32367 30583
rect 32309 30543 32367 30549
rect 1104 30490 38272 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 38272 30490
rect 1104 30416 38272 30438
rect 3513 30379 3571 30385
rect 3513 30345 3525 30379
rect 3559 30376 3571 30379
rect 4062 30376 4068 30388
rect 3559 30348 4068 30376
rect 3559 30345 3571 30348
rect 3513 30339 3571 30345
rect 4062 30336 4068 30348
rect 4120 30336 4126 30388
rect 4430 30336 4436 30388
rect 4488 30336 4494 30388
rect 4522 30336 4528 30388
rect 4580 30376 4586 30388
rect 4580 30348 4936 30376
rect 4580 30336 4586 30348
rect 4908 30317 4936 30348
rect 7282 30336 7288 30388
rect 7340 30376 7346 30388
rect 8113 30379 8171 30385
rect 8113 30376 8125 30379
rect 7340 30348 8125 30376
rect 7340 30336 7346 30348
rect 8113 30345 8125 30348
rect 8159 30345 8171 30379
rect 8113 30339 8171 30345
rect 8938 30336 8944 30388
rect 8996 30336 9002 30388
rect 13446 30336 13452 30388
rect 13504 30336 13510 30388
rect 20533 30379 20591 30385
rect 20533 30376 20545 30379
rect 19996 30348 20545 30376
rect 4893 30311 4951 30317
rect 3344 30280 4660 30308
rect 3344 30252 3372 30280
rect 4632 30252 4660 30280
rect 4893 30277 4905 30311
rect 4939 30277 4951 30311
rect 4893 30271 4951 30277
rect 4985 30311 5043 30317
rect 4985 30277 4997 30311
rect 5031 30308 5043 30311
rect 5258 30308 5264 30320
rect 5031 30280 5264 30308
rect 5031 30277 5043 30280
rect 4985 30271 5043 30277
rect 5258 30268 5264 30280
rect 5316 30268 5322 30320
rect 3326 30200 3332 30252
rect 3384 30200 3390 30252
rect 3418 30200 3424 30252
rect 3476 30200 3482 30252
rect 3510 30200 3516 30252
rect 3568 30200 3574 30252
rect 4525 30243 4583 30249
rect 4525 30209 4537 30243
rect 4571 30209 4583 30243
rect 4525 30203 4583 30209
rect 3237 30175 3295 30181
rect 3237 30141 3249 30175
rect 3283 30141 3295 30175
rect 3237 30135 3295 30141
rect 3252 30104 3280 30135
rect 3602 30132 3608 30184
rect 3660 30132 3666 30184
rect 4540 30172 4568 30203
rect 4614 30200 4620 30252
rect 4672 30200 4678 30252
rect 4765 30243 4823 30249
rect 4765 30209 4777 30243
rect 4811 30240 4823 30243
rect 5121 30243 5179 30249
rect 4811 30212 5028 30240
rect 4811 30209 4823 30212
rect 4765 30203 4823 30209
rect 5000 30184 5028 30212
rect 5121 30209 5133 30243
rect 5167 30240 5179 30243
rect 5442 30240 5448 30252
rect 5167 30212 5448 30240
rect 5167 30209 5179 30212
rect 5121 30203 5179 30209
rect 4540 30144 4844 30172
rect 4816 30116 4844 30144
rect 4982 30132 4988 30184
rect 5040 30132 5046 30184
rect 4706 30104 4712 30116
rect 3252 30076 4712 30104
rect 4706 30064 4712 30076
rect 4764 30064 4770 30116
rect 4798 30064 4804 30116
rect 4856 30064 4862 30116
rect 5138 30104 5166 30203
rect 5442 30200 5448 30212
rect 5500 30200 5506 30252
rect 8297 30243 8355 30249
rect 8297 30209 8309 30243
rect 8343 30240 8355 30243
rect 8956 30240 8984 30336
rect 8343 30212 8984 30240
rect 8343 30209 8355 30212
rect 8297 30203 8355 30209
rect 13262 30200 13268 30252
rect 13320 30200 13326 30252
rect 13464 30249 13492 30336
rect 13538 30268 13544 30320
rect 13596 30308 13602 30320
rect 13596 30280 14228 30308
rect 13596 30268 13602 30280
rect 13357 30243 13415 30249
rect 13357 30209 13369 30243
rect 13403 30209 13415 30243
rect 13357 30203 13415 30209
rect 13449 30243 13507 30249
rect 13449 30209 13461 30243
rect 13495 30209 13507 30243
rect 13449 30203 13507 30209
rect 13633 30243 13691 30249
rect 13633 30209 13645 30243
rect 13679 30240 13691 30243
rect 13814 30240 13820 30252
rect 13679 30212 13820 30240
rect 13679 30209 13691 30212
rect 13633 30203 13691 30209
rect 6546 30132 6552 30184
rect 6604 30132 6610 30184
rect 13372 30172 13400 30203
rect 13814 30200 13820 30212
rect 13872 30240 13878 30252
rect 14090 30240 14096 30252
rect 13872 30212 14096 30240
rect 13872 30200 13878 30212
rect 14090 30200 14096 30212
rect 14148 30200 14154 30252
rect 14200 30240 14228 30280
rect 17678 30268 17684 30320
rect 17736 30308 17742 30320
rect 19996 30317 20024 30348
rect 20533 30345 20545 30348
rect 20579 30376 20591 30379
rect 27985 30379 28043 30385
rect 20579 30348 24900 30376
rect 20579 30345 20591 30348
rect 20533 30339 20591 30345
rect 19981 30311 20039 30317
rect 19981 30308 19993 30311
rect 17736 30280 19993 30308
rect 17736 30268 17742 30280
rect 19981 30277 19993 30280
rect 20027 30277 20039 30311
rect 19981 30271 20039 30277
rect 20197 30311 20255 30317
rect 20197 30277 20209 30311
rect 20243 30308 20255 30311
rect 20717 30311 20775 30317
rect 20717 30308 20729 30311
rect 20243 30280 20729 30308
rect 20243 30277 20255 30280
rect 20197 30271 20255 30277
rect 20717 30277 20729 30280
rect 20763 30308 20775 30311
rect 20990 30308 20996 30320
rect 20763 30280 20996 30308
rect 20763 30277 20775 30280
rect 20717 30271 20775 30277
rect 20990 30268 20996 30280
rect 21048 30308 21054 30320
rect 21910 30308 21916 30320
rect 21048 30280 21916 30308
rect 21048 30268 21054 30280
rect 21910 30268 21916 30280
rect 21968 30268 21974 30320
rect 22738 30268 22744 30320
rect 22796 30308 22802 30320
rect 23293 30311 23351 30317
rect 23293 30308 23305 30311
rect 22796 30280 23305 30308
rect 22796 30268 22802 30280
rect 23293 30277 23305 30280
rect 23339 30308 23351 30311
rect 23382 30308 23388 30320
rect 23339 30280 23388 30308
rect 23339 30277 23351 30280
rect 23293 30271 23351 30277
rect 23382 30268 23388 30280
rect 23440 30268 23446 30320
rect 23676 30280 24532 30308
rect 19610 30240 19616 30252
rect 14200 30212 19616 30240
rect 19610 30200 19616 30212
rect 19668 30240 19674 30252
rect 20070 30240 20076 30252
rect 19668 30212 20076 30240
rect 19668 30200 19674 30212
rect 20070 30200 20076 30212
rect 20128 30200 20134 30252
rect 20441 30243 20499 30249
rect 20441 30240 20453 30243
rect 20180 30212 20453 30240
rect 13372 30144 13676 30172
rect 4908 30076 5166 30104
rect 5261 30107 5319 30113
rect 3970 29996 3976 30048
rect 4028 30036 4034 30048
rect 4249 30039 4307 30045
rect 4249 30036 4261 30039
rect 4028 30008 4261 30036
rect 4028 29996 4034 30008
rect 4249 30005 4261 30008
rect 4295 30005 4307 30039
rect 4249 29999 4307 30005
rect 4338 29996 4344 30048
rect 4396 30036 4402 30048
rect 4908 30036 4936 30076
rect 5261 30073 5273 30107
rect 5307 30104 5319 30107
rect 6564 30104 6592 30132
rect 5307 30076 6592 30104
rect 5307 30073 5319 30076
rect 5261 30067 5319 30073
rect 13648 30048 13676 30144
rect 13722 30064 13728 30116
rect 13780 30104 13786 30116
rect 19886 30104 19892 30116
rect 13780 30076 19892 30104
rect 13780 30064 13786 30076
rect 19886 30064 19892 30076
rect 19944 30064 19950 30116
rect 4396 30008 4936 30036
rect 4396 29996 4402 30008
rect 4982 29996 4988 30048
rect 5040 30036 5046 30048
rect 10594 30036 10600 30048
rect 5040 30008 10600 30036
rect 5040 29996 5046 30008
rect 10594 29996 10600 30008
rect 10652 29996 10658 30048
rect 12618 29996 12624 30048
rect 12676 30036 12682 30048
rect 12989 30039 13047 30045
rect 12989 30036 13001 30039
rect 12676 30008 13001 30036
rect 12676 29996 12682 30008
rect 12989 30005 13001 30008
rect 13035 30005 13047 30039
rect 12989 29999 13047 30005
rect 13630 29996 13636 30048
rect 13688 29996 13694 30048
rect 15654 29996 15660 30048
rect 15712 30036 15718 30048
rect 20180 30045 20208 30212
rect 20441 30209 20453 30212
rect 20487 30209 20499 30243
rect 20441 30203 20499 30209
rect 23109 30243 23167 30249
rect 23109 30209 23121 30243
rect 23155 30240 23167 30243
rect 23474 30240 23480 30252
rect 23155 30212 23480 30240
rect 23155 30209 23167 30212
rect 23109 30203 23167 30209
rect 23474 30200 23480 30212
rect 23532 30240 23538 30252
rect 23676 30240 23704 30280
rect 23532 30212 23704 30240
rect 23532 30200 23538 30212
rect 23750 30200 23756 30252
rect 23808 30200 23814 30252
rect 24213 30243 24271 30249
rect 24213 30240 24225 30243
rect 24044 30212 24225 30240
rect 23566 30132 23572 30184
rect 23624 30172 23630 30184
rect 23661 30175 23719 30181
rect 23661 30172 23673 30175
rect 23624 30144 23673 30172
rect 23624 30132 23630 30144
rect 23661 30141 23673 30144
rect 23707 30141 23719 30175
rect 23661 30135 23719 30141
rect 23842 30132 23848 30184
rect 23900 30132 23906 30184
rect 23937 30175 23995 30181
rect 23937 30141 23949 30175
rect 23983 30141 23995 30175
rect 23937 30135 23995 30141
rect 23474 30064 23480 30116
rect 23532 30104 23538 30116
rect 23952 30104 23980 30135
rect 23532 30076 23980 30104
rect 23532 30064 23538 30076
rect 24044 30048 24072 30212
rect 24213 30209 24225 30212
rect 24259 30209 24271 30243
rect 24213 30203 24271 30209
rect 24397 30243 24455 30249
rect 24397 30209 24409 30243
rect 24443 30209 24455 30243
rect 24397 30203 24455 30209
rect 24121 30175 24179 30181
rect 24121 30141 24133 30175
rect 24167 30172 24179 30175
rect 24412 30172 24440 30203
rect 24167 30144 24440 30172
rect 24504 30172 24532 30280
rect 24872 30252 24900 30348
rect 27985 30345 27997 30379
rect 28031 30376 28043 30379
rect 28074 30376 28080 30388
rect 28031 30348 28080 30376
rect 28031 30345 28043 30348
rect 27985 30339 28043 30345
rect 28074 30336 28080 30348
rect 28132 30376 28138 30388
rect 28534 30376 28540 30388
rect 28132 30348 28540 30376
rect 28132 30336 28138 30348
rect 28534 30336 28540 30348
rect 28592 30336 28598 30388
rect 28626 30336 28632 30388
rect 28684 30376 28690 30388
rect 37550 30376 37556 30388
rect 28684 30348 37556 30376
rect 28684 30336 28690 30348
rect 37550 30336 37556 30348
rect 37608 30336 37614 30388
rect 27617 30311 27675 30317
rect 27617 30277 27629 30311
rect 27663 30308 27675 30311
rect 27706 30308 27712 30320
rect 27663 30280 27712 30308
rect 27663 30277 27675 30280
rect 27617 30271 27675 30277
rect 27706 30268 27712 30280
rect 27764 30268 27770 30320
rect 28166 30308 28172 30320
rect 28092 30280 28172 30308
rect 24854 30200 24860 30252
rect 24912 30200 24918 30252
rect 26418 30200 26424 30252
rect 26476 30240 26482 30252
rect 28092 30249 28120 30280
rect 28166 30268 28172 30280
rect 28224 30268 28230 30320
rect 29641 30311 29699 30317
rect 29641 30277 29653 30311
rect 29687 30308 29699 30311
rect 30190 30308 30196 30320
rect 29687 30280 30196 30308
rect 29687 30277 29699 30280
rect 29641 30271 29699 30277
rect 30190 30268 30196 30280
rect 30248 30308 30254 30320
rect 30248 30280 30512 30308
rect 30248 30268 30254 30280
rect 27801 30243 27859 30249
rect 27801 30240 27813 30243
rect 26476 30212 27813 30240
rect 26476 30200 26482 30212
rect 27801 30209 27813 30212
rect 27847 30209 27859 30243
rect 27801 30203 27859 30209
rect 28077 30243 28135 30249
rect 28077 30209 28089 30243
rect 28123 30209 28135 30243
rect 28077 30203 28135 30209
rect 27816 30172 27844 30203
rect 28258 30200 28264 30252
rect 28316 30200 28322 30252
rect 29549 30243 29607 30249
rect 29549 30209 29561 30243
rect 29595 30240 29607 30243
rect 29733 30243 29791 30249
rect 29595 30212 29684 30240
rect 29595 30209 29607 30212
rect 29549 30203 29607 30209
rect 29656 30184 29684 30212
rect 29733 30209 29745 30243
rect 29779 30209 29791 30243
rect 29733 30203 29791 30209
rect 28169 30175 28227 30181
rect 28169 30172 28181 30175
rect 24504 30144 27614 30172
rect 27816 30144 28181 30172
rect 24167 30141 24179 30144
rect 24121 30135 24179 30141
rect 24489 30107 24547 30113
rect 24489 30073 24501 30107
rect 24535 30073 24547 30107
rect 27586 30104 27614 30144
rect 28169 30141 28181 30144
rect 28215 30141 28227 30175
rect 28169 30135 28227 30141
rect 29638 30132 29644 30184
rect 29696 30132 29702 30184
rect 29748 30104 29776 30203
rect 29914 30200 29920 30252
rect 29972 30240 29978 30252
rect 30009 30243 30067 30249
rect 30009 30240 30021 30243
rect 29972 30212 30021 30240
rect 29972 30200 29978 30212
rect 30009 30209 30021 30212
rect 30055 30209 30067 30243
rect 30009 30203 30067 30209
rect 30285 30243 30343 30249
rect 30285 30209 30297 30243
rect 30331 30240 30343 30243
rect 30374 30240 30380 30252
rect 30331 30212 30380 30240
rect 30331 30209 30343 30212
rect 30285 30203 30343 30209
rect 30024 30172 30052 30203
rect 30374 30200 30380 30212
rect 30432 30200 30438 30252
rect 30484 30249 30512 30280
rect 31386 30268 31392 30320
rect 31444 30308 31450 30320
rect 34606 30308 34612 30320
rect 31444 30280 34612 30308
rect 31444 30268 31450 30280
rect 34606 30268 34612 30280
rect 34664 30268 34670 30320
rect 30469 30243 30527 30249
rect 30469 30209 30481 30243
rect 30515 30209 30527 30243
rect 30745 30243 30803 30249
rect 30745 30240 30757 30243
rect 30469 30203 30527 30209
rect 30668 30212 30757 30240
rect 30561 30175 30619 30181
rect 30561 30172 30573 30175
rect 30024 30144 30573 30172
rect 30561 30141 30573 30144
rect 30607 30141 30619 30175
rect 30561 30135 30619 30141
rect 30668 30104 30696 30212
rect 30745 30209 30757 30212
rect 30791 30209 30803 30243
rect 30745 30203 30803 30209
rect 32766 30200 32772 30252
rect 32824 30200 32830 30252
rect 30926 30132 30932 30184
rect 30984 30132 30990 30184
rect 32674 30132 32680 30184
rect 32732 30132 32738 30184
rect 33597 30175 33655 30181
rect 33597 30141 33609 30175
rect 33643 30172 33655 30175
rect 33643 30144 37228 30172
rect 33643 30141 33655 30144
rect 33597 30135 33655 30141
rect 27586 30076 28212 30104
rect 24489 30067 24547 30073
rect 20165 30039 20223 30045
rect 20165 30036 20177 30039
rect 15712 30008 20177 30036
rect 15712 29996 15718 30008
rect 20165 30005 20177 30008
rect 20211 30005 20223 30039
rect 20165 29999 20223 30005
rect 20346 29996 20352 30048
rect 20404 29996 20410 30048
rect 20714 29996 20720 30048
rect 20772 29996 20778 30048
rect 24026 29996 24032 30048
rect 24084 29996 24090 30048
rect 24118 29996 24124 30048
rect 24176 30036 24182 30048
rect 24504 30036 24532 30067
rect 28184 30048 28212 30076
rect 29472 30076 30696 30104
rect 29472 30048 29500 30076
rect 24176 30008 24532 30036
rect 24176 29996 24182 30008
rect 28166 29996 28172 30048
rect 28224 29996 28230 30048
rect 29454 29996 29460 30048
rect 29512 29996 29518 30048
rect 29638 29996 29644 30048
rect 29696 30036 29702 30048
rect 29825 30039 29883 30045
rect 29825 30036 29837 30039
rect 29696 30008 29837 30036
rect 29696 29996 29702 30008
rect 29825 30005 29837 30008
rect 29871 30005 29883 30039
rect 29825 29999 29883 30005
rect 29914 29996 29920 30048
rect 29972 30036 29978 30048
rect 30944 30036 30972 30132
rect 37200 30048 37228 30144
rect 29972 30008 30972 30036
rect 29972 29996 29978 30008
rect 37182 29996 37188 30048
rect 37240 29996 37246 30048
rect 1104 29946 38272 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38272 29946
rect 1104 29872 38272 29894
rect 12802 29832 12808 29844
rect 2746 29804 12808 29832
rect 1397 29699 1455 29705
rect 1397 29665 1409 29699
rect 1443 29696 1455 29699
rect 1762 29696 1768 29708
rect 1443 29668 1768 29696
rect 1443 29665 1455 29668
rect 1397 29659 1455 29665
rect 1762 29656 1768 29668
rect 1820 29656 1826 29708
rect 2746 29696 2774 29804
rect 12802 29792 12808 29804
rect 12860 29792 12866 29844
rect 14553 29835 14611 29841
rect 14553 29801 14565 29835
rect 14599 29832 14611 29835
rect 20257 29835 20315 29841
rect 14599 29804 19334 29832
rect 14599 29801 14611 29804
rect 14553 29795 14611 29801
rect 3145 29767 3203 29773
rect 3145 29733 3157 29767
rect 3191 29764 3203 29767
rect 3602 29764 3608 29776
rect 3191 29736 3608 29764
rect 3191 29733 3203 29736
rect 3145 29727 3203 29733
rect 3602 29724 3608 29736
rect 3660 29724 3666 29776
rect 4798 29724 4804 29776
rect 4856 29724 4862 29776
rect 4982 29724 4988 29776
rect 5040 29764 5046 29776
rect 5077 29767 5135 29773
rect 5077 29764 5089 29767
rect 5040 29736 5089 29764
rect 5040 29724 5046 29736
rect 5077 29733 5089 29736
rect 5123 29733 5135 29767
rect 5077 29727 5135 29733
rect 10137 29767 10195 29773
rect 10137 29733 10149 29767
rect 10183 29733 10195 29767
rect 10137 29727 10195 29733
rect 2700 29668 2774 29696
rect 2700 29640 2728 29668
rect 2682 29588 2688 29640
rect 2740 29588 2746 29640
rect 2774 29588 2780 29640
rect 2832 29588 2838 29640
rect 4522 29588 4528 29640
rect 4580 29628 4586 29640
rect 4816 29628 4844 29724
rect 7009 29699 7067 29705
rect 7009 29665 7021 29699
rect 7055 29696 7067 29699
rect 8018 29696 8024 29708
rect 7055 29668 8024 29696
rect 7055 29665 7067 29668
rect 7009 29659 7067 29665
rect 8018 29656 8024 29668
rect 8076 29656 8082 29708
rect 4985 29631 5043 29637
rect 4985 29628 4997 29631
rect 4580 29600 4997 29628
rect 4580 29588 4586 29600
rect 4985 29597 4997 29600
rect 5031 29597 5043 29631
rect 4985 29591 5043 29597
rect 5169 29631 5227 29637
rect 5169 29597 5181 29631
rect 5215 29597 5227 29631
rect 5169 29591 5227 29597
rect 9861 29631 9919 29637
rect 9861 29597 9873 29631
rect 9907 29628 9919 29631
rect 10152 29628 10180 29727
rect 12066 29724 12072 29776
rect 12124 29764 12130 29776
rect 12342 29764 12348 29776
rect 12124 29736 12348 29764
rect 12124 29724 12130 29736
rect 12342 29724 12348 29736
rect 12400 29724 12406 29776
rect 12710 29724 12716 29776
rect 12768 29764 12774 29776
rect 12768 29736 13400 29764
rect 12768 29724 12774 29736
rect 13372 29708 13400 29736
rect 15102 29724 15108 29776
rect 15160 29724 15166 29776
rect 15565 29767 15623 29773
rect 15565 29764 15577 29767
rect 15212 29736 15577 29764
rect 10686 29656 10692 29708
rect 10744 29696 10750 29708
rect 10870 29696 10876 29708
rect 10744 29668 10876 29696
rect 10744 29656 10750 29668
rect 10870 29656 10876 29668
rect 10928 29656 10934 29708
rect 12805 29699 12863 29705
rect 12805 29665 12817 29699
rect 12851 29696 12863 29699
rect 13170 29696 13176 29708
rect 12851 29668 13176 29696
rect 12851 29665 12863 29668
rect 12805 29659 12863 29665
rect 9907 29600 10180 29628
rect 9907 29597 9919 29600
rect 9861 29591 9919 29597
rect 1670 29520 1676 29572
rect 1728 29520 1734 29572
rect 2792 29492 2820 29588
rect 4338 29520 4344 29572
rect 4396 29560 4402 29572
rect 4706 29560 4712 29572
rect 4396 29532 4712 29560
rect 4396 29520 4402 29532
rect 4706 29520 4712 29532
rect 4764 29560 4770 29572
rect 5184 29560 5212 29591
rect 11146 29588 11152 29640
rect 11204 29628 11210 29640
rect 11425 29631 11483 29637
rect 11425 29628 11437 29631
rect 11204 29600 11437 29628
rect 11204 29588 11210 29600
rect 11425 29597 11437 29600
rect 11471 29597 11483 29631
rect 11425 29591 11483 29597
rect 4764 29532 5212 29560
rect 4764 29520 4770 29532
rect 7282 29520 7288 29572
rect 7340 29520 7346 29572
rect 10505 29563 10563 29569
rect 7392 29532 7774 29560
rect 7392 29492 7420 29532
rect 2792 29464 7420 29492
rect 7668 29492 7696 29532
rect 10505 29529 10517 29563
rect 10551 29560 10563 29563
rect 10870 29560 10876 29572
rect 10551 29532 10876 29560
rect 10551 29529 10563 29532
rect 10505 29523 10563 29529
rect 10870 29520 10876 29532
rect 10928 29560 10934 29572
rect 11609 29563 11667 29569
rect 11609 29560 11621 29563
rect 10928 29532 11621 29560
rect 10928 29520 10934 29532
rect 11609 29529 11621 29532
rect 11655 29560 11667 29563
rect 12710 29560 12716 29572
rect 11655 29532 12716 29560
rect 11655 29529 11667 29532
rect 11609 29523 11667 29529
rect 12710 29520 12716 29532
rect 12768 29520 12774 29572
rect 12820 29560 12848 29659
rect 13170 29656 13176 29668
rect 13228 29656 13234 29708
rect 13354 29656 13360 29708
rect 13412 29696 13418 29708
rect 13722 29696 13728 29708
rect 13412 29668 13728 29696
rect 13412 29656 13418 29668
rect 13722 29656 13728 29668
rect 13780 29656 13786 29708
rect 14369 29699 14427 29705
rect 14369 29665 14381 29699
rect 14415 29696 14427 29699
rect 15120 29696 15148 29724
rect 15212 29705 15240 29736
rect 15565 29733 15577 29736
rect 15611 29733 15623 29767
rect 15565 29727 15623 29733
rect 15838 29724 15844 29776
rect 15896 29764 15902 29776
rect 16577 29767 16635 29773
rect 15896 29736 16160 29764
rect 15896 29724 15902 29736
rect 16132 29708 16160 29736
rect 16577 29733 16589 29767
rect 16623 29764 16635 29767
rect 18138 29764 18144 29776
rect 16623 29736 18144 29764
rect 16623 29733 16635 29736
rect 16577 29727 16635 29733
rect 18138 29724 18144 29736
rect 18196 29724 18202 29776
rect 14415 29668 15148 29696
rect 15197 29699 15255 29705
rect 14415 29665 14427 29668
rect 14369 29659 14427 29665
rect 15197 29665 15209 29699
rect 15243 29665 15255 29699
rect 15197 29659 15255 29665
rect 15473 29699 15531 29705
rect 15473 29665 15485 29699
rect 15519 29696 15531 29699
rect 15654 29696 15660 29708
rect 15519 29668 15660 29696
rect 15519 29665 15531 29668
rect 15473 29659 15531 29665
rect 15654 29656 15660 29668
rect 15712 29656 15718 29708
rect 15930 29656 15936 29708
rect 15988 29696 15994 29708
rect 16025 29699 16083 29705
rect 16025 29696 16037 29699
rect 15988 29668 16037 29696
rect 15988 29656 15994 29668
rect 16025 29665 16037 29668
rect 16071 29665 16083 29699
rect 16025 29659 16083 29665
rect 16114 29656 16120 29708
rect 16172 29656 16178 29708
rect 19306 29696 19334 29804
rect 20257 29801 20269 29835
rect 20303 29832 20315 29835
rect 20346 29832 20352 29844
rect 20303 29804 20352 29832
rect 20303 29801 20315 29804
rect 20257 29795 20315 29801
rect 20346 29792 20352 29804
rect 20404 29792 20410 29844
rect 20625 29835 20683 29841
rect 20625 29801 20637 29835
rect 20671 29832 20683 29835
rect 20714 29832 20720 29844
rect 20671 29804 20720 29832
rect 20671 29801 20683 29804
rect 20625 29795 20683 29801
rect 20088 29736 20576 29764
rect 20088 29705 20116 29736
rect 20548 29705 20576 29736
rect 20073 29699 20131 29705
rect 20073 29696 20085 29699
rect 19306 29668 20085 29696
rect 20073 29665 20085 29668
rect 20119 29665 20131 29699
rect 20073 29659 20131 29665
rect 20533 29699 20591 29705
rect 20533 29665 20545 29699
rect 20579 29665 20591 29699
rect 20533 29659 20591 29665
rect 12894 29588 12900 29640
rect 12952 29628 12958 29640
rect 13081 29631 13139 29637
rect 13081 29628 13093 29631
rect 12952 29600 13093 29628
rect 12952 29588 12958 29600
rect 13081 29597 13093 29600
rect 13127 29597 13139 29631
rect 13081 29591 13139 29597
rect 13262 29588 13268 29640
rect 13320 29628 13326 29640
rect 14277 29631 14335 29637
rect 14277 29628 14289 29631
rect 13320 29600 14289 29628
rect 13320 29588 13326 29600
rect 14277 29597 14289 29600
rect 14323 29597 14335 29631
rect 14277 29591 14335 29597
rect 15105 29631 15163 29637
rect 15105 29597 15117 29631
rect 15151 29628 15163 29631
rect 15838 29628 15844 29640
rect 15151 29600 15844 29628
rect 15151 29597 15163 29600
rect 15105 29591 15163 29597
rect 12989 29563 13047 29569
rect 12820 29532 12940 29560
rect 12912 29504 12940 29532
rect 12989 29529 13001 29563
rect 13035 29560 13047 29563
rect 14182 29560 14188 29572
rect 13035 29532 14188 29560
rect 13035 29529 13047 29532
rect 12989 29523 13047 29529
rect 14182 29520 14188 29532
rect 14240 29520 14246 29572
rect 8294 29492 8300 29504
rect 7668 29464 8300 29492
rect 8294 29452 8300 29464
rect 8352 29452 8358 29504
rect 8754 29452 8760 29504
rect 8812 29452 8818 29504
rect 9674 29452 9680 29504
rect 9732 29452 9738 29504
rect 10597 29495 10655 29501
rect 10597 29461 10609 29495
rect 10643 29492 10655 29495
rect 11514 29492 11520 29504
rect 10643 29464 11520 29492
rect 10643 29461 10655 29464
rect 10597 29455 10655 29461
rect 11514 29452 11520 29464
rect 11572 29452 11578 29504
rect 11790 29452 11796 29504
rect 11848 29452 11854 29504
rect 12894 29452 12900 29504
rect 12952 29452 12958 29504
rect 13446 29452 13452 29504
rect 13504 29452 13510 29504
rect 14292 29492 14320 29591
rect 15838 29588 15844 29600
rect 15896 29628 15902 29640
rect 16393 29631 16451 29637
rect 16393 29628 16405 29631
rect 15896 29600 16405 29628
rect 15896 29588 15902 29600
rect 16393 29597 16405 29600
rect 16439 29597 16451 29631
rect 16393 29591 16451 29597
rect 16577 29631 16635 29637
rect 16577 29597 16589 29631
rect 16623 29628 16635 29631
rect 17218 29628 17224 29640
rect 16623 29600 17224 29628
rect 16623 29597 16635 29600
rect 16577 29591 16635 29597
rect 15933 29563 15991 29569
rect 15933 29529 15945 29563
rect 15979 29560 15991 29563
rect 16592 29560 16620 29591
rect 17218 29588 17224 29600
rect 17276 29588 17282 29640
rect 20349 29631 20407 29637
rect 20349 29597 20361 29631
rect 20395 29597 20407 29631
rect 20349 29591 20407 29597
rect 15979 29532 16620 29560
rect 20364 29560 20392 29591
rect 20438 29588 20444 29640
rect 20496 29588 20502 29640
rect 20640 29560 20668 29795
rect 20714 29792 20720 29804
rect 20772 29792 20778 29844
rect 23382 29792 23388 29844
rect 23440 29792 23446 29844
rect 23753 29835 23811 29841
rect 23753 29801 23765 29835
rect 23799 29832 23811 29835
rect 24026 29832 24032 29844
rect 23799 29804 24032 29832
rect 23799 29801 23811 29804
rect 23753 29795 23811 29801
rect 24026 29792 24032 29804
rect 24084 29792 24090 29844
rect 26602 29792 26608 29844
rect 26660 29832 26666 29844
rect 27154 29832 27160 29844
rect 26660 29804 27160 29832
rect 26660 29792 26666 29804
rect 27154 29792 27160 29804
rect 27212 29832 27218 29844
rect 27212 29804 28580 29832
rect 27212 29792 27218 29804
rect 20898 29724 20904 29776
rect 20956 29764 20962 29776
rect 21453 29767 21511 29773
rect 20956 29736 21312 29764
rect 20956 29724 20962 29736
rect 21284 29696 21312 29736
rect 21453 29733 21465 29767
rect 21499 29764 21511 29767
rect 22186 29764 22192 29776
rect 21499 29736 22192 29764
rect 21499 29733 21511 29736
rect 21453 29727 21511 29733
rect 22186 29724 22192 29736
rect 22244 29724 22250 29776
rect 23400 29696 23428 29792
rect 28552 29776 28580 29804
rect 28920 29804 30972 29832
rect 28920 29776 28948 29804
rect 26050 29724 26056 29776
rect 26108 29764 26114 29776
rect 28353 29767 28411 29773
rect 28353 29764 28365 29767
rect 26108 29736 28365 29764
rect 26108 29724 26114 29736
rect 28353 29733 28365 29736
rect 28399 29733 28411 29767
rect 28353 29727 28411 29733
rect 28534 29724 28540 29776
rect 28592 29724 28598 29776
rect 28902 29724 28908 29776
rect 28960 29724 28966 29776
rect 30944 29764 30972 29804
rect 31018 29792 31024 29844
rect 31076 29792 31082 29844
rect 34149 29835 34207 29841
rect 34149 29801 34161 29835
rect 34195 29832 34207 29835
rect 34790 29832 34796 29844
rect 34195 29804 34796 29832
rect 34195 29801 34207 29804
rect 34149 29795 34207 29801
rect 34790 29792 34796 29804
rect 34848 29792 34854 29844
rect 34241 29767 34299 29773
rect 30944 29736 34192 29764
rect 28000 29696 28212 29704
rect 20364 29532 20668 29560
rect 20732 29668 21220 29696
rect 21284 29668 21588 29696
rect 23400 29668 24440 29696
rect 15979 29529 15991 29532
rect 15933 29523 15991 29529
rect 15562 29492 15568 29504
rect 14292 29464 15568 29492
rect 15562 29452 15568 29464
rect 15620 29492 15626 29504
rect 16206 29492 16212 29504
rect 15620 29464 16212 29492
rect 15620 29452 15626 29464
rect 16206 29452 16212 29464
rect 16264 29452 16270 29504
rect 20073 29495 20131 29501
rect 20073 29461 20085 29495
rect 20119 29492 20131 29495
rect 20732 29492 20760 29668
rect 21192 29640 21220 29668
rect 20990 29588 20996 29640
rect 21048 29628 21054 29640
rect 21085 29631 21143 29637
rect 21085 29628 21097 29631
rect 21048 29600 21097 29628
rect 21048 29588 21054 29600
rect 21085 29597 21097 29600
rect 21131 29597 21143 29631
rect 21085 29591 21143 29597
rect 21174 29588 21180 29640
rect 21232 29588 21238 29640
rect 21453 29631 21511 29637
rect 21453 29597 21465 29631
rect 21499 29597 21511 29631
rect 21453 29591 21511 29597
rect 21266 29560 21272 29572
rect 20824 29532 21272 29560
rect 20824 29501 20852 29532
rect 21266 29520 21272 29532
rect 21324 29520 21330 29572
rect 21468 29504 21496 29591
rect 21560 29560 21588 29668
rect 23474 29588 23480 29640
rect 23532 29588 23538 29640
rect 23750 29588 23756 29640
rect 23808 29588 23814 29640
rect 24412 29637 24440 29668
rect 28000 29676 28304 29696
rect 24578 29637 24584 29640
rect 24397 29631 24455 29637
rect 24397 29597 24409 29631
rect 24443 29597 24455 29631
rect 24574 29628 24584 29637
rect 24539 29600 24584 29628
rect 24397 29591 24455 29597
rect 24574 29591 24584 29600
rect 24578 29588 24584 29591
rect 24636 29588 24642 29640
rect 26418 29588 26424 29640
rect 26476 29588 26482 29640
rect 26602 29588 26608 29640
rect 26660 29588 26666 29640
rect 26697 29631 26755 29637
rect 26697 29597 26709 29631
rect 26743 29628 26755 29631
rect 26881 29631 26939 29637
rect 26881 29628 26893 29631
rect 26743 29600 26893 29628
rect 26743 29597 26755 29600
rect 26697 29591 26755 29597
rect 26881 29597 26893 29600
rect 26927 29597 26939 29631
rect 26881 29591 26939 29597
rect 26970 29588 26976 29640
rect 27028 29588 27034 29640
rect 28000 29560 28028 29676
rect 28184 29668 28304 29676
rect 28074 29588 28080 29640
rect 28132 29637 28138 29640
rect 28276 29637 28304 29668
rect 28810 29656 28816 29708
rect 28868 29705 28874 29708
rect 28868 29659 28877 29705
rect 31662 29696 31668 29708
rect 30852 29668 31668 29696
rect 28868 29656 28874 29659
rect 30852 29640 30880 29668
rect 31662 29656 31668 29668
rect 31720 29696 31726 29708
rect 31720 29668 31800 29696
rect 31720 29656 31726 29668
rect 28132 29631 28158 29637
rect 28146 29597 28158 29631
rect 28132 29591 28158 29597
rect 28261 29631 28319 29637
rect 28261 29597 28273 29631
rect 28307 29597 28319 29631
rect 28261 29591 28319 29597
rect 28132 29588 28138 29591
rect 28534 29588 28540 29640
rect 28592 29588 28598 29640
rect 28718 29588 28724 29640
rect 28776 29588 28782 29640
rect 28902 29588 28908 29640
rect 28960 29588 28966 29640
rect 29089 29631 29147 29637
rect 29089 29597 29101 29631
rect 29135 29597 29147 29631
rect 29089 29591 29147 29597
rect 29104 29560 29132 29591
rect 30374 29588 30380 29640
rect 30432 29628 30438 29640
rect 30834 29628 30840 29640
rect 30432 29600 30840 29628
rect 30432 29588 30438 29600
rect 30834 29588 30840 29600
rect 30892 29588 30898 29640
rect 31772 29637 31800 29668
rect 31021 29631 31079 29637
rect 31021 29597 31033 29631
rect 31067 29597 31079 29631
rect 31021 29591 31079 29597
rect 31757 29631 31815 29637
rect 31757 29597 31769 29631
rect 31803 29597 31815 29631
rect 31757 29591 31815 29597
rect 21560 29532 28028 29560
rect 28276 29532 29132 29560
rect 20119 29464 20760 29492
rect 20809 29495 20867 29501
rect 20119 29461 20131 29464
rect 20073 29455 20131 29461
rect 20809 29461 20821 29495
rect 20855 29461 20867 29495
rect 20809 29455 20867 29461
rect 20990 29452 20996 29504
rect 21048 29452 21054 29504
rect 21450 29452 21456 29504
rect 21508 29452 21514 29504
rect 23569 29495 23627 29501
rect 23569 29461 23581 29495
rect 23615 29492 23627 29495
rect 23842 29492 23848 29504
rect 23615 29464 23848 29492
rect 23615 29461 23627 29464
rect 23569 29455 23627 29461
rect 23842 29452 23848 29464
rect 23900 29492 23906 29504
rect 24489 29495 24547 29501
rect 24489 29492 24501 29495
rect 23900 29464 24501 29492
rect 23900 29452 23906 29464
rect 24489 29461 24501 29464
rect 24535 29492 24547 29495
rect 24762 29492 24768 29504
rect 24535 29464 24768 29492
rect 24535 29461 24547 29464
rect 24489 29455 24547 29461
rect 24762 29452 24768 29464
rect 24820 29452 24826 29504
rect 26234 29452 26240 29504
rect 26292 29452 26298 29504
rect 27338 29452 27344 29504
rect 27396 29492 27402 29504
rect 28074 29492 28080 29504
rect 27396 29464 28080 29492
rect 27396 29452 27402 29464
rect 28074 29452 28080 29464
rect 28132 29452 28138 29504
rect 28276 29501 28304 29532
rect 30006 29520 30012 29572
rect 30064 29560 30070 29572
rect 31036 29560 31064 29591
rect 32030 29588 32036 29640
rect 32088 29588 32094 29640
rect 33778 29588 33784 29640
rect 33836 29588 33842 29640
rect 33962 29588 33968 29640
rect 34020 29588 34026 29640
rect 34057 29631 34115 29637
rect 34057 29597 34069 29631
rect 34103 29597 34115 29631
rect 34164 29628 34192 29736
rect 34241 29733 34253 29767
rect 34287 29764 34299 29767
rect 34330 29764 34336 29776
rect 34287 29736 34336 29764
rect 34287 29733 34299 29736
rect 34241 29727 34299 29733
rect 34330 29724 34336 29736
rect 34388 29724 34394 29776
rect 36725 29767 36783 29773
rect 36725 29733 36737 29767
rect 36771 29733 36783 29767
rect 36725 29727 36783 29733
rect 36446 29656 36452 29708
rect 36504 29656 36510 29708
rect 36740 29696 36768 29727
rect 36740 29668 37504 29696
rect 34333 29631 34391 29637
rect 34333 29628 34345 29631
rect 34164 29600 34345 29628
rect 34057 29591 34115 29597
rect 34333 29597 34345 29600
rect 34379 29628 34391 29631
rect 34422 29628 34428 29640
rect 34379 29600 34428 29628
rect 34379 29597 34391 29600
rect 34333 29591 34391 29597
rect 31478 29560 31484 29572
rect 30064 29532 31484 29560
rect 30064 29520 30070 29532
rect 31478 29520 31484 29532
rect 31536 29520 31542 29572
rect 34072 29560 34100 29591
rect 34422 29588 34428 29600
rect 34480 29588 34486 29640
rect 36354 29588 36360 29640
rect 36412 29588 36418 29640
rect 37182 29588 37188 29640
rect 37240 29588 37246 29640
rect 37476 29637 37504 29668
rect 37461 29631 37519 29637
rect 37461 29597 37473 29631
rect 37507 29597 37519 29631
rect 37461 29591 37519 29597
rect 34072 29532 35020 29560
rect 34992 29504 35020 29532
rect 28261 29495 28319 29501
rect 28261 29461 28273 29495
rect 28307 29461 28319 29495
rect 28261 29455 28319 29461
rect 31938 29452 31944 29504
rect 31996 29492 32002 29504
rect 32033 29495 32091 29501
rect 32033 29492 32045 29495
rect 31996 29464 32045 29492
rect 31996 29452 32002 29464
rect 32033 29461 32045 29464
rect 32079 29492 32091 29495
rect 32766 29492 32772 29504
rect 32079 29464 32772 29492
rect 32079 29461 32091 29464
rect 32033 29455 32091 29461
rect 32766 29452 32772 29464
rect 32824 29452 32830 29504
rect 34974 29452 34980 29504
rect 35032 29452 35038 29504
rect 36814 29452 36820 29504
rect 36872 29452 36878 29504
rect 1104 29402 38272 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 38272 29402
rect 1104 29328 38272 29350
rect 1670 29248 1676 29300
rect 1728 29288 1734 29300
rect 1857 29291 1915 29297
rect 1857 29288 1869 29291
rect 1728 29260 1869 29288
rect 1728 29248 1734 29260
rect 1857 29257 1869 29260
rect 1903 29257 1915 29291
rect 1857 29251 1915 29257
rect 3605 29291 3663 29297
rect 3605 29257 3617 29291
rect 3651 29288 3663 29291
rect 3970 29288 3976 29300
rect 3651 29260 3976 29288
rect 3651 29257 3663 29260
rect 3605 29251 3663 29257
rect 3970 29248 3976 29260
rect 4028 29248 4034 29300
rect 4522 29248 4528 29300
rect 4580 29248 4586 29300
rect 5074 29248 5080 29300
rect 5132 29288 5138 29300
rect 5169 29291 5227 29297
rect 5169 29288 5181 29291
rect 5132 29260 5181 29288
rect 5132 29248 5138 29260
rect 5169 29257 5181 29260
rect 5215 29257 5227 29291
rect 5169 29251 5227 29257
rect 7282 29248 7288 29300
rect 7340 29288 7346 29300
rect 8021 29291 8079 29297
rect 8021 29288 8033 29291
rect 7340 29260 8033 29288
rect 7340 29248 7346 29260
rect 8021 29257 8033 29260
rect 8067 29257 8079 29291
rect 8021 29251 8079 29257
rect 8772 29260 10824 29288
rect 4540 29161 4568 29248
rect 8772 29232 8800 29260
rect 7469 29223 7527 29229
rect 5092 29192 6868 29220
rect 2041 29155 2099 29161
rect 2041 29121 2053 29155
rect 2087 29152 2099 29155
rect 3697 29155 3755 29161
rect 2087 29124 2774 29152
rect 2087 29121 2099 29124
rect 2041 29115 2099 29121
rect 2746 29016 2774 29124
rect 3697 29121 3709 29155
rect 3743 29152 3755 29155
rect 4525 29155 4583 29161
rect 3743 29124 4476 29152
rect 3743 29121 3755 29124
rect 3697 29115 3755 29121
rect 3881 29087 3939 29093
rect 3881 29053 3893 29087
rect 3927 29053 3939 29087
rect 3881 29047 3939 29053
rect 3237 29019 3295 29025
rect 3237 29016 3249 29019
rect 2746 28988 3249 29016
rect 3237 28985 3249 28988
rect 3283 28985 3295 29019
rect 3896 29016 3924 29047
rect 4338 29044 4344 29096
rect 4396 29044 4402 29096
rect 4448 29084 4476 29124
rect 4525 29121 4537 29155
rect 4571 29121 4583 29155
rect 4525 29115 4583 29121
rect 4798 29112 4804 29164
rect 4856 29161 4862 29164
rect 4856 29155 4883 29161
rect 4871 29121 4883 29155
rect 4856 29115 4883 29121
rect 4856 29112 4862 29115
rect 4982 29112 4988 29164
rect 5040 29112 5046 29164
rect 5092 29161 5120 29192
rect 6840 29164 6868 29192
rect 7469 29189 7481 29223
rect 7515 29220 7527 29223
rect 8754 29220 8760 29232
rect 7515 29192 8760 29220
rect 7515 29189 7527 29192
rect 7469 29183 7527 29189
rect 8754 29180 8760 29192
rect 8812 29180 8818 29232
rect 9401 29223 9459 29229
rect 9401 29189 9413 29223
rect 9447 29220 9459 29223
rect 9674 29220 9680 29232
rect 9447 29192 9680 29220
rect 9447 29189 9459 29192
rect 9401 29183 9459 29189
rect 9674 29180 9680 29192
rect 9732 29180 9738 29232
rect 9858 29180 9864 29232
rect 9916 29180 9922 29232
rect 5077 29155 5135 29161
rect 5077 29121 5089 29155
rect 5123 29121 5135 29155
rect 5077 29115 5135 29121
rect 5092 29084 5120 29115
rect 5258 29112 5264 29164
rect 5316 29112 5322 29164
rect 6822 29112 6828 29164
rect 6880 29112 6886 29164
rect 7561 29155 7619 29161
rect 7561 29121 7573 29155
rect 7607 29121 7619 29155
rect 8205 29155 8263 29161
rect 8205 29152 8217 29155
rect 7561 29115 7619 29121
rect 7944 29124 8217 29152
rect 4448 29056 5120 29084
rect 6914 29044 6920 29096
rect 6972 29084 6978 29096
rect 7282 29084 7288 29096
rect 6972 29056 7288 29084
rect 6972 29044 6978 29056
rect 7282 29044 7288 29056
rect 7340 29044 7346 29096
rect 4614 29016 4620 29028
rect 3896 28988 4620 29016
rect 3237 28979 3295 28985
rect 4614 28976 4620 28988
rect 4672 29016 4678 29028
rect 4982 29016 4988 29028
rect 4672 28988 4988 29016
rect 4672 28976 4678 28988
rect 4982 28976 4988 28988
rect 5040 28976 5046 29028
rect 7576 29016 7604 29115
rect 7944 29025 7972 29124
rect 8205 29121 8217 29124
rect 8251 29121 8263 29155
rect 8205 29115 8263 29121
rect 8018 29044 8024 29096
rect 8076 29084 8082 29096
rect 9125 29087 9183 29093
rect 9125 29084 9137 29087
rect 8076 29056 9137 29084
rect 8076 29044 8082 29056
rect 9125 29053 9137 29056
rect 9171 29053 9183 29087
rect 9125 29047 9183 29053
rect 6196 28988 7604 29016
rect 7929 29019 7987 29025
rect 6196 28960 6224 28988
rect 7929 28985 7941 29019
rect 7975 28985 7987 29019
rect 10796 29016 10824 29260
rect 10870 29248 10876 29300
rect 10928 29248 10934 29300
rect 11514 29248 11520 29300
rect 11572 29248 11578 29300
rect 11790 29248 11796 29300
rect 11848 29248 11854 29300
rect 12158 29248 12164 29300
rect 12216 29288 12222 29300
rect 12216 29260 12480 29288
rect 12216 29248 12222 29260
rect 10888 29220 10916 29248
rect 11808 29220 11836 29248
rect 10888 29192 11376 29220
rect 11146 29112 11152 29164
rect 11204 29112 11210 29164
rect 11348 29161 11376 29192
rect 11716 29192 11836 29220
rect 11716 29161 11744 29192
rect 11882 29180 11888 29232
rect 11940 29220 11946 29232
rect 12250 29220 12256 29232
rect 11940 29192 12256 29220
rect 11940 29180 11946 29192
rect 12250 29180 12256 29192
rect 12308 29180 12314 29232
rect 12342 29180 12348 29232
rect 12400 29180 12406 29232
rect 11333 29155 11391 29161
rect 11333 29121 11345 29155
rect 11379 29121 11391 29155
rect 11333 29115 11391 29121
rect 11701 29155 11759 29161
rect 11701 29121 11713 29155
rect 11747 29121 11759 29155
rect 11701 29115 11759 29121
rect 11790 29112 11796 29164
rect 11848 29112 11854 29164
rect 12023 29155 12081 29161
rect 12023 29121 12035 29155
rect 12069 29152 12081 29155
rect 12360 29152 12388 29180
rect 12452 29161 12480 29260
rect 12544 29260 12756 29288
rect 12069 29124 12388 29152
rect 12437 29155 12495 29161
rect 12069 29121 12081 29124
rect 12023 29115 12081 29121
rect 12437 29121 12449 29155
rect 12483 29121 12495 29155
rect 12437 29115 12495 29121
rect 11241 29087 11299 29093
rect 11241 29053 11253 29087
rect 11287 29084 11299 29087
rect 11808 29084 11836 29112
rect 11287 29056 11836 29084
rect 12161 29087 12219 29093
rect 11287 29053 11299 29056
rect 11241 29047 11299 29053
rect 12161 29053 12173 29087
rect 12207 29084 12219 29087
rect 12544 29084 12572 29260
rect 12728 29229 12756 29260
rect 12802 29248 12808 29300
rect 12860 29288 12866 29300
rect 13081 29291 13139 29297
rect 13081 29288 13093 29291
rect 12860 29260 13093 29288
rect 12860 29248 12866 29260
rect 13081 29257 13093 29260
rect 13127 29257 13139 29291
rect 13081 29251 13139 29257
rect 13446 29248 13452 29300
rect 13504 29248 13510 29300
rect 14182 29248 14188 29300
rect 14240 29248 14246 29300
rect 15930 29248 15936 29300
rect 15988 29248 15994 29300
rect 21177 29291 21235 29297
rect 21177 29257 21189 29291
rect 21223 29257 21235 29291
rect 21177 29251 21235 29257
rect 24397 29291 24455 29297
rect 24397 29257 24409 29291
rect 24443 29257 24455 29291
rect 26050 29288 26056 29300
rect 24397 29251 24455 29257
rect 24504 29260 26056 29288
rect 12713 29223 12771 29229
rect 12713 29189 12725 29223
rect 12759 29189 12771 29223
rect 13354 29220 13360 29232
rect 12713 29183 12771 29189
rect 12820 29192 13360 29220
rect 12820 29161 12848 29192
rect 13354 29180 13360 29192
rect 13412 29180 13418 29232
rect 12621 29155 12679 29161
rect 12621 29121 12633 29155
rect 12667 29152 12679 29155
rect 12805 29155 12863 29161
rect 12667 29124 12756 29152
rect 12667 29121 12679 29124
rect 12621 29115 12679 29121
rect 12207 29056 12572 29084
rect 12728 29084 12756 29124
rect 12805 29121 12817 29155
rect 12851 29121 12863 29155
rect 12805 29115 12863 29121
rect 13265 29155 13323 29161
rect 13265 29121 13277 29155
rect 13311 29152 13323 29155
rect 13464 29152 13492 29248
rect 13311 29124 13492 29152
rect 13311 29121 13323 29124
rect 13265 29115 13323 29121
rect 13354 29084 13360 29096
rect 12728 29056 13360 29084
rect 12207 29053 12219 29056
rect 12161 29047 12219 29053
rect 12176 29016 12204 29047
rect 13354 29044 13360 29056
rect 13412 29044 13418 29096
rect 13449 29087 13507 29093
rect 13449 29053 13461 29087
rect 13495 29084 13507 29087
rect 13814 29084 13820 29096
rect 13495 29056 13820 29084
rect 13495 29053 13507 29056
rect 13449 29047 13507 29053
rect 13814 29044 13820 29056
rect 13872 29044 13878 29096
rect 14200 29084 14228 29248
rect 15948 29220 15976 29248
rect 15856 29192 15976 29220
rect 18509 29223 18567 29229
rect 15856 29161 15884 29192
rect 18509 29189 18521 29223
rect 18555 29220 18567 29223
rect 20898 29220 20904 29232
rect 18555 29192 20904 29220
rect 18555 29189 18567 29192
rect 18509 29183 18567 29189
rect 20898 29180 20904 29192
rect 20956 29180 20962 29232
rect 15841 29155 15899 29161
rect 15841 29121 15853 29155
rect 15887 29121 15899 29155
rect 15841 29115 15899 29121
rect 15930 29112 15936 29164
rect 15988 29112 15994 29164
rect 16114 29112 16120 29164
rect 16172 29112 16178 29164
rect 17862 29112 17868 29164
rect 17920 29112 17926 29164
rect 17954 29112 17960 29164
rect 18012 29112 18018 29164
rect 18138 29112 18144 29164
rect 18196 29112 18202 29164
rect 19518 29112 19524 29164
rect 19576 29152 19582 29164
rect 20809 29155 20867 29161
rect 20809 29152 20821 29155
rect 19576 29124 20821 29152
rect 19576 29112 19582 29124
rect 20809 29121 20821 29124
rect 20855 29121 20867 29155
rect 21192 29152 21220 29251
rect 21266 29180 21272 29232
rect 21324 29180 21330 29232
rect 21450 29180 21456 29232
rect 21508 29229 21514 29232
rect 21508 29223 21527 29229
rect 21515 29189 21527 29223
rect 24412 29220 24440 29251
rect 21508 29183 21527 29189
rect 21560 29192 24440 29220
rect 21508 29180 21514 29183
rect 21468 29152 21496 29180
rect 21192 29124 21496 29152
rect 20809 29115 20867 29121
rect 20901 29087 20959 29093
rect 14200 29056 20852 29084
rect 20824 29028 20852 29056
rect 20901 29053 20913 29087
rect 20947 29084 20959 29087
rect 21560 29084 21588 29192
rect 21726 29112 21732 29164
rect 21784 29152 21790 29164
rect 22005 29155 22063 29161
rect 22005 29152 22017 29155
rect 21784 29124 22017 29152
rect 21784 29112 21790 29124
rect 22005 29121 22017 29124
rect 22051 29121 22063 29155
rect 22005 29115 22063 29121
rect 23937 29155 23995 29161
rect 23937 29121 23949 29155
rect 23983 29121 23995 29155
rect 24504 29152 24532 29260
rect 26050 29248 26056 29260
rect 26108 29248 26114 29300
rect 26329 29291 26387 29297
rect 26329 29257 26341 29291
rect 26375 29288 26387 29291
rect 26786 29288 26792 29300
rect 26375 29260 26792 29288
rect 26375 29257 26387 29260
rect 26329 29251 26387 29257
rect 26786 29248 26792 29260
rect 26844 29288 26850 29300
rect 27522 29288 27528 29300
rect 26844 29260 27528 29288
rect 26844 29248 26850 29260
rect 27522 29248 27528 29260
rect 27580 29248 27586 29300
rect 27801 29291 27859 29297
rect 27801 29257 27813 29291
rect 27847 29288 27859 29291
rect 27890 29288 27896 29300
rect 27847 29260 27896 29288
rect 27847 29257 27859 29260
rect 27801 29251 27859 29257
rect 27890 29248 27896 29260
rect 27948 29248 27954 29300
rect 28258 29248 28264 29300
rect 28316 29248 28322 29300
rect 28353 29291 28411 29297
rect 28353 29257 28365 29291
rect 28399 29288 28411 29291
rect 33042 29288 33048 29300
rect 28399 29260 33048 29288
rect 28399 29257 28411 29260
rect 28353 29251 28411 29257
rect 26418 29220 26424 29232
rect 25976 29192 26424 29220
rect 25976 29161 26004 29192
rect 26418 29180 26424 29192
rect 26476 29220 26482 29232
rect 31389 29223 31447 29229
rect 31389 29220 31401 29223
rect 26476 29192 28120 29220
rect 26476 29180 26482 29192
rect 23937 29115 23995 29121
rect 24044 29124 24532 29152
rect 24765 29155 24823 29161
rect 20947 29056 21588 29084
rect 20947 29053 20959 29056
rect 20901 29047 20959 29053
rect 21910 29044 21916 29096
rect 21968 29044 21974 29096
rect 10796 28988 12204 29016
rect 7929 28979 7987 28985
rect 12250 28976 12256 29028
rect 12308 29016 12314 29028
rect 12802 29016 12808 29028
rect 12308 28988 12808 29016
rect 12308 28976 12314 28988
rect 12802 28976 12808 28988
rect 12860 28976 12866 29028
rect 12989 29019 13047 29025
rect 12989 28985 13001 29019
rect 13035 29016 13047 29019
rect 15102 29016 15108 29028
rect 13035 28988 15108 29016
rect 13035 28985 13047 28988
rect 12989 28979 13047 28985
rect 15102 28976 15108 28988
rect 15160 28976 15166 29028
rect 16117 29019 16175 29025
rect 16117 28985 16129 29019
rect 16163 29016 16175 29019
rect 17126 29016 17132 29028
rect 16163 28988 17132 29016
rect 16163 28985 16175 28988
rect 16117 28979 16175 28985
rect 17126 28976 17132 28988
rect 17184 28976 17190 29028
rect 19426 28976 19432 29028
rect 19484 29016 19490 29028
rect 19886 29016 19892 29028
rect 19484 28988 19892 29016
rect 19484 28976 19490 28988
rect 19886 28976 19892 28988
rect 19944 28976 19950 29028
rect 20806 28976 20812 29028
rect 20864 29016 20870 29028
rect 20990 29016 20996 29028
rect 20864 28988 20996 29016
rect 20864 28976 20870 28988
rect 20990 28976 20996 28988
rect 21048 28976 21054 29028
rect 21637 29019 21695 29025
rect 21637 28985 21649 29019
rect 21683 29016 21695 29019
rect 22094 29016 22100 29028
rect 21683 28988 22100 29016
rect 21683 28985 21695 28988
rect 21637 28979 21695 28985
rect 22094 28976 22100 28988
rect 22152 28976 22158 29028
rect 23382 28976 23388 29028
rect 23440 29016 23446 29028
rect 23952 29016 23980 29115
rect 24044 29093 24072 29124
rect 24765 29121 24777 29155
rect 24811 29121 24823 29155
rect 24765 29115 24823 29121
rect 25961 29155 26019 29161
rect 25961 29121 25973 29155
rect 26007 29121 26019 29155
rect 25961 29115 26019 29121
rect 24029 29087 24087 29093
rect 24029 29053 24041 29087
rect 24075 29053 24087 29087
rect 24029 29047 24087 29053
rect 24118 29044 24124 29096
rect 24176 29044 24182 29096
rect 24673 29087 24731 29093
rect 24673 29084 24685 29087
rect 24320 29056 24685 29084
rect 24136 29016 24164 29044
rect 24320 29025 24348 29056
rect 24673 29053 24685 29056
rect 24719 29053 24731 29087
rect 24673 29047 24731 29053
rect 23440 28988 24164 29016
rect 24305 29019 24363 29025
rect 23440 28976 23446 28988
rect 24305 28985 24317 29019
rect 24351 28985 24363 29019
rect 24780 29016 24808 29115
rect 26142 29112 26148 29164
rect 26200 29152 26206 29164
rect 26200 29124 26832 29152
rect 26200 29112 26206 29124
rect 26053 29087 26111 29093
rect 26053 29053 26065 29087
rect 26099 29084 26111 29087
rect 26234 29084 26240 29096
rect 26099 29056 26240 29084
rect 26099 29053 26111 29056
rect 26053 29047 26111 29053
rect 26234 29044 26240 29056
rect 26292 29044 26298 29096
rect 26804 29084 26832 29124
rect 26878 29112 26884 29164
rect 26936 29152 26942 29164
rect 27157 29155 27215 29161
rect 27157 29152 27169 29155
rect 26936 29124 27169 29152
rect 26936 29112 26942 29124
rect 27157 29121 27169 29124
rect 27203 29121 27215 29155
rect 27157 29115 27215 29121
rect 27433 29155 27491 29161
rect 27433 29121 27445 29155
rect 27479 29121 27491 29155
rect 27433 29115 27491 29121
rect 27341 29087 27399 29093
rect 27341 29084 27353 29087
rect 26804 29056 27353 29084
rect 27341 29053 27353 29056
rect 27387 29053 27399 29087
rect 27341 29047 27399 29053
rect 26973 29019 27031 29025
rect 26973 29016 26985 29019
rect 24780 28988 26985 29016
rect 24305 28979 24363 28985
rect 26973 28985 26985 28988
rect 27019 28985 27031 29019
rect 27448 29016 27476 29115
rect 27522 29112 27528 29164
rect 27580 29112 27586 29164
rect 27614 29112 27620 29164
rect 27672 29152 27678 29164
rect 27709 29155 27767 29161
rect 27709 29152 27721 29155
rect 27672 29124 27721 29152
rect 27672 29112 27678 29124
rect 27709 29121 27721 29124
rect 27755 29121 27767 29155
rect 27709 29115 27767 29121
rect 28092 29093 28120 29192
rect 28467 29192 31401 29220
rect 28467 29161 28495 29192
rect 31389 29189 31401 29192
rect 31435 29189 31447 29223
rect 31389 29183 31447 29189
rect 28445 29155 28503 29161
rect 28445 29121 28457 29155
rect 28491 29121 28503 29155
rect 28445 29115 28503 29121
rect 28537 29155 28595 29161
rect 28537 29121 28549 29155
rect 28583 29121 28595 29155
rect 28537 29115 28595 29121
rect 27985 29087 28043 29093
rect 27985 29053 27997 29087
rect 28031 29053 28043 29087
rect 27985 29047 28043 29053
rect 28077 29087 28135 29093
rect 28077 29053 28089 29087
rect 28123 29084 28135 29087
rect 28558 29084 28586 29115
rect 28626 29112 28632 29164
rect 28684 29152 28690 29164
rect 28721 29155 28779 29161
rect 28721 29152 28733 29155
rect 28684 29124 28733 29152
rect 28684 29112 28690 29124
rect 28721 29121 28733 29124
rect 28767 29121 28779 29155
rect 28721 29115 28779 29121
rect 28994 29112 29000 29164
rect 29052 29112 29058 29164
rect 29457 29155 29515 29161
rect 29457 29121 29469 29155
rect 29503 29152 29515 29155
rect 29638 29152 29644 29164
rect 29503 29124 29644 29152
rect 29503 29121 29515 29124
rect 29457 29115 29515 29121
rect 29638 29112 29644 29124
rect 29696 29112 29702 29164
rect 30006 29112 30012 29164
rect 30064 29112 30070 29164
rect 30098 29112 30104 29164
rect 30156 29152 30162 29164
rect 31297 29155 31355 29161
rect 31297 29152 31309 29155
rect 30156 29124 31309 29152
rect 30156 29112 30162 29124
rect 31297 29121 31309 29124
rect 31343 29121 31355 29155
rect 31297 29115 31355 29121
rect 31481 29155 31539 29161
rect 31481 29121 31493 29155
rect 31527 29152 31539 29155
rect 31938 29152 31944 29164
rect 31527 29124 31944 29152
rect 31527 29121 31539 29124
rect 31481 29115 31539 29121
rect 31938 29112 31944 29124
rect 31996 29112 32002 29164
rect 32140 29161 32168 29260
rect 33042 29248 33048 29260
rect 33100 29248 33106 29300
rect 34701 29291 34759 29297
rect 34701 29257 34713 29291
rect 34747 29288 34759 29291
rect 36354 29288 36360 29300
rect 34747 29260 36360 29288
rect 34747 29257 34759 29260
rect 34701 29251 34759 29257
rect 36354 29248 36360 29260
rect 36412 29248 36418 29300
rect 33413 29223 33471 29229
rect 32416 29192 33364 29220
rect 32125 29155 32183 29161
rect 32125 29121 32137 29155
rect 32171 29121 32183 29155
rect 32125 29115 32183 29121
rect 28123 29056 28586 29084
rect 29365 29087 29423 29093
rect 28123 29053 28135 29056
rect 28077 29047 28135 29053
rect 29365 29053 29377 29087
rect 29411 29084 29423 29087
rect 29917 29087 29975 29093
rect 29917 29084 29929 29087
rect 29411 29056 29929 29084
rect 29411 29053 29423 29056
rect 29365 29047 29423 29053
rect 29917 29053 29929 29056
rect 29963 29053 29975 29087
rect 29917 29047 29975 29053
rect 30193 29087 30251 29093
rect 30193 29053 30205 29087
rect 30239 29053 30251 29087
rect 30193 29047 30251 29053
rect 26973 28979 27031 28985
rect 27080 28988 27476 29016
rect 4706 28908 4712 28960
rect 4764 28908 4770 28960
rect 6178 28908 6184 28960
rect 6236 28908 6242 28960
rect 18506 28908 18512 28960
rect 18564 28908 18570 28960
rect 21266 28908 21272 28960
rect 21324 28948 21330 28960
rect 21453 28951 21511 28957
rect 21453 28948 21465 28951
rect 21324 28920 21465 28948
rect 21324 28908 21330 28920
rect 21453 28917 21465 28920
rect 21499 28917 21511 28951
rect 21453 28911 21511 28917
rect 22278 28908 22284 28960
rect 22336 28908 22342 28960
rect 25406 28908 25412 28960
rect 25464 28948 25470 28960
rect 27080 28948 27108 28988
rect 25464 28920 27108 28948
rect 27448 28948 27476 28988
rect 27522 28976 27528 29028
rect 27580 29016 27586 29028
rect 28000 29016 28028 29047
rect 27580 28988 28028 29016
rect 27580 28976 27586 28988
rect 28258 28976 28264 29028
rect 28316 29016 28322 29028
rect 28534 29016 28540 29028
rect 28316 28988 28540 29016
rect 28316 28976 28322 28988
rect 28534 28976 28540 28988
rect 28592 28976 28598 29028
rect 28721 29019 28779 29025
rect 28721 28985 28733 29019
rect 28767 29016 28779 29019
rect 29380 29016 29408 29047
rect 28767 28988 29408 29016
rect 29641 29019 29699 29025
rect 28767 28985 28779 28988
rect 28721 28979 28779 28985
rect 29641 28985 29653 29019
rect 29687 29016 29699 29019
rect 30208 29016 30236 29047
rect 31662 29044 31668 29096
rect 31720 29084 31726 29096
rect 32217 29087 32275 29093
rect 32217 29084 32229 29087
rect 31720 29056 32229 29084
rect 31720 29044 31726 29056
rect 32217 29053 32229 29056
rect 32263 29053 32275 29087
rect 32217 29047 32275 29053
rect 29687 28988 30236 29016
rect 29687 28985 29699 28988
rect 29641 28979 29699 28985
rect 31018 28976 31024 29028
rect 31076 29016 31082 29028
rect 32416 29016 32444 29192
rect 32861 29155 32919 29161
rect 32861 29152 32873 29155
rect 32508 29124 32873 29152
rect 32508 29025 32536 29124
rect 32861 29121 32873 29124
rect 32907 29121 32919 29155
rect 32861 29115 32919 29121
rect 33134 29112 33140 29164
rect 33192 29112 33198 29164
rect 33336 29161 33364 29192
rect 33413 29189 33425 29223
rect 33459 29220 33471 29223
rect 34974 29220 34980 29232
rect 33459 29192 34008 29220
rect 33459 29189 33471 29192
rect 33413 29183 33471 29189
rect 33321 29155 33379 29161
rect 33321 29121 33333 29155
rect 33367 29121 33379 29155
rect 33321 29115 33379 29121
rect 33502 29112 33508 29164
rect 33560 29112 33566 29164
rect 33980 29161 34008 29192
rect 34348 29192 34980 29220
rect 33965 29155 34023 29161
rect 33965 29121 33977 29155
rect 34011 29121 34023 29155
rect 33965 29115 34023 29121
rect 34146 29112 34152 29164
rect 34204 29112 34210 29164
rect 34250 29155 34308 29161
rect 34250 29121 34262 29155
rect 34296 29152 34308 29155
rect 34348 29152 34376 29192
rect 34974 29180 34980 29192
rect 35032 29180 35038 29232
rect 35345 29223 35403 29229
rect 35345 29189 35357 29223
rect 35391 29220 35403 29223
rect 36265 29223 36323 29229
rect 36265 29220 36277 29223
rect 35391 29192 36277 29220
rect 35391 29189 35403 29192
rect 35345 29183 35403 29189
rect 36265 29189 36277 29192
rect 36311 29189 36323 29223
rect 36265 29183 36323 29189
rect 34296 29124 34376 29152
rect 34296 29121 34308 29124
rect 34250 29115 34308 29121
rect 34422 29112 34428 29164
rect 34480 29152 34486 29164
rect 34517 29155 34575 29161
rect 34517 29152 34529 29155
rect 34480 29124 34529 29152
rect 34480 29112 34486 29124
rect 34517 29121 34529 29124
rect 34563 29152 34575 29155
rect 34790 29152 34796 29164
rect 34563 29124 34796 29152
rect 34563 29121 34575 29124
rect 34517 29115 34575 29121
rect 34790 29112 34796 29124
rect 34848 29112 34854 29164
rect 35158 29112 35164 29164
rect 35216 29152 35222 29164
rect 35526 29152 35532 29164
rect 35216 29124 35532 29152
rect 35216 29112 35222 29124
rect 35526 29112 35532 29124
rect 35584 29112 35590 29164
rect 35621 29155 35679 29161
rect 35621 29121 35633 29155
rect 35667 29121 35679 29155
rect 35621 29115 35679 29121
rect 33229 29087 33287 29093
rect 33229 29053 33241 29087
rect 33275 29084 33287 29087
rect 34330 29084 34336 29096
rect 33275 29056 34336 29084
rect 33275 29053 33287 29056
rect 33229 29047 33287 29053
rect 34330 29044 34336 29056
rect 34388 29044 34394 29096
rect 35636 29084 35664 29115
rect 35986 29112 35992 29164
rect 36044 29112 36050 29164
rect 36170 29112 36176 29164
rect 36228 29112 36234 29164
rect 36354 29112 36360 29164
rect 36412 29112 36418 29164
rect 35452 29056 35664 29084
rect 36004 29084 36032 29112
rect 36081 29087 36139 29093
rect 36081 29084 36093 29087
rect 36004 29056 36093 29084
rect 35452 29028 35480 29056
rect 36081 29053 36093 29056
rect 36127 29084 36139 29087
rect 36722 29084 36728 29096
rect 36127 29056 36728 29084
rect 36127 29053 36139 29056
rect 36081 29047 36139 29053
rect 36722 29044 36728 29056
rect 36780 29044 36786 29096
rect 31076 28988 32444 29016
rect 32493 29019 32551 29025
rect 31076 28976 31082 28988
rect 32493 28985 32505 29019
rect 32539 28985 32551 29019
rect 32493 28979 32551 28985
rect 35434 28976 35440 29028
rect 35492 28976 35498 29028
rect 28074 28948 28080 28960
rect 27448 28920 28080 28948
rect 25464 28908 25470 28920
rect 28074 28908 28080 28920
rect 28132 28908 28138 28960
rect 28810 28908 28816 28960
rect 28868 28948 28874 28960
rect 29733 28951 29791 28957
rect 29733 28948 29745 28951
rect 28868 28920 29745 28948
rect 28868 28908 28874 28920
rect 29733 28917 29745 28920
rect 29779 28917 29791 28951
rect 29733 28911 29791 28917
rect 32030 28908 32036 28960
rect 32088 28948 32094 28960
rect 32125 28951 32183 28957
rect 32125 28948 32137 28951
rect 32088 28920 32137 28948
rect 32088 28908 32094 28920
rect 32125 28917 32137 28920
rect 32171 28917 32183 28951
rect 32125 28911 32183 28917
rect 34422 28908 34428 28960
rect 34480 28948 34486 28960
rect 35713 28951 35771 28957
rect 35713 28948 35725 28951
rect 34480 28920 35725 28948
rect 34480 28908 34486 28920
rect 35713 28917 35725 28920
rect 35759 28917 35771 28951
rect 35713 28911 35771 28917
rect 35802 28908 35808 28960
rect 35860 28948 35866 28960
rect 36722 28948 36728 28960
rect 35860 28920 36728 28948
rect 35860 28908 35866 28920
rect 36722 28908 36728 28920
rect 36780 28908 36786 28960
rect 1104 28858 38272 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38272 28858
rect 1104 28784 38272 28806
rect 3510 28704 3516 28756
rect 3568 28744 3574 28756
rect 3605 28747 3663 28753
rect 3605 28744 3617 28747
rect 3568 28716 3617 28744
rect 3568 28704 3574 28716
rect 3605 28713 3617 28716
rect 3651 28713 3663 28747
rect 3605 28707 3663 28713
rect 1762 28568 1768 28620
rect 1820 28608 1826 28620
rect 1857 28611 1915 28617
rect 1857 28608 1869 28611
rect 1820 28580 1869 28608
rect 1820 28568 1826 28580
rect 1857 28577 1869 28580
rect 1903 28608 1915 28611
rect 2130 28608 2136 28620
rect 1903 28580 2136 28608
rect 1903 28577 1915 28580
rect 1857 28571 1915 28577
rect 2130 28568 2136 28580
rect 2188 28568 2194 28620
rect 3620 28608 3648 28707
rect 4614 28704 4620 28756
rect 4672 28704 4678 28756
rect 5258 28704 5264 28756
rect 5316 28704 5322 28756
rect 6822 28704 6828 28756
rect 6880 28704 6886 28756
rect 15933 28747 15991 28753
rect 15933 28713 15945 28747
rect 15979 28744 15991 28747
rect 16114 28744 16120 28756
rect 15979 28716 16120 28744
rect 15979 28713 15991 28716
rect 15933 28707 15991 28713
rect 16114 28704 16120 28716
rect 16172 28704 16178 28756
rect 17589 28747 17647 28753
rect 17589 28713 17601 28747
rect 17635 28744 17647 28747
rect 21726 28744 21732 28756
rect 17635 28716 21732 28744
rect 17635 28713 17647 28716
rect 17589 28707 17647 28713
rect 21726 28704 21732 28716
rect 21784 28704 21790 28756
rect 22186 28704 22192 28756
rect 22244 28704 22250 28756
rect 24854 28704 24860 28756
rect 24912 28744 24918 28756
rect 26142 28744 26148 28756
rect 24912 28716 26148 28744
rect 24912 28704 24918 28716
rect 26142 28704 26148 28716
rect 26200 28704 26206 28756
rect 27157 28747 27215 28753
rect 27157 28713 27169 28747
rect 27203 28744 27215 28747
rect 27430 28744 27436 28756
rect 27203 28716 27436 28744
rect 27203 28713 27215 28716
rect 27157 28707 27215 28713
rect 27430 28704 27436 28716
rect 27488 28704 27494 28756
rect 27893 28747 27951 28753
rect 27893 28713 27905 28747
rect 27939 28744 27951 28747
rect 28166 28744 28172 28756
rect 27939 28716 28172 28744
rect 27939 28713 27951 28716
rect 27893 28707 27951 28713
rect 28166 28704 28172 28716
rect 28224 28744 28230 28756
rect 28810 28744 28816 28756
rect 28224 28716 28816 28744
rect 28224 28704 28230 28716
rect 28810 28704 28816 28716
rect 28868 28704 28874 28756
rect 29086 28704 29092 28756
rect 29144 28744 29150 28756
rect 29549 28747 29607 28753
rect 29549 28744 29561 28747
rect 29144 28716 29561 28744
rect 29144 28704 29150 28716
rect 29549 28713 29561 28716
rect 29595 28713 29607 28747
rect 29549 28707 29607 28713
rect 29917 28747 29975 28753
rect 29917 28713 29929 28747
rect 29963 28713 29975 28747
rect 29917 28707 29975 28713
rect 30944 28716 31432 28744
rect 3789 28611 3847 28617
rect 3789 28608 3801 28611
rect 3620 28580 3801 28608
rect 3789 28577 3801 28580
rect 3835 28577 3847 28611
rect 5276 28608 5304 28704
rect 6733 28679 6791 28685
rect 6733 28645 6745 28679
rect 6779 28676 6791 28679
rect 6779 28648 7328 28676
rect 6779 28645 6791 28648
rect 6733 28639 6791 28645
rect 3789 28571 3847 28577
rect 4816 28580 5304 28608
rect 5721 28611 5779 28617
rect 4816 28549 4844 28580
rect 5721 28577 5733 28611
rect 5767 28608 5779 28611
rect 5905 28611 5963 28617
rect 5767 28580 5856 28608
rect 5767 28577 5779 28580
rect 5721 28571 5779 28577
rect 4433 28543 4491 28549
rect 4433 28509 4445 28543
rect 4479 28540 4491 28543
rect 4525 28543 4583 28549
rect 4525 28540 4537 28543
rect 4479 28512 4537 28540
rect 4479 28509 4491 28512
rect 4433 28503 4491 28509
rect 4525 28509 4537 28512
rect 4571 28509 4583 28543
rect 4525 28503 4583 28509
rect 4801 28543 4859 28549
rect 4801 28509 4813 28543
rect 4847 28509 4859 28543
rect 4801 28503 4859 28509
rect 4982 28500 4988 28552
rect 5040 28540 5046 28552
rect 5261 28543 5319 28549
rect 5261 28540 5273 28543
rect 5040 28512 5273 28540
rect 5040 28500 5046 28512
rect 5261 28509 5273 28512
rect 5307 28509 5319 28543
rect 5261 28503 5319 28509
rect 5353 28543 5411 28549
rect 5353 28509 5365 28543
rect 5399 28509 5411 28543
rect 5353 28503 5411 28509
rect 2133 28475 2191 28481
rect 2133 28441 2145 28475
rect 2179 28441 2191 28475
rect 2133 28435 2191 28441
rect 2148 28404 2176 28435
rect 2774 28432 2780 28484
rect 2832 28432 2838 28484
rect 3528 28444 5028 28472
rect 3528 28404 3556 28444
rect 5000 28413 5028 28444
rect 2148 28376 3556 28404
rect 4985 28407 5043 28413
rect 4985 28373 4997 28407
rect 5031 28373 5043 28407
rect 5368 28404 5396 28503
rect 5534 28500 5540 28552
rect 5592 28500 5598 28552
rect 5629 28543 5687 28549
rect 5629 28509 5641 28543
rect 5675 28540 5687 28543
rect 5828 28540 5856 28580
rect 5905 28577 5917 28611
rect 5951 28608 5963 28611
rect 6822 28608 6828 28620
rect 5951 28580 6224 28608
rect 5951 28577 5963 28580
rect 5905 28571 5963 28577
rect 6196 28552 6224 28580
rect 6288 28580 6828 28608
rect 5675 28512 5856 28540
rect 5675 28509 5687 28512
rect 5629 28503 5687 28509
rect 5828 28484 5856 28512
rect 5997 28543 6055 28549
rect 5997 28509 6009 28543
rect 6043 28509 6055 28543
rect 5997 28503 6055 28509
rect 5810 28432 5816 28484
rect 5868 28432 5874 28484
rect 6012 28472 6040 28503
rect 6086 28500 6092 28552
rect 6144 28500 6150 28552
rect 6178 28500 6184 28552
rect 6236 28500 6242 28552
rect 6288 28472 6316 28580
rect 6822 28568 6828 28580
rect 6880 28608 6886 28620
rect 7300 28617 7328 28648
rect 17218 28636 17224 28688
rect 17276 28636 17282 28688
rect 17681 28679 17739 28685
rect 17681 28645 17693 28679
rect 17727 28676 17739 28679
rect 18046 28676 18052 28688
rect 17727 28648 18052 28676
rect 17727 28645 17739 28648
rect 17681 28639 17739 28645
rect 7101 28611 7159 28617
rect 7101 28608 7113 28611
rect 6880 28580 7113 28608
rect 6880 28568 6886 28580
rect 7101 28577 7113 28580
rect 7147 28577 7159 28611
rect 7101 28571 7159 28577
rect 7285 28611 7343 28617
rect 7285 28577 7297 28611
rect 7331 28577 7343 28611
rect 15565 28611 15623 28617
rect 15565 28608 15577 28611
rect 7285 28571 7343 28577
rect 15488 28580 15577 28608
rect 6362 28500 6368 28552
rect 6420 28540 6426 28552
rect 7009 28543 7067 28549
rect 7009 28540 7021 28543
rect 6420 28512 7021 28540
rect 6420 28500 6426 28512
rect 7009 28509 7021 28512
rect 7055 28509 7067 28543
rect 7009 28503 7067 28509
rect 7193 28543 7251 28549
rect 7193 28509 7205 28543
rect 7239 28540 7251 28543
rect 7374 28540 7380 28552
rect 7239 28512 7380 28540
rect 7239 28509 7251 28512
rect 7193 28503 7251 28509
rect 7374 28500 7380 28512
rect 7432 28500 7438 28552
rect 12710 28500 12716 28552
rect 12768 28540 12774 28552
rect 12989 28543 13047 28549
rect 12989 28540 13001 28543
rect 12768 28512 13001 28540
rect 12768 28500 12774 28512
rect 12989 28509 13001 28512
rect 13035 28509 13047 28543
rect 12989 28503 13047 28509
rect 15102 28500 15108 28552
rect 15160 28540 15166 28552
rect 15488 28549 15516 28580
rect 15565 28577 15577 28580
rect 15611 28608 15623 28611
rect 17236 28608 17264 28636
rect 15611 28580 17264 28608
rect 15611 28577 15623 28580
rect 15565 28571 15623 28577
rect 16040 28549 16068 28580
rect 17310 28568 17316 28620
rect 17368 28568 17374 28620
rect 15289 28543 15347 28549
rect 15289 28540 15301 28543
rect 15160 28512 15301 28540
rect 15160 28500 15166 28512
rect 15289 28509 15301 28512
rect 15335 28509 15347 28543
rect 15289 28503 15347 28509
rect 15473 28543 15531 28549
rect 15473 28509 15485 28543
rect 15519 28509 15531 28543
rect 15473 28503 15531 28509
rect 15749 28543 15807 28549
rect 15749 28509 15761 28543
rect 15795 28509 15807 28543
rect 15749 28503 15807 28509
rect 16025 28543 16083 28549
rect 16025 28509 16037 28543
rect 16071 28509 16083 28543
rect 16025 28503 16083 28509
rect 16117 28543 16175 28549
rect 16117 28509 16129 28543
rect 16163 28540 16175 28543
rect 16301 28543 16359 28549
rect 16301 28540 16313 28543
rect 16163 28512 16313 28540
rect 16163 28509 16175 28512
rect 16117 28503 16175 28509
rect 16301 28509 16313 28512
rect 16347 28509 16359 28543
rect 16301 28503 16359 28509
rect 16485 28543 16543 28549
rect 16485 28509 16497 28543
rect 16531 28509 16543 28543
rect 16485 28503 16543 28509
rect 6012 28444 6316 28472
rect 6574 28475 6632 28481
rect 6574 28441 6586 28475
rect 6620 28472 6632 28475
rect 6730 28472 6736 28484
rect 6620 28444 6736 28472
rect 6620 28441 6632 28444
rect 6574 28435 6632 28441
rect 6730 28432 6736 28444
rect 6788 28432 6794 28484
rect 12805 28475 12863 28481
rect 12805 28441 12817 28475
rect 12851 28472 12863 28475
rect 12894 28472 12900 28484
rect 12851 28444 12900 28472
rect 12851 28441 12863 28444
rect 12805 28435 12863 28441
rect 12894 28432 12900 28444
rect 12952 28432 12958 28484
rect 15304 28472 15332 28503
rect 15764 28472 15792 28503
rect 16500 28472 16528 28503
rect 17126 28500 17132 28552
rect 17184 28500 17190 28552
rect 17221 28543 17279 28549
rect 17221 28509 17233 28543
rect 17267 28540 17279 28543
rect 17696 28540 17724 28639
rect 18046 28636 18052 28648
rect 18104 28636 18110 28688
rect 19794 28676 19800 28688
rect 18432 28648 19800 28676
rect 17770 28568 17776 28620
rect 17828 28568 17834 28620
rect 17267 28512 17724 28540
rect 18049 28543 18107 28549
rect 17267 28509 17279 28512
rect 17221 28503 17279 28509
rect 18049 28509 18061 28543
rect 18095 28540 18107 28543
rect 18432 28540 18460 28648
rect 19794 28636 19800 28648
rect 19852 28636 19858 28688
rect 22094 28636 22100 28688
rect 22152 28676 22158 28688
rect 22649 28679 22707 28685
rect 22649 28676 22661 28679
rect 22152 28648 22661 28676
rect 22152 28636 22158 28648
rect 22649 28645 22661 28648
rect 22695 28645 22707 28679
rect 22649 28639 22707 28645
rect 23474 28636 23480 28688
rect 23532 28676 23538 28688
rect 24946 28676 24952 28688
rect 23532 28648 24952 28676
rect 23532 28636 23538 28648
rect 24946 28636 24952 28648
rect 25004 28636 25010 28688
rect 29932 28676 29960 28707
rect 30944 28676 30972 28716
rect 29932 28648 30972 28676
rect 18616 28580 19472 28608
rect 18095 28512 18460 28540
rect 18095 28509 18107 28512
rect 18049 28503 18107 28509
rect 18506 28500 18512 28552
rect 18564 28500 18570 28552
rect 15304 28444 16528 28472
rect 17144 28472 17172 28500
rect 18616 28472 18644 28580
rect 19444 28549 19472 28580
rect 19536 28580 20116 28608
rect 19536 28549 19564 28580
rect 18877 28543 18935 28549
rect 18877 28509 18889 28543
rect 18923 28540 18935 28543
rect 19429 28543 19487 28549
rect 18923 28512 19012 28540
rect 18923 28509 18935 28512
rect 18877 28503 18935 28509
rect 18984 28484 19012 28512
rect 19429 28509 19441 28543
rect 19475 28509 19487 28543
rect 19429 28503 19487 28509
rect 19521 28543 19579 28549
rect 19521 28509 19533 28543
rect 19567 28509 19579 28543
rect 19521 28503 19579 28509
rect 19705 28543 19763 28549
rect 19705 28509 19717 28543
rect 19751 28509 19763 28543
rect 19705 28503 19763 28509
rect 17144 28444 18644 28472
rect 18966 28432 18972 28484
rect 19024 28432 19030 28484
rect 19058 28432 19064 28484
rect 19116 28472 19122 28484
rect 19720 28472 19748 28503
rect 19794 28500 19800 28552
rect 19852 28500 19858 28552
rect 19886 28500 19892 28552
rect 19944 28500 19950 28552
rect 19978 28500 19984 28552
rect 20036 28500 20042 28552
rect 20088 28549 20116 28580
rect 22112 28549 22140 28636
rect 22189 28611 22247 28617
rect 22189 28577 22201 28611
rect 22235 28608 22247 28611
rect 22278 28608 22284 28620
rect 22235 28580 22284 28608
rect 22235 28577 22247 28580
rect 22189 28571 22247 28577
rect 22278 28568 22284 28580
rect 22336 28608 22342 28620
rect 22833 28611 22891 28617
rect 22833 28608 22845 28611
rect 22336 28580 22845 28608
rect 22336 28568 22342 28580
rect 22833 28577 22845 28580
rect 22879 28577 22891 28611
rect 27249 28611 27307 28617
rect 27249 28608 27261 28611
rect 22833 28571 22891 28577
rect 24872 28580 27261 28608
rect 20073 28543 20131 28549
rect 20073 28509 20085 28543
rect 20119 28540 20131 28543
rect 22102 28543 22160 28549
rect 20119 28512 20392 28540
rect 20119 28509 20131 28512
rect 20073 28503 20131 28509
rect 19996 28472 20024 28500
rect 19116 28444 19380 28472
rect 19720 28444 20024 28472
rect 19116 28432 19122 28444
rect 5626 28404 5632 28416
rect 5368 28376 5632 28404
rect 4985 28367 5043 28373
rect 5626 28364 5632 28376
rect 5684 28364 5690 28416
rect 5721 28407 5779 28413
rect 5721 28373 5733 28407
rect 5767 28404 5779 28407
rect 6365 28407 6423 28413
rect 6365 28404 6377 28407
rect 5767 28376 6377 28404
rect 5767 28373 5779 28376
rect 5721 28367 5779 28373
rect 6365 28373 6377 28376
rect 6411 28373 6423 28407
rect 6365 28367 6423 28373
rect 6454 28364 6460 28416
rect 6512 28364 6518 28416
rect 13170 28364 13176 28416
rect 13228 28364 13234 28416
rect 15378 28364 15384 28416
rect 15436 28364 15442 28416
rect 16393 28407 16451 28413
rect 16393 28373 16405 28407
rect 16439 28404 16451 28407
rect 17954 28404 17960 28416
rect 16439 28376 17960 28404
rect 16439 28373 16451 28376
rect 16393 28367 16451 28373
rect 17954 28364 17960 28376
rect 18012 28364 18018 28416
rect 19242 28364 19248 28416
rect 19300 28364 19306 28416
rect 19352 28404 19380 28444
rect 20364 28416 20392 28512
rect 22102 28509 22114 28543
rect 22148 28509 22160 28543
rect 22557 28543 22615 28549
rect 22557 28540 22569 28543
rect 22102 28503 22160 28509
rect 22204 28512 22569 28540
rect 22204 28484 22232 28512
rect 22557 28509 22569 28512
rect 22603 28509 22615 28543
rect 22557 28503 22615 28509
rect 23842 28500 23848 28552
rect 23900 28540 23906 28552
rect 24673 28543 24731 28549
rect 24673 28540 24685 28543
rect 23900 28512 24685 28540
rect 23900 28500 23906 28512
rect 24673 28509 24685 28512
rect 24719 28509 24731 28543
rect 24673 28503 24731 28509
rect 24762 28500 24768 28552
rect 24820 28500 24826 28552
rect 24872 28549 24900 28580
rect 27249 28577 27261 28580
rect 27295 28577 27307 28611
rect 27249 28571 27307 28577
rect 30009 28611 30067 28617
rect 30009 28577 30021 28611
rect 30055 28608 30067 28611
rect 30098 28608 30104 28620
rect 30055 28580 30104 28608
rect 30055 28577 30067 28580
rect 30009 28571 30067 28577
rect 30098 28568 30104 28580
rect 30156 28568 30162 28620
rect 30834 28568 30840 28620
rect 30892 28568 30898 28620
rect 31404 28608 31432 28716
rect 31570 28704 31576 28756
rect 31628 28744 31634 28756
rect 31665 28747 31723 28753
rect 31665 28744 31677 28747
rect 31628 28716 31677 28744
rect 31628 28704 31634 28716
rect 31665 28713 31677 28716
rect 31711 28713 31723 28747
rect 31665 28707 31723 28713
rect 32030 28704 32036 28756
rect 32088 28704 32094 28756
rect 32490 28704 32496 28756
rect 32548 28744 32554 28756
rect 32769 28747 32827 28753
rect 32769 28744 32781 28747
rect 32548 28716 32781 28744
rect 32548 28704 32554 28716
rect 32769 28713 32781 28716
rect 32815 28713 32827 28747
rect 32769 28707 32827 28713
rect 33042 28704 33048 28756
rect 33100 28704 33106 28756
rect 35618 28704 35624 28756
rect 35676 28744 35682 28756
rect 36262 28744 36268 28756
rect 35676 28716 36268 28744
rect 35676 28704 35682 28716
rect 36262 28704 36268 28716
rect 36320 28704 36326 28756
rect 36354 28704 36360 28756
rect 36412 28744 36418 28756
rect 36449 28747 36507 28753
rect 36449 28744 36461 28747
rect 36412 28716 36461 28744
rect 36412 28704 36418 28716
rect 36449 28713 36461 28716
rect 36495 28713 36507 28747
rect 36449 28707 36507 28713
rect 36722 28704 36728 28756
rect 36780 28744 36786 28756
rect 36780 28716 36952 28744
rect 36780 28704 36786 28716
rect 31481 28679 31539 28685
rect 31481 28645 31493 28679
rect 31527 28676 31539 28679
rect 32048 28676 32076 28704
rect 31527 28648 32076 28676
rect 32585 28679 32643 28685
rect 31527 28645 31539 28648
rect 31481 28639 31539 28645
rect 32585 28645 32597 28679
rect 32631 28676 32643 28679
rect 33134 28676 33140 28688
rect 32631 28648 33140 28676
rect 32631 28645 32643 28648
rect 32585 28639 32643 28645
rect 32600 28608 32628 28639
rect 33134 28636 33140 28648
rect 33192 28636 33198 28688
rect 35434 28636 35440 28688
rect 35492 28636 35498 28688
rect 35526 28636 35532 28688
rect 35584 28676 35590 28688
rect 35713 28679 35771 28685
rect 35713 28676 35725 28679
rect 35584 28648 35725 28676
rect 35584 28636 35590 28648
rect 35713 28645 35725 28648
rect 35759 28645 35771 28679
rect 35713 28639 35771 28645
rect 36081 28679 36139 28685
rect 36081 28645 36093 28679
rect 36127 28676 36139 28679
rect 36127 28648 36492 28676
rect 36127 28645 36139 28648
rect 36081 28639 36139 28645
rect 31404 28580 32628 28608
rect 24857 28543 24915 28549
rect 24857 28509 24869 28543
rect 24903 28509 24915 28543
rect 24857 28503 24915 28509
rect 25041 28543 25099 28549
rect 25041 28509 25053 28543
rect 25087 28509 25099 28543
rect 25041 28503 25099 28509
rect 22186 28432 22192 28484
rect 22244 28432 22250 28484
rect 23014 28432 23020 28484
rect 23072 28472 23078 28484
rect 25056 28472 25084 28503
rect 26694 28500 26700 28552
rect 26752 28500 26758 28552
rect 26786 28500 26792 28552
rect 26844 28500 26850 28552
rect 26970 28500 26976 28552
rect 27028 28500 27034 28552
rect 27525 28543 27583 28549
rect 27525 28509 27537 28543
rect 27571 28509 27583 28543
rect 27525 28503 27583 28509
rect 27709 28543 27767 28549
rect 27709 28509 27721 28543
rect 27755 28540 27767 28543
rect 27798 28540 27804 28552
rect 27755 28512 27804 28540
rect 27755 28509 27767 28512
rect 27709 28503 27767 28509
rect 23072 28444 25084 28472
rect 27540 28472 27568 28503
rect 27798 28500 27804 28512
rect 27856 28500 27862 28552
rect 27985 28543 28043 28549
rect 27985 28509 27997 28543
rect 28031 28540 28043 28543
rect 28442 28540 28448 28552
rect 28031 28512 28448 28540
rect 28031 28509 28043 28512
rect 27985 28503 28043 28509
rect 28442 28500 28448 28512
rect 28500 28500 28506 28552
rect 29730 28500 29736 28552
rect 29788 28500 29794 28552
rect 30650 28500 30656 28552
rect 30708 28500 30714 28552
rect 30742 28500 30748 28552
rect 30800 28500 30806 28552
rect 30929 28543 30987 28549
rect 30929 28509 30941 28543
rect 30975 28542 30987 28543
rect 30975 28514 31064 28542
rect 30975 28509 30987 28514
rect 30929 28503 30987 28509
rect 30668 28472 30696 28500
rect 31036 28472 31064 28514
rect 31110 28500 31116 28552
rect 31168 28500 31174 28552
rect 31772 28549 31800 28580
rect 32766 28568 32772 28620
rect 32824 28608 32830 28620
rect 32861 28611 32919 28617
rect 32861 28608 32873 28611
rect 32824 28580 32873 28608
rect 32824 28568 32830 28580
rect 32861 28577 32873 28580
rect 32907 28608 32919 28611
rect 36262 28608 36268 28620
rect 32907 28580 36268 28608
rect 32907 28577 32919 28580
rect 32861 28571 32919 28577
rect 36262 28568 36268 28580
rect 36320 28568 36326 28620
rect 36464 28608 36492 28648
rect 36654 28648 36860 28676
rect 36654 28608 36682 28648
rect 36464 28580 36682 28608
rect 36722 28568 36728 28620
rect 36780 28568 36786 28620
rect 31297 28543 31355 28549
rect 31297 28509 31309 28543
rect 31343 28509 31355 28543
rect 31297 28503 31355 28509
rect 31573 28543 31631 28549
rect 31573 28509 31585 28543
rect 31619 28509 31631 28543
rect 31573 28503 31631 28509
rect 31757 28543 31815 28549
rect 31757 28509 31769 28543
rect 31803 28509 31815 28543
rect 31757 28503 31815 28509
rect 31312 28472 31340 28503
rect 27540 28444 28672 28472
rect 30668 28444 31340 28472
rect 23072 28432 23078 28444
rect 28644 28416 28672 28444
rect 19981 28407 20039 28413
rect 19981 28404 19993 28407
rect 19352 28376 19993 28404
rect 19981 28373 19993 28376
rect 20027 28373 20039 28407
rect 19981 28367 20039 28373
rect 20346 28364 20352 28416
rect 20404 28364 20410 28416
rect 22462 28364 22468 28416
rect 22520 28364 22526 28416
rect 22830 28364 22836 28416
rect 22888 28364 22894 28416
rect 24394 28364 24400 28416
rect 24452 28364 24458 28416
rect 26050 28364 26056 28416
rect 26108 28404 26114 28416
rect 27617 28407 27675 28413
rect 27617 28404 27629 28407
rect 26108 28376 27629 28404
rect 26108 28364 26114 28376
rect 27617 28373 27629 28376
rect 27663 28373 27675 28407
rect 27617 28367 27675 28373
rect 28626 28364 28632 28416
rect 28684 28364 28690 28416
rect 30926 28364 30932 28416
rect 30984 28404 30990 28416
rect 31588 28404 31616 28503
rect 32490 28500 32496 28552
rect 32548 28500 32554 28552
rect 32953 28543 33011 28549
rect 32953 28509 32965 28543
rect 32999 28540 33011 28543
rect 33042 28540 33048 28552
rect 32999 28512 33048 28540
rect 32999 28509 33011 28512
rect 32953 28503 33011 28509
rect 33042 28500 33048 28512
rect 33100 28500 33106 28552
rect 33229 28543 33287 28549
rect 33229 28509 33241 28543
rect 33275 28509 33287 28543
rect 33229 28503 33287 28509
rect 32508 28472 32536 28500
rect 33244 28472 33272 28503
rect 35802 28500 35808 28552
rect 35860 28500 35866 28552
rect 35894 28500 35900 28552
rect 35952 28500 35958 28552
rect 35986 28500 35992 28552
rect 36044 28500 36050 28552
rect 36173 28543 36231 28549
rect 36173 28518 36185 28543
rect 36096 28509 36185 28518
rect 36219 28509 36231 28543
rect 36280 28540 36308 28568
rect 36832 28549 36860 28648
rect 36924 28549 36952 28716
rect 36357 28543 36415 28549
rect 36357 28540 36369 28543
rect 36280 28512 36369 28540
rect 36096 28503 36231 28509
rect 36357 28509 36369 28512
rect 36403 28509 36415 28543
rect 36633 28543 36691 28549
rect 36633 28540 36645 28543
rect 36357 28503 36415 28509
rect 36556 28512 36645 28540
rect 32508 28444 33272 28472
rect 33318 28432 33324 28484
rect 33376 28472 33382 28484
rect 34422 28472 34428 28484
rect 33376 28444 34428 28472
rect 33376 28432 33382 28444
rect 34422 28432 34428 28444
rect 34480 28472 34486 28484
rect 35161 28475 35219 28481
rect 35161 28472 35173 28475
rect 34480 28444 35173 28472
rect 34480 28432 34486 28444
rect 35161 28441 35173 28444
rect 35207 28441 35219 28475
rect 35161 28435 35219 28441
rect 35250 28432 35256 28484
rect 35308 28472 35314 28484
rect 35618 28472 35624 28484
rect 35308 28444 35624 28472
rect 35308 28432 35314 28444
rect 35618 28432 35624 28444
rect 35676 28432 35682 28484
rect 35820 28472 35848 28500
rect 36096 28490 36215 28503
rect 36096 28472 36124 28490
rect 36556 28472 36584 28512
rect 36633 28509 36645 28512
rect 36679 28509 36691 28543
rect 36633 28503 36691 28509
rect 36817 28543 36875 28549
rect 36817 28509 36829 28543
rect 36863 28509 36875 28543
rect 36817 28503 36875 28509
rect 36909 28543 36967 28549
rect 36909 28509 36921 28543
rect 36955 28509 36967 28543
rect 36909 28503 36967 28509
rect 35820 28444 36124 28472
rect 36464 28444 36584 28472
rect 36832 28472 36860 28503
rect 37090 28500 37096 28552
rect 37148 28500 37154 28552
rect 37108 28472 37136 28500
rect 36832 28444 37136 28472
rect 36464 28416 36492 28444
rect 30984 28376 31616 28404
rect 30984 28364 30990 28376
rect 35894 28364 35900 28416
rect 35952 28404 35958 28416
rect 36446 28404 36452 28416
rect 35952 28376 36452 28404
rect 35952 28364 35958 28376
rect 36446 28364 36452 28376
rect 36504 28364 36510 28416
rect 1104 28314 38272 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 38272 28314
rect 1104 28240 38272 28262
rect 5810 28160 5816 28212
rect 5868 28200 5874 28212
rect 6457 28203 6515 28209
rect 6457 28200 6469 28203
rect 5868 28172 6469 28200
rect 5868 28160 5874 28172
rect 6457 28169 6469 28172
rect 6503 28169 6515 28203
rect 6457 28163 6515 28169
rect 9030 28160 9036 28212
rect 9088 28200 9094 28212
rect 12618 28200 12624 28212
rect 9088 28172 12624 28200
rect 9088 28160 9094 28172
rect 12618 28160 12624 28172
rect 12676 28160 12682 28212
rect 13170 28160 13176 28212
rect 13228 28160 13234 28212
rect 15378 28160 15384 28212
rect 15436 28160 15442 28212
rect 15749 28203 15807 28209
rect 15749 28169 15761 28203
rect 15795 28200 15807 28203
rect 15930 28200 15936 28212
rect 15795 28172 15936 28200
rect 15795 28169 15807 28172
rect 15749 28163 15807 28169
rect 15930 28160 15936 28172
rect 15988 28160 15994 28212
rect 17589 28203 17647 28209
rect 17589 28169 17601 28203
rect 17635 28200 17647 28203
rect 17770 28200 17776 28212
rect 17635 28172 17776 28200
rect 17635 28169 17647 28172
rect 17589 28163 17647 28169
rect 17770 28160 17776 28172
rect 17828 28160 17834 28212
rect 17862 28160 17868 28212
rect 17920 28200 17926 28212
rect 17920 28172 18184 28200
rect 17920 28160 17926 28172
rect 4706 28092 4712 28144
rect 4764 28092 4770 28144
rect 8294 28092 8300 28144
rect 8352 28132 8358 28144
rect 8570 28132 8576 28144
rect 8352 28104 8576 28132
rect 8352 28092 8358 28104
rect 8570 28092 8576 28104
rect 8628 28132 8634 28144
rect 13188 28132 13216 28160
rect 8628 28104 8786 28132
rect 13188 28104 13768 28132
rect 8628 28092 8634 28104
rect 1949 28067 2007 28073
rect 1949 28033 1961 28067
rect 1995 28064 2007 28067
rect 2682 28064 2688 28076
rect 1995 28036 2688 28064
rect 1995 28033 2007 28036
rect 1949 28027 2007 28033
rect 2682 28024 2688 28036
rect 2740 28024 2746 28076
rect 6365 28067 6423 28073
rect 6365 28033 6377 28067
rect 6411 28033 6423 28067
rect 6365 28027 6423 28033
rect 6549 28067 6607 28073
rect 6549 28033 6561 28067
rect 6595 28064 6607 28067
rect 7374 28064 7380 28076
rect 6595 28036 7380 28064
rect 6595 28033 6607 28036
rect 6549 28027 6607 28033
rect 1762 27820 1768 27872
rect 1820 27820 1826 27872
rect 4985 27863 5043 27869
rect 4985 27829 4997 27863
rect 5031 27860 5043 27863
rect 5258 27860 5264 27872
rect 5031 27832 5264 27860
rect 5031 27829 5043 27832
rect 4985 27823 5043 27829
rect 5258 27820 5264 27832
rect 5316 27820 5322 27872
rect 6086 27820 6092 27872
rect 6144 27860 6150 27872
rect 6380 27860 6408 28027
rect 7374 28024 7380 28036
rect 7432 28024 7438 28076
rect 11698 28024 11704 28076
rect 11756 28024 11762 28076
rect 13541 28067 13599 28073
rect 13541 28033 13553 28067
rect 13587 28033 13599 28067
rect 13541 28027 13599 28033
rect 8018 27956 8024 28008
rect 8076 27956 8082 28008
rect 8294 27956 8300 28008
rect 8352 27956 8358 28008
rect 8938 27956 8944 28008
rect 8996 27996 9002 28008
rect 8996 27968 9904 27996
rect 8996 27956 9002 27968
rect 6822 27860 6828 27872
rect 6144 27832 6828 27860
rect 6144 27820 6150 27832
rect 6822 27820 6828 27832
rect 6880 27860 6886 27872
rect 9582 27860 9588 27872
rect 6880 27832 9588 27860
rect 6880 27820 6886 27832
rect 9582 27820 9588 27832
rect 9640 27820 9646 27872
rect 9766 27820 9772 27872
rect 9824 27820 9830 27872
rect 9876 27860 9904 27968
rect 11790 27956 11796 28008
rect 11848 27956 11854 28008
rect 13556 27996 13584 28027
rect 13630 28024 13636 28076
rect 13688 28024 13694 28076
rect 13740 28073 13768 28104
rect 13725 28067 13783 28073
rect 13725 28033 13737 28067
rect 13771 28033 13783 28067
rect 13725 28027 13783 28033
rect 13814 28024 13820 28076
rect 13872 28064 13878 28076
rect 13909 28067 13967 28073
rect 13909 28064 13921 28067
rect 13872 28036 13921 28064
rect 13872 28024 13878 28036
rect 13909 28033 13921 28036
rect 13955 28064 13967 28067
rect 14458 28064 14464 28076
rect 13955 28036 14464 28064
rect 13955 28033 13967 28036
rect 13909 28027 13967 28033
rect 14458 28024 14464 28036
rect 14516 28024 14522 28076
rect 15396 28064 15424 28160
rect 17880 28132 17908 28160
rect 17236 28104 17908 28132
rect 18156 28132 18184 28172
rect 19058 28160 19064 28212
rect 19116 28160 19122 28212
rect 19242 28160 19248 28212
rect 19300 28160 19306 28212
rect 19886 28160 19892 28212
rect 19944 28160 19950 28212
rect 24121 28203 24179 28209
rect 22388 28172 23152 28200
rect 19076 28132 19104 28160
rect 18156 28104 19104 28132
rect 15657 28067 15715 28073
rect 15657 28064 15669 28067
rect 15396 28036 15669 28064
rect 15657 28033 15669 28036
rect 15703 28033 15715 28067
rect 15657 28027 15715 28033
rect 15841 28067 15899 28073
rect 15841 28033 15853 28067
rect 15887 28064 15899 28067
rect 16114 28064 16120 28076
rect 15887 28036 16120 28064
rect 15887 28033 15899 28036
rect 15841 28027 15899 28033
rect 16114 28024 16120 28036
rect 16172 28024 16178 28076
rect 17236 28073 17264 28104
rect 17221 28067 17279 28073
rect 17221 28033 17233 28067
rect 17267 28033 17279 28067
rect 17221 28027 17279 28033
rect 17865 28067 17923 28073
rect 17865 28033 17877 28067
rect 17911 28064 17923 28067
rect 17954 28064 17960 28076
rect 17911 28036 17960 28064
rect 17911 28033 17923 28036
rect 17865 28027 17923 28033
rect 17954 28024 17960 28036
rect 18012 28024 18018 28076
rect 18156 28073 18184 28104
rect 18141 28067 18199 28073
rect 18141 28033 18153 28067
rect 18187 28033 18199 28067
rect 18141 28027 18199 28033
rect 18506 28024 18512 28076
rect 18564 28064 18570 28076
rect 19260 28073 19288 28160
rect 22388 28141 22416 28172
rect 23124 28141 23152 28172
rect 24121 28169 24133 28203
rect 24167 28200 24179 28203
rect 24302 28200 24308 28212
rect 24167 28172 24308 28200
rect 24167 28169 24179 28172
rect 24121 28163 24179 28169
rect 24302 28160 24308 28172
rect 24360 28160 24366 28212
rect 24394 28160 24400 28212
rect 24452 28160 24458 28212
rect 26053 28203 26111 28209
rect 26053 28169 26065 28203
rect 26099 28200 26111 28203
rect 27338 28200 27344 28212
rect 26099 28172 27344 28200
rect 26099 28169 26111 28172
rect 26053 28163 26111 28169
rect 27338 28160 27344 28172
rect 27396 28160 27402 28212
rect 30742 28160 30748 28212
rect 30800 28200 30806 28212
rect 31110 28200 31116 28212
rect 30800 28172 31116 28200
rect 30800 28160 30806 28172
rect 31110 28160 31116 28172
rect 31168 28160 31174 28212
rect 32769 28203 32827 28209
rect 32769 28169 32781 28203
rect 32815 28200 32827 28203
rect 33778 28200 33784 28212
rect 32815 28172 33784 28200
rect 32815 28169 32827 28172
rect 32769 28163 32827 28169
rect 33778 28160 33784 28172
rect 33836 28160 33842 28212
rect 34146 28160 34152 28212
rect 34204 28160 34210 28212
rect 35897 28203 35955 28209
rect 35897 28169 35909 28203
rect 35943 28200 35955 28203
rect 35986 28200 35992 28212
rect 35943 28172 35992 28200
rect 35943 28169 35955 28172
rect 35897 28163 35955 28169
rect 35986 28160 35992 28172
rect 36044 28200 36050 28212
rect 36722 28200 36728 28212
rect 36044 28172 36728 28200
rect 36044 28160 36050 28172
rect 22373 28135 22431 28141
rect 22373 28101 22385 28135
rect 22419 28101 22431 28135
rect 23109 28135 23167 28141
rect 22373 28095 22431 28101
rect 22603 28101 22661 28107
rect 19061 28067 19119 28073
rect 19061 28064 19073 28067
rect 18564 28036 19073 28064
rect 18564 28024 18570 28036
rect 19061 28033 19073 28036
rect 19107 28033 19119 28067
rect 19061 28027 19119 28033
rect 19245 28067 19303 28073
rect 19245 28033 19257 28067
rect 19291 28033 19303 28067
rect 19245 28027 19303 28033
rect 19521 28067 19579 28073
rect 19521 28033 19533 28067
rect 19567 28033 19579 28067
rect 19521 28027 19579 28033
rect 19797 28067 19855 28073
rect 19797 28033 19809 28067
rect 19843 28033 19855 28067
rect 19797 28027 19855 28033
rect 15010 27996 15016 28008
rect 13556 27968 15016 27996
rect 15010 27956 15016 27968
rect 15068 27956 15074 28008
rect 17126 27956 17132 28008
rect 17184 27956 17190 28008
rect 18325 27999 18383 28005
rect 18325 27965 18337 27999
rect 18371 27996 18383 27999
rect 18966 27996 18972 28008
rect 18371 27968 18972 27996
rect 18371 27965 18383 27968
rect 18325 27959 18383 27965
rect 18966 27956 18972 27968
rect 19024 27996 19030 28008
rect 19429 27999 19487 28005
rect 19429 27996 19441 27999
rect 19024 27968 19441 27996
rect 19024 27956 19030 27968
rect 19429 27965 19441 27968
rect 19475 27965 19487 27999
rect 19429 27959 19487 27965
rect 12069 27931 12127 27937
rect 12069 27897 12081 27931
rect 12115 27928 12127 27931
rect 12526 27928 12532 27940
rect 12115 27900 12532 27928
rect 12115 27897 12127 27900
rect 12069 27891 12127 27897
rect 12526 27888 12532 27900
rect 12584 27888 12590 27940
rect 17957 27931 18015 27937
rect 17957 27897 17969 27931
rect 18003 27928 18015 27931
rect 18138 27928 18144 27940
rect 18003 27900 18144 27928
rect 18003 27897 18015 27900
rect 17957 27891 18015 27897
rect 18138 27888 18144 27900
rect 18196 27888 18202 27940
rect 19334 27888 19340 27940
rect 19392 27888 19398 27940
rect 13265 27863 13323 27869
rect 13265 27860 13277 27863
rect 9876 27832 13277 27860
rect 13265 27829 13277 27832
rect 13311 27829 13323 27863
rect 19536 27860 19564 28027
rect 19812 27996 19840 28027
rect 19886 28024 19892 28076
rect 19944 28064 19950 28076
rect 22278 28064 22284 28076
rect 19944 28036 22284 28064
rect 19944 28024 19950 28036
rect 22278 28024 22284 28036
rect 22336 28024 22342 28076
rect 22603 28067 22615 28101
rect 22649 28067 22661 28101
rect 23109 28101 23121 28135
rect 23155 28132 23167 28135
rect 23155 28104 24164 28132
rect 23155 28101 23167 28104
rect 23109 28095 23167 28101
rect 22603 28064 22661 28067
rect 22830 28064 22836 28076
rect 22603 28061 22836 28064
rect 22604 28036 22836 28061
rect 22830 28024 22836 28036
rect 22888 28024 22894 28076
rect 22925 28067 22983 28073
rect 22925 28033 22937 28067
rect 22971 28033 22983 28067
rect 22925 28027 22983 28033
rect 23937 28067 23995 28073
rect 23937 28033 23949 28067
rect 23983 28033 23995 28067
rect 23937 28027 23995 28033
rect 19978 27996 19984 28008
rect 19812 27968 19984 27996
rect 19978 27956 19984 27968
rect 20036 27956 20042 28008
rect 22462 27956 22468 28008
rect 22520 27996 22526 28008
rect 22940 27996 22968 28027
rect 22520 27968 22968 27996
rect 22520 27956 22526 27968
rect 19705 27931 19763 27937
rect 19705 27897 19717 27931
rect 19751 27928 19763 27931
rect 23952 27928 23980 28027
rect 24136 27996 24164 28104
rect 24213 28067 24271 28073
rect 24213 28033 24225 28067
rect 24259 28064 24271 28067
rect 24412 28064 24440 28160
rect 27065 28135 27123 28141
rect 24780 28104 24992 28132
rect 24780 28073 24808 28104
rect 24964 28076 24992 28104
rect 27065 28101 27077 28135
rect 27111 28132 27123 28135
rect 27246 28132 27252 28144
rect 27111 28104 27252 28132
rect 27111 28101 27123 28104
rect 27065 28095 27123 28101
rect 27246 28092 27252 28104
rect 27304 28092 27310 28144
rect 34164 28132 34192 28160
rect 32968 28104 34008 28132
rect 34164 28104 34560 28132
rect 32968 28076 32996 28104
rect 24259 28036 24440 28064
rect 24765 28067 24823 28073
rect 24259 28033 24271 28036
rect 24213 28027 24271 28033
rect 24765 28033 24777 28067
rect 24811 28033 24823 28067
rect 24765 28027 24823 28033
rect 24854 28024 24860 28076
rect 24912 28024 24918 28076
rect 24946 28024 24952 28076
rect 25004 28024 25010 28076
rect 25590 28024 25596 28076
rect 25648 28024 25654 28076
rect 25866 28024 25872 28076
rect 25924 28024 25930 28076
rect 26602 28024 26608 28076
rect 26660 28064 26666 28076
rect 26786 28064 26792 28076
rect 26660 28036 26792 28064
rect 26660 28024 26666 28036
rect 26786 28024 26792 28036
rect 26844 28064 26850 28076
rect 26973 28067 27031 28073
rect 26973 28064 26985 28067
rect 26844 28036 26985 28064
rect 26844 28024 26850 28036
rect 26973 28033 26985 28036
rect 27019 28033 27031 28067
rect 26973 28027 27031 28033
rect 27154 28024 27160 28076
rect 27212 28064 27218 28076
rect 28534 28064 28540 28076
rect 27212 28036 28540 28064
rect 27212 28024 27218 28036
rect 28534 28024 28540 28036
rect 28592 28024 28598 28076
rect 32122 28024 32128 28076
rect 32180 28024 32186 28076
rect 32309 28067 32367 28073
rect 32309 28033 32321 28067
rect 32355 28033 32367 28067
rect 32309 28027 32367 28033
rect 32324 27996 32352 28027
rect 32398 28024 32404 28076
rect 32456 28024 32462 28076
rect 32493 28067 32551 28073
rect 32493 28033 32505 28067
rect 32539 28064 32551 28067
rect 32766 28064 32772 28076
rect 32539 28036 32772 28064
rect 32539 28033 32551 28036
rect 32493 28027 32551 28033
rect 32766 28024 32772 28036
rect 32824 28024 32830 28076
rect 32861 28067 32919 28073
rect 32861 28033 32873 28067
rect 32907 28064 32919 28067
rect 32950 28064 32956 28076
rect 32907 28036 32956 28064
rect 32907 28033 32919 28036
rect 32861 28027 32919 28033
rect 32950 28024 32956 28036
rect 33008 28024 33014 28076
rect 33045 28067 33103 28073
rect 33045 28033 33057 28067
rect 33091 28064 33103 28067
rect 33318 28064 33324 28076
rect 33091 28036 33324 28064
rect 33091 28033 33103 28036
rect 33045 28027 33103 28033
rect 33318 28024 33324 28036
rect 33376 28064 33382 28076
rect 33505 28067 33563 28073
rect 33505 28064 33517 28067
rect 33376 28036 33517 28064
rect 33376 28024 33382 28036
rect 33505 28033 33517 28036
rect 33551 28033 33563 28067
rect 33505 28027 33563 28033
rect 32582 27996 32588 28008
rect 24136 27968 31754 27996
rect 32324 27968 32588 27996
rect 19751 27900 23980 27928
rect 24857 27931 24915 27937
rect 19751 27897 19763 27900
rect 19705 27891 19763 27897
rect 24857 27897 24869 27931
rect 24903 27928 24915 27931
rect 25406 27928 25412 27940
rect 24903 27900 25412 27928
rect 24903 27897 24915 27900
rect 24857 27891 24915 27897
rect 25406 27888 25412 27900
rect 25464 27888 25470 27940
rect 25685 27931 25743 27937
rect 25685 27897 25697 27931
rect 25731 27897 25743 27931
rect 25685 27891 25743 27897
rect 22370 27860 22376 27872
rect 19536 27832 22376 27860
rect 13265 27823 13323 27829
rect 22370 27820 22376 27832
rect 22428 27820 22434 27872
rect 22462 27820 22468 27872
rect 22520 27860 22526 27872
rect 22557 27863 22615 27869
rect 22557 27860 22569 27863
rect 22520 27832 22569 27860
rect 22520 27820 22526 27832
rect 22557 27829 22569 27832
rect 22603 27829 22615 27863
rect 22557 27823 22615 27829
rect 22738 27820 22744 27872
rect 22796 27820 22802 27872
rect 23106 27820 23112 27872
rect 23164 27820 23170 27872
rect 23934 27820 23940 27872
rect 23992 27820 23998 27872
rect 25130 27820 25136 27872
rect 25188 27860 25194 27872
rect 25700 27860 25728 27891
rect 25774 27888 25780 27940
rect 25832 27888 25838 27940
rect 31726 27928 31754 27968
rect 32582 27956 32588 27968
rect 32640 27956 32646 28008
rect 33520 27996 33548 28027
rect 33594 28024 33600 28076
rect 33652 28064 33658 28076
rect 33870 28064 33876 28076
rect 33652 28036 33876 28064
rect 33652 28024 33658 28036
rect 33870 28024 33876 28036
rect 33928 28024 33934 28076
rect 33980 28064 34008 28104
rect 33980 28036 34192 28064
rect 34164 27996 34192 28036
rect 34422 28024 34428 28076
rect 34480 28024 34486 28076
rect 34532 28073 34560 28104
rect 34517 28067 34575 28073
rect 34517 28033 34529 28067
rect 34563 28033 34575 28067
rect 34517 28027 34575 28033
rect 34698 28024 34704 28076
rect 34756 28064 34762 28076
rect 35069 28067 35127 28073
rect 35069 28064 35081 28067
rect 34756 28036 35081 28064
rect 34756 28024 34762 28036
rect 35069 28033 35081 28036
rect 35115 28033 35127 28067
rect 35069 28027 35127 28033
rect 35250 28024 35256 28076
rect 35308 28064 35314 28076
rect 36188 28073 36216 28172
rect 36722 28160 36728 28172
rect 36780 28160 36786 28212
rect 35989 28067 36047 28073
rect 35989 28064 36001 28067
rect 35308 28036 36001 28064
rect 35308 28024 35314 28036
rect 35989 28033 36001 28036
rect 36035 28033 36047 28067
rect 35989 28027 36047 28033
rect 36173 28067 36231 28073
rect 36173 28033 36185 28067
rect 36219 28033 36231 28067
rect 36173 28027 36231 28033
rect 35434 27996 35440 28008
rect 33520 27968 34100 27996
rect 34164 27968 35440 27996
rect 33873 27931 33931 27937
rect 33873 27928 33885 27931
rect 31726 27900 33885 27928
rect 33873 27897 33885 27900
rect 33919 27897 33931 27931
rect 34072 27928 34100 27968
rect 35434 27956 35440 27968
rect 35492 27956 35498 28008
rect 35713 27931 35771 27937
rect 35713 27928 35725 27931
rect 34072 27900 35725 27928
rect 33873 27891 33931 27897
rect 35713 27897 35725 27900
rect 35759 27897 35771 27931
rect 35713 27891 35771 27897
rect 36265 27931 36323 27937
rect 36265 27897 36277 27931
rect 36311 27928 36323 27931
rect 36722 27928 36728 27940
rect 36311 27900 36728 27928
rect 36311 27897 36323 27900
rect 36265 27891 36323 27897
rect 36722 27888 36728 27900
rect 36780 27888 36786 27940
rect 26786 27860 26792 27872
rect 25188 27832 26792 27860
rect 25188 27820 25194 27832
rect 26786 27820 26792 27832
rect 26844 27820 26850 27872
rect 32490 27820 32496 27872
rect 32548 27860 32554 27872
rect 32861 27863 32919 27869
rect 32861 27860 32873 27863
rect 32548 27832 32873 27860
rect 32548 27820 32554 27832
rect 32861 27829 32873 27832
rect 32907 27829 32919 27863
rect 32861 27823 32919 27829
rect 1104 27770 38272 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38272 27770
rect 1104 27696 38272 27718
rect 4798 27616 4804 27668
rect 4856 27656 4862 27668
rect 4893 27659 4951 27665
rect 4893 27656 4905 27659
rect 4856 27628 4905 27656
rect 4856 27616 4862 27628
rect 4893 27625 4905 27628
rect 4939 27625 4951 27659
rect 4893 27619 4951 27625
rect 5534 27616 5540 27668
rect 5592 27656 5598 27668
rect 6365 27659 6423 27665
rect 6365 27656 6377 27659
rect 5592 27628 6377 27656
rect 5592 27616 5598 27628
rect 6365 27625 6377 27628
rect 6411 27625 6423 27659
rect 6914 27656 6920 27668
rect 6365 27619 6423 27625
rect 6656 27628 6920 27656
rect 4154 27548 4160 27600
rect 4212 27588 4218 27600
rect 6656 27588 6684 27628
rect 6914 27616 6920 27628
rect 6972 27616 6978 27668
rect 7006 27616 7012 27668
rect 7064 27656 7070 27668
rect 7193 27659 7251 27665
rect 7193 27656 7205 27659
rect 7064 27628 7205 27656
rect 7064 27616 7070 27628
rect 7193 27625 7205 27628
rect 7239 27625 7251 27659
rect 7193 27619 7251 27625
rect 8294 27616 8300 27668
rect 8352 27616 8358 27668
rect 8570 27616 8576 27668
rect 8628 27656 8634 27668
rect 9858 27656 9864 27668
rect 8628 27628 9864 27656
rect 8628 27616 8634 27628
rect 9858 27616 9864 27628
rect 9916 27616 9922 27668
rect 12544 27628 14964 27656
rect 4212 27560 6684 27588
rect 6733 27591 6791 27597
rect 4212 27548 4218 27560
rect 6733 27557 6745 27591
rect 6779 27588 6791 27591
rect 7098 27588 7104 27600
rect 6779 27560 7104 27588
rect 6779 27557 6791 27560
rect 6733 27551 6791 27557
rect 7098 27548 7104 27560
rect 7156 27548 7162 27600
rect 7282 27548 7288 27600
rect 7340 27588 7346 27600
rect 9766 27588 9772 27600
rect 7340 27560 7788 27588
rect 7340 27548 7346 27560
rect 6641 27523 6699 27529
rect 6641 27489 6653 27523
rect 6687 27520 6699 27523
rect 7760 27520 7788 27560
rect 9416 27560 9772 27588
rect 9416 27529 9444 27560
rect 9766 27548 9772 27560
rect 9824 27588 9830 27600
rect 12544 27588 12572 27628
rect 9824 27560 12572 27588
rect 9824 27548 9830 27560
rect 9401 27523 9459 27529
rect 6687 27492 7696 27520
rect 7760 27492 9352 27520
rect 6687 27489 6699 27492
rect 6641 27483 6699 27489
rect 7668 27464 7696 27492
rect 4893 27455 4951 27461
rect 4893 27452 4905 27455
rect 4632 27424 4905 27452
rect 4632 27328 4660 27424
rect 4893 27421 4905 27424
rect 4939 27421 4951 27455
rect 4893 27415 4951 27421
rect 5077 27455 5135 27461
rect 5077 27421 5089 27455
rect 5123 27452 5135 27455
rect 6549 27455 6607 27461
rect 5123 27424 5304 27452
rect 5123 27421 5135 27424
rect 5077 27415 5135 27421
rect 5276 27328 5304 27424
rect 6549 27421 6561 27455
rect 6595 27421 6607 27455
rect 6549 27415 6607 27421
rect 6825 27455 6883 27461
rect 6825 27421 6837 27455
rect 6871 27421 6883 27455
rect 6825 27415 6883 27421
rect 4614 27276 4620 27328
rect 4672 27276 4678 27328
rect 4706 27276 4712 27328
rect 4764 27276 4770 27328
rect 5258 27276 5264 27328
rect 5316 27276 5322 27328
rect 6564 27316 6592 27415
rect 6840 27384 6868 27415
rect 6914 27412 6920 27464
rect 6972 27452 6978 27464
rect 7101 27455 7159 27461
rect 7101 27452 7113 27455
rect 6972 27424 7113 27452
rect 6972 27412 6978 27424
rect 7101 27421 7113 27424
rect 7147 27421 7159 27455
rect 7101 27415 7159 27421
rect 7650 27412 7656 27464
rect 7708 27412 7714 27464
rect 8481 27455 8539 27461
rect 8481 27421 8493 27455
rect 8527 27452 8539 27455
rect 9324 27452 9352 27492
rect 9401 27489 9413 27523
rect 9447 27489 9459 27523
rect 9401 27483 9459 27489
rect 9493 27523 9551 27529
rect 9493 27489 9505 27523
rect 9539 27489 9551 27523
rect 9493 27483 9551 27489
rect 9508 27452 9536 27483
rect 9674 27480 9680 27532
rect 9732 27520 9738 27532
rect 10686 27520 10692 27532
rect 9732 27492 10692 27520
rect 9732 27480 9738 27492
rect 10686 27480 10692 27492
rect 10744 27520 10750 27532
rect 11885 27523 11943 27529
rect 11885 27520 11897 27523
rect 10744 27492 11897 27520
rect 10744 27480 10750 27492
rect 11885 27489 11897 27492
rect 11931 27489 11943 27523
rect 12544 27520 12572 27560
rect 12710 27548 12716 27600
rect 12768 27548 12774 27600
rect 13078 27548 13084 27600
rect 13136 27588 13142 27600
rect 13265 27591 13323 27597
rect 13265 27588 13277 27591
rect 13136 27560 13277 27588
rect 13136 27548 13142 27560
rect 13265 27557 13277 27560
rect 13311 27557 13323 27591
rect 14826 27588 14832 27600
rect 13265 27551 13323 27557
rect 13372 27560 14832 27588
rect 11885 27483 11943 27489
rect 12452 27492 12572 27520
rect 8527 27424 8984 27452
rect 9324 27424 9536 27452
rect 11057 27455 11115 27461
rect 8527 27421 8539 27424
rect 8481 27415 8539 27421
rect 8202 27384 8208 27396
rect 6840 27356 8208 27384
rect 8202 27344 8208 27356
rect 8260 27344 8266 27396
rect 7282 27316 7288 27328
rect 6564 27288 7288 27316
rect 7282 27276 7288 27288
rect 7340 27276 7346 27328
rect 7558 27276 7564 27328
rect 7616 27276 7622 27328
rect 8956 27325 8984 27424
rect 11057 27421 11069 27455
rect 11103 27452 11115 27455
rect 11103 27424 11376 27452
rect 11103 27421 11115 27424
rect 11057 27415 11115 27421
rect 8941 27319 8999 27325
rect 8941 27285 8953 27319
rect 8987 27285 8999 27319
rect 8941 27279 8999 27285
rect 9309 27319 9367 27325
rect 9309 27285 9321 27319
rect 9355 27316 9367 27319
rect 9582 27316 9588 27328
rect 9355 27288 9588 27316
rect 9355 27285 9367 27288
rect 9309 27279 9367 27285
rect 9582 27276 9588 27288
rect 9640 27276 9646 27328
rect 11238 27276 11244 27328
rect 11296 27276 11302 27328
rect 11348 27325 11376 27424
rect 12342 27412 12348 27464
rect 12400 27412 12406 27464
rect 12452 27461 12480 27492
rect 12437 27455 12495 27461
rect 12437 27421 12449 27455
rect 12483 27421 12495 27455
rect 12437 27415 12495 27421
rect 12526 27412 12532 27464
rect 12584 27412 12590 27464
rect 12720 27461 12748 27548
rect 13372 27520 13400 27560
rect 14826 27548 14832 27560
rect 14884 27548 14890 27600
rect 12820 27492 13400 27520
rect 13449 27523 13507 27529
rect 12693 27455 12751 27461
rect 12693 27421 12705 27455
rect 12739 27421 12751 27455
rect 12693 27415 12751 27421
rect 11698 27344 11704 27396
rect 11756 27384 11762 27396
rect 12820 27393 12848 27492
rect 13449 27489 13461 27523
rect 13495 27520 13507 27523
rect 14936 27520 14964 27628
rect 15010 27616 15016 27668
rect 15068 27616 15074 27668
rect 19334 27616 19340 27668
rect 19392 27656 19398 27668
rect 19429 27659 19487 27665
rect 19429 27656 19441 27659
rect 19392 27628 19441 27656
rect 19392 27616 19398 27628
rect 19429 27625 19441 27628
rect 19475 27625 19487 27659
rect 19429 27619 19487 27625
rect 19978 27616 19984 27668
rect 20036 27616 20042 27668
rect 20346 27616 20352 27668
rect 20404 27616 20410 27668
rect 22370 27616 22376 27668
rect 22428 27656 22434 27668
rect 25406 27656 25412 27668
rect 22428 27628 25412 27656
rect 22428 27616 22434 27628
rect 25406 27616 25412 27628
rect 25464 27616 25470 27668
rect 36633 27659 36691 27665
rect 29196 27628 29592 27656
rect 15028 27588 15056 27616
rect 15749 27591 15807 27597
rect 15749 27588 15761 27591
rect 15028 27560 15761 27588
rect 15749 27557 15761 27560
rect 15795 27557 15807 27591
rect 15749 27551 15807 27557
rect 16390 27548 16396 27600
rect 16448 27588 16454 27600
rect 19518 27588 19524 27600
rect 16448 27560 19524 27588
rect 16448 27548 16454 27560
rect 19518 27548 19524 27560
rect 19576 27548 19582 27600
rect 23014 27588 23020 27600
rect 22388 27560 23020 27588
rect 13495 27492 14412 27520
rect 14936 27492 19564 27520
rect 13495 27489 13507 27492
rect 13449 27483 13507 27489
rect 12989 27455 13047 27461
rect 12989 27421 13001 27455
rect 13035 27452 13047 27455
rect 13464 27452 13492 27483
rect 14384 27464 14412 27492
rect 19536 27464 19564 27492
rect 19904 27492 20208 27520
rect 19904 27464 19932 27492
rect 13035 27424 13492 27452
rect 13541 27455 13599 27461
rect 13035 27421 13047 27424
rect 12989 27415 13047 27421
rect 13541 27421 13553 27455
rect 13587 27452 13599 27455
rect 13587 27424 14320 27452
rect 13587 27421 13599 27424
rect 13541 27415 13599 27421
rect 12805 27387 12863 27393
rect 11756 27356 12434 27384
rect 11756 27344 11762 27356
rect 11333 27319 11391 27325
rect 11333 27285 11345 27319
rect 11379 27285 11391 27319
rect 11333 27279 11391 27285
rect 11793 27319 11851 27325
rect 11793 27285 11805 27319
rect 11839 27316 11851 27319
rect 12161 27319 12219 27325
rect 12161 27316 12173 27319
rect 11839 27288 12173 27316
rect 11839 27285 11851 27288
rect 11793 27279 11851 27285
rect 12161 27285 12173 27288
rect 12207 27285 12219 27319
rect 12406 27316 12434 27356
rect 12805 27353 12817 27387
rect 12851 27353 12863 27387
rect 13262 27384 13268 27396
rect 12805 27347 12863 27353
rect 13096 27356 13268 27384
rect 13096 27316 13124 27356
rect 13262 27344 13268 27356
rect 13320 27384 13326 27396
rect 13817 27387 13875 27393
rect 13817 27384 13829 27387
rect 13320 27356 13829 27384
rect 13320 27344 13326 27356
rect 13817 27353 13829 27356
rect 13863 27353 13875 27387
rect 13817 27347 13875 27353
rect 13909 27387 13967 27393
rect 13909 27353 13921 27387
rect 13955 27384 13967 27387
rect 14090 27384 14096 27396
rect 13955 27356 14096 27384
rect 13955 27353 13967 27356
rect 13909 27347 13967 27353
rect 14090 27344 14096 27356
rect 14148 27344 14154 27396
rect 14292 27384 14320 27424
rect 14366 27412 14372 27464
rect 14424 27412 14430 27464
rect 14826 27412 14832 27464
rect 14884 27412 14890 27464
rect 15654 27412 15660 27464
rect 15712 27452 15718 27464
rect 15933 27455 15991 27461
rect 15933 27452 15945 27455
rect 15712 27424 15945 27452
rect 15712 27412 15718 27424
rect 15933 27421 15945 27424
rect 15979 27421 15991 27455
rect 15933 27415 15991 27421
rect 16117 27455 16175 27461
rect 16117 27421 16129 27455
rect 16163 27452 16175 27455
rect 17678 27452 17684 27464
rect 16163 27424 17684 27452
rect 16163 27421 16175 27424
rect 16117 27415 16175 27421
rect 17678 27412 17684 27424
rect 17736 27412 17742 27464
rect 19429 27455 19487 27461
rect 19429 27421 19441 27455
rect 19475 27421 19487 27455
rect 19429 27415 19487 27421
rect 17494 27384 17500 27396
rect 14292 27356 17500 27384
rect 17494 27344 17500 27356
rect 17552 27344 17558 27396
rect 18690 27384 18696 27396
rect 17604 27356 18696 27384
rect 12406 27288 13124 27316
rect 12161 27279 12219 27285
rect 13170 27276 13176 27328
rect 13228 27276 13234 27328
rect 14182 27276 14188 27328
rect 14240 27276 14246 27328
rect 15378 27276 15384 27328
rect 15436 27316 15442 27328
rect 17604 27316 17632 27356
rect 18690 27344 18696 27356
rect 18748 27344 18754 27396
rect 19242 27344 19248 27396
rect 19300 27384 19306 27396
rect 19444 27384 19472 27415
rect 19518 27412 19524 27464
rect 19576 27412 19582 27464
rect 19613 27455 19671 27461
rect 19613 27421 19625 27455
rect 19659 27452 19671 27455
rect 19797 27455 19855 27461
rect 19797 27452 19809 27455
rect 19659 27424 19809 27452
rect 19659 27421 19671 27424
rect 19613 27415 19671 27421
rect 19797 27421 19809 27424
rect 19843 27421 19855 27455
rect 19797 27415 19855 27421
rect 19886 27412 19892 27464
rect 19944 27412 19950 27464
rect 20180 27461 20208 27492
rect 19981 27455 20039 27461
rect 19981 27421 19993 27455
rect 20027 27421 20039 27455
rect 19981 27415 20039 27421
rect 20165 27455 20223 27461
rect 20165 27421 20177 27455
rect 20211 27452 20223 27455
rect 20257 27455 20315 27461
rect 20257 27452 20269 27455
rect 20211 27424 20269 27452
rect 20211 27421 20223 27424
rect 20165 27415 20223 27421
rect 20257 27421 20269 27424
rect 20303 27421 20315 27455
rect 20257 27415 20315 27421
rect 20441 27455 20499 27461
rect 20441 27421 20453 27455
rect 20487 27421 20499 27455
rect 20441 27415 20499 27421
rect 19996 27384 20024 27415
rect 20456 27384 20484 27415
rect 22186 27412 22192 27464
rect 22244 27452 22250 27464
rect 22388 27461 22416 27560
rect 23014 27548 23020 27560
rect 23072 27548 23078 27600
rect 23106 27548 23112 27600
rect 23164 27548 23170 27600
rect 24394 27548 24400 27600
rect 24452 27588 24458 27600
rect 25958 27588 25964 27600
rect 24452 27560 25964 27588
rect 24452 27548 24458 27560
rect 25958 27548 25964 27560
rect 26016 27548 26022 27600
rect 27341 27591 27399 27597
rect 27341 27557 27353 27591
rect 27387 27588 27399 27591
rect 27522 27588 27528 27600
rect 27387 27560 27528 27588
rect 27387 27557 27399 27560
rect 27341 27551 27399 27557
rect 27522 27548 27528 27560
rect 27580 27548 27586 27600
rect 27798 27548 27804 27600
rect 27856 27588 27862 27600
rect 29196 27588 29224 27628
rect 27856 27560 29224 27588
rect 29273 27591 29331 27597
rect 27856 27548 27862 27560
rect 29273 27557 29285 27591
rect 29319 27588 29331 27591
rect 29454 27588 29460 27600
rect 29319 27560 29460 27588
rect 29319 27557 29331 27560
rect 29273 27551 29331 27557
rect 29454 27548 29460 27560
rect 29512 27548 29518 27600
rect 29564 27588 29592 27628
rect 36633 27625 36645 27659
rect 36679 27656 36691 27659
rect 36679 27628 36952 27656
rect 36679 27625 36691 27628
rect 36633 27619 36691 27625
rect 36924 27588 36952 27628
rect 29564 27560 31754 27588
rect 36924 27560 37320 27588
rect 23124 27520 23152 27548
rect 29730 27520 29736 27532
rect 22572 27492 23152 27520
rect 25240 27492 28488 27520
rect 22572 27461 22600 27492
rect 22373 27455 22431 27461
rect 22373 27452 22385 27455
rect 22244 27424 22385 27452
rect 22244 27412 22250 27424
rect 22373 27421 22385 27424
rect 22419 27421 22431 27455
rect 22373 27415 22431 27421
rect 22557 27455 22615 27461
rect 22557 27421 22569 27455
rect 22603 27421 22615 27455
rect 22557 27415 22615 27421
rect 22738 27412 22744 27464
rect 22796 27412 22802 27464
rect 22830 27412 22836 27464
rect 22888 27452 22894 27464
rect 25130 27452 25136 27464
rect 22888 27424 25136 27452
rect 22888 27412 22894 27424
rect 25130 27412 25136 27424
rect 25188 27412 25194 27464
rect 25240 27396 25268 27492
rect 27154 27412 27160 27464
rect 27212 27452 27218 27464
rect 27249 27455 27307 27461
rect 27249 27452 27261 27455
rect 27212 27424 27261 27452
rect 27212 27412 27218 27424
rect 27249 27421 27261 27424
rect 27295 27421 27307 27455
rect 27249 27415 27307 27421
rect 27430 27412 27436 27464
rect 27488 27412 27494 27464
rect 22925 27387 22983 27393
rect 22925 27384 22937 27387
rect 19300 27356 20484 27384
rect 22066 27356 22937 27384
rect 19300 27344 19306 27356
rect 15436 27288 17632 27316
rect 15436 27276 15442 27288
rect 17678 27276 17684 27328
rect 17736 27316 17742 27328
rect 22066 27316 22094 27356
rect 22925 27353 22937 27356
rect 22971 27353 22983 27387
rect 22925 27347 22983 27353
rect 23017 27387 23075 27393
rect 23017 27353 23029 27387
rect 23063 27384 23075 27387
rect 23106 27384 23112 27396
rect 23063 27356 23112 27384
rect 23063 27353 23075 27356
rect 23017 27347 23075 27353
rect 23106 27344 23112 27356
rect 23164 27344 23170 27396
rect 25222 27344 25228 27396
rect 25280 27344 25286 27396
rect 28460 27384 28488 27492
rect 28736 27492 29736 27520
rect 28736 27464 28764 27492
rect 29730 27480 29736 27492
rect 29788 27520 29794 27532
rect 30101 27523 30159 27529
rect 30101 27520 30113 27523
rect 29788 27492 30113 27520
rect 29788 27480 29794 27492
rect 30101 27489 30113 27492
rect 30147 27489 30159 27523
rect 31726 27520 31754 27560
rect 32858 27520 32864 27532
rect 31726 27492 32864 27520
rect 30101 27483 30159 27489
rect 32858 27480 32864 27492
rect 32916 27480 32922 27532
rect 37090 27520 37096 27532
rect 36648 27492 37096 27520
rect 28718 27412 28724 27464
rect 28776 27412 28782 27464
rect 29181 27455 29239 27461
rect 29181 27421 29193 27455
rect 29227 27421 29239 27455
rect 29181 27415 29239 27421
rect 29196 27384 29224 27415
rect 29362 27412 29368 27464
rect 29420 27452 29426 27464
rect 29549 27455 29607 27461
rect 29549 27452 29561 27455
rect 29420 27424 29561 27452
rect 29420 27412 29426 27424
rect 29549 27421 29561 27424
rect 29595 27421 29607 27455
rect 29549 27415 29607 27421
rect 29825 27455 29883 27461
rect 29825 27421 29837 27455
rect 29871 27452 29883 27455
rect 29914 27452 29920 27464
rect 29871 27424 29920 27452
rect 29871 27421 29883 27424
rect 29825 27415 29883 27421
rect 29638 27384 29644 27396
rect 28460 27356 29644 27384
rect 29638 27344 29644 27356
rect 29696 27344 29702 27396
rect 17736 27288 22094 27316
rect 17736 27276 17742 27288
rect 22278 27276 22284 27328
rect 22336 27316 22342 27328
rect 24578 27316 24584 27328
rect 22336 27288 24584 27316
rect 22336 27276 22342 27288
rect 24578 27276 24584 27288
rect 24636 27316 24642 27328
rect 28902 27316 28908 27328
rect 24636 27288 28908 27316
rect 24636 27276 24642 27288
rect 28902 27276 28908 27288
rect 28960 27276 28966 27328
rect 29546 27276 29552 27328
rect 29604 27316 29610 27328
rect 29840 27316 29868 27415
rect 29914 27412 29920 27424
rect 29972 27412 29978 27464
rect 30285 27455 30343 27461
rect 30285 27421 30297 27455
rect 30331 27452 30343 27455
rect 30374 27452 30380 27464
rect 30331 27424 30380 27452
rect 30331 27421 30343 27424
rect 30285 27415 30343 27421
rect 30374 27412 30380 27424
rect 30432 27412 30438 27464
rect 30561 27455 30619 27461
rect 30561 27421 30573 27455
rect 30607 27452 30619 27455
rect 30607 27424 30972 27452
rect 30607 27421 30619 27424
rect 30561 27415 30619 27421
rect 30006 27344 30012 27396
rect 30064 27384 30070 27396
rect 30469 27387 30527 27393
rect 30469 27384 30481 27387
rect 30064 27356 30481 27384
rect 30064 27344 30070 27356
rect 30469 27353 30481 27356
rect 30515 27353 30527 27387
rect 30469 27347 30527 27353
rect 30944 27328 30972 27424
rect 34514 27412 34520 27464
rect 34572 27452 34578 27464
rect 34701 27455 34759 27461
rect 34701 27452 34713 27455
rect 34572 27424 34713 27452
rect 34572 27412 34578 27424
rect 34701 27421 34713 27424
rect 34747 27452 34759 27455
rect 34790 27452 34796 27464
rect 34747 27424 34796 27452
rect 34747 27421 34759 27424
rect 34701 27415 34759 27421
rect 34790 27412 34796 27424
rect 34848 27412 34854 27464
rect 34882 27412 34888 27464
rect 34940 27412 34946 27464
rect 36446 27412 36452 27464
rect 36504 27412 36510 27464
rect 36648 27461 36676 27492
rect 37090 27480 37096 27492
rect 37148 27480 37154 27532
rect 37292 27529 37320 27560
rect 37277 27523 37335 27529
rect 37277 27489 37289 27523
rect 37323 27489 37335 27523
rect 37277 27483 37335 27489
rect 36633 27455 36691 27461
rect 36633 27421 36645 27455
rect 36679 27421 36691 27455
rect 36633 27415 36691 27421
rect 36814 27412 36820 27464
rect 36872 27454 36878 27464
rect 37369 27455 37427 27461
rect 36872 27452 36952 27454
rect 37369 27452 37381 27455
rect 36872 27426 37381 27452
rect 36872 27412 36878 27426
rect 36924 27424 37381 27426
rect 37369 27421 37381 27424
rect 37415 27421 37427 27455
rect 37369 27415 37427 27421
rect 34422 27344 34428 27396
rect 34480 27384 34486 27396
rect 36725 27387 36783 27393
rect 36725 27384 36737 27387
rect 34480 27356 36737 27384
rect 34480 27344 34486 27356
rect 36725 27353 36737 27356
rect 36771 27353 36783 27387
rect 36725 27347 36783 27353
rect 29604 27288 29868 27316
rect 29604 27276 29610 27288
rect 30926 27276 30932 27328
rect 30984 27276 30990 27328
rect 34330 27276 34336 27328
rect 34388 27316 34394 27328
rect 34793 27319 34851 27325
rect 34793 27316 34805 27319
rect 34388 27288 34805 27316
rect 34388 27276 34394 27288
rect 34793 27285 34805 27288
rect 34839 27285 34851 27319
rect 34793 27279 34851 27285
rect 1104 27226 38272 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 38272 27226
rect 1104 27152 38272 27174
rect 2774 27072 2780 27124
rect 2832 27072 2838 27124
rect 5626 27072 5632 27124
rect 5684 27072 5690 27124
rect 7101 27115 7159 27121
rect 7101 27112 7113 27115
rect 5828 27084 7113 27112
rect 2792 27044 2820 27072
rect 2792 27016 2898 27044
rect 2130 26936 2136 26988
rect 2188 26936 2194 26988
rect 3970 26936 3976 26988
rect 4028 26936 4034 26988
rect 4709 26979 4767 26985
rect 4709 26945 4721 26979
rect 4755 26976 4767 26979
rect 4798 26976 4804 26988
rect 4755 26948 4804 26976
rect 4755 26945 4767 26948
rect 4709 26939 4767 26945
rect 2409 26911 2467 26917
rect 2409 26877 2421 26911
rect 2455 26908 2467 26911
rect 3418 26908 3424 26920
rect 2455 26880 3424 26908
rect 2455 26877 2467 26880
rect 2409 26871 2467 26877
rect 3418 26868 3424 26880
rect 3476 26868 3482 26920
rect 3881 26911 3939 26917
rect 3881 26877 3893 26911
rect 3927 26908 3939 26911
rect 4724 26908 4752 26939
rect 4798 26936 4804 26948
rect 4856 26976 4862 26988
rect 5828 26985 5856 27084
rect 7101 27081 7113 27084
rect 7147 27081 7159 27115
rect 7101 27075 7159 27081
rect 7208 27084 7972 27112
rect 6914 27044 6920 27056
rect 6589 27016 6920 27044
rect 4985 26979 5043 26985
rect 4985 26976 4997 26979
rect 4856 26948 4997 26976
rect 4856 26936 4862 26948
rect 4985 26945 4997 26948
rect 5031 26945 5043 26979
rect 4985 26939 5043 26945
rect 5353 26979 5411 26985
rect 5353 26945 5365 26979
rect 5399 26945 5411 26979
rect 5353 26939 5411 26945
rect 5813 26979 5871 26985
rect 5813 26945 5825 26979
rect 5859 26945 5871 26979
rect 5813 26939 5871 26945
rect 3927 26880 4752 26908
rect 3927 26877 3939 26880
rect 3881 26871 3939 26877
rect 5368 26840 5396 26939
rect 5902 26936 5908 26988
rect 5960 26936 5966 26988
rect 6086 26936 6092 26988
rect 6144 26936 6150 26988
rect 6178 26936 6184 26988
rect 6236 26936 6242 26988
rect 6589 26985 6617 27016
rect 6914 27004 6920 27016
rect 6972 27004 6978 27056
rect 6552 26979 6617 26985
rect 6552 26945 6564 26979
rect 6598 26946 6617 26979
rect 7009 26979 7067 26985
rect 7009 26976 7021 26979
rect 6932 26948 7021 26976
rect 6598 26945 6610 26946
rect 6552 26939 6610 26945
rect 6932 26920 6960 26948
rect 7009 26945 7021 26948
rect 7055 26945 7067 26979
rect 7009 26939 7067 26945
rect 7208 26920 7236 27084
rect 7558 27004 7564 27056
rect 7616 27044 7622 27056
rect 7616 27016 7788 27044
rect 7616 27004 7622 27016
rect 7282 26936 7288 26988
rect 7340 26976 7346 26988
rect 7340 26948 7604 26976
rect 7340 26936 7346 26948
rect 5534 26868 5540 26920
rect 5592 26868 5598 26920
rect 6638 26868 6644 26920
rect 6696 26868 6702 26920
rect 6914 26868 6920 26920
rect 6972 26868 6978 26920
rect 7190 26868 7196 26920
rect 7248 26908 7254 26920
rect 7377 26911 7435 26917
rect 7377 26908 7389 26911
rect 7248 26880 7389 26908
rect 7248 26868 7254 26880
rect 7377 26877 7389 26880
rect 7423 26877 7435 26911
rect 7576 26908 7604 26948
rect 7650 26936 7656 26988
rect 7708 26936 7714 26988
rect 7760 26985 7788 27016
rect 7745 26979 7803 26985
rect 7745 26945 7757 26979
rect 7791 26945 7803 26979
rect 7745 26939 7803 26945
rect 7837 26979 7895 26985
rect 7837 26945 7849 26979
rect 7883 26945 7895 26979
rect 7944 26976 7972 27084
rect 8202 27072 8208 27124
rect 8260 27072 8266 27124
rect 8849 27115 8907 27121
rect 8849 27081 8861 27115
rect 8895 27081 8907 27115
rect 8849 27075 8907 27081
rect 8864 27044 8892 27075
rect 12434 27072 12440 27124
rect 12492 27112 12498 27124
rect 14277 27115 14335 27121
rect 14277 27112 14289 27115
rect 12492 27084 14289 27112
rect 12492 27072 12498 27084
rect 14277 27081 14289 27084
rect 14323 27081 14335 27115
rect 14277 27075 14335 27081
rect 15289 27115 15347 27121
rect 15289 27081 15301 27115
rect 15335 27112 15347 27115
rect 15746 27112 15752 27124
rect 15335 27084 15752 27112
rect 15335 27081 15347 27084
rect 15289 27075 15347 27081
rect 15746 27072 15752 27084
rect 15804 27072 15810 27124
rect 17494 27112 17500 27124
rect 17420 27084 17500 27112
rect 9217 27047 9275 27053
rect 9217 27044 9229 27047
rect 8864 27016 9229 27044
rect 9217 27013 9229 27016
rect 9263 27013 9275 27047
rect 9217 27007 9275 27013
rect 9858 27004 9864 27056
rect 9916 27004 9922 27056
rect 12986 27004 12992 27056
rect 13044 27004 13050 27056
rect 13630 27004 13636 27056
rect 13688 27044 13694 27056
rect 14090 27044 14096 27056
rect 13688 27016 14096 27044
rect 13688 27004 13694 27016
rect 14090 27004 14096 27016
rect 14148 27004 14154 27056
rect 8021 26979 8079 26985
rect 8021 26976 8033 26979
rect 7944 26948 8033 26976
rect 7837 26939 7895 26945
rect 8021 26945 8033 26948
rect 8067 26945 8079 26979
rect 8021 26939 8079 26945
rect 7852 26908 7880 26939
rect 8662 26936 8668 26988
rect 8720 26936 8726 26988
rect 15378 26936 15384 26988
rect 15436 26936 15442 26988
rect 16390 26936 16396 26988
rect 16448 26936 16454 26988
rect 16942 26936 16948 26988
rect 17000 26976 17006 26988
rect 17420 26985 17448 27084
rect 17494 27072 17500 27084
rect 17552 27072 17558 27124
rect 18046 27072 18052 27124
rect 18104 27072 18110 27124
rect 19242 27072 19248 27124
rect 19300 27072 19306 27124
rect 19426 27072 19432 27124
rect 19484 27112 19490 27124
rect 22554 27112 22560 27124
rect 19484 27084 22560 27112
rect 19484 27072 19490 27084
rect 22554 27072 22560 27084
rect 22612 27112 22618 27124
rect 25130 27112 25136 27124
rect 22612 27084 25136 27112
rect 22612 27072 22618 27084
rect 25130 27072 25136 27084
rect 25188 27072 25194 27124
rect 25222 27072 25228 27124
rect 25280 27072 25286 27124
rect 25590 27072 25596 27124
rect 25648 27112 25654 27124
rect 26145 27115 26203 27121
rect 26145 27112 26157 27115
rect 25648 27084 26157 27112
rect 25648 27072 25654 27084
rect 26145 27081 26157 27084
rect 26191 27081 26203 27115
rect 26145 27075 26203 27081
rect 27062 27072 27068 27124
rect 27120 27072 27126 27124
rect 27246 27072 27252 27124
rect 27304 27072 27310 27124
rect 27430 27072 27436 27124
rect 27488 27112 27494 27124
rect 27617 27115 27675 27121
rect 27617 27112 27629 27115
rect 27488 27084 27629 27112
rect 27488 27072 27494 27084
rect 27617 27081 27629 27084
rect 27663 27081 27675 27115
rect 27617 27075 27675 27081
rect 28350 27072 28356 27124
rect 28408 27072 28414 27124
rect 30837 27115 30895 27121
rect 29764 27084 30788 27112
rect 17221 26979 17279 26985
rect 17221 26976 17233 26979
rect 17000 26948 17233 26976
rect 17000 26936 17006 26948
rect 17221 26945 17233 26948
rect 17267 26945 17279 26979
rect 17221 26939 17279 26945
rect 17405 26979 17463 26985
rect 17405 26945 17417 26979
rect 17451 26945 17463 26979
rect 17405 26939 17463 26945
rect 17497 26979 17555 26985
rect 17497 26945 17509 26979
rect 17543 26945 17555 26979
rect 17497 26939 17555 26945
rect 17681 26979 17739 26985
rect 17681 26945 17693 26979
rect 17727 26976 17739 26979
rect 18064 26976 18092 27072
rect 25685 27047 25743 27053
rect 17727 26948 18092 26976
rect 18708 27016 24992 27044
rect 17727 26945 17739 26948
rect 17681 26939 17739 26945
rect 7576 26880 7880 26908
rect 8941 26911 8999 26917
rect 7377 26871 7435 26877
rect 8941 26877 8953 26911
rect 8987 26877 8999 26911
rect 8941 26871 8999 26877
rect 4632 26812 5396 26840
rect 5552 26840 5580 26868
rect 8018 26840 8024 26852
rect 5552 26812 8024 26840
rect 4632 26784 4660 26812
rect 8018 26800 8024 26812
rect 8076 26840 8082 26852
rect 8956 26840 8984 26871
rect 12802 26868 12808 26920
rect 12860 26908 12866 26920
rect 14182 26908 14188 26920
rect 12860 26880 14188 26908
rect 12860 26868 12866 26880
rect 14182 26868 14188 26880
rect 14240 26908 14246 26920
rect 15473 26911 15531 26917
rect 15473 26908 15485 26911
rect 14240 26880 15485 26908
rect 14240 26868 14246 26880
rect 15473 26877 15485 26880
rect 15519 26877 15531 26911
rect 17512 26908 17540 26939
rect 18506 26908 18512 26920
rect 17512 26880 18512 26908
rect 15473 26871 15531 26877
rect 18506 26868 18512 26880
rect 18564 26868 18570 26920
rect 8076 26812 8984 26840
rect 10689 26843 10747 26849
rect 8076 26800 8082 26812
rect 10689 26809 10701 26843
rect 10735 26840 10747 26843
rect 18708 26840 18736 27016
rect 19426 26936 19432 26988
rect 19484 26936 19490 26988
rect 19518 26936 19524 26988
rect 19576 26936 19582 26988
rect 19610 26936 19616 26988
rect 19668 26936 19674 26988
rect 19794 26936 19800 26988
rect 19852 26936 19858 26988
rect 20622 26976 20628 26988
rect 19904 26948 20628 26976
rect 18782 26868 18788 26920
rect 18840 26908 18846 26920
rect 19904 26908 19932 26948
rect 20622 26936 20628 26948
rect 20680 26936 20686 26988
rect 20714 26936 20720 26988
rect 20772 26936 20778 26988
rect 22922 26936 22928 26988
rect 22980 26936 22986 26988
rect 23014 26936 23020 26988
rect 23072 26976 23078 26988
rect 23109 26979 23167 26985
rect 23109 26976 23121 26979
rect 23072 26948 23121 26976
rect 23072 26936 23078 26948
rect 23109 26945 23121 26948
rect 23155 26945 23167 26979
rect 23109 26939 23167 26945
rect 24489 26979 24547 26985
rect 24489 26945 24501 26979
rect 24535 26945 24547 26979
rect 24489 26939 24547 26945
rect 18840 26880 19932 26908
rect 18840 26868 18846 26880
rect 20070 26868 20076 26920
rect 20128 26908 20134 26920
rect 20809 26911 20867 26917
rect 20809 26908 20821 26911
rect 20128 26880 20821 26908
rect 20128 26868 20134 26880
rect 20809 26877 20821 26880
rect 20855 26908 20867 26911
rect 24504 26908 24532 26939
rect 24578 26936 24584 26988
rect 24636 26936 24642 26988
rect 24762 26976 24768 26988
rect 24688 26948 24768 26976
rect 24688 26908 24716 26948
rect 24762 26936 24768 26948
rect 24820 26936 24826 26988
rect 24857 26979 24915 26985
rect 24857 26945 24869 26979
rect 24903 26945 24915 26979
rect 24857 26939 24915 26945
rect 20855 26880 21956 26908
rect 24504 26880 24716 26908
rect 20855 26877 20867 26880
rect 20809 26871 20867 26877
rect 10735 26812 18736 26840
rect 10735 26809 10747 26812
rect 10689 26803 10747 26809
rect 4062 26732 4068 26784
rect 4120 26732 4126 26784
rect 4614 26732 4620 26784
rect 4672 26732 4678 26784
rect 4798 26732 4804 26784
rect 4856 26732 4862 26784
rect 5258 26732 5264 26784
rect 5316 26732 5322 26784
rect 5902 26732 5908 26784
rect 5960 26772 5966 26784
rect 6365 26775 6423 26781
rect 6365 26772 6377 26775
rect 5960 26744 6377 26772
rect 5960 26732 5966 26744
rect 6365 26741 6377 26744
rect 6411 26741 6423 26775
rect 6365 26735 6423 26741
rect 6822 26732 6828 26784
rect 6880 26732 6886 26784
rect 7282 26732 7288 26784
rect 7340 26732 7346 26784
rect 7650 26732 7656 26784
rect 7708 26772 7714 26784
rect 8202 26772 8208 26784
rect 7708 26744 8208 26772
rect 7708 26732 7714 26744
rect 8202 26732 8208 26744
rect 8260 26772 8266 26784
rect 9306 26772 9312 26784
rect 8260 26744 9312 26772
rect 8260 26732 8266 26744
rect 9306 26732 9312 26744
rect 9364 26732 9370 26784
rect 9398 26732 9404 26784
rect 9456 26772 9462 26784
rect 10704 26772 10732 26803
rect 9456 26744 10732 26772
rect 9456 26732 9462 26744
rect 14918 26732 14924 26784
rect 14976 26732 14982 26784
rect 16298 26732 16304 26784
rect 16356 26732 16362 26784
rect 17313 26775 17371 26781
rect 17313 26741 17325 26775
rect 17359 26772 17371 26775
rect 17770 26772 17776 26784
rect 17359 26744 17776 26772
rect 17359 26741 17371 26744
rect 17313 26735 17371 26741
rect 17770 26732 17776 26744
rect 17828 26732 17834 26784
rect 20990 26732 20996 26784
rect 21048 26732 21054 26784
rect 21928 26772 21956 26880
rect 23017 26843 23075 26849
rect 23017 26809 23029 26843
rect 23063 26840 23075 26843
rect 23106 26840 23112 26852
rect 23063 26812 23112 26840
rect 23063 26809 23075 26812
rect 23017 26803 23075 26809
rect 23106 26800 23112 26812
rect 23164 26800 23170 26852
rect 24118 26772 24124 26784
rect 21928 26744 24124 26772
rect 24118 26732 24124 26744
rect 24176 26732 24182 26784
rect 24688 26772 24716 26880
rect 24872 26840 24900 26939
rect 24964 26908 24992 27016
rect 25685 27013 25697 27047
rect 25731 27044 25743 27047
rect 25866 27044 25872 27056
rect 25731 27016 25872 27044
rect 25731 27013 25743 27016
rect 25685 27007 25743 27013
rect 25866 27004 25872 27016
rect 25924 27004 25930 27056
rect 27080 27044 27108 27072
rect 26620 27016 27108 27044
rect 27264 27044 27292 27072
rect 28718 27044 28724 27056
rect 27264 27016 27384 27044
rect 26620 26988 26648 27016
rect 25041 26979 25099 26985
rect 25041 26945 25053 26979
rect 25087 26976 25099 26979
rect 25130 26976 25136 26988
rect 25087 26948 25136 26976
rect 25087 26945 25099 26948
rect 25041 26939 25099 26945
rect 25130 26936 25136 26948
rect 25188 26936 25194 26988
rect 25222 26936 25228 26988
rect 25280 26936 25286 26988
rect 25501 26979 25559 26985
rect 25501 26945 25513 26979
rect 25547 26976 25559 26979
rect 25777 26979 25835 26985
rect 25777 26976 25789 26979
rect 25547 26948 25789 26976
rect 25547 26945 25559 26948
rect 25501 26939 25559 26945
rect 25777 26945 25789 26948
rect 25823 26945 25835 26979
rect 25777 26939 25835 26945
rect 25248 26908 25276 26936
rect 24964 26880 25276 26908
rect 25317 26911 25375 26917
rect 25317 26877 25329 26911
rect 25363 26877 25375 26911
rect 25792 26908 25820 26939
rect 25958 26936 25964 26988
rect 26016 26936 26022 26988
rect 26602 26936 26608 26988
rect 26660 26936 26666 26988
rect 26786 26936 26792 26988
rect 26844 26936 26850 26988
rect 27065 26979 27123 26985
rect 27065 26945 27077 26979
rect 27111 26945 27123 26979
rect 27065 26939 27123 26945
rect 27157 26979 27215 26985
rect 27157 26945 27169 26979
rect 27203 26976 27215 26979
rect 27246 26976 27252 26988
rect 27203 26948 27252 26976
rect 27203 26945 27215 26948
rect 27157 26939 27215 26945
rect 26697 26911 26755 26917
rect 25792 26880 26188 26908
rect 25317 26871 25375 26877
rect 25130 26840 25136 26852
rect 24872 26812 25136 26840
rect 25130 26800 25136 26812
rect 25188 26800 25194 26852
rect 25222 26772 25228 26784
rect 24688 26744 25228 26772
rect 25222 26732 25228 26744
rect 25280 26732 25286 26784
rect 25332 26772 25360 26871
rect 26160 26784 26188 26880
rect 26697 26877 26709 26911
rect 26743 26908 26755 26911
rect 27080 26908 27108 26939
rect 27246 26936 27252 26948
rect 27304 26936 27310 26988
rect 27356 26985 27384 27016
rect 27448 27016 28724 27044
rect 27448 26985 27476 27016
rect 28718 27004 28724 27016
rect 28776 27004 28782 27056
rect 29764 27044 29792 27084
rect 28828 27016 29792 27044
rect 27341 26979 27399 26985
rect 27341 26945 27353 26979
rect 27387 26945 27399 26979
rect 27341 26939 27399 26945
rect 27433 26979 27491 26985
rect 27433 26945 27445 26979
rect 27479 26945 27491 26979
rect 27433 26939 27491 26945
rect 26743 26880 27108 26908
rect 27356 26908 27384 26939
rect 27706 26936 27712 26988
rect 27764 26936 27770 26988
rect 27890 26936 27896 26988
rect 27948 26936 27954 26988
rect 27982 26936 27988 26988
rect 28040 26936 28046 26988
rect 28077 26979 28135 26985
rect 28077 26945 28089 26979
rect 28123 26945 28135 26979
rect 28077 26939 28135 26945
rect 28092 26908 28120 26939
rect 27356 26880 28120 26908
rect 26743 26877 26755 26880
rect 26697 26871 26755 26877
rect 27080 26840 27108 26880
rect 27154 26840 27160 26852
rect 27080 26812 27160 26840
rect 27154 26800 27160 26812
rect 27212 26800 27218 26852
rect 27982 26800 27988 26852
rect 28040 26840 28046 26852
rect 28828 26840 28856 27016
rect 29178 26936 29184 26988
rect 29236 26976 29242 26988
rect 29764 26985 29792 27016
rect 30006 27004 30012 27056
rect 30064 27004 30070 27056
rect 30101 27047 30159 27053
rect 30101 27013 30113 27047
rect 30147 27044 30159 27047
rect 30760 27044 30788 27084
rect 30837 27081 30849 27115
rect 30883 27112 30895 27115
rect 31294 27112 31300 27124
rect 30883 27084 31300 27112
rect 30883 27081 30895 27084
rect 30837 27075 30895 27081
rect 31294 27072 31300 27084
rect 31352 27072 31358 27124
rect 31757 27115 31815 27121
rect 31757 27081 31769 27115
rect 31803 27112 31815 27115
rect 32122 27112 32128 27124
rect 31803 27084 32128 27112
rect 31803 27081 31815 27084
rect 31757 27075 31815 27081
rect 32122 27072 32128 27084
rect 32180 27072 32186 27124
rect 34882 27072 34888 27124
rect 34940 27112 34946 27124
rect 36265 27115 36323 27121
rect 34940 27084 35480 27112
rect 34940 27072 34946 27084
rect 32953 27047 33011 27053
rect 30147 27016 30420 27044
rect 30760 27016 31340 27044
rect 30147 27013 30159 27016
rect 30101 27007 30159 27013
rect 29365 26979 29423 26985
rect 29365 26976 29377 26979
rect 29236 26948 29377 26976
rect 29236 26936 29242 26948
rect 29365 26945 29377 26948
rect 29411 26945 29423 26979
rect 29365 26939 29423 26945
rect 29549 26979 29607 26985
rect 29549 26945 29561 26979
rect 29595 26945 29607 26979
rect 29549 26939 29607 26945
rect 29733 26979 29792 26985
rect 29733 26945 29745 26979
rect 29779 26948 29792 26979
rect 29917 26979 29975 26985
rect 29779 26945 29791 26948
rect 29733 26939 29791 26945
rect 29917 26945 29929 26979
rect 29963 26976 29975 26979
rect 30024 26976 30052 27004
rect 29963 26948 30052 26976
rect 29963 26945 29975 26948
rect 29917 26939 29975 26945
rect 29564 26908 29592 26939
rect 30190 26936 30196 26988
rect 30248 26936 30254 26988
rect 30392 26985 30420 27016
rect 30377 26979 30435 26985
rect 30377 26945 30389 26979
rect 30423 26945 30435 26979
rect 30377 26939 30435 26945
rect 30466 26936 30472 26988
rect 30524 26936 30530 26988
rect 30561 26979 30619 26985
rect 30561 26945 30573 26979
rect 30607 26945 30619 26979
rect 30561 26939 30619 26945
rect 28040 26812 28856 26840
rect 28920 26880 29592 26908
rect 28040 26800 28046 26812
rect 25866 26772 25872 26784
rect 25332 26744 25872 26772
rect 25866 26732 25872 26744
rect 25924 26732 25930 26784
rect 26142 26732 26148 26784
rect 26200 26732 26206 26784
rect 27430 26732 27436 26784
rect 27488 26772 27494 26784
rect 28920 26772 28948 26880
rect 27488 26744 28948 26772
rect 29564 26772 29592 26880
rect 29641 26911 29699 26917
rect 29641 26877 29653 26911
rect 29687 26877 29699 26911
rect 29641 26871 29699 26877
rect 29656 26840 29684 26871
rect 30282 26868 30288 26920
rect 30340 26908 30346 26920
rect 30576 26908 30604 26939
rect 30926 26936 30932 26988
rect 30984 26976 30990 26988
rect 31312 26985 31340 27016
rect 32953 27013 32965 27047
rect 32999 27044 33011 27047
rect 33965 27047 34023 27053
rect 32999 27016 33732 27044
rect 32999 27013 33011 27016
rect 32953 27007 33011 27013
rect 31113 26979 31171 26985
rect 31113 26976 31125 26979
rect 30984 26948 31125 26976
rect 30984 26936 30990 26948
rect 31113 26945 31125 26948
rect 31159 26945 31171 26979
rect 31113 26939 31171 26945
rect 31297 26979 31355 26985
rect 31297 26945 31309 26979
rect 31343 26945 31355 26979
rect 31297 26939 31355 26945
rect 30340 26880 30604 26908
rect 30340 26868 30346 26880
rect 30742 26840 30748 26852
rect 29656 26812 30748 26840
rect 30576 26784 30604 26812
rect 30742 26800 30748 26812
rect 30800 26800 30806 26852
rect 31312 26840 31340 26939
rect 31570 26936 31576 26988
rect 31628 26936 31634 26988
rect 32398 26936 32404 26988
rect 32456 26976 32462 26988
rect 33137 26979 33195 26985
rect 33137 26976 33149 26979
rect 32456 26948 33149 26976
rect 32456 26936 32462 26948
rect 32784 26920 32812 26948
rect 33137 26945 33149 26948
rect 33183 26945 33195 26979
rect 33137 26939 33195 26945
rect 33226 26936 33232 26988
rect 33284 26936 33290 26988
rect 33704 26985 33732 27016
rect 33965 27013 33977 27047
rect 34011 27044 34023 27047
rect 34422 27044 34428 27056
rect 34011 27016 34428 27044
rect 34011 27013 34023 27016
rect 33965 27007 34023 27013
rect 34422 27004 34428 27016
rect 34480 27004 34486 27056
rect 35069 27047 35127 27053
rect 35069 27044 35081 27047
rect 34624 27016 35081 27044
rect 33689 26979 33747 26985
rect 33689 26945 33701 26979
rect 33735 26945 33747 26979
rect 33689 26939 33747 26945
rect 33778 26936 33784 26988
rect 33836 26936 33842 26988
rect 34054 26936 34060 26988
rect 34112 26936 34118 26988
rect 34195 26979 34253 26985
rect 34195 26945 34207 26979
rect 34241 26976 34253 26979
rect 34624 26976 34652 27016
rect 35069 27013 35081 27016
rect 35115 27013 35127 27047
rect 35069 27007 35127 27013
rect 35452 26988 35480 27084
rect 36265 27081 36277 27115
rect 36311 27112 36323 27115
rect 36538 27112 36544 27124
rect 36311 27084 36544 27112
rect 36311 27081 36323 27084
rect 36265 27075 36323 27081
rect 36538 27072 36544 27084
rect 36596 27112 36602 27124
rect 36596 27084 36860 27112
rect 36596 27072 36602 27084
rect 36081 27047 36139 27053
rect 36081 27013 36093 27047
rect 36127 27044 36139 27047
rect 36170 27044 36176 27056
rect 36127 27016 36176 27044
rect 36127 27013 36139 27016
rect 36081 27007 36139 27013
rect 36170 27004 36176 27016
rect 36228 27044 36234 27056
rect 36630 27044 36636 27056
rect 36228 27016 36636 27044
rect 36228 27004 36234 27016
rect 36630 27004 36636 27016
rect 36688 27004 36694 27056
rect 36722 27004 36728 27056
rect 36780 27004 36786 27056
rect 36832 26988 36860 27084
rect 34241 26948 34652 26976
rect 34241 26945 34253 26948
rect 34195 26939 34253 26945
rect 34698 26936 34704 26988
rect 34756 26936 34762 26988
rect 34977 26979 35035 26985
rect 34977 26945 34989 26979
rect 35023 26976 35035 26979
rect 35253 26979 35311 26985
rect 35023 26948 35204 26976
rect 35023 26945 35035 26948
rect 34977 26939 35035 26945
rect 32766 26868 32772 26920
rect 32824 26868 32830 26920
rect 32950 26868 32956 26920
rect 33008 26868 33014 26920
rect 34072 26908 34100 26936
rect 34072 26880 35020 26908
rect 34333 26843 34391 26849
rect 31312 26812 33180 26840
rect 33152 26784 33180 26812
rect 34333 26809 34345 26843
rect 34379 26840 34391 26843
rect 34885 26843 34943 26849
rect 34885 26840 34897 26843
rect 34379 26812 34897 26840
rect 34379 26809 34391 26812
rect 34333 26803 34391 26809
rect 34885 26809 34897 26812
rect 34931 26809 34943 26843
rect 34885 26803 34943 26809
rect 30374 26772 30380 26784
rect 29564 26744 30380 26772
rect 27488 26732 27494 26744
rect 30374 26732 30380 26744
rect 30432 26732 30438 26784
rect 30558 26732 30564 26784
rect 30616 26732 30622 26784
rect 33134 26732 33140 26784
rect 33192 26732 33198 26784
rect 33410 26732 33416 26784
rect 33468 26772 33474 26784
rect 34517 26775 34575 26781
rect 34517 26772 34529 26775
rect 33468 26744 34529 26772
rect 33468 26732 33474 26744
rect 34517 26741 34529 26744
rect 34563 26741 34575 26775
rect 34992 26772 35020 26880
rect 35176 26840 35204 26948
rect 35253 26945 35265 26979
rect 35299 26976 35311 26979
rect 35342 26976 35348 26988
rect 35299 26948 35348 26976
rect 35299 26945 35311 26948
rect 35253 26939 35311 26945
rect 35342 26936 35348 26948
rect 35400 26936 35406 26988
rect 35434 26936 35440 26988
rect 35492 26976 35498 26988
rect 35621 26979 35679 26985
rect 35621 26976 35633 26979
rect 35492 26948 35633 26976
rect 35492 26936 35498 26948
rect 35621 26945 35633 26948
rect 35667 26945 35679 26979
rect 35621 26939 35679 26945
rect 35805 26979 35863 26985
rect 35805 26945 35817 26979
rect 35851 26976 35863 26979
rect 36357 26979 36415 26985
rect 35851 26948 35885 26976
rect 35851 26945 35863 26948
rect 35805 26939 35863 26945
rect 36357 26945 36369 26979
rect 36403 26976 36415 26979
rect 36541 26979 36599 26985
rect 36541 26976 36553 26979
rect 36403 26948 36553 26976
rect 36403 26945 36415 26948
rect 36357 26939 36415 26945
rect 36541 26945 36553 26948
rect 36587 26945 36599 26979
rect 36541 26939 36599 26945
rect 35529 26911 35587 26917
rect 35529 26877 35541 26911
rect 35575 26908 35587 26911
rect 35820 26908 35848 26939
rect 36814 26936 36820 26988
rect 36872 26936 36878 26988
rect 36909 26979 36967 26985
rect 36909 26945 36921 26979
rect 36955 26976 36967 26979
rect 36955 26948 37044 26976
rect 36955 26945 36967 26948
rect 36909 26939 36967 26945
rect 35986 26908 35992 26920
rect 35575 26880 35992 26908
rect 35575 26877 35587 26880
rect 35529 26871 35587 26877
rect 35986 26868 35992 26880
rect 36044 26868 36050 26920
rect 36081 26843 36139 26849
rect 36081 26840 36093 26843
rect 35176 26812 36093 26840
rect 36081 26809 36093 26812
rect 36127 26809 36139 26843
rect 36081 26803 36139 26809
rect 37016 26784 37044 26948
rect 35713 26775 35771 26781
rect 35713 26772 35725 26775
rect 34992 26744 35725 26772
rect 34517 26735 34575 26741
rect 35713 26741 35725 26744
rect 35759 26741 35771 26775
rect 35713 26735 35771 26741
rect 36998 26732 37004 26784
rect 37056 26732 37062 26784
rect 1104 26682 38272 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38272 26682
rect 1104 26608 38272 26630
rect 2130 26568 2136 26580
rect 1412 26540 2136 26568
rect 1412 26444 1440 26540
rect 2130 26528 2136 26540
rect 2188 26568 2194 26580
rect 5534 26568 5540 26580
rect 2188 26540 5540 26568
rect 2188 26528 2194 26540
rect 5534 26528 5540 26540
rect 5592 26528 5598 26580
rect 6822 26528 6828 26580
rect 6880 26568 6886 26580
rect 7193 26571 7251 26577
rect 7193 26568 7205 26571
rect 6880 26540 7205 26568
rect 6880 26528 6886 26540
rect 7193 26537 7205 26540
rect 7239 26537 7251 26571
rect 7193 26531 7251 26537
rect 7282 26528 7288 26580
rect 7340 26568 7346 26580
rect 7561 26571 7619 26577
rect 7561 26568 7573 26571
rect 7340 26540 7573 26568
rect 7340 26528 7346 26540
rect 7561 26537 7573 26540
rect 7607 26537 7619 26571
rect 7561 26531 7619 26537
rect 8662 26528 8668 26580
rect 8720 26568 8726 26580
rect 9033 26571 9091 26577
rect 9033 26568 9045 26571
rect 8720 26540 9045 26568
rect 8720 26528 8726 26540
rect 9033 26537 9045 26540
rect 9079 26537 9091 26571
rect 9033 26531 9091 26537
rect 9140 26540 9628 26568
rect 3605 26503 3663 26509
rect 3605 26500 3617 26503
rect 2746 26472 3617 26500
rect 1394 26392 1400 26444
rect 1452 26392 1458 26444
rect 1673 26435 1731 26441
rect 1673 26401 1685 26435
rect 1719 26432 1731 26435
rect 2746 26432 2774 26472
rect 3605 26469 3617 26472
rect 3651 26500 3663 26503
rect 3970 26500 3976 26512
rect 3651 26472 3976 26500
rect 3651 26469 3663 26472
rect 3605 26463 3663 26469
rect 3970 26460 3976 26472
rect 4028 26460 4034 26512
rect 4798 26460 4804 26512
rect 4856 26460 4862 26512
rect 9140 26500 9168 26540
rect 5000 26472 9168 26500
rect 1719 26404 2774 26432
rect 3145 26435 3203 26441
rect 1719 26401 1731 26404
rect 1673 26395 1731 26401
rect 3145 26401 3157 26435
rect 3191 26432 3203 26435
rect 4341 26435 4399 26441
rect 4341 26432 4353 26435
rect 3191 26404 4353 26432
rect 3191 26401 3203 26404
rect 3145 26395 3203 26401
rect 4341 26401 4353 26404
rect 4387 26432 4399 26435
rect 4614 26432 4620 26444
rect 4387 26404 4620 26432
rect 4387 26401 4399 26404
rect 4341 26395 4399 26401
rect 4614 26392 4620 26404
rect 4672 26392 4678 26444
rect 2774 26324 2780 26376
rect 2832 26324 2838 26376
rect 3421 26367 3479 26373
rect 3421 26333 3433 26367
rect 3467 26333 3479 26367
rect 3421 26327 3479 26333
rect 3605 26367 3663 26373
rect 3605 26333 3617 26367
rect 3651 26364 3663 26367
rect 4816 26364 4844 26460
rect 4893 26367 4951 26373
rect 4893 26364 4905 26367
rect 3651 26336 4476 26364
rect 4816 26336 4905 26364
rect 3651 26333 3663 26336
rect 3605 26327 3663 26333
rect 3436 26296 3464 26327
rect 3789 26299 3847 26305
rect 3789 26296 3801 26299
rect 3436 26268 3801 26296
rect 3789 26265 3801 26268
rect 3835 26265 3847 26299
rect 3789 26259 3847 26265
rect 4448 26228 4476 26336
rect 4893 26333 4905 26336
rect 4939 26333 4951 26367
rect 4893 26327 4951 26333
rect 4522 26256 4528 26308
rect 4580 26296 4586 26308
rect 5000 26296 5028 26472
rect 9398 26460 9404 26512
rect 9456 26460 9462 26512
rect 7006 26392 7012 26444
rect 7064 26392 7070 26444
rect 8018 26392 8024 26444
rect 8076 26392 8082 26444
rect 9416 26432 9444 26460
rect 9493 26435 9551 26441
rect 9493 26432 9505 26435
rect 9416 26404 9505 26432
rect 9493 26401 9505 26404
rect 9539 26401 9551 26435
rect 9600 26432 9628 26540
rect 11238 26528 11244 26580
rect 11296 26528 11302 26580
rect 13170 26528 13176 26580
rect 13228 26528 13234 26580
rect 13262 26528 13268 26580
rect 13320 26528 13326 26580
rect 15562 26528 15568 26580
rect 15620 26568 15626 26580
rect 15841 26571 15899 26577
rect 15841 26568 15853 26571
rect 15620 26540 15853 26568
rect 15620 26528 15626 26540
rect 15841 26537 15853 26540
rect 15887 26537 15899 26571
rect 19334 26568 19340 26580
rect 15841 26531 15899 26537
rect 16224 26540 19340 26568
rect 9677 26435 9735 26441
rect 9677 26432 9689 26435
rect 9600 26404 9689 26432
rect 9493 26395 9551 26401
rect 9677 26401 9689 26404
rect 9723 26432 9735 26435
rect 10410 26432 10416 26444
rect 9723 26404 10416 26432
rect 9723 26401 9735 26404
rect 9677 26395 9735 26401
rect 10410 26392 10416 26404
rect 10468 26392 10474 26444
rect 11256 26432 11284 26528
rect 11793 26435 11851 26441
rect 11793 26432 11805 26435
rect 11256 26404 11805 26432
rect 11793 26401 11805 26404
rect 11839 26401 11851 26435
rect 11793 26395 11851 26401
rect 12250 26392 12256 26444
rect 12308 26432 12314 26444
rect 12434 26432 12440 26444
rect 12308 26404 12440 26432
rect 12308 26392 12314 26404
rect 12434 26392 12440 26404
rect 12492 26392 12498 26444
rect 7024 26364 7052 26392
rect 7101 26367 7159 26373
rect 7101 26364 7113 26367
rect 7024 26336 7113 26364
rect 7101 26333 7113 26336
rect 7147 26333 7159 26367
rect 7101 26327 7159 26333
rect 7466 26324 7472 26376
rect 7524 26324 7530 26376
rect 8036 26364 8064 26392
rect 11517 26367 11575 26373
rect 11517 26364 11529 26367
rect 8036 26336 11529 26364
rect 11517 26333 11529 26336
rect 11563 26333 11575 26367
rect 13188 26364 13216 26528
rect 14090 26460 14096 26512
rect 14148 26500 14154 26512
rect 16224 26500 16252 26540
rect 19334 26528 19340 26540
rect 19392 26568 19398 26580
rect 20622 26568 20628 26580
rect 19392 26540 20628 26568
rect 19392 26528 19398 26540
rect 20622 26528 20628 26540
rect 20680 26528 20686 26580
rect 20990 26528 20996 26580
rect 21048 26528 21054 26580
rect 22557 26571 22615 26577
rect 21468 26540 22508 26568
rect 14148 26472 16252 26500
rect 16301 26503 16359 26509
rect 14148 26460 14154 26472
rect 14384 26441 14412 26472
rect 16301 26469 16313 26503
rect 16347 26500 16359 26503
rect 16850 26500 16856 26512
rect 16347 26472 16856 26500
rect 16347 26469 16359 26472
rect 16301 26463 16359 26469
rect 16850 26460 16856 26472
rect 16908 26460 16914 26512
rect 16942 26460 16948 26512
rect 17000 26500 17006 26512
rect 17037 26503 17095 26509
rect 17037 26500 17049 26503
rect 17000 26472 17049 26500
rect 17000 26460 17006 26472
rect 17037 26469 17049 26472
rect 17083 26500 17095 26503
rect 17083 26472 17264 26500
rect 17083 26469 17095 26472
rect 17037 26463 17095 26469
rect 14369 26435 14427 26441
rect 14369 26401 14381 26435
rect 14415 26401 14427 26435
rect 14369 26395 14427 26401
rect 15194 26392 15200 26444
rect 15252 26432 15258 26444
rect 15933 26435 15991 26441
rect 15933 26432 15945 26435
rect 15252 26404 15945 26432
rect 15252 26392 15258 26404
rect 15933 26401 15945 26404
rect 15979 26432 15991 26435
rect 16022 26432 16028 26444
rect 15979 26404 16028 26432
rect 15979 26401 15991 26404
rect 15933 26395 15991 26401
rect 16022 26392 16028 26404
rect 16080 26392 16086 26444
rect 17236 26441 17264 26472
rect 17310 26460 17316 26512
rect 17368 26500 17374 26512
rect 18233 26503 18291 26509
rect 18233 26500 18245 26503
rect 17368 26472 18245 26500
rect 17368 26460 17374 26472
rect 18233 26469 18245 26472
rect 18279 26469 18291 26503
rect 18233 26463 18291 26469
rect 17221 26435 17279 26441
rect 17221 26401 17233 26435
rect 17267 26401 17279 26435
rect 17221 26395 17279 26401
rect 18322 26392 18328 26444
rect 18380 26392 18386 26444
rect 21008 26432 21036 26528
rect 21269 26435 21327 26441
rect 21269 26432 21281 26435
rect 21008 26404 21281 26432
rect 21269 26401 21281 26404
rect 21315 26401 21327 26435
rect 21269 26395 21327 26401
rect 14093 26367 14151 26373
rect 14093 26364 14105 26367
rect 13188 26336 14105 26364
rect 11517 26327 11575 26333
rect 14093 26333 14105 26336
rect 14139 26333 14151 26367
rect 14093 26327 14151 26333
rect 15010 26324 15016 26376
rect 15068 26364 15074 26376
rect 16117 26367 16175 26373
rect 16117 26364 16129 26367
rect 15068 26336 16129 26364
rect 15068 26324 15074 26336
rect 16117 26333 16129 26336
rect 16163 26333 16175 26367
rect 16117 26327 16175 26333
rect 16298 26324 16304 26376
rect 16356 26324 16362 26376
rect 16945 26367 17003 26373
rect 16945 26333 16957 26367
rect 16991 26364 17003 26367
rect 17034 26364 17040 26376
rect 16991 26336 17040 26364
rect 16991 26333 17003 26336
rect 16945 26327 17003 26333
rect 17034 26324 17040 26336
rect 17092 26324 17098 26376
rect 17129 26367 17187 26373
rect 17129 26333 17141 26367
rect 17175 26333 17187 26367
rect 17129 26327 17187 26333
rect 4580 26268 5028 26296
rect 7009 26299 7067 26305
rect 4580 26256 4586 26268
rect 7009 26265 7021 26299
rect 7055 26296 7067 26299
rect 7484 26296 7512 26324
rect 7926 26296 7932 26308
rect 7055 26268 7932 26296
rect 7055 26265 7067 26268
rect 7009 26259 7067 26265
rect 7926 26256 7932 26268
rect 7984 26256 7990 26308
rect 9324 26268 9536 26296
rect 5258 26228 5264 26240
rect 4448 26200 5264 26228
rect 5258 26188 5264 26200
rect 5316 26188 5322 26240
rect 6822 26188 6828 26240
rect 6880 26228 6886 26240
rect 9324 26228 9352 26268
rect 6880 26200 9352 26228
rect 6880 26188 6886 26200
rect 9398 26188 9404 26240
rect 9456 26188 9462 26240
rect 9508 26228 9536 26268
rect 9858 26256 9864 26308
rect 9916 26296 9922 26308
rect 12250 26296 12256 26308
rect 9916 26268 12256 26296
rect 9916 26256 9922 26268
rect 12250 26256 12256 26268
rect 12308 26256 12314 26308
rect 15841 26299 15899 26305
rect 15841 26265 15853 26299
rect 15887 26296 15899 26299
rect 16316 26296 16344 26324
rect 15887 26268 16344 26296
rect 15887 26265 15899 26268
rect 15841 26259 15899 26265
rect 16482 26256 16488 26308
rect 16540 26296 16546 26308
rect 17144 26296 17172 26327
rect 17586 26324 17592 26376
rect 17644 26324 17650 26376
rect 17681 26367 17739 26373
rect 17681 26333 17693 26367
rect 17727 26364 17739 26367
rect 18046 26364 18052 26376
rect 17727 26336 18052 26364
rect 17727 26333 17739 26336
rect 17681 26327 17739 26333
rect 18046 26324 18052 26336
rect 18104 26364 18110 26376
rect 18141 26367 18199 26373
rect 18141 26364 18153 26367
rect 18104 26336 18153 26364
rect 18104 26324 18110 26336
rect 18141 26333 18153 26336
rect 18187 26333 18199 26367
rect 18141 26327 18199 26333
rect 18417 26367 18475 26373
rect 18417 26333 18429 26367
rect 18463 26364 18475 26367
rect 18506 26364 18512 26376
rect 18463 26336 18512 26364
rect 18463 26333 18475 26336
rect 18417 26327 18475 26333
rect 18506 26324 18512 26336
rect 18564 26324 18570 26376
rect 21358 26324 21364 26376
rect 21416 26324 21422 26376
rect 16540 26268 20668 26296
rect 16540 26256 16546 26268
rect 17494 26228 17500 26240
rect 9508 26200 17500 26228
rect 17494 26188 17500 26200
rect 17552 26188 17558 26240
rect 17862 26188 17868 26240
rect 17920 26188 17926 26240
rect 17957 26231 18015 26237
rect 17957 26197 17969 26231
rect 18003 26228 18015 26231
rect 18046 26228 18052 26240
rect 18003 26200 18052 26228
rect 18003 26197 18015 26200
rect 17957 26191 18015 26197
rect 18046 26188 18052 26200
rect 18104 26188 18110 26240
rect 20640 26228 20668 26268
rect 20714 26256 20720 26308
rect 20772 26296 20778 26308
rect 21468 26296 21496 26540
rect 21729 26503 21787 26509
rect 21729 26469 21741 26503
rect 21775 26500 21787 26503
rect 22480 26500 22508 26540
rect 22557 26537 22569 26571
rect 22603 26568 22615 26571
rect 22922 26568 22928 26580
rect 22603 26540 22928 26568
rect 22603 26537 22615 26540
rect 22557 26531 22615 26537
rect 22922 26528 22928 26540
rect 22980 26528 22986 26580
rect 24394 26568 24400 26580
rect 23032 26540 24400 26568
rect 23032 26500 23060 26540
rect 24394 26528 24400 26540
rect 24452 26528 24458 26580
rect 24949 26571 25007 26577
rect 24949 26537 24961 26571
rect 24995 26568 25007 26571
rect 25498 26568 25504 26580
rect 24995 26540 25504 26568
rect 24995 26537 25007 26540
rect 24949 26531 25007 26537
rect 25498 26528 25504 26540
rect 25556 26528 25562 26580
rect 25608 26540 27184 26568
rect 21775 26472 22094 26500
rect 22480 26472 23060 26500
rect 21775 26469 21787 26472
rect 21729 26463 21787 26469
rect 22066 26432 22094 26472
rect 23290 26460 23296 26512
rect 23348 26500 23354 26512
rect 23348 26472 23796 26500
rect 23348 26460 23354 26472
rect 22189 26435 22247 26441
rect 22189 26432 22201 26435
rect 22066 26404 22201 26432
rect 22189 26401 22201 26404
rect 22235 26401 22247 26435
rect 22189 26395 22247 26401
rect 23474 26392 23480 26444
rect 23532 26432 23538 26444
rect 23532 26404 23618 26432
rect 23532 26392 23538 26404
rect 22370 26373 22376 26376
rect 22359 26367 22376 26373
rect 22359 26333 22371 26367
rect 22428 26364 22434 26376
rect 23590 26373 23618 26404
rect 23768 26373 23796 26472
rect 23842 26460 23848 26512
rect 23900 26500 23906 26512
rect 24762 26500 24768 26512
rect 23900 26472 24768 26500
rect 23900 26460 23906 26472
rect 24762 26460 24768 26472
rect 24820 26460 24826 26512
rect 25608 26500 25636 26540
rect 26326 26500 26332 26512
rect 25148 26472 25636 26500
rect 25976 26472 26332 26500
rect 23860 26404 25084 26432
rect 23860 26376 23888 26404
rect 25056 26376 25084 26404
rect 23569 26367 23627 26373
rect 22428 26336 22876 26364
rect 22359 26327 22376 26333
rect 22370 26324 22376 26327
rect 22428 26324 22434 26336
rect 22186 26296 22192 26308
rect 20772 26268 21496 26296
rect 21560 26268 22192 26296
rect 20772 26256 20778 26268
rect 21560 26228 21588 26268
rect 22186 26256 22192 26268
rect 22244 26256 22250 26308
rect 22848 26296 22876 26336
rect 23569 26333 23581 26367
rect 23615 26333 23627 26367
rect 23569 26327 23627 26333
rect 23753 26367 23811 26373
rect 23753 26333 23765 26367
rect 23799 26333 23811 26367
rect 23753 26327 23811 26333
rect 23842 26324 23848 26376
rect 23900 26324 23906 26376
rect 23937 26367 23995 26373
rect 23937 26333 23949 26367
rect 23983 26364 23995 26367
rect 23983 26336 24348 26364
rect 23983 26333 23995 26336
rect 23937 26327 23995 26333
rect 23952 26296 23980 26327
rect 22848 26268 23980 26296
rect 24210 26256 24216 26308
rect 24268 26256 24274 26308
rect 24320 26296 24348 26336
rect 25038 26324 25044 26376
rect 25096 26324 25102 26376
rect 25148 26296 25176 26472
rect 25406 26392 25412 26444
rect 25464 26432 25470 26444
rect 25501 26435 25559 26441
rect 25501 26432 25513 26435
rect 25464 26404 25513 26432
rect 25464 26392 25470 26404
rect 25501 26401 25513 26404
rect 25547 26401 25559 26435
rect 25501 26395 25559 26401
rect 25314 26324 25320 26376
rect 25372 26324 25378 26376
rect 25976 26373 26004 26472
rect 26326 26460 26332 26472
rect 26384 26500 26390 26512
rect 26878 26500 26884 26512
rect 26384 26472 26884 26500
rect 26384 26460 26390 26472
rect 26878 26460 26884 26472
rect 26936 26460 26942 26512
rect 26697 26435 26755 26441
rect 26697 26401 26709 26435
rect 26743 26432 26755 26435
rect 27156 26432 27184 26540
rect 27706 26528 27712 26580
rect 27764 26528 27770 26580
rect 27801 26571 27859 26577
rect 27801 26537 27813 26571
rect 27847 26568 27859 26571
rect 27890 26568 27896 26580
rect 27847 26540 27896 26568
rect 27847 26537 27859 26540
rect 27801 26531 27859 26537
rect 27890 26528 27896 26540
rect 27948 26528 27954 26580
rect 28997 26571 29055 26577
rect 28184 26540 28948 26568
rect 27724 26500 27752 26528
rect 28077 26503 28135 26509
rect 28077 26500 28089 26503
rect 27724 26472 28089 26500
rect 28077 26469 28089 26472
rect 28123 26469 28135 26503
rect 28077 26463 28135 26469
rect 28184 26432 28212 26540
rect 28920 26500 28948 26540
rect 28997 26537 29009 26571
rect 29043 26568 29055 26571
rect 29178 26568 29184 26580
rect 29043 26540 29184 26568
rect 29043 26537 29055 26540
rect 28997 26531 29055 26537
rect 29178 26528 29184 26540
rect 29236 26528 29242 26580
rect 29638 26528 29644 26580
rect 29696 26568 29702 26580
rect 29733 26571 29791 26577
rect 29733 26568 29745 26571
rect 29696 26540 29745 26568
rect 29696 26528 29702 26540
rect 29733 26537 29745 26540
rect 29779 26537 29791 26571
rect 29733 26531 29791 26537
rect 29917 26571 29975 26577
rect 29917 26537 29929 26571
rect 29963 26568 29975 26571
rect 30282 26568 30288 26580
rect 29963 26540 30288 26568
rect 29963 26537 29975 26540
rect 29917 26531 29975 26537
rect 30282 26528 30288 26540
rect 30340 26528 30346 26580
rect 32950 26528 32956 26580
rect 33008 26528 33014 26580
rect 33410 26568 33416 26580
rect 33152 26540 33416 26568
rect 33152 26500 33180 26540
rect 33410 26528 33416 26540
rect 33468 26528 33474 26580
rect 34698 26568 34704 26580
rect 34440 26540 34704 26568
rect 34440 26509 34468 26540
rect 34698 26528 34704 26540
rect 34756 26528 34762 26580
rect 35161 26571 35219 26577
rect 35161 26537 35173 26571
rect 35207 26568 35219 26571
rect 35434 26568 35440 26580
rect 35207 26540 35440 26568
rect 35207 26537 35219 26540
rect 35161 26531 35219 26537
rect 35434 26528 35440 26540
rect 35492 26528 35498 26580
rect 36814 26528 36820 26580
rect 36872 26528 36878 26580
rect 36998 26528 37004 26580
rect 37056 26528 37062 26580
rect 26743 26404 27108 26432
rect 27156 26404 28212 26432
rect 28368 26472 28856 26500
rect 28920 26472 33180 26500
rect 34425 26503 34483 26509
rect 26743 26401 26755 26404
rect 26697 26395 26755 26401
rect 25961 26367 26019 26373
rect 25961 26333 25973 26367
rect 26007 26333 26019 26367
rect 25961 26327 26019 26333
rect 26142 26324 26148 26376
rect 26200 26324 26206 26376
rect 26605 26367 26663 26373
rect 26605 26333 26617 26367
rect 26651 26333 26663 26367
rect 26605 26327 26663 26333
rect 26789 26367 26847 26373
rect 26789 26333 26801 26367
rect 26835 26364 26847 26367
rect 26878 26364 26884 26376
rect 26835 26336 26884 26364
rect 26835 26333 26847 26336
rect 26789 26327 26847 26333
rect 24320 26268 25176 26296
rect 25409 26299 25467 26305
rect 25409 26265 25421 26299
rect 25455 26296 25467 26299
rect 25682 26296 25688 26308
rect 25455 26268 25688 26296
rect 25455 26265 25467 26268
rect 25409 26259 25467 26265
rect 25682 26256 25688 26268
rect 25740 26256 25746 26308
rect 26053 26299 26111 26305
rect 26053 26265 26065 26299
rect 26099 26296 26111 26299
rect 26620 26296 26648 26327
rect 26878 26324 26884 26336
rect 26936 26324 26942 26376
rect 27080 26373 27108 26404
rect 27065 26367 27123 26373
rect 27065 26333 27077 26367
rect 27111 26333 27123 26367
rect 27065 26327 27123 26333
rect 27154 26324 27160 26376
rect 27212 26364 27218 26376
rect 27249 26367 27307 26373
rect 27249 26364 27261 26367
rect 27212 26336 27261 26364
rect 27212 26324 27218 26336
rect 27249 26333 27261 26336
rect 27295 26333 27307 26367
rect 27249 26327 27307 26333
rect 27338 26324 27344 26376
rect 27396 26324 27402 26376
rect 27430 26324 27436 26376
rect 27488 26324 27494 26376
rect 27617 26367 27675 26373
rect 27617 26333 27629 26367
rect 27663 26364 27675 26367
rect 28166 26364 28172 26376
rect 27663 26336 28172 26364
rect 27663 26333 27675 26336
rect 27617 26327 27675 26333
rect 28166 26324 28172 26336
rect 28224 26324 28230 26376
rect 27890 26296 27896 26308
rect 26099 26268 26556 26296
rect 26620 26268 27896 26296
rect 26099 26265 26111 26268
rect 26053 26259 26111 26265
rect 20640 26200 21588 26228
rect 26528 26228 26556 26268
rect 27890 26256 27896 26268
rect 27948 26296 27954 26308
rect 28368 26296 28396 26472
rect 28534 26392 28540 26444
rect 28592 26432 28598 26444
rect 28629 26435 28687 26441
rect 28629 26432 28641 26435
rect 28592 26404 28641 26432
rect 28592 26392 28598 26404
rect 28629 26401 28641 26404
rect 28675 26432 28687 26435
rect 28718 26432 28724 26444
rect 28675 26404 28724 26432
rect 28675 26401 28687 26404
rect 28629 26395 28687 26401
rect 28718 26392 28724 26404
rect 28776 26392 28782 26444
rect 28828 26432 28856 26472
rect 34425 26469 34437 26503
rect 34471 26469 34483 26503
rect 36722 26500 36728 26512
rect 34425 26463 34483 26469
rect 36188 26472 36728 26500
rect 31110 26432 31116 26444
rect 28828 26404 31116 26432
rect 28902 26324 28908 26376
rect 28960 26366 28966 26376
rect 29104 26373 29132 26404
rect 31110 26392 31116 26404
rect 31168 26392 31174 26444
rect 32490 26392 32496 26444
rect 32548 26392 32554 26444
rect 32585 26435 32643 26441
rect 32585 26401 32597 26435
rect 32631 26432 32643 26435
rect 32631 26404 33088 26432
rect 32631 26401 32643 26404
rect 32585 26395 32643 26401
rect 29089 26367 29147 26373
rect 28960 26338 29003 26366
rect 28960 26324 28966 26338
rect 29089 26333 29101 26367
rect 29135 26333 29147 26367
rect 29089 26327 29147 26333
rect 29380 26336 29684 26364
rect 29380 26308 29408 26336
rect 27948 26268 28396 26296
rect 28445 26299 28503 26305
rect 27948 26256 27954 26268
rect 28445 26265 28457 26299
rect 28491 26296 28503 26299
rect 28491 26268 28994 26296
rect 28491 26265 28503 26268
rect 28445 26259 28503 26265
rect 27246 26228 27252 26240
rect 26528 26200 27252 26228
rect 27246 26188 27252 26200
rect 27304 26188 27310 26240
rect 28534 26188 28540 26240
rect 28592 26188 28598 26240
rect 28966 26228 28994 26268
rect 29362 26256 29368 26308
rect 29420 26256 29426 26308
rect 29546 26256 29552 26308
rect 29604 26256 29610 26308
rect 29656 26296 29684 26336
rect 32214 26324 32220 26376
rect 32272 26324 32278 26376
rect 32401 26367 32459 26373
rect 32401 26333 32413 26367
rect 32447 26333 32459 26367
rect 32401 26327 32459 26333
rect 32769 26367 32827 26373
rect 32769 26333 32781 26367
rect 32815 26364 32827 26367
rect 32950 26364 32956 26376
rect 32815 26336 32956 26364
rect 32815 26333 32827 26336
rect 32769 26327 32827 26333
rect 29749 26299 29807 26305
rect 29749 26296 29761 26299
rect 29656 26268 29761 26296
rect 29749 26265 29761 26268
rect 29795 26265 29807 26299
rect 29749 26259 29807 26265
rect 32306 26256 32312 26308
rect 32364 26296 32370 26308
rect 32416 26296 32444 26327
rect 32950 26324 32956 26336
rect 33008 26324 33014 26376
rect 33060 26364 33088 26404
rect 33226 26392 33232 26444
rect 33284 26432 33290 26444
rect 36188 26441 36216 26472
rect 36722 26460 36728 26472
rect 36780 26460 36786 26512
rect 34793 26435 34851 26441
rect 34793 26432 34805 26435
rect 33284 26404 34805 26432
rect 33284 26392 33290 26404
rect 34793 26401 34805 26404
rect 34839 26432 34851 26435
rect 36173 26435 36231 26441
rect 36173 26432 36185 26435
rect 34839 26404 36185 26432
rect 34839 26401 34851 26404
rect 34793 26395 34851 26401
rect 36173 26401 36185 26404
rect 36219 26401 36231 26435
rect 36173 26395 36231 26401
rect 36541 26435 36599 26441
rect 36541 26401 36553 26435
rect 36587 26432 36599 26435
rect 36587 26404 37136 26432
rect 36587 26401 36599 26404
rect 36541 26395 36599 26401
rect 33134 26364 33140 26376
rect 33060 26336 33140 26364
rect 33134 26324 33140 26336
rect 33192 26364 33198 26376
rect 33410 26364 33416 26376
rect 33192 26336 33416 26364
rect 33192 26324 33198 26336
rect 33410 26324 33416 26336
rect 33468 26324 33474 26376
rect 34330 26324 34336 26376
rect 34388 26364 34394 26376
rect 34517 26367 34575 26373
rect 34517 26364 34529 26367
rect 34388 26336 34529 26364
rect 34388 26324 34394 26336
rect 34517 26333 34529 26336
rect 34563 26333 34575 26367
rect 34517 26327 34575 26333
rect 34885 26367 34943 26373
rect 34885 26333 34897 26367
rect 34931 26333 34943 26367
rect 34885 26327 34943 26333
rect 36633 26367 36691 26373
rect 36633 26333 36645 26367
rect 36679 26364 36691 26367
rect 36722 26364 36728 26376
rect 36679 26336 36728 26364
rect 36679 26333 36691 26336
rect 36633 26327 36691 26333
rect 32364 26268 32444 26296
rect 32364 26256 32370 26268
rect 34238 26256 34244 26308
rect 34296 26296 34302 26308
rect 34900 26296 34928 26327
rect 36722 26324 36728 26336
rect 36780 26364 36786 26376
rect 37108 26373 37136 26404
rect 36909 26367 36967 26373
rect 36909 26364 36921 26367
rect 36780 26336 36921 26364
rect 36780 26324 36786 26336
rect 36909 26333 36921 26336
rect 36955 26333 36967 26367
rect 36909 26327 36967 26333
rect 37093 26367 37151 26373
rect 37093 26333 37105 26367
rect 37139 26364 37151 26367
rect 37139 26336 37228 26364
rect 37139 26333 37151 26336
rect 37093 26327 37151 26333
rect 34296 26268 34928 26296
rect 34296 26256 34302 26268
rect 37200 26240 37228 26336
rect 29178 26228 29184 26240
rect 28966 26200 29184 26228
rect 29178 26188 29184 26200
rect 29236 26188 29242 26240
rect 31202 26188 31208 26240
rect 31260 26228 31266 26240
rect 34330 26228 34336 26240
rect 31260 26200 34336 26228
rect 31260 26188 31266 26200
rect 34330 26188 34336 26200
rect 34388 26188 34394 26240
rect 37182 26188 37188 26240
rect 37240 26188 37246 26240
rect 1104 26138 38272 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 38272 26138
rect 1104 26064 38272 26086
rect 3418 25984 3424 26036
rect 3476 25984 3482 26036
rect 5629 26027 5687 26033
rect 5629 25993 5641 26027
rect 5675 25993 5687 26027
rect 5629 25987 5687 25993
rect 1762 25916 1768 25968
rect 1820 25916 1826 25968
rect 4522 25956 4528 25968
rect 3344 25928 4528 25956
rect 3344 25900 3372 25928
rect 4522 25916 4528 25928
rect 4580 25916 4586 25968
rect 5644 25956 5672 25987
rect 5718 25984 5724 26036
rect 5776 26024 5782 26036
rect 6641 26027 6699 26033
rect 6641 26024 6653 26027
rect 5776 25996 6653 26024
rect 5776 25984 5782 25996
rect 6641 25993 6653 25996
rect 6687 26024 6699 26027
rect 6914 26024 6920 26036
rect 6687 25996 6920 26024
rect 6687 25993 6699 25996
rect 6641 25987 6699 25993
rect 6914 25984 6920 25996
rect 6972 25984 6978 26036
rect 9674 26024 9680 26036
rect 7024 25996 9680 26024
rect 7024 25956 7052 25996
rect 9674 25984 9680 25996
rect 9732 25984 9738 26036
rect 14093 26027 14151 26033
rect 14093 25993 14105 26027
rect 14139 26024 14151 26027
rect 14642 26024 14648 26036
rect 14139 25996 14648 26024
rect 14139 25993 14151 25996
rect 14093 25987 14151 25993
rect 14642 25984 14648 25996
rect 14700 25984 14706 26036
rect 14752 25996 19932 26024
rect 5644 25928 7052 25956
rect 7101 25959 7159 25965
rect 7101 25925 7113 25959
rect 7147 25956 7159 25959
rect 7282 25956 7288 25968
rect 7147 25928 7288 25956
rect 7147 25925 7159 25928
rect 7101 25919 7159 25925
rect 7282 25916 7288 25928
rect 7340 25916 7346 25968
rect 13354 25916 13360 25968
rect 13412 25916 13418 25968
rect 13464 25928 14688 25956
rect 934 25848 940 25900
rect 992 25888 998 25900
rect 1397 25891 1455 25897
rect 1397 25888 1409 25891
rect 992 25860 1409 25888
rect 992 25848 998 25860
rect 1397 25857 1409 25860
rect 1443 25857 1455 25891
rect 1397 25851 1455 25857
rect 3326 25848 3332 25900
rect 3384 25848 3390 25900
rect 3513 25891 3571 25897
rect 3513 25857 3525 25891
rect 3559 25888 3571 25891
rect 4154 25888 4160 25900
rect 3559 25860 4160 25888
rect 3559 25857 3571 25860
rect 3513 25851 3571 25857
rect 4154 25848 4160 25860
rect 4212 25848 4218 25900
rect 4614 25848 4620 25900
rect 4672 25848 4678 25900
rect 5258 25848 5264 25900
rect 5316 25888 5322 25900
rect 5629 25891 5687 25897
rect 5629 25888 5641 25891
rect 5316 25860 5641 25888
rect 5316 25848 5322 25860
rect 5629 25857 5641 25860
rect 5675 25857 5687 25891
rect 5629 25851 5687 25857
rect 5644 25820 5672 25851
rect 6362 25848 6368 25900
rect 6420 25848 6426 25900
rect 7742 25888 7748 25900
rect 6472 25860 7748 25888
rect 6472 25820 6500 25860
rect 7742 25848 7748 25860
rect 7800 25848 7806 25900
rect 13170 25897 13176 25900
rect 13168 25851 13176 25897
rect 13170 25848 13176 25851
rect 13228 25848 13234 25900
rect 13265 25891 13323 25897
rect 13265 25857 13277 25891
rect 13311 25888 13323 25891
rect 13464 25888 13492 25928
rect 13311 25860 13492 25888
rect 13311 25857 13323 25860
rect 13265 25851 13323 25857
rect 13538 25848 13544 25900
rect 13596 25848 13602 25900
rect 13817 25891 13875 25897
rect 13817 25857 13829 25891
rect 13863 25888 13875 25891
rect 14182 25888 14188 25900
rect 13863 25860 14188 25888
rect 13863 25857 13875 25860
rect 13817 25851 13875 25857
rect 14182 25848 14188 25860
rect 14240 25848 14246 25900
rect 14369 25891 14427 25897
rect 14369 25857 14381 25891
rect 14415 25888 14427 25891
rect 14458 25888 14464 25900
rect 14415 25860 14464 25888
rect 14415 25857 14427 25860
rect 14369 25851 14427 25857
rect 14458 25848 14464 25860
rect 14516 25848 14522 25900
rect 5644 25792 6500 25820
rect 6549 25823 6607 25829
rect 6549 25789 6561 25823
rect 6595 25820 6607 25823
rect 6638 25820 6644 25832
rect 6595 25792 6644 25820
rect 6595 25789 6607 25792
rect 6549 25783 6607 25789
rect 6638 25780 6644 25792
rect 6696 25780 6702 25832
rect 13725 25823 13783 25829
rect 13725 25820 13737 25823
rect 6748 25792 13737 25820
rect 4798 25712 4804 25764
rect 4856 25752 4862 25764
rect 5442 25752 5448 25764
rect 4856 25724 5448 25752
rect 4856 25712 4862 25724
rect 5442 25712 5448 25724
rect 5500 25752 5506 25764
rect 6748 25752 6776 25792
rect 13725 25789 13737 25792
rect 13771 25789 13783 25823
rect 14660 25820 14688 25928
rect 14752 25900 14780 25996
rect 14826 25916 14832 25968
rect 14884 25956 14890 25968
rect 16025 25959 16083 25965
rect 16025 25956 16037 25959
rect 14884 25928 16037 25956
rect 14884 25916 14890 25928
rect 16025 25925 16037 25928
rect 16071 25925 16083 25959
rect 16025 25919 16083 25925
rect 16117 25959 16175 25965
rect 16117 25925 16129 25959
rect 16163 25956 16175 25959
rect 16206 25956 16212 25968
rect 16163 25928 16212 25956
rect 16163 25925 16175 25928
rect 16117 25919 16175 25925
rect 14734 25897 14740 25900
rect 14732 25851 14740 25897
rect 14734 25848 14740 25851
rect 14792 25848 14798 25900
rect 14844 25820 14872 25916
rect 14921 25891 14979 25897
rect 14921 25857 14933 25891
rect 14967 25857 14979 25891
rect 14921 25851 14979 25857
rect 15105 25891 15163 25897
rect 15105 25857 15117 25891
rect 15151 25888 15163 25891
rect 15562 25888 15568 25900
rect 15151 25860 15568 25888
rect 15151 25857 15163 25860
rect 15105 25851 15163 25857
rect 14660 25792 14872 25820
rect 14936 25820 14964 25851
rect 15562 25848 15568 25860
rect 15620 25848 15626 25900
rect 15928 25891 15986 25897
rect 15928 25857 15940 25891
rect 15974 25857 15986 25891
rect 15928 25851 15986 25857
rect 14936 25792 15884 25820
rect 13725 25783 13783 25789
rect 5500 25724 6776 25752
rect 7101 25755 7159 25761
rect 5500 25712 5506 25724
rect 7101 25721 7113 25755
rect 7147 25752 7159 25755
rect 7282 25752 7288 25764
rect 7147 25724 7288 25752
rect 7147 25721 7159 25724
rect 7101 25715 7159 25721
rect 7282 25712 7288 25724
rect 7340 25752 7346 25764
rect 15102 25752 15108 25764
rect 7340 25724 15108 25752
rect 7340 25712 7346 25724
rect 15102 25712 15108 25724
rect 15160 25712 15166 25764
rect 9674 25644 9680 25696
rect 9732 25684 9738 25696
rect 12989 25687 13047 25693
rect 12989 25684 13001 25687
rect 9732 25656 13001 25684
rect 9732 25644 9738 25656
rect 12989 25653 13001 25656
rect 13035 25653 13047 25687
rect 12989 25647 13047 25653
rect 14550 25644 14556 25696
rect 14608 25644 14614 25696
rect 14734 25644 14740 25696
rect 14792 25684 14798 25696
rect 15286 25684 15292 25696
rect 14792 25656 15292 25684
rect 14792 25644 14798 25656
rect 15286 25644 15292 25656
rect 15344 25684 15350 25696
rect 15654 25684 15660 25696
rect 15344 25656 15660 25684
rect 15344 25644 15350 25656
rect 15654 25644 15660 25656
rect 15712 25644 15718 25696
rect 15746 25644 15752 25696
rect 15804 25644 15810 25696
rect 15856 25684 15884 25792
rect 15948 25752 15976 25851
rect 16040 25820 16068 25919
rect 16206 25916 16212 25928
rect 16264 25916 16270 25968
rect 16390 25916 16396 25968
rect 16448 25956 16454 25968
rect 19702 25956 19708 25968
rect 16448 25928 17724 25956
rect 16448 25916 16454 25928
rect 16301 25891 16359 25897
rect 16301 25857 16313 25891
rect 16347 25888 16359 25891
rect 16574 25888 16580 25900
rect 16347 25860 16580 25888
rect 16347 25857 16359 25860
rect 16301 25851 16359 25857
rect 16574 25848 16580 25860
rect 16632 25888 16638 25900
rect 17586 25888 17592 25900
rect 16632 25860 17592 25888
rect 16632 25848 16638 25860
rect 17586 25848 17592 25860
rect 17644 25848 17650 25900
rect 16482 25820 16488 25832
rect 16040 25792 16488 25820
rect 16482 25780 16488 25792
rect 16540 25780 16546 25832
rect 17696 25820 17724 25928
rect 19536 25928 19708 25956
rect 19242 25848 19248 25900
rect 19300 25848 19306 25900
rect 19334 25848 19340 25900
rect 19392 25848 19398 25900
rect 19450 25897 19508 25903
rect 19450 25894 19462 25897
rect 19444 25863 19462 25894
rect 19496 25888 19508 25897
rect 19536 25888 19564 25928
rect 19702 25916 19708 25928
rect 19760 25916 19766 25968
rect 19904 25956 19932 25996
rect 20622 25984 20628 26036
rect 20680 26024 20686 26036
rect 23842 26024 23848 26036
rect 20680 25996 23848 26024
rect 20680 25984 20686 25996
rect 23842 25984 23848 25996
rect 23900 25984 23906 26036
rect 26326 25984 26332 26036
rect 26384 25984 26390 26036
rect 28166 25984 28172 26036
rect 28224 26024 28230 26036
rect 29086 26024 29092 26036
rect 28224 25996 29092 26024
rect 28224 25984 28230 25996
rect 29086 25984 29092 25996
rect 29144 25984 29150 26036
rect 30101 26027 30159 26033
rect 30101 25993 30113 26027
rect 30147 26024 30159 26027
rect 30190 26024 30196 26036
rect 30147 25996 30196 26024
rect 30147 25993 30159 25996
rect 30101 25987 30159 25993
rect 30190 25984 30196 25996
rect 30248 25984 30254 26036
rect 31849 26027 31907 26033
rect 31849 25993 31861 26027
rect 31895 26024 31907 26027
rect 32214 26024 32220 26036
rect 31895 25996 32220 26024
rect 31895 25993 31907 25996
rect 31849 25987 31907 25993
rect 32214 25984 32220 25996
rect 32272 25984 32278 26036
rect 32582 25984 32588 26036
rect 32640 26024 32646 26036
rect 32640 25996 32812 26024
rect 32640 25984 32646 25996
rect 19904 25928 22416 25956
rect 19904 25897 19932 25928
rect 22388 25900 22416 25928
rect 23198 25916 23204 25968
rect 23256 25956 23262 25968
rect 23860 25956 23888 25984
rect 23256 25928 23704 25956
rect 23256 25916 23262 25928
rect 19496 25863 19564 25888
rect 19444 25860 19564 25863
rect 19613 25891 19671 25897
rect 19450 25857 19508 25860
rect 19613 25857 19625 25891
rect 19659 25857 19671 25891
rect 19613 25851 19671 25857
rect 19889 25891 19947 25897
rect 19889 25857 19901 25891
rect 19935 25857 19947 25891
rect 19889 25851 19947 25857
rect 19981 25891 20039 25897
rect 19981 25857 19993 25891
rect 20027 25888 20039 25891
rect 20070 25888 20076 25900
rect 20027 25860 20076 25888
rect 20027 25857 20039 25860
rect 19981 25851 20039 25857
rect 19628 25820 19656 25851
rect 20070 25848 20076 25860
rect 20128 25848 20134 25900
rect 20162 25848 20168 25900
rect 20220 25848 20226 25900
rect 22370 25848 22376 25900
rect 22428 25848 22434 25900
rect 23474 25848 23480 25900
rect 23532 25848 23538 25900
rect 23676 25897 23704 25928
rect 23768 25928 23888 25956
rect 23768 25897 23796 25928
rect 23661 25891 23719 25897
rect 23661 25857 23673 25891
rect 23707 25857 23719 25891
rect 23661 25851 23719 25857
rect 23753 25891 23811 25897
rect 23753 25857 23765 25891
rect 23799 25857 23811 25891
rect 23753 25851 23811 25857
rect 23845 25891 23903 25897
rect 23845 25857 23857 25891
rect 23891 25857 23903 25891
rect 23845 25851 23903 25857
rect 23492 25820 23520 25848
rect 17696 25792 23520 25820
rect 17126 25752 17132 25764
rect 15948 25724 17132 25752
rect 17126 25712 17132 25724
rect 17184 25752 17190 25764
rect 17184 25724 19656 25752
rect 17184 25712 17190 25724
rect 17310 25684 17316 25696
rect 15856 25656 17316 25684
rect 17310 25644 17316 25656
rect 17368 25644 17374 25696
rect 17402 25644 17408 25696
rect 17460 25684 17466 25696
rect 18782 25684 18788 25696
rect 17460 25656 18788 25684
rect 17460 25644 17466 25656
rect 18782 25644 18788 25656
rect 18840 25644 18846 25696
rect 18966 25644 18972 25696
rect 19024 25644 19030 25696
rect 19628 25684 19656 25724
rect 19702 25712 19708 25764
rect 19760 25712 19766 25764
rect 23860 25752 23888 25851
rect 26142 25848 26148 25900
rect 26200 25848 26206 25900
rect 26344 25897 26372 25984
rect 29178 25916 29184 25968
rect 29236 25956 29242 25968
rect 29641 25959 29699 25965
rect 29641 25956 29653 25959
rect 29236 25928 29653 25956
rect 29236 25916 29242 25928
rect 29641 25925 29653 25928
rect 29687 25956 29699 25959
rect 30282 25956 30288 25968
rect 29687 25928 30288 25956
rect 29687 25925 29699 25928
rect 29641 25919 29699 25925
rect 30282 25916 30288 25928
rect 30340 25956 30346 25968
rect 30745 25959 30803 25965
rect 30745 25956 30757 25959
rect 30340 25928 30757 25956
rect 30340 25916 30346 25928
rect 30745 25925 30757 25928
rect 30791 25925 30803 25959
rect 30745 25919 30803 25925
rect 30929 25959 30987 25965
rect 30929 25925 30941 25959
rect 30975 25956 30987 25959
rect 31018 25956 31024 25968
rect 30975 25928 31024 25956
rect 30975 25925 30987 25928
rect 30929 25919 30987 25925
rect 31018 25916 31024 25928
rect 31076 25916 31082 25968
rect 31113 25959 31171 25965
rect 31113 25925 31125 25959
rect 31159 25956 31171 25959
rect 32784 25956 32812 25996
rect 32950 25984 32956 26036
rect 33008 26024 33014 26036
rect 33045 26027 33103 26033
rect 33045 26024 33057 26027
rect 33008 25996 33057 26024
rect 33008 25984 33014 25996
rect 33045 25993 33057 25996
rect 33091 25993 33103 26027
rect 33045 25987 33103 25993
rect 32861 25959 32919 25965
rect 32861 25956 32873 25959
rect 31159 25928 32168 25956
rect 31159 25925 31171 25928
rect 31113 25919 31171 25925
rect 26329 25891 26387 25897
rect 26329 25857 26341 25891
rect 26375 25857 26387 25891
rect 26329 25851 26387 25857
rect 28534 25848 28540 25900
rect 28592 25888 28598 25900
rect 29733 25891 29791 25897
rect 29733 25888 29745 25891
rect 28592 25860 29745 25888
rect 28592 25848 28598 25860
rect 29733 25857 29745 25860
rect 29779 25857 29791 25891
rect 29733 25851 29791 25857
rect 30374 25848 30380 25900
rect 30432 25888 30438 25900
rect 30834 25888 30840 25900
rect 30432 25860 30840 25888
rect 30432 25848 30438 25860
rect 30834 25848 30840 25860
rect 30892 25848 30898 25900
rect 31202 25848 31208 25900
rect 31260 25848 31266 25900
rect 31386 25848 31392 25900
rect 31444 25848 31450 25900
rect 31478 25848 31484 25900
rect 31536 25848 31542 25900
rect 32140 25897 32168 25928
rect 32232 25928 32720 25956
rect 32784 25928 32873 25956
rect 32232 25900 32260 25928
rect 31573 25891 31631 25897
rect 31573 25857 31585 25891
rect 31619 25857 31631 25891
rect 31573 25851 31631 25857
rect 32125 25891 32183 25897
rect 32125 25857 32137 25891
rect 32171 25857 32183 25891
rect 32125 25851 32183 25857
rect 24854 25780 24860 25832
rect 24912 25820 24918 25832
rect 26160 25820 26188 25848
rect 24912 25792 26188 25820
rect 24912 25780 24918 25792
rect 29086 25780 29092 25832
rect 29144 25820 29150 25832
rect 29457 25823 29515 25829
rect 29457 25820 29469 25823
rect 29144 25792 29469 25820
rect 29144 25780 29150 25792
rect 29457 25789 29469 25792
rect 29503 25820 29515 25823
rect 29546 25820 29552 25832
rect 29503 25792 29552 25820
rect 29503 25789 29515 25792
rect 29457 25783 29515 25789
rect 29546 25780 29552 25792
rect 29604 25780 29610 25832
rect 30558 25780 30564 25832
rect 30616 25820 30622 25832
rect 31588 25820 31616 25851
rect 32214 25848 32220 25900
rect 32272 25848 32278 25900
rect 32306 25848 32312 25900
rect 32364 25848 32370 25900
rect 32692 25897 32720 25928
rect 32861 25925 32873 25928
rect 32907 25925 32919 25959
rect 32861 25919 32919 25925
rect 32677 25891 32735 25897
rect 32677 25857 32689 25891
rect 32723 25857 32735 25891
rect 32953 25891 33011 25897
rect 32953 25888 32965 25891
rect 32677 25851 32735 25857
rect 32876 25860 32965 25888
rect 30616 25792 31616 25820
rect 30616 25780 30622 25792
rect 31294 25752 31300 25764
rect 22066 25724 31300 25752
rect 19889 25687 19947 25693
rect 19889 25684 19901 25687
rect 19628 25656 19901 25684
rect 19889 25653 19901 25656
rect 19935 25684 19947 25687
rect 19978 25684 19984 25696
rect 19935 25656 19984 25684
rect 19935 25653 19947 25656
rect 19889 25647 19947 25653
rect 19978 25644 19984 25656
rect 20036 25684 20042 25696
rect 22066 25684 22094 25724
rect 31294 25712 31300 25724
rect 31352 25712 31358 25764
rect 20036 25656 22094 25684
rect 20036 25644 20042 25656
rect 24118 25644 24124 25696
rect 24176 25644 24182 25696
rect 26237 25687 26295 25693
rect 26237 25653 26249 25687
rect 26283 25684 26295 25687
rect 27062 25684 27068 25696
rect 26283 25656 27068 25684
rect 26283 25653 26295 25656
rect 26237 25647 26295 25653
rect 27062 25644 27068 25656
rect 27120 25644 27126 25696
rect 31588 25684 31616 25792
rect 31938 25712 31944 25764
rect 31996 25752 32002 25764
rect 32324 25752 32352 25848
rect 32876 25832 32904 25860
rect 32953 25857 32965 25860
rect 32999 25857 33011 25891
rect 32953 25851 33011 25857
rect 33137 25891 33195 25897
rect 33137 25857 33149 25891
rect 33183 25888 33195 25891
rect 33183 25860 33272 25888
rect 33183 25857 33195 25860
rect 33137 25851 33195 25857
rect 33244 25832 33272 25860
rect 32401 25823 32459 25829
rect 32401 25789 32413 25823
rect 32447 25789 32459 25823
rect 32401 25783 32459 25789
rect 31996 25724 32352 25752
rect 31996 25712 32002 25724
rect 32416 25684 32444 25783
rect 32490 25780 32496 25832
rect 32548 25780 32554 25832
rect 32858 25780 32864 25832
rect 32916 25780 32922 25832
rect 33226 25780 33232 25832
rect 33284 25780 33290 25832
rect 31588 25656 32444 25684
rect 1104 25594 38272 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38272 25594
rect 1104 25520 38272 25542
rect 7282 25440 7288 25492
rect 7340 25440 7346 25492
rect 14734 25480 14740 25492
rect 7392 25452 8708 25480
rect 1394 25304 1400 25356
rect 1452 25304 1458 25356
rect 3145 25347 3203 25353
rect 3145 25313 3157 25347
rect 3191 25344 3203 25347
rect 4341 25347 4399 25353
rect 4341 25344 4353 25347
rect 3191 25316 4353 25344
rect 3191 25313 3203 25316
rect 3145 25307 3203 25313
rect 4341 25313 4353 25316
rect 4387 25344 4399 25347
rect 4522 25344 4528 25356
rect 4387 25316 4528 25344
rect 4387 25313 4399 25316
rect 4341 25307 4399 25313
rect 4522 25304 4528 25316
rect 4580 25304 4586 25356
rect 7300 25353 7328 25440
rect 7285 25347 7343 25353
rect 6656 25316 6960 25344
rect 2774 25236 2780 25288
rect 2832 25236 2838 25288
rect 4617 25279 4675 25285
rect 4617 25245 4629 25279
rect 4663 25276 4675 25279
rect 4706 25276 4712 25288
rect 4663 25248 4712 25276
rect 4663 25245 4675 25248
rect 4617 25239 4675 25245
rect 4706 25236 4712 25248
rect 4764 25236 4770 25288
rect 6656 25285 6684 25316
rect 6932 25288 6960 25316
rect 7285 25313 7297 25347
rect 7331 25313 7343 25347
rect 7285 25307 7343 25313
rect 6641 25279 6699 25285
rect 6641 25245 6653 25279
rect 6687 25245 6699 25279
rect 6641 25239 6699 25245
rect 6822 25236 6828 25288
rect 6880 25236 6886 25288
rect 6914 25236 6920 25288
rect 6972 25276 6978 25288
rect 7101 25279 7159 25285
rect 7101 25276 7113 25279
rect 6972 25248 7113 25276
rect 6972 25236 6978 25248
rect 7101 25245 7113 25248
rect 7147 25245 7159 25279
rect 7101 25239 7159 25245
rect 1670 25168 1676 25220
rect 1728 25168 1734 25220
rect 4985 25211 5043 25217
rect 4985 25177 4997 25211
rect 5031 25208 5043 25211
rect 5442 25208 5448 25220
rect 5031 25180 5448 25208
rect 5031 25177 5043 25180
rect 4985 25171 5043 25177
rect 5442 25168 5448 25180
rect 5500 25208 5506 25220
rect 7392 25208 7420 25452
rect 7929 25415 7987 25421
rect 7929 25381 7941 25415
rect 7975 25412 7987 25415
rect 8294 25412 8300 25424
rect 7975 25384 8300 25412
rect 7975 25381 7987 25384
rect 7929 25375 7987 25381
rect 8294 25372 8300 25384
rect 8352 25372 8358 25424
rect 8680 25353 8708 25452
rect 13464 25452 14740 25480
rect 9677 25415 9735 25421
rect 9677 25381 9689 25415
rect 9723 25412 9735 25415
rect 9766 25412 9772 25424
rect 9723 25384 9772 25412
rect 9723 25381 9735 25384
rect 9677 25375 9735 25381
rect 9766 25372 9772 25384
rect 9824 25372 9830 25424
rect 8665 25347 8723 25353
rect 5500 25180 7420 25208
rect 7668 25316 8248 25344
rect 5500 25168 5506 25180
rect 3786 25100 3792 25152
rect 3844 25100 3850 25152
rect 5810 25100 5816 25152
rect 5868 25140 5874 25152
rect 6454 25140 6460 25152
rect 5868 25112 6460 25140
rect 5868 25100 5874 25112
rect 6454 25100 6460 25112
rect 6512 25100 6518 25152
rect 6917 25143 6975 25149
rect 6917 25109 6929 25143
rect 6963 25140 6975 25143
rect 7668 25140 7696 25316
rect 8220 25288 8248 25316
rect 8665 25313 8677 25347
rect 8711 25344 8723 25347
rect 9033 25347 9091 25353
rect 9033 25344 9045 25347
rect 8711 25316 9045 25344
rect 8711 25313 8723 25316
rect 8665 25307 8723 25313
rect 9033 25313 9045 25316
rect 9079 25313 9091 25347
rect 9033 25307 9091 25313
rect 10410 25304 10416 25356
rect 10468 25304 10474 25356
rect 10597 25347 10655 25353
rect 10597 25313 10609 25347
rect 10643 25344 10655 25347
rect 12894 25344 12900 25356
rect 10643 25316 12900 25344
rect 10643 25313 10655 25316
rect 10597 25307 10655 25313
rect 12894 25304 12900 25316
rect 12952 25304 12958 25356
rect 7745 25279 7803 25285
rect 7745 25245 7757 25279
rect 7791 25276 7803 25279
rect 7791 25248 8064 25276
rect 7791 25245 7803 25248
rect 7745 25239 7803 25245
rect 8036 25149 8064 25248
rect 8202 25236 8208 25288
rect 8260 25276 8266 25288
rect 8389 25279 8447 25285
rect 8389 25276 8401 25279
rect 8260 25248 8401 25276
rect 8260 25236 8266 25248
rect 8389 25245 8401 25248
rect 8435 25245 8447 25279
rect 8389 25239 8447 25245
rect 9490 25236 9496 25288
rect 9548 25276 9554 25288
rect 11149 25279 11207 25285
rect 11149 25276 11161 25279
rect 9548 25248 11161 25276
rect 9548 25236 9554 25248
rect 11149 25245 11161 25248
rect 11195 25245 11207 25279
rect 11149 25239 11207 25245
rect 12434 25236 12440 25288
rect 12492 25276 12498 25288
rect 13081 25279 13139 25285
rect 13081 25276 13093 25279
rect 12492 25248 13093 25276
rect 12492 25236 12498 25248
rect 13081 25245 13093 25248
rect 13127 25245 13139 25279
rect 13464 25276 13492 25452
rect 14734 25440 14740 25452
rect 14792 25440 14798 25492
rect 14826 25440 14832 25492
rect 14884 25440 14890 25492
rect 14918 25440 14924 25492
rect 14976 25480 14982 25492
rect 17402 25480 17408 25492
rect 14976 25452 17408 25480
rect 14976 25440 14982 25452
rect 17402 25440 17408 25452
rect 17460 25440 17466 25492
rect 17681 25483 17739 25489
rect 17681 25449 17693 25483
rect 17727 25449 17739 25483
rect 17681 25443 17739 25449
rect 14844 25412 14872 25440
rect 14384 25384 14872 25412
rect 15657 25415 15715 25421
rect 13633 25279 13691 25285
rect 13633 25276 13645 25279
rect 13464 25248 13645 25276
rect 13081 25239 13139 25245
rect 13633 25245 13645 25248
rect 13679 25245 13691 25279
rect 13633 25239 13691 25245
rect 14274 25236 14280 25288
rect 14332 25236 14338 25288
rect 14384 25285 14412 25384
rect 15657 25381 15669 25415
rect 15703 25412 15715 25415
rect 16206 25412 16212 25424
rect 15703 25384 16212 25412
rect 15703 25381 15715 25384
rect 15657 25375 15715 25381
rect 16206 25372 16212 25384
rect 16264 25372 16270 25424
rect 17221 25415 17279 25421
rect 17221 25381 17233 25415
rect 17267 25412 17279 25415
rect 17310 25412 17316 25424
rect 17267 25384 17316 25412
rect 17267 25381 17279 25384
rect 17221 25375 17279 25381
rect 17310 25372 17316 25384
rect 17368 25372 17374 25424
rect 17696 25412 17724 25443
rect 17954 25440 17960 25492
rect 18012 25440 18018 25492
rect 18046 25440 18052 25492
rect 18104 25440 18110 25492
rect 18690 25440 18696 25492
rect 18748 25440 18754 25492
rect 19702 25480 19708 25492
rect 18800 25452 19708 25480
rect 18064 25412 18092 25440
rect 18325 25415 18383 25421
rect 18325 25412 18337 25415
rect 17696 25384 18092 25412
rect 18156 25384 18337 25412
rect 14734 25344 14740 25356
rect 14660 25316 14740 25344
rect 14660 25285 14688 25316
rect 14734 25304 14740 25316
rect 14792 25344 14798 25356
rect 15562 25344 15568 25356
rect 14792 25316 15568 25344
rect 14792 25304 14798 25316
rect 15562 25304 15568 25316
rect 15620 25344 15626 25356
rect 17589 25347 17647 25353
rect 15620 25316 16252 25344
rect 15620 25304 15626 25316
rect 14369 25279 14427 25285
rect 14369 25245 14381 25279
rect 14415 25245 14427 25279
rect 14369 25239 14427 25245
rect 14645 25279 14703 25285
rect 14645 25245 14657 25279
rect 14691 25245 14703 25279
rect 14645 25239 14703 25245
rect 15010 25236 15016 25288
rect 15068 25236 15074 25288
rect 15838 25285 15844 25288
rect 15836 25276 15844 25285
rect 15799 25248 15844 25276
rect 15836 25239 15844 25248
rect 15838 25236 15844 25239
rect 15896 25236 15902 25288
rect 16022 25236 16028 25288
rect 16080 25236 16086 25288
rect 16224 25285 16252 25316
rect 17589 25313 17601 25347
rect 17635 25344 17647 25347
rect 18156 25344 18184 25384
rect 18325 25381 18337 25384
rect 18371 25381 18383 25415
rect 18325 25375 18383 25381
rect 18800 25344 18828 25452
rect 19702 25440 19708 25452
rect 19760 25440 19766 25492
rect 20809 25483 20867 25489
rect 20809 25449 20821 25483
rect 20855 25480 20867 25483
rect 21358 25480 21364 25492
rect 20855 25452 21364 25480
rect 20855 25449 20867 25452
rect 20809 25443 20867 25449
rect 21358 25440 21364 25452
rect 21416 25440 21422 25492
rect 25409 25483 25467 25489
rect 25409 25449 25421 25483
rect 25455 25480 25467 25483
rect 26326 25480 26332 25492
rect 25455 25452 26332 25480
rect 25455 25449 25467 25452
rect 25409 25443 25467 25449
rect 26326 25440 26332 25452
rect 26384 25440 26390 25492
rect 30282 25440 30288 25492
rect 30340 25480 30346 25492
rect 30561 25483 30619 25489
rect 30561 25480 30573 25483
rect 30340 25452 30573 25480
rect 30340 25440 30346 25452
rect 30561 25449 30573 25452
rect 30607 25449 30619 25483
rect 30561 25443 30619 25449
rect 31021 25483 31079 25489
rect 31021 25449 31033 25483
rect 31067 25480 31079 25483
rect 31386 25480 31392 25492
rect 31067 25452 31392 25480
rect 31067 25449 31079 25452
rect 31021 25443 31079 25449
rect 31386 25440 31392 25452
rect 31444 25440 31450 25492
rect 33042 25440 33048 25492
rect 33100 25440 33106 25492
rect 36722 25440 36728 25492
rect 36780 25440 36786 25492
rect 37182 25440 37188 25492
rect 37240 25440 37246 25492
rect 19058 25372 19064 25424
rect 19116 25412 19122 25424
rect 22186 25412 22192 25424
rect 19116 25384 22192 25412
rect 19116 25372 19122 25384
rect 22186 25372 22192 25384
rect 22244 25372 22250 25424
rect 32858 25412 32864 25424
rect 26896 25384 32864 25412
rect 17635 25316 18184 25344
rect 18248 25316 18828 25344
rect 17635 25313 17647 25316
rect 17589 25307 17647 25313
rect 16209 25279 16267 25285
rect 16209 25245 16221 25279
rect 16255 25276 16267 25279
rect 16574 25276 16580 25288
rect 16255 25248 16580 25276
rect 16255 25245 16267 25248
rect 16209 25239 16267 25245
rect 16574 25236 16580 25248
rect 16632 25236 16638 25288
rect 17034 25236 17040 25288
rect 17092 25276 17098 25288
rect 17405 25279 17463 25285
rect 17405 25276 17417 25279
rect 17092 25248 17417 25276
rect 17092 25236 17098 25248
rect 17405 25245 17417 25248
rect 17451 25276 17463 25279
rect 17494 25276 17500 25288
rect 17451 25248 17500 25276
rect 17451 25245 17463 25248
rect 17405 25239 17463 25245
rect 17494 25236 17500 25248
rect 17552 25236 17558 25288
rect 17957 25279 18015 25285
rect 17604 25248 17908 25276
rect 9217 25211 9275 25217
rect 9217 25177 9229 25211
rect 9263 25208 9275 25211
rect 9858 25208 9864 25220
rect 9263 25180 9864 25208
rect 9263 25177 9275 25180
rect 9217 25171 9275 25177
rect 9858 25168 9864 25180
rect 9916 25168 9922 25220
rect 10689 25211 10747 25217
rect 10689 25177 10701 25211
rect 10735 25208 10747 25211
rect 10735 25180 11192 25208
rect 10735 25177 10747 25180
rect 10689 25171 10747 25177
rect 6963 25112 7696 25140
rect 8021 25143 8079 25149
rect 6963 25109 6975 25112
rect 6917 25103 6975 25109
rect 8021 25109 8033 25143
rect 8067 25109 8079 25143
rect 8021 25103 8079 25109
rect 8481 25143 8539 25149
rect 8481 25109 8493 25143
rect 8527 25140 8539 25143
rect 9030 25140 9036 25152
rect 8527 25112 9036 25140
rect 8527 25109 8539 25112
rect 8481 25103 8539 25109
rect 9030 25100 9036 25112
rect 9088 25100 9094 25152
rect 9309 25143 9367 25149
rect 9309 25109 9321 25143
rect 9355 25140 9367 25143
rect 9582 25140 9588 25152
rect 9355 25112 9588 25140
rect 9355 25109 9367 25112
rect 9309 25103 9367 25109
rect 9582 25100 9588 25112
rect 9640 25140 9646 25152
rect 10704 25140 10732 25171
rect 9640 25112 10732 25140
rect 9640 25100 9646 25112
rect 11054 25100 11060 25152
rect 11112 25100 11118 25152
rect 11164 25140 11192 25180
rect 11422 25168 11428 25220
rect 11480 25168 11486 25220
rect 13446 25168 13452 25220
rect 13504 25208 13510 25220
rect 14461 25211 14519 25217
rect 13504 25180 14412 25208
rect 13504 25168 13510 25180
rect 11606 25140 11612 25152
rect 11164 25112 11612 25140
rect 11606 25100 11612 25112
rect 11664 25100 11670 25152
rect 14090 25100 14096 25152
rect 14148 25100 14154 25152
rect 14384 25140 14412 25180
rect 14461 25177 14473 25211
rect 14507 25208 14519 25211
rect 15028 25208 15056 25236
rect 14507 25180 15056 25208
rect 15933 25211 15991 25217
rect 14507 25177 14519 25180
rect 14461 25171 14519 25177
rect 15933 25177 15945 25211
rect 15979 25208 15991 25211
rect 16482 25208 16488 25220
rect 15979 25180 16488 25208
rect 15979 25177 15991 25180
rect 15933 25171 15991 25177
rect 16482 25168 16488 25180
rect 16540 25168 16546 25220
rect 17604 25140 17632 25248
rect 17681 25211 17739 25217
rect 17681 25177 17693 25211
rect 17727 25208 17739 25211
rect 17727 25180 17816 25208
rect 17727 25177 17739 25180
rect 17681 25171 17739 25177
rect 17788 25149 17816 25180
rect 14384 25112 17632 25140
rect 17773 25143 17831 25149
rect 17773 25109 17785 25143
rect 17819 25109 17831 25143
rect 17880 25140 17908 25248
rect 17957 25245 17969 25279
rect 18003 25245 18015 25279
rect 17957 25239 18015 25245
rect 17972 25208 18000 25239
rect 18046 25236 18052 25288
rect 18104 25236 18110 25288
rect 18138 25236 18144 25288
rect 18196 25236 18202 25288
rect 18248 25285 18276 25316
rect 19978 25304 19984 25356
rect 20036 25304 20042 25356
rect 20257 25347 20315 25353
rect 20257 25313 20269 25347
rect 20303 25344 20315 25347
rect 20441 25347 20499 25353
rect 20441 25344 20453 25347
rect 20303 25316 20453 25344
rect 20303 25313 20315 25316
rect 20257 25307 20315 25313
rect 20441 25313 20453 25316
rect 20487 25313 20499 25347
rect 20441 25307 20499 25313
rect 21910 25304 21916 25356
rect 21968 25344 21974 25356
rect 26896 25344 26924 25384
rect 32858 25372 32864 25384
rect 32916 25372 32922 25424
rect 21968 25316 26924 25344
rect 30484 25316 32904 25344
rect 21968 25304 21974 25316
rect 30484 25288 30512 25316
rect 18233 25279 18291 25285
rect 18233 25245 18245 25279
rect 18279 25245 18291 25279
rect 18233 25239 18291 25245
rect 18509 25279 18567 25285
rect 18509 25245 18521 25279
rect 18555 25245 18567 25279
rect 18509 25239 18567 25245
rect 18785 25279 18843 25285
rect 18785 25245 18797 25279
rect 18831 25276 18843 25279
rect 18831 25248 19334 25276
rect 18831 25245 18843 25248
rect 18785 25239 18843 25245
rect 18156 25208 18184 25236
rect 17972 25180 18184 25208
rect 18524 25152 18552 25239
rect 18506 25140 18512 25152
rect 17880 25112 18512 25140
rect 17773 25103 17831 25109
rect 18506 25100 18512 25112
rect 18564 25100 18570 25152
rect 19306 25140 19334 25248
rect 19886 25236 19892 25288
rect 19944 25236 19950 25288
rect 20530 25236 20536 25288
rect 20588 25236 20594 25288
rect 23750 25276 23756 25288
rect 20640 25248 23756 25276
rect 19904 25208 19932 25236
rect 20640 25208 20668 25248
rect 23750 25236 23756 25248
rect 23808 25276 23814 25288
rect 24670 25276 24676 25288
rect 23808 25248 24676 25276
rect 23808 25236 23814 25248
rect 24670 25236 24676 25248
rect 24728 25236 24734 25288
rect 25038 25236 25044 25288
rect 25096 25236 25102 25288
rect 25225 25279 25283 25285
rect 25225 25245 25237 25279
rect 25271 25276 25283 25279
rect 25271 25248 25360 25276
rect 25271 25245 25283 25248
rect 25225 25239 25283 25245
rect 19904 25180 20668 25208
rect 20806 25168 20812 25220
rect 20864 25208 20870 25220
rect 23198 25208 23204 25220
rect 20864 25180 23204 25208
rect 20864 25168 20870 25180
rect 23198 25168 23204 25180
rect 23256 25168 23262 25220
rect 20824 25140 20852 25168
rect 25332 25152 25360 25248
rect 26694 25236 26700 25288
rect 26752 25236 26758 25288
rect 27246 25236 27252 25288
rect 27304 25236 27310 25288
rect 27338 25236 27344 25288
rect 27396 25276 27402 25288
rect 27433 25279 27491 25285
rect 27433 25276 27445 25279
rect 27396 25248 27445 25276
rect 27396 25236 27402 25248
rect 27433 25245 27445 25248
rect 27479 25245 27491 25279
rect 27433 25239 27491 25245
rect 26712 25208 26740 25236
rect 27448 25208 27476 25239
rect 30466 25236 30472 25288
rect 30524 25236 30530 25288
rect 30742 25236 30748 25288
rect 30800 25236 30806 25288
rect 30834 25236 30840 25288
rect 30892 25236 30898 25288
rect 31110 25236 31116 25288
rect 31168 25276 31174 25288
rect 31757 25279 31815 25285
rect 31757 25276 31769 25279
rect 31168 25248 31769 25276
rect 31168 25236 31174 25248
rect 31757 25245 31769 25248
rect 31803 25276 31815 25279
rect 32582 25276 32588 25288
rect 31803 25248 32588 25276
rect 31803 25245 31815 25248
rect 31757 25239 31815 25245
rect 32582 25236 32588 25248
rect 32640 25236 32646 25288
rect 30374 25208 30380 25220
rect 26712 25180 30380 25208
rect 30374 25168 30380 25180
rect 30432 25208 30438 25220
rect 32122 25208 32128 25220
rect 30432 25180 32128 25208
rect 30432 25168 30438 25180
rect 32122 25168 32128 25180
rect 32180 25168 32186 25220
rect 32876 25208 32904 25316
rect 32968 25316 33548 25344
rect 32968 25288 32996 25316
rect 32950 25236 32956 25288
rect 33008 25236 33014 25288
rect 33318 25236 33324 25288
rect 33376 25236 33382 25288
rect 33520 25285 33548 25316
rect 36446 25304 36452 25356
rect 36504 25344 36510 25356
rect 36909 25347 36967 25353
rect 36909 25344 36921 25347
rect 36504 25316 36921 25344
rect 36504 25304 36510 25316
rect 33413 25279 33471 25285
rect 33413 25245 33425 25279
rect 33459 25245 33471 25279
rect 33413 25239 33471 25245
rect 33505 25279 33563 25285
rect 33505 25245 33517 25279
rect 33551 25245 33563 25279
rect 33505 25239 33563 25245
rect 33226 25208 33232 25220
rect 32876 25180 33232 25208
rect 33226 25168 33232 25180
rect 33284 25168 33290 25220
rect 33428 25208 33456 25239
rect 33686 25236 33692 25288
rect 33744 25236 33750 25288
rect 36556 25285 36584 25316
rect 36909 25313 36921 25316
rect 36955 25313 36967 25347
rect 36909 25307 36967 25313
rect 36265 25279 36323 25285
rect 36265 25245 36277 25279
rect 36311 25245 36323 25279
rect 36265 25239 36323 25245
rect 36541 25279 36599 25285
rect 36541 25245 36553 25279
rect 36587 25245 36599 25279
rect 36541 25239 36599 25245
rect 36817 25279 36875 25285
rect 36817 25245 36829 25279
rect 36863 25245 36875 25279
rect 36817 25239 36875 25245
rect 36280 25208 36308 25239
rect 36832 25208 36860 25239
rect 36998 25236 37004 25288
rect 37056 25276 37062 25288
rect 37093 25279 37151 25285
rect 37093 25276 37105 25279
rect 37056 25248 37105 25276
rect 37056 25236 37062 25248
rect 37093 25245 37105 25248
rect 37139 25245 37151 25279
rect 37277 25279 37335 25285
rect 37277 25276 37289 25279
rect 37093 25239 37151 25245
rect 37200 25248 37289 25276
rect 37200 25208 37228 25248
rect 37277 25245 37289 25248
rect 37323 25245 37335 25279
rect 37277 25239 37335 25245
rect 33428 25180 33824 25208
rect 36280 25180 36768 25208
rect 36832 25180 37228 25208
rect 33796 25152 33824 25180
rect 36740 25152 36768 25180
rect 37200 25152 37228 25180
rect 19306 25112 20852 25140
rect 22002 25100 22008 25152
rect 22060 25140 22066 25152
rect 22094 25140 22100 25152
rect 22060 25112 22100 25140
rect 22060 25100 22066 25112
rect 22094 25100 22100 25112
rect 22152 25100 22158 25152
rect 25314 25100 25320 25152
rect 25372 25100 25378 25152
rect 27341 25143 27399 25149
rect 27341 25109 27353 25143
rect 27387 25140 27399 25143
rect 27614 25140 27620 25152
rect 27387 25112 27620 25140
rect 27387 25109 27399 25112
rect 27341 25103 27399 25109
rect 27614 25100 27620 25112
rect 27672 25100 27678 25152
rect 31478 25100 31484 25152
rect 31536 25140 31542 25152
rect 31849 25143 31907 25149
rect 31849 25140 31861 25143
rect 31536 25112 31861 25140
rect 31536 25100 31542 25112
rect 31849 25109 31861 25112
rect 31895 25140 31907 25143
rect 32490 25140 32496 25152
rect 31895 25112 32496 25140
rect 31895 25109 31907 25112
rect 31849 25103 31907 25109
rect 32490 25100 32496 25112
rect 32548 25140 32554 25152
rect 33502 25140 33508 25152
rect 32548 25112 33508 25140
rect 32548 25100 32554 25112
rect 33502 25100 33508 25112
rect 33560 25100 33566 25152
rect 33778 25100 33784 25152
rect 33836 25100 33842 25152
rect 36357 25143 36415 25149
rect 36357 25109 36369 25143
rect 36403 25140 36415 25143
rect 36630 25140 36636 25152
rect 36403 25112 36636 25140
rect 36403 25109 36415 25112
rect 36357 25103 36415 25109
rect 36630 25100 36636 25112
rect 36688 25100 36694 25152
rect 36722 25100 36728 25152
rect 36780 25100 36786 25152
rect 37182 25100 37188 25152
rect 37240 25100 37246 25152
rect 1104 25050 38272 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 38272 25050
rect 1104 24976 38272 24998
rect 1670 24896 1676 24948
rect 1728 24936 1734 24948
rect 2501 24939 2559 24945
rect 2501 24936 2513 24939
rect 1728 24908 2513 24936
rect 1728 24896 1734 24908
rect 2501 24905 2513 24908
rect 2547 24905 2559 24939
rect 2501 24899 2559 24905
rect 2774 24896 2780 24948
rect 2832 24936 2838 24948
rect 2869 24939 2927 24945
rect 2869 24936 2881 24939
rect 2832 24908 2881 24936
rect 2832 24896 2838 24908
rect 2869 24905 2881 24908
rect 2915 24936 2927 24939
rect 3786 24936 3792 24948
rect 2915 24908 3792 24936
rect 2915 24905 2927 24908
rect 2869 24899 2927 24905
rect 3786 24896 3792 24908
rect 3844 24896 3850 24948
rect 4065 24939 4123 24945
rect 4065 24905 4077 24939
rect 4111 24936 4123 24939
rect 4798 24936 4804 24948
rect 4111 24908 4804 24936
rect 4111 24905 4123 24908
rect 4065 24899 4123 24905
rect 4798 24896 4804 24908
rect 4856 24896 4862 24948
rect 8110 24896 8116 24948
rect 8168 24936 8174 24948
rect 8168 24908 10456 24936
rect 8168 24896 8174 24908
rect 10428 24880 10456 24908
rect 11054 24896 11060 24948
rect 11112 24896 11118 24948
rect 11422 24896 11428 24948
rect 11480 24936 11486 24948
rect 11517 24939 11575 24945
rect 11517 24936 11529 24939
rect 11480 24908 11529 24936
rect 11480 24896 11486 24908
rect 11517 24905 11529 24908
rect 11563 24905 11575 24939
rect 11517 24899 11575 24905
rect 11606 24896 11612 24948
rect 11664 24936 11670 24948
rect 11885 24939 11943 24945
rect 11885 24936 11897 24939
rect 11664 24908 11897 24936
rect 11664 24896 11670 24908
rect 11885 24905 11897 24908
rect 11931 24905 11943 24939
rect 11885 24899 11943 24905
rect 14274 24896 14280 24948
rect 14332 24936 14338 24948
rect 14918 24936 14924 24948
rect 14332 24908 14924 24936
rect 14332 24896 14338 24908
rect 14918 24896 14924 24908
rect 14976 24896 14982 24948
rect 15838 24896 15844 24948
rect 15896 24936 15902 24948
rect 19889 24939 19947 24945
rect 15896 24908 18092 24936
rect 15896 24896 15902 24908
rect 7944 24840 8786 24868
rect 2685 24803 2743 24809
rect 2685 24769 2697 24803
rect 2731 24769 2743 24803
rect 2685 24763 2743 24769
rect 2700 24732 2728 24763
rect 2958 24760 2964 24812
rect 3016 24760 3022 24812
rect 4433 24803 4491 24809
rect 4433 24769 4445 24803
rect 4479 24800 4491 24803
rect 4614 24800 4620 24812
rect 4479 24772 4620 24800
rect 4479 24769 4491 24772
rect 4433 24763 4491 24769
rect 4614 24760 4620 24772
rect 4672 24760 4678 24812
rect 4709 24803 4767 24809
rect 4709 24769 4721 24803
rect 4755 24800 4767 24803
rect 4798 24800 4804 24812
rect 4755 24772 4804 24800
rect 4755 24769 4767 24772
rect 4709 24763 4767 24769
rect 4798 24760 4804 24772
rect 4856 24760 4862 24812
rect 5353 24803 5411 24809
rect 5353 24769 5365 24803
rect 5399 24800 5411 24803
rect 6825 24803 6883 24809
rect 6825 24800 6837 24803
rect 5399 24772 6837 24800
rect 5399 24769 5411 24772
rect 5353 24763 5411 24769
rect 6825 24769 6837 24772
rect 6871 24800 6883 24803
rect 6914 24800 6920 24812
rect 6871 24772 6920 24800
rect 6871 24769 6883 24772
rect 6825 24763 6883 24769
rect 6914 24760 6920 24772
rect 6972 24800 6978 24812
rect 7285 24803 7343 24809
rect 7285 24800 7297 24803
rect 6972 24772 7297 24800
rect 6972 24760 6978 24772
rect 7285 24769 7297 24772
rect 7331 24800 7343 24803
rect 7331 24772 7604 24800
rect 7331 24769 7343 24772
rect 7285 24763 7343 24769
rect 7576 24744 7604 24772
rect 7650 24760 7656 24812
rect 7708 24800 7714 24812
rect 7944 24800 7972 24840
rect 10410 24828 10416 24880
rect 10468 24828 10474 24880
rect 7708 24772 7972 24800
rect 7708 24760 7714 24772
rect 8018 24760 8024 24812
rect 8076 24760 8082 24812
rect 11072 24800 11100 24896
rect 14093 24871 14151 24877
rect 14093 24837 14105 24871
rect 14139 24868 14151 24871
rect 14642 24868 14648 24880
rect 14139 24840 14648 24868
rect 14139 24837 14151 24840
rect 14093 24831 14151 24837
rect 14642 24828 14648 24840
rect 14700 24828 14706 24880
rect 14752 24840 15332 24868
rect 11701 24803 11759 24809
rect 11701 24800 11713 24803
rect 11072 24772 11713 24800
rect 11701 24769 11713 24772
rect 11747 24769 11759 24803
rect 11701 24763 11759 24769
rect 12069 24803 12127 24809
rect 12069 24769 12081 24803
rect 12115 24769 12127 24803
rect 12069 24763 12127 24769
rect 13817 24803 13875 24809
rect 13817 24769 13829 24803
rect 13863 24769 13875 24803
rect 13817 24763 13875 24769
rect 4341 24735 4399 24741
rect 4341 24732 4353 24735
rect 2700 24704 4353 24732
rect 4341 24701 4353 24704
rect 4387 24732 4399 24735
rect 4525 24735 4583 24741
rect 4525 24732 4537 24735
rect 4387 24704 4537 24732
rect 4387 24701 4399 24704
rect 4341 24695 4399 24701
rect 4525 24701 4537 24704
rect 4571 24701 4583 24735
rect 4525 24695 4583 24701
rect 4893 24735 4951 24741
rect 4893 24701 4905 24735
rect 4939 24732 4951 24735
rect 4939 24704 5028 24732
rect 4939 24701 4951 24704
rect 4893 24695 4951 24701
rect 3694 24556 3700 24608
rect 3752 24596 3758 24608
rect 4249 24599 4307 24605
rect 4249 24596 4261 24599
rect 3752 24568 4261 24596
rect 3752 24556 3758 24568
rect 4249 24565 4261 24568
rect 4295 24565 4307 24599
rect 5000 24596 5028 24704
rect 5534 24692 5540 24744
rect 5592 24732 5598 24744
rect 6546 24732 6552 24744
rect 5592 24704 6552 24732
rect 5592 24692 5598 24704
rect 6546 24692 6552 24704
rect 6604 24692 6610 24744
rect 6638 24692 6644 24744
rect 6696 24692 6702 24744
rect 7009 24735 7067 24741
rect 7009 24701 7021 24735
rect 7055 24732 7067 24735
rect 7098 24732 7104 24744
rect 7055 24704 7104 24732
rect 7055 24701 7067 24704
rect 7009 24695 7067 24701
rect 7098 24692 7104 24704
rect 7156 24692 7162 24744
rect 7466 24692 7472 24744
rect 7524 24692 7530 24744
rect 7558 24692 7564 24744
rect 7616 24692 7622 24744
rect 5169 24667 5227 24673
rect 5169 24633 5181 24667
rect 5215 24664 5227 24667
rect 5350 24664 5356 24676
rect 5215 24636 5356 24664
rect 5215 24633 5227 24636
rect 5169 24627 5227 24633
rect 5350 24624 5356 24636
rect 5408 24624 5414 24676
rect 6822 24624 6828 24676
rect 6880 24664 6886 24676
rect 8036 24664 8064 24760
rect 8294 24692 8300 24744
rect 8352 24692 8358 24744
rect 9030 24692 9036 24744
rect 9088 24732 9094 24744
rect 10045 24735 10103 24741
rect 10045 24732 10057 24735
rect 9088 24704 10057 24732
rect 9088 24692 9094 24704
rect 10045 24701 10057 24704
rect 10091 24732 10103 24735
rect 10410 24732 10416 24744
rect 10091 24704 10416 24732
rect 10091 24701 10103 24704
rect 10045 24695 10103 24701
rect 10410 24692 10416 24704
rect 10468 24692 10474 24744
rect 11882 24692 11888 24744
rect 11940 24732 11946 24744
rect 12084 24732 12112 24763
rect 11940 24704 12112 24732
rect 12253 24735 12311 24741
rect 11940 24692 11946 24704
rect 12253 24701 12265 24735
rect 12299 24732 12311 24735
rect 13630 24732 13636 24744
rect 12299 24704 13636 24732
rect 12299 24701 12311 24704
rect 12253 24695 12311 24701
rect 13630 24692 13636 24704
rect 13688 24692 13694 24744
rect 11900 24664 11928 24692
rect 6880 24636 8064 24664
rect 9324 24636 11928 24664
rect 6880 24624 6886 24636
rect 5258 24596 5264 24608
rect 5000 24568 5264 24596
rect 4249 24559 4307 24565
rect 5258 24556 5264 24568
rect 5316 24556 5322 24608
rect 5902 24556 5908 24608
rect 5960 24596 5966 24608
rect 6178 24596 6184 24608
rect 5960 24568 6184 24596
rect 5960 24556 5966 24568
rect 6178 24556 6184 24568
rect 6236 24596 6242 24608
rect 7101 24599 7159 24605
rect 7101 24596 7113 24599
rect 6236 24568 7113 24596
rect 6236 24556 6242 24568
rect 7101 24565 7113 24568
rect 7147 24565 7159 24599
rect 7101 24559 7159 24565
rect 7558 24556 7564 24608
rect 7616 24596 7622 24608
rect 9324 24596 9352 24636
rect 12158 24624 12164 24676
rect 12216 24664 12222 24676
rect 13832 24664 13860 24763
rect 13998 24760 14004 24812
rect 14056 24800 14062 24812
rect 14056 24772 14136 24800
rect 14056 24760 14062 24772
rect 14108 24732 14136 24772
rect 14182 24760 14188 24812
rect 14240 24809 14246 24812
rect 14752 24809 14780 24840
rect 14240 24803 14295 24809
rect 14240 24769 14249 24803
rect 14283 24800 14295 24803
rect 14737 24803 14795 24809
rect 14737 24800 14749 24803
rect 14283 24772 14749 24800
rect 14283 24769 14295 24772
rect 14240 24763 14295 24769
rect 14737 24769 14749 24772
rect 14783 24769 14795 24803
rect 14737 24763 14795 24769
rect 14240 24760 14246 24763
rect 14826 24760 14832 24812
rect 14884 24760 14890 24812
rect 14921 24803 14979 24809
rect 14921 24769 14933 24803
rect 14967 24769 14979 24803
rect 14921 24763 14979 24769
rect 15105 24804 15163 24809
rect 15194 24804 15200 24812
rect 15105 24803 15200 24804
rect 15105 24769 15117 24803
rect 15151 24776 15200 24803
rect 15151 24769 15163 24776
rect 15105 24763 15163 24769
rect 14936 24732 14964 24763
rect 15194 24760 15200 24776
rect 15252 24760 15258 24812
rect 15304 24800 15332 24840
rect 15654 24828 15660 24880
rect 15712 24868 15718 24880
rect 16206 24868 16212 24880
rect 15712 24840 16212 24868
rect 15712 24828 15718 24840
rect 16206 24828 16212 24840
rect 16264 24828 16270 24880
rect 16945 24871 17003 24877
rect 16945 24837 16957 24871
rect 16991 24868 17003 24871
rect 17126 24868 17132 24880
rect 16991 24840 17132 24868
rect 16991 24837 17003 24840
rect 16945 24831 17003 24837
rect 17126 24828 17132 24840
rect 17184 24828 17190 24880
rect 17310 24828 17316 24880
rect 17368 24868 17374 24880
rect 17862 24868 17868 24880
rect 17368 24840 17868 24868
rect 17368 24828 17374 24840
rect 17862 24828 17868 24840
rect 17920 24828 17926 24880
rect 16850 24800 16856 24812
rect 15304 24772 16856 24800
rect 16850 24760 16856 24772
rect 16908 24760 16914 24812
rect 17037 24803 17095 24809
rect 17037 24769 17049 24803
rect 17083 24769 17095 24803
rect 17037 24763 17095 24769
rect 17221 24803 17279 24809
rect 17221 24769 17233 24803
rect 17267 24800 17279 24803
rect 17402 24800 17408 24812
rect 17267 24772 17408 24800
rect 17267 24769 17279 24772
rect 17221 24763 17279 24769
rect 14108 24704 14964 24732
rect 12216 24636 13860 24664
rect 14936 24664 14964 24704
rect 17052 24664 17080 24763
rect 17402 24760 17408 24772
rect 17460 24760 17466 24812
rect 18064 24744 18092 24908
rect 19889 24905 19901 24939
rect 19935 24936 19947 24939
rect 20530 24936 20536 24948
rect 19935 24908 20536 24936
rect 19935 24905 19947 24908
rect 19889 24899 19947 24905
rect 20530 24896 20536 24908
rect 20588 24896 20594 24948
rect 22186 24896 22192 24948
rect 22244 24936 22250 24948
rect 22830 24936 22836 24948
rect 22244 24908 22836 24936
rect 22244 24896 22250 24908
rect 22830 24896 22836 24908
rect 22888 24896 22894 24948
rect 27893 24939 27951 24945
rect 27893 24905 27905 24939
rect 27939 24936 27951 24939
rect 28166 24936 28172 24948
rect 27939 24908 28172 24936
rect 27939 24905 27951 24908
rect 27893 24899 27951 24905
rect 28166 24896 28172 24908
rect 28224 24896 28230 24948
rect 28534 24896 28540 24948
rect 28592 24936 28598 24948
rect 28994 24936 29000 24948
rect 28592 24908 29000 24936
rect 28592 24896 28598 24908
rect 28994 24896 29000 24908
rect 29052 24896 29058 24948
rect 30282 24896 30288 24948
rect 30340 24936 30346 24948
rect 30340 24908 31708 24936
rect 30340 24896 30346 24908
rect 18690 24828 18696 24880
rect 18748 24868 18754 24880
rect 23382 24868 23388 24880
rect 18748 24840 23388 24868
rect 18748 24828 18754 24840
rect 18138 24760 18144 24812
rect 18196 24800 18202 24812
rect 18601 24803 18659 24809
rect 18601 24800 18613 24803
rect 18196 24772 18613 24800
rect 18196 24760 18202 24772
rect 18601 24769 18613 24772
rect 18647 24800 18659 24803
rect 18782 24800 18788 24812
rect 18647 24772 18788 24800
rect 18647 24769 18659 24772
rect 18601 24763 18659 24769
rect 18782 24760 18788 24772
rect 18840 24760 18846 24812
rect 19334 24760 19340 24812
rect 19392 24800 19398 24812
rect 19521 24803 19579 24809
rect 19521 24800 19533 24803
rect 19392 24772 19533 24800
rect 19392 24760 19398 24772
rect 19521 24769 19533 24772
rect 19567 24800 19579 24803
rect 20162 24800 20168 24812
rect 19567 24772 20168 24800
rect 19567 24769 19579 24772
rect 19521 24763 19579 24769
rect 20162 24760 20168 24772
rect 20220 24800 20226 24812
rect 21174 24800 21180 24812
rect 20220 24772 21180 24800
rect 20220 24760 20226 24772
rect 21174 24760 21180 24772
rect 21232 24800 21238 24812
rect 22002 24800 22008 24812
rect 21232 24772 22008 24800
rect 21232 24760 21238 24772
rect 22002 24760 22008 24772
rect 22060 24760 22066 24812
rect 22281 24803 22339 24809
rect 22281 24769 22293 24803
rect 22327 24800 22339 24803
rect 22833 24803 22891 24809
rect 22327 24772 22784 24800
rect 22327 24769 22339 24772
rect 22281 24763 22339 24769
rect 18046 24692 18052 24744
rect 18104 24732 18110 24744
rect 18690 24732 18696 24744
rect 18104 24704 18696 24732
rect 18104 24692 18110 24704
rect 18690 24692 18696 24704
rect 18748 24692 18754 24744
rect 18969 24735 19027 24741
rect 18969 24701 18981 24735
rect 19015 24732 19027 24735
rect 19429 24735 19487 24741
rect 19429 24732 19441 24735
rect 19015 24704 19441 24732
rect 19015 24701 19027 24704
rect 18969 24695 19027 24701
rect 19429 24701 19441 24704
rect 19475 24701 19487 24735
rect 19429 24695 19487 24701
rect 20806 24692 20812 24744
rect 20864 24732 20870 24744
rect 22373 24735 22431 24741
rect 20864 24704 22232 24732
rect 20864 24692 20870 24704
rect 21358 24664 21364 24676
rect 14936 24636 21364 24664
rect 12216 24624 12222 24636
rect 21358 24624 21364 24636
rect 21416 24624 21422 24676
rect 22204 24664 22232 24704
rect 22373 24701 22385 24735
rect 22419 24701 22431 24735
rect 22756 24732 22784 24772
rect 22833 24769 22845 24803
rect 22879 24800 22891 24803
rect 22922 24800 22928 24812
rect 22879 24772 22928 24800
rect 22879 24769 22891 24772
rect 22833 24763 22891 24769
rect 22922 24760 22928 24772
rect 22980 24760 22986 24812
rect 23032 24809 23060 24840
rect 23382 24828 23388 24840
rect 23440 24828 23446 24880
rect 23842 24868 23848 24880
rect 23803 24840 23848 24868
rect 23842 24828 23848 24840
rect 23900 24868 23906 24880
rect 23900 24840 24348 24868
rect 23900 24828 23906 24840
rect 23017 24803 23075 24809
rect 23017 24769 23029 24803
rect 23063 24769 23075 24803
rect 23017 24763 23075 24769
rect 23106 24760 23112 24812
rect 23164 24760 23170 24812
rect 23201 24803 23259 24809
rect 23201 24769 23213 24803
rect 23247 24800 23259 24803
rect 23247 24772 23520 24800
rect 23247 24769 23259 24772
rect 23201 24763 23259 24769
rect 23382 24732 23388 24744
rect 22756 24704 23388 24732
rect 22373 24695 22431 24701
rect 22388 24664 22416 24695
rect 23382 24692 23388 24704
rect 23440 24692 23446 24744
rect 23492 24664 23520 24772
rect 23566 24760 23572 24812
rect 23624 24800 23630 24812
rect 23661 24803 23719 24809
rect 23661 24800 23673 24803
rect 23624 24772 23673 24800
rect 23624 24760 23630 24772
rect 23661 24769 23673 24772
rect 23707 24769 23719 24803
rect 23661 24763 23719 24769
rect 23676 24732 23704 24763
rect 23750 24760 23756 24812
rect 23808 24760 23814 24812
rect 24026 24760 24032 24812
rect 24084 24760 24090 24812
rect 24118 24760 24124 24812
rect 24176 24760 24182 24812
rect 24320 24809 24348 24840
rect 26418 24828 26424 24880
rect 26476 24868 26482 24880
rect 28074 24868 28080 24880
rect 26476 24840 27292 24868
rect 26476 24828 26482 24840
rect 24305 24803 24363 24809
rect 24305 24769 24317 24803
rect 24351 24769 24363 24803
rect 24305 24763 24363 24769
rect 24394 24760 24400 24812
rect 24452 24760 24458 24812
rect 24494 24803 24552 24809
rect 24494 24769 24506 24803
rect 24540 24769 24552 24803
rect 24494 24763 24552 24769
rect 24509 24732 24537 24763
rect 24854 24760 24860 24812
rect 24912 24800 24918 24812
rect 24949 24803 25007 24809
rect 24949 24800 24961 24803
rect 24912 24772 24961 24800
rect 24912 24760 24918 24772
rect 24949 24769 24961 24772
rect 24995 24769 25007 24803
rect 24949 24763 25007 24769
rect 25866 24760 25872 24812
rect 25924 24800 25930 24812
rect 25924 24772 26654 24800
rect 25924 24760 25930 24772
rect 23676 24704 24537 24732
rect 24670 24692 24676 24744
rect 24728 24741 24734 24744
rect 24728 24735 24748 24741
rect 24736 24701 24748 24735
rect 24728 24695 24748 24701
rect 24728 24692 24734 24695
rect 26234 24692 26240 24744
rect 26292 24692 26298 24744
rect 26418 24692 26424 24744
rect 26476 24692 26482 24744
rect 26252 24664 26280 24692
rect 22204 24636 22416 24664
rect 22480 24636 26280 24664
rect 26626 24664 26654 24772
rect 26970 24760 26976 24812
rect 27028 24760 27034 24812
rect 27154 24760 27160 24812
rect 27212 24760 27218 24812
rect 27264 24809 27292 24840
rect 27724 24840 28080 24868
rect 27249 24803 27307 24809
rect 27249 24769 27261 24803
rect 27295 24769 27307 24803
rect 27249 24763 27307 24769
rect 27430 24760 27436 24812
rect 27488 24760 27494 24812
rect 27522 24760 27528 24812
rect 27580 24760 27586 24812
rect 27617 24803 27675 24809
rect 27617 24769 27629 24803
rect 27663 24800 27675 24803
rect 27724 24800 27752 24840
rect 28074 24828 28080 24840
rect 28132 24828 28138 24880
rect 28629 24871 28687 24877
rect 28629 24837 28641 24871
rect 28675 24868 28687 24871
rect 28675 24840 28994 24868
rect 28675 24837 28687 24840
rect 28629 24831 28687 24837
rect 28966 24800 28994 24840
rect 30558 24828 30564 24880
rect 30616 24828 30622 24880
rect 31680 24868 31708 24908
rect 31754 24896 31760 24948
rect 31812 24936 31818 24948
rect 32214 24936 32220 24948
rect 31812 24908 32220 24936
rect 31812 24896 31818 24908
rect 32214 24896 32220 24908
rect 32272 24896 32278 24948
rect 33686 24896 33692 24948
rect 33744 24936 33750 24948
rect 34057 24939 34115 24945
rect 34057 24936 34069 24939
rect 33744 24908 34069 24936
rect 33744 24896 33750 24908
rect 34057 24905 34069 24908
rect 34103 24905 34115 24939
rect 34057 24899 34115 24905
rect 33704 24868 33732 24896
rect 31680 24840 31754 24868
rect 27663 24772 27752 24800
rect 27816 24772 28764 24800
rect 28966 24772 29224 24800
rect 27663 24769 27675 24772
rect 27617 24763 27675 24769
rect 27816 24664 27844 24772
rect 28736 24744 28764 24772
rect 29196 24744 29224 24772
rect 29270 24760 29276 24812
rect 29328 24800 29334 24812
rect 29917 24803 29975 24809
rect 29917 24800 29929 24803
rect 29328 24772 29929 24800
rect 29328 24760 29334 24772
rect 29917 24769 29929 24772
rect 29963 24800 29975 24803
rect 30193 24803 30251 24809
rect 30193 24800 30205 24803
rect 29963 24772 30205 24800
rect 29963 24769 29975 24772
rect 29917 24763 29975 24769
rect 30193 24769 30205 24772
rect 30239 24769 30251 24803
rect 30193 24763 30251 24769
rect 30377 24803 30435 24809
rect 30377 24769 30389 24803
rect 30423 24769 30435 24803
rect 31726 24800 31754 24840
rect 33428 24840 33732 24868
rect 32030 24800 32036 24812
rect 31726 24772 32036 24800
rect 30377 24763 30435 24769
rect 27893 24735 27951 24741
rect 27893 24701 27905 24735
rect 27939 24701 27951 24735
rect 27893 24695 27951 24701
rect 26626 24636 27844 24664
rect 27908 24664 27936 24695
rect 28718 24692 28724 24744
rect 28776 24692 28782 24744
rect 29178 24692 29184 24744
rect 29236 24692 29242 24744
rect 29733 24735 29791 24741
rect 29733 24701 29745 24735
rect 29779 24732 29791 24735
rect 30392 24732 30420 24763
rect 32030 24760 32036 24772
rect 32088 24760 32094 24812
rect 33428 24809 33456 24840
rect 33229 24803 33287 24809
rect 33229 24769 33241 24803
rect 33275 24769 33287 24803
rect 33229 24763 33287 24769
rect 33413 24803 33471 24809
rect 33413 24769 33425 24803
rect 33459 24769 33471 24803
rect 33413 24763 33471 24769
rect 33597 24803 33655 24809
rect 33597 24769 33609 24803
rect 33643 24800 33655 24803
rect 33962 24800 33968 24812
rect 33643 24772 33968 24800
rect 33643 24769 33655 24772
rect 33597 24763 33655 24769
rect 29779 24704 30420 24732
rect 33244 24732 33272 24763
rect 33962 24760 33968 24772
rect 34020 24760 34026 24812
rect 34072 24732 34100 24899
rect 34440 24840 36492 24868
rect 34440 24812 34468 24840
rect 34422 24760 34428 24812
rect 34480 24760 34486 24812
rect 36170 24760 36176 24812
rect 36228 24800 36234 24812
rect 36464 24809 36492 24840
rect 36357 24803 36415 24809
rect 36357 24800 36369 24803
rect 36228 24772 36369 24800
rect 36228 24760 36234 24772
rect 36357 24769 36369 24772
rect 36403 24769 36415 24803
rect 36357 24763 36415 24769
rect 36449 24803 36507 24809
rect 36449 24769 36461 24803
rect 36495 24800 36507 24803
rect 36495 24772 36952 24800
rect 36495 24769 36507 24772
rect 36449 24763 36507 24769
rect 36924 24744 36952 24772
rect 34149 24735 34207 24741
rect 34149 24732 34161 24735
rect 33244 24704 33456 24732
rect 34072 24704 34161 24732
rect 29779 24701 29791 24704
rect 29733 24695 29791 24701
rect 28169 24667 28227 24673
rect 28169 24664 28181 24667
rect 27908 24636 28181 24664
rect 7616 24568 9352 24596
rect 7616 24556 7622 24568
rect 13814 24556 13820 24608
rect 13872 24596 13878 24608
rect 14369 24599 14427 24605
rect 14369 24596 14381 24599
rect 13872 24568 14381 24596
rect 13872 24556 13878 24568
rect 14369 24565 14381 24568
rect 14415 24565 14427 24599
rect 14369 24559 14427 24565
rect 14553 24599 14611 24605
rect 14553 24565 14565 24599
rect 14599 24596 14611 24599
rect 15010 24596 15016 24608
rect 14599 24568 15016 24596
rect 14599 24565 14611 24568
rect 14553 24559 14611 24565
rect 15010 24556 15016 24568
rect 15068 24556 15074 24608
rect 16669 24599 16727 24605
rect 16669 24565 16681 24599
rect 16715 24596 16727 24599
rect 17126 24596 17132 24608
rect 16715 24568 17132 24596
rect 16715 24565 16727 24568
rect 16669 24559 16727 24565
rect 17126 24556 17132 24568
rect 17184 24556 17190 24608
rect 18506 24556 18512 24608
rect 18564 24596 18570 24608
rect 19886 24596 19892 24608
rect 18564 24568 19892 24596
rect 18564 24556 18570 24568
rect 19886 24556 19892 24568
rect 19944 24556 19950 24608
rect 21634 24556 21640 24608
rect 21692 24596 21698 24608
rect 21821 24599 21879 24605
rect 21821 24596 21833 24599
rect 21692 24568 21833 24596
rect 21692 24556 21698 24568
rect 21821 24565 21833 24568
rect 21867 24565 21879 24599
rect 21821 24559 21879 24565
rect 22002 24556 22008 24608
rect 22060 24596 22066 24608
rect 22480 24596 22508 24636
rect 28169 24633 28181 24636
rect 28215 24633 28227 24667
rect 28169 24627 28227 24633
rect 29932 24608 29960 24704
rect 33428 24676 33456 24704
rect 34149 24701 34161 24704
rect 34195 24701 34207 24735
rect 34149 24695 34207 24701
rect 36541 24735 36599 24741
rect 36541 24701 36553 24735
rect 36587 24701 36599 24735
rect 36541 24695 36599 24701
rect 36633 24735 36691 24741
rect 36633 24701 36645 24735
rect 36679 24732 36691 24735
rect 36722 24732 36728 24744
rect 36679 24704 36728 24732
rect 36679 24701 36691 24704
rect 36633 24695 36691 24701
rect 30742 24624 30748 24676
rect 30800 24664 30806 24676
rect 31386 24664 31392 24676
rect 30800 24636 31392 24664
rect 30800 24624 30806 24636
rect 31386 24624 31392 24636
rect 31444 24664 31450 24676
rect 31444 24636 33364 24664
rect 31444 24624 31450 24636
rect 22060 24568 22508 24596
rect 22060 24556 22066 24568
rect 23106 24556 23112 24608
rect 23164 24596 23170 24608
rect 23385 24599 23443 24605
rect 23385 24596 23397 24599
rect 23164 24568 23397 24596
rect 23164 24556 23170 24568
rect 23385 24565 23397 24568
rect 23431 24565 23443 24599
rect 23385 24559 23443 24565
rect 23474 24556 23480 24608
rect 23532 24556 23538 24608
rect 24394 24556 24400 24608
rect 24452 24596 24458 24608
rect 25130 24596 25136 24608
rect 24452 24568 25136 24596
rect 24452 24556 24458 24568
rect 25130 24556 25136 24568
rect 25188 24556 25194 24608
rect 27062 24556 27068 24608
rect 27120 24596 27126 24608
rect 27709 24599 27767 24605
rect 27709 24596 27721 24599
rect 27120 24568 27721 24596
rect 27120 24556 27126 24568
rect 27709 24565 27721 24568
rect 27755 24565 27767 24599
rect 27709 24559 27767 24565
rect 29914 24556 29920 24608
rect 29972 24556 29978 24608
rect 30101 24599 30159 24605
rect 30101 24565 30113 24599
rect 30147 24596 30159 24599
rect 31018 24596 31024 24608
rect 30147 24568 31024 24596
rect 30147 24565 30159 24568
rect 30101 24559 30159 24565
rect 31018 24556 31024 24568
rect 31076 24556 31082 24608
rect 31294 24556 31300 24608
rect 31352 24596 31358 24608
rect 33042 24596 33048 24608
rect 31352 24568 33048 24596
rect 31352 24556 31358 24568
rect 33042 24556 33048 24568
rect 33100 24556 33106 24608
rect 33226 24556 33232 24608
rect 33284 24556 33290 24608
rect 33336 24596 33364 24636
rect 33410 24624 33416 24676
rect 33468 24624 33474 24676
rect 34333 24667 34391 24673
rect 34333 24664 34345 24667
rect 33796 24636 34345 24664
rect 33796 24608 33824 24636
rect 34333 24633 34345 24636
rect 34379 24633 34391 24667
rect 36556 24664 36584 24695
rect 36722 24692 36728 24704
rect 36780 24692 36786 24744
rect 36906 24692 36912 24744
rect 36964 24692 36970 24744
rect 36556 24636 36676 24664
rect 34333 24627 34391 24633
rect 36648 24608 36676 24636
rect 33689 24599 33747 24605
rect 33689 24596 33701 24599
rect 33336 24568 33701 24596
rect 33689 24565 33701 24568
rect 33735 24565 33747 24599
rect 33689 24559 33747 24565
rect 33778 24556 33784 24608
rect 33836 24556 33842 24608
rect 34238 24556 34244 24608
rect 34296 24556 34302 24608
rect 36630 24556 36636 24608
rect 36688 24556 36694 24608
rect 36814 24556 36820 24608
rect 36872 24556 36878 24608
rect 1104 24506 38272 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38272 24506
rect 1104 24432 38272 24454
rect 4706 24352 4712 24404
rect 4764 24352 4770 24404
rect 6549 24395 6607 24401
rect 6549 24361 6561 24395
rect 6595 24392 6607 24395
rect 6730 24392 6736 24404
rect 6595 24364 6736 24392
rect 6595 24361 6607 24364
rect 6549 24355 6607 24361
rect 6730 24352 6736 24364
rect 6788 24352 6794 24404
rect 6914 24352 6920 24404
rect 6972 24352 6978 24404
rect 9766 24392 9772 24404
rect 9232 24364 9772 24392
rect 2958 24216 2964 24268
rect 3016 24256 3022 24268
rect 3694 24256 3700 24268
rect 3016 24228 3700 24256
rect 3016 24216 3022 24228
rect 3694 24216 3700 24228
rect 3752 24216 3758 24268
rect 4525 24259 4583 24265
rect 4525 24225 4537 24259
rect 4571 24256 4583 24259
rect 4614 24256 4620 24268
rect 4571 24228 4620 24256
rect 4571 24225 4583 24228
rect 4525 24219 4583 24225
rect 4614 24216 4620 24228
rect 4672 24216 4678 24268
rect 4724 24256 4752 24352
rect 5537 24259 5595 24265
rect 4724 24228 4844 24256
rect 2685 24191 2743 24197
rect 2685 24157 2697 24191
rect 2731 24188 2743 24191
rect 2774 24188 2780 24200
rect 2731 24160 2780 24188
rect 2731 24157 2743 24160
rect 2685 24151 2743 24157
rect 2774 24148 2780 24160
rect 2832 24148 2838 24200
rect 3786 24148 3792 24200
rect 3844 24148 3850 24200
rect 3970 24148 3976 24200
rect 4028 24188 4034 24200
rect 4709 24191 4767 24197
rect 4709 24188 4721 24191
rect 4028 24160 4721 24188
rect 4028 24148 4034 24160
rect 4709 24157 4721 24160
rect 4755 24157 4767 24191
rect 4709 24151 4767 24157
rect 2314 24012 2320 24064
rect 2372 24012 2378 24064
rect 2777 24055 2835 24061
rect 2777 24021 2789 24055
rect 2823 24052 2835 24055
rect 3988 24052 4016 24148
rect 4816 24120 4844 24228
rect 5537 24225 5549 24259
rect 5583 24256 5595 24259
rect 6932 24256 6960 24352
rect 5583 24228 5672 24256
rect 5583 24225 5595 24228
rect 5537 24219 5595 24225
rect 5644 24200 5672 24228
rect 5736 24228 6960 24256
rect 5077 24191 5135 24197
rect 5077 24157 5089 24191
rect 5123 24188 5135 24191
rect 5123 24160 5304 24188
rect 5123 24157 5135 24160
rect 5077 24151 5135 24157
rect 4816 24092 5028 24120
rect 2823 24024 4016 24052
rect 4433 24055 4491 24061
rect 2823 24021 2835 24024
rect 2777 24015 2835 24021
rect 4433 24021 4445 24055
rect 4479 24052 4491 24055
rect 4798 24052 4804 24064
rect 4479 24024 4804 24052
rect 4479 24021 4491 24024
rect 4433 24015 4491 24021
rect 4798 24012 4804 24024
rect 4856 24012 4862 24064
rect 5000 24061 5028 24092
rect 5276 24064 5304 24160
rect 5626 24148 5632 24200
rect 5684 24148 5690 24200
rect 5736 24197 5764 24228
rect 5721 24191 5779 24197
rect 5721 24157 5733 24191
rect 5767 24157 5779 24191
rect 5721 24151 5779 24157
rect 5905 24191 5963 24197
rect 5905 24157 5917 24191
rect 5951 24188 5963 24191
rect 6086 24188 6092 24200
rect 5951 24160 6092 24188
rect 5951 24157 5963 24160
rect 5905 24151 5963 24157
rect 6086 24148 6092 24160
rect 6144 24188 6150 24200
rect 6638 24188 6644 24200
rect 6144 24160 6644 24188
rect 6144 24148 6150 24160
rect 6638 24148 6644 24160
rect 6696 24148 6702 24200
rect 6748 24197 6776 24228
rect 6733 24191 6791 24197
rect 6733 24157 6745 24191
rect 6779 24157 6791 24191
rect 6733 24151 6791 24157
rect 6914 24148 6920 24200
rect 6972 24148 6978 24200
rect 9232 24197 9260 24364
rect 9766 24352 9772 24364
rect 9824 24352 9830 24404
rect 11882 24352 11888 24404
rect 11940 24352 11946 24404
rect 12158 24352 12164 24404
rect 12216 24352 12222 24404
rect 12710 24352 12716 24404
rect 12768 24392 12774 24404
rect 12768 24364 16068 24392
rect 12768 24352 12774 24364
rect 11974 24284 11980 24336
rect 12032 24284 12038 24336
rect 12176 24256 12204 24352
rect 12342 24284 12348 24336
rect 12400 24324 12406 24336
rect 16040 24333 16068 24364
rect 16206 24352 16212 24404
rect 16264 24392 16270 24404
rect 19058 24392 19064 24404
rect 16264 24364 19064 24392
rect 16264 24352 16270 24364
rect 19058 24352 19064 24364
rect 19116 24352 19122 24404
rect 19702 24352 19708 24404
rect 19760 24392 19766 24404
rect 25409 24395 25467 24401
rect 19760 24364 24348 24392
rect 19760 24352 19766 24364
rect 15105 24327 15163 24333
rect 15105 24324 15117 24327
rect 12400 24296 15117 24324
rect 12400 24284 12406 24296
rect 15105 24293 15117 24296
rect 15151 24293 15163 24327
rect 15105 24287 15163 24293
rect 16025 24327 16083 24333
rect 16025 24293 16037 24327
rect 16071 24293 16083 24327
rect 16025 24287 16083 24293
rect 17586 24284 17592 24336
rect 17644 24324 17650 24336
rect 17644 24296 21680 24324
rect 17644 24284 17650 24296
rect 9324 24228 12204 24256
rect 13265 24259 13323 24265
rect 9217 24191 9275 24197
rect 9217 24157 9229 24191
rect 9263 24157 9275 24191
rect 9217 24151 9275 24157
rect 5534 24080 5540 24132
rect 5592 24120 5598 24132
rect 5994 24120 6000 24132
rect 5592 24092 6000 24120
rect 5592 24080 5598 24092
rect 5994 24080 6000 24092
rect 6052 24120 6058 24132
rect 9324 24120 9352 24228
rect 13265 24225 13277 24259
rect 13311 24256 13323 24259
rect 13722 24256 13728 24268
rect 13311 24228 13728 24256
rect 13311 24225 13323 24228
rect 13265 24219 13323 24225
rect 13722 24216 13728 24228
rect 13780 24256 13786 24268
rect 13780 24228 14136 24256
rect 13780 24216 13786 24228
rect 9490 24148 9496 24200
rect 9548 24148 9554 24200
rect 12342 24148 12348 24200
rect 12400 24148 12406 24200
rect 13173 24191 13231 24197
rect 13173 24157 13185 24191
rect 13219 24157 13231 24191
rect 13173 24151 13231 24157
rect 9769 24123 9827 24129
rect 9769 24120 9781 24123
rect 6052 24092 9352 24120
rect 9416 24092 9781 24120
rect 6052 24080 6058 24092
rect 4985 24055 5043 24061
rect 4985 24021 4997 24055
rect 5031 24021 5043 24055
rect 4985 24015 5043 24021
rect 5258 24012 5264 24064
rect 5316 24012 5322 24064
rect 6638 24012 6644 24064
rect 6696 24052 6702 24064
rect 7190 24052 7196 24064
rect 6696 24024 7196 24052
rect 6696 24012 6702 24024
rect 7190 24012 7196 24024
rect 7248 24012 7254 24064
rect 9416 24061 9444 24092
rect 9769 24089 9781 24092
rect 9815 24089 9827 24123
rect 9769 24083 9827 24089
rect 10226 24080 10232 24132
rect 10284 24080 10290 24132
rect 13188 24120 13216 24151
rect 13446 24148 13452 24200
rect 13504 24148 13510 24200
rect 13538 24148 13544 24200
rect 13596 24188 13602 24200
rect 14108 24197 14136 24228
rect 14366 24216 14372 24268
rect 14424 24256 14430 24268
rect 14461 24259 14519 24265
rect 14461 24256 14473 24259
rect 14424 24228 14473 24256
rect 14424 24216 14430 24228
rect 14461 24225 14473 24228
rect 14507 24225 14519 24259
rect 14461 24219 14519 24225
rect 14734 24216 14740 24268
rect 14792 24216 14798 24268
rect 15488 24228 16436 24256
rect 13633 24191 13691 24197
rect 13633 24188 13645 24191
rect 13596 24160 13645 24188
rect 13596 24148 13602 24160
rect 13633 24157 13645 24160
rect 13679 24188 13691 24191
rect 14093 24191 14151 24197
rect 13679 24160 14044 24188
rect 13679 24157 13691 24160
rect 13633 24151 13691 24157
rect 14016 24120 14044 24160
rect 14093 24157 14105 24191
rect 14139 24157 14151 24191
rect 14752 24188 14780 24216
rect 14093 24151 14151 24157
rect 14200 24160 14780 24188
rect 14200 24120 14228 24160
rect 15378 24148 15384 24200
rect 15436 24148 15442 24200
rect 15488 24197 15516 24228
rect 16408 24200 16436 24228
rect 16850 24216 16856 24268
rect 16908 24256 16914 24268
rect 20990 24256 20996 24268
rect 16908 24228 20996 24256
rect 16908 24216 16914 24228
rect 20990 24216 20996 24228
rect 21048 24256 21054 24268
rect 21652 24256 21680 24296
rect 21818 24284 21824 24336
rect 21876 24284 21882 24336
rect 22094 24284 22100 24336
rect 22152 24324 22158 24336
rect 22152 24296 22416 24324
rect 22152 24284 22158 24296
rect 22388 24265 22416 24296
rect 23014 24284 23020 24336
rect 23072 24284 23078 24336
rect 23658 24284 23664 24336
rect 23716 24284 23722 24336
rect 22373 24259 22431 24265
rect 21048 24228 21588 24256
rect 21652 24228 22094 24256
rect 21048 24216 21054 24228
rect 15473 24191 15531 24197
rect 15473 24157 15485 24191
rect 15519 24157 15531 24191
rect 15473 24151 15531 24157
rect 15565 24191 15623 24197
rect 15565 24157 15577 24191
rect 15611 24157 15623 24191
rect 15565 24151 15623 24157
rect 15749 24191 15807 24197
rect 15749 24157 15761 24191
rect 15795 24188 15807 24191
rect 16022 24188 16028 24200
rect 15795 24160 16028 24188
rect 15795 24157 15807 24160
rect 15749 24151 15807 24157
rect 11072 24092 13216 24120
rect 13556 24092 13768 24120
rect 14016 24092 14228 24120
rect 14277 24123 14335 24129
rect 9401 24055 9459 24061
rect 9401 24021 9413 24055
rect 9447 24021 9459 24055
rect 9401 24015 9459 24021
rect 9582 24012 9588 24064
rect 9640 24052 9646 24064
rect 11072 24052 11100 24092
rect 9640 24024 11100 24052
rect 11241 24055 11299 24061
rect 9640 24012 9646 24024
rect 11241 24021 11253 24055
rect 11287 24052 11299 24055
rect 11514 24052 11520 24064
rect 11287 24024 11520 24052
rect 11287 24021 11299 24024
rect 11241 24015 11299 24021
rect 11514 24012 11520 24024
rect 11572 24012 11578 24064
rect 11606 24012 11612 24064
rect 11664 24052 11670 24064
rect 13556 24052 13584 24092
rect 11664 24024 13584 24052
rect 13740 24052 13768 24092
rect 14277 24089 14289 24123
rect 14323 24120 14335 24123
rect 14642 24120 14648 24132
rect 14323 24092 14648 24120
rect 14323 24089 14335 24092
rect 14277 24083 14335 24089
rect 14642 24080 14648 24092
rect 14700 24080 14706 24132
rect 15580 24120 15608 24151
rect 16022 24148 16028 24160
rect 16080 24148 16086 24200
rect 16390 24148 16396 24200
rect 16448 24148 16454 24200
rect 16758 24148 16764 24200
rect 16816 24148 16822 24200
rect 18690 24148 18696 24200
rect 18748 24188 18754 24200
rect 18748 24160 20300 24188
rect 18748 24148 18754 24160
rect 20162 24120 20168 24132
rect 15580 24092 20168 24120
rect 20162 24080 20168 24092
rect 20220 24080 20226 24132
rect 20272 24120 20300 24160
rect 20714 24148 20720 24200
rect 20772 24188 20778 24200
rect 21269 24191 21327 24197
rect 21269 24188 21281 24191
rect 20772 24160 21281 24188
rect 20772 24148 20778 24160
rect 21269 24157 21281 24160
rect 21315 24157 21327 24191
rect 21269 24151 21327 24157
rect 21358 24148 21364 24200
rect 21416 24188 21422 24200
rect 21453 24191 21511 24197
rect 21453 24188 21465 24191
rect 21416 24160 21465 24188
rect 21416 24148 21422 24160
rect 21453 24157 21465 24160
rect 21499 24157 21511 24191
rect 21560 24188 21588 24228
rect 21642 24191 21700 24197
rect 21642 24188 21654 24191
rect 21560 24160 21654 24188
rect 21453 24151 21511 24157
rect 21642 24157 21654 24160
rect 21688 24157 21700 24191
rect 21642 24151 21700 24157
rect 21545 24123 21603 24129
rect 21545 24120 21557 24123
rect 20272 24092 21557 24120
rect 21545 24089 21557 24092
rect 21591 24089 21603 24123
rect 22066 24120 22094 24228
rect 22373 24225 22385 24259
rect 22419 24225 22431 24259
rect 22373 24219 22431 24225
rect 22554 24216 22560 24268
rect 22612 24265 22618 24268
rect 22612 24259 22631 24265
rect 22619 24225 22631 24259
rect 23032 24256 23060 24284
rect 24320 24256 24348 24364
rect 25409 24361 25421 24395
rect 25455 24392 25467 24395
rect 25866 24392 25872 24404
rect 25455 24364 25872 24392
rect 25455 24361 25467 24364
rect 25409 24355 25467 24361
rect 25866 24352 25872 24364
rect 25924 24352 25930 24404
rect 26602 24352 26608 24404
rect 26660 24392 26666 24404
rect 26789 24395 26847 24401
rect 26789 24392 26801 24395
rect 26660 24364 26801 24392
rect 26660 24352 26666 24364
rect 26789 24361 26801 24364
rect 26835 24361 26847 24395
rect 26789 24355 26847 24361
rect 27065 24395 27123 24401
rect 27065 24361 27077 24395
rect 27111 24392 27123 24395
rect 27430 24392 27436 24404
rect 27111 24364 27436 24392
rect 27111 24361 27123 24364
rect 27065 24355 27123 24361
rect 26804 24256 26832 24355
rect 27430 24352 27436 24364
rect 27488 24352 27494 24404
rect 27522 24352 27528 24404
rect 27580 24392 27586 24404
rect 27709 24395 27767 24401
rect 27709 24392 27721 24395
rect 27580 24364 27721 24392
rect 27580 24352 27586 24364
rect 27709 24361 27721 24364
rect 27755 24361 27767 24395
rect 27709 24355 27767 24361
rect 28626 24352 28632 24404
rect 28684 24352 28690 24404
rect 28994 24352 29000 24404
rect 29052 24392 29058 24404
rect 29089 24395 29147 24401
rect 29089 24392 29101 24395
rect 29052 24364 29101 24392
rect 29052 24352 29058 24364
rect 29089 24361 29101 24364
rect 29135 24361 29147 24395
rect 29089 24355 29147 24361
rect 31021 24395 31079 24401
rect 31021 24361 31033 24395
rect 31067 24392 31079 24395
rect 31570 24392 31576 24404
rect 31067 24364 31576 24392
rect 31067 24361 31079 24364
rect 31021 24355 31079 24361
rect 31570 24352 31576 24364
rect 31628 24352 31634 24404
rect 33134 24352 33140 24404
rect 33192 24352 33198 24404
rect 34885 24395 34943 24401
rect 34885 24361 34897 24395
rect 34931 24392 34943 24395
rect 34931 24364 35296 24392
rect 34931 24361 34943 24364
rect 34885 24355 34943 24361
rect 27614 24284 27620 24336
rect 27672 24284 27678 24336
rect 29730 24324 29736 24336
rect 28460 24296 29736 24324
rect 23032 24228 23428 24256
rect 22612 24219 22631 24225
rect 22612 24216 22618 24219
rect 22278 24148 22284 24200
rect 22336 24148 22342 24200
rect 22922 24188 22928 24200
rect 22664 24160 22928 24188
rect 22664 24120 22692 24160
rect 22922 24148 22928 24160
rect 22980 24188 22986 24200
rect 23109 24191 23167 24197
rect 23109 24188 23121 24191
rect 22980 24160 23121 24188
rect 22980 24148 22986 24160
rect 23109 24157 23121 24160
rect 23155 24157 23167 24191
rect 23109 24151 23167 24157
rect 23198 24148 23204 24200
rect 23256 24188 23262 24200
rect 23400 24197 23428 24228
rect 24320 24228 26372 24256
rect 26804 24228 27384 24256
rect 23293 24191 23351 24197
rect 23293 24188 23305 24191
rect 23256 24160 23305 24188
rect 23256 24148 23262 24160
rect 23293 24157 23305 24160
rect 23339 24157 23351 24191
rect 23293 24151 23351 24157
rect 23385 24191 23443 24197
rect 23385 24157 23397 24191
rect 23431 24157 23443 24191
rect 23385 24151 23443 24157
rect 23529 24191 23587 24197
rect 23529 24157 23541 24191
rect 23575 24188 23587 24191
rect 24210 24188 24216 24200
rect 23575 24160 24216 24188
rect 23575 24157 23587 24160
rect 23529 24151 23587 24157
rect 24210 24148 24216 24160
rect 24268 24148 24274 24200
rect 24320 24188 24348 24228
rect 24489 24191 24547 24197
rect 24489 24188 24501 24191
rect 24320 24160 24501 24188
rect 24489 24157 24501 24160
rect 24535 24157 24547 24191
rect 24489 24151 24547 24157
rect 24857 24191 24915 24197
rect 24857 24157 24869 24191
rect 24903 24157 24915 24191
rect 24857 24151 24915 24157
rect 22066 24092 22692 24120
rect 21545 24083 21603 24089
rect 20622 24052 20628 24064
rect 13740 24024 20628 24052
rect 11664 24012 11670 24024
rect 20622 24012 20628 24024
rect 20680 24012 20686 24064
rect 21560 24052 21588 24083
rect 22830 24080 22836 24132
rect 22888 24080 22894 24132
rect 23017 24123 23075 24129
rect 23017 24089 23029 24123
rect 23063 24089 23075 24123
rect 24872 24120 24900 24151
rect 25038 24148 25044 24200
rect 25096 24148 25102 24200
rect 25314 24148 25320 24200
rect 25372 24148 25378 24200
rect 25590 24148 25596 24200
rect 25648 24188 25654 24200
rect 26053 24191 26111 24197
rect 26053 24188 26065 24191
rect 25648 24160 26065 24188
rect 25648 24148 25654 24160
rect 26053 24157 26065 24160
rect 26099 24188 26111 24191
rect 26142 24188 26148 24200
rect 26099 24160 26148 24188
rect 26099 24157 26111 24160
rect 26053 24151 26111 24157
rect 26142 24148 26148 24160
rect 26200 24148 26206 24200
rect 26344 24197 26372 24228
rect 27356 24197 27384 24228
rect 27632 24197 27660 24284
rect 27890 24216 27896 24268
rect 27948 24256 27954 24268
rect 27948 24228 28396 24256
rect 27948 24216 27954 24228
rect 26329 24191 26387 24197
rect 26329 24157 26341 24191
rect 26375 24157 26387 24191
rect 26329 24151 26387 24157
rect 27249 24191 27307 24197
rect 27249 24157 27261 24191
rect 27295 24157 27307 24191
rect 27249 24151 27307 24157
rect 27341 24191 27399 24197
rect 27341 24157 27353 24191
rect 27387 24157 27399 24191
rect 27341 24151 27399 24157
rect 27525 24191 27583 24197
rect 27525 24157 27537 24191
rect 27571 24157 27583 24191
rect 27525 24151 27583 24157
rect 27617 24191 27675 24197
rect 27617 24157 27629 24191
rect 27663 24157 27675 24191
rect 27617 24151 27675 24157
rect 25056 24120 25084 24148
rect 25608 24120 25636 24148
rect 24872 24092 24992 24120
rect 25056 24092 25636 24120
rect 26513 24123 26571 24129
rect 23017 24083 23075 24089
rect 21634 24052 21640 24064
rect 21560 24024 21640 24052
rect 21634 24012 21640 24024
rect 21692 24012 21698 24064
rect 22462 24012 22468 24064
rect 22520 24012 22526 24064
rect 23032 24052 23060 24083
rect 24854 24052 24860 24064
rect 23032 24024 24860 24052
rect 24854 24012 24860 24024
rect 24912 24012 24918 24064
rect 24964 24052 24992 24092
rect 26513 24089 26525 24123
rect 26559 24120 26571 24123
rect 26697 24123 26755 24129
rect 26697 24120 26709 24123
rect 26559 24092 26709 24120
rect 26559 24089 26571 24092
rect 26513 24083 26571 24089
rect 26697 24089 26709 24092
rect 26743 24089 26755 24123
rect 27264 24120 27292 24151
rect 27264 24092 27476 24120
rect 26697 24083 26755 24089
rect 27448 24064 27476 24092
rect 25774 24052 25780 24064
rect 24964 24024 25780 24052
rect 25774 24012 25780 24024
rect 25832 24012 25838 24064
rect 27430 24012 27436 24064
rect 27488 24012 27494 24064
rect 27540 24052 27568 24151
rect 27798 24148 27804 24200
rect 27856 24188 27862 24200
rect 27982 24188 27988 24200
rect 27856 24160 27988 24188
rect 27856 24148 27862 24160
rect 27982 24148 27988 24160
rect 28040 24148 28046 24200
rect 28077 24191 28135 24197
rect 28077 24157 28089 24191
rect 28123 24157 28135 24191
rect 28077 24151 28135 24157
rect 28093 24120 28121 24151
rect 28166 24148 28172 24200
rect 28224 24148 28230 24200
rect 28368 24197 28396 24228
rect 28460 24197 28488 24296
rect 29730 24284 29736 24296
rect 29788 24284 29794 24336
rect 32214 24284 32220 24336
rect 32272 24324 32278 24336
rect 32272 24296 35020 24324
rect 32272 24284 32278 24296
rect 28810 24216 28816 24268
rect 28868 24256 28874 24268
rect 28868 24228 29224 24256
rect 28868 24216 28874 24228
rect 28353 24191 28411 24197
rect 28353 24157 28365 24191
rect 28399 24157 28411 24191
rect 28353 24151 28411 24157
rect 28445 24191 28503 24197
rect 28445 24157 28457 24191
rect 28491 24157 28503 24191
rect 28445 24151 28503 24157
rect 28460 24120 28488 24151
rect 28718 24148 28724 24200
rect 28776 24148 28782 24200
rect 28902 24148 28908 24200
rect 28960 24148 28966 24200
rect 29196 24197 29224 24228
rect 31386 24216 31392 24268
rect 31444 24256 31450 24268
rect 31757 24259 31815 24265
rect 31757 24256 31769 24259
rect 31444 24228 31769 24256
rect 31444 24216 31450 24228
rect 31757 24225 31769 24228
rect 31803 24225 31815 24259
rect 31757 24219 31815 24225
rect 32861 24201 32919 24207
rect 32861 24200 32873 24201
rect 32907 24200 32919 24201
rect 28997 24191 29055 24197
rect 28997 24157 29009 24191
rect 29043 24157 29055 24191
rect 28997 24151 29055 24157
rect 29181 24191 29239 24197
rect 29181 24157 29193 24191
rect 29227 24157 29239 24191
rect 29181 24151 29239 24157
rect 28093 24092 28488 24120
rect 28629 24123 28687 24129
rect 28629 24089 28641 24123
rect 28675 24120 28687 24123
rect 29012 24120 29040 24151
rect 30098 24148 30104 24200
rect 30156 24148 30162 24200
rect 30466 24148 30472 24200
rect 30524 24148 30530 24200
rect 30834 24148 30840 24200
rect 30892 24148 30898 24200
rect 31941 24191 31999 24197
rect 31941 24157 31953 24191
rect 31987 24188 31999 24191
rect 32030 24188 32036 24200
rect 31987 24160 32036 24188
rect 31987 24157 31999 24160
rect 31941 24151 31999 24157
rect 32030 24148 32036 24160
rect 32088 24148 32094 24200
rect 32122 24148 32128 24200
rect 32180 24188 32186 24200
rect 32858 24188 32864 24200
rect 32180 24160 32864 24188
rect 32916 24198 32922 24200
rect 32916 24170 32951 24198
rect 33689 24191 33747 24197
rect 32180 24148 32186 24160
rect 32858 24148 32864 24160
rect 32916 24148 32922 24170
rect 33689 24157 33701 24191
rect 33735 24157 33747 24191
rect 33689 24151 33747 24157
rect 29638 24120 29644 24132
rect 28675 24092 28856 24120
rect 29012 24092 29644 24120
rect 28675 24089 28687 24092
rect 28629 24083 28687 24089
rect 27614 24052 27620 24064
rect 27540 24024 27620 24052
rect 27614 24012 27620 24024
rect 27672 24012 27678 24064
rect 28828 24061 28856 24092
rect 29638 24080 29644 24092
rect 29696 24120 29702 24132
rect 30116 24120 30144 24148
rect 29696 24092 30144 24120
rect 29696 24080 29702 24092
rect 30558 24080 30564 24132
rect 30616 24120 30622 24132
rect 30653 24123 30711 24129
rect 30653 24120 30665 24123
rect 30616 24092 30665 24120
rect 30616 24080 30622 24092
rect 30653 24089 30665 24092
rect 30699 24089 30711 24123
rect 30653 24083 30711 24089
rect 30742 24080 30748 24132
rect 30800 24080 30806 24132
rect 31864 24092 32536 24120
rect 28813 24055 28871 24061
rect 28813 24021 28825 24055
rect 28859 24052 28871 24055
rect 28902 24052 28908 24064
rect 28859 24024 28908 24052
rect 28859 24021 28871 24024
rect 28813 24015 28871 24021
rect 28902 24012 28908 24024
rect 28960 24012 28966 24064
rect 29822 24012 29828 24064
rect 29880 24052 29886 24064
rect 31864 24052 31892 24092
rect 29880 24024 31892 24052
rect 29880 24012 29886 24024
rect 31938 24012 31944 24064
rect 31996 24052 32002 24064
rect 32033 24055 32091 24061
rect 32033 24052 32045 24055
rect 31996 24024 32045 24052
rect 31996 24012 32002 24024
rect 32033 24021 32045 24024
rect 32079 24021 32091 24055
rect 32033 24015 32091 24021
rect 32398 24012 32404 24064
rect 32456 24012 32462 24064
rect 32508 24052 32536 24092
rect 33042 24080 33048 24132
rect 33100 24080 33106 24132
rect 33137 24123 33195 24129
rect 33137 24089 33149 24123
rect 33183 24120 33195 24123
rect 33318 24120 33324 24132
rect 33183 24092 33324 24120
rect 33183 24089 33195 24092
rect 33137 24083 33195 24089
rect 33318 24080 33324 24092
rect 33376 24120 33382 24132
rect 33704 24120 33732 24151
rect 33778 24148 33784 24200
rect 33836 24188 33842 24200
rect 33965 24191 34023 24197
rect 33965 24188 33977 24191
rect 33836 24160 33977 24188
rect 33836 24148 33842 24160
rect 33965 24157 33977 24160
rect 34011 24157 34023 24191
rect 33965 24151 34023 24157
rect 34422 24148 34428 24200
rect 34480 24148 34486 24200
rect 34606 24148 34612 24200
rect 34664 24188 34670 24200
rect 34701 24191 34759 24197
rect 34701 24188 34713 24191
rect 34664 24160 34713 24188
rect 34664 24148 34670 24160
rect 34701 24157 34713 24160
rect 34747 24157 34759 24191
rect 34701 24151 34759 24157
rect 34882 24148 34888 24200
rect 34940 24148 34946 24200
rect 34992 24188 35020 24296
rect 35268 24256 35296 24364
rect 35621 24327 35679 24333
rect 35621 24293 35633 24327
rect 35667 24324 35679 24327
rect 36262 24324 36268 24336
rect 35667 24296 36268 24324
rect 35667 24293 35679 24296
rect 35621 24287 35679 24293
rect 36262 24284 36268 24296
rect 36320 24284 36326 24336
rect 35713 24259 35771 24265
rect 35713 24256 35725 24259
rect 35268 24228 35725 24256
rect 35713 24225 35725 24228
rect 35759 24225 35771 24259
rect 35713 24219 35771 24225
rect 35158 24188 35164 24200
rect 35216 24197 35222 24200
rect 35216 24191 35249 24197
rect 34992 24160 35164 24188
rect 35158 24148 35164 24160
rect 35237 24157 35249 24191
rect 35216 24151 35249 24157
rect 35216 24148 35222 24151
rect 36078 24148 36084 24200
rect 36136 24188 36142 24200
rect 36998 24198 37004 24200
rect 36541 24191 36599 24197
rect 36541 24188 36553 24191
rect 36136 24160 36553 24188
rect 36136 24148 36142 24160
rect 36541 24157 36553 24160
rect 36587 24188 36599 24191
rect 36832 24188 37004 24198
rect 36587 24170 37004 24188
rect 36587 24160 36860 24170
rect 36587 24157 36599 24160
rect 36541 24151 36599 24157
rect 36998 24148 37004 24170
rect 37056 24148 37062 24200
rect 37182 24148 37188 24200
rect 37240 24148 37246 24200
rect 34440 24120 34468 24148
rect 36912 24132 36964 24138
rect 33376 24092 34468 24120
rect 34517 24123 34575 24129
rect 33376 24080 33382 24092
rect 34517 24089 34529 24123
rect 34563 24120 34575 24123
rect 34563 24092 35296 24120
rect 34563 24089 34575 24092
rect 34517 24083 34575 24089
rect 32766 24052 32772 24064
rect 32508 24024 32772 24052
rect 32766 24012 32772 24024
rect 32824 24052 32830 24064
rect 32953 24055 33011 24061
rect 32953 24052 32965 24055
rect 32824 24024 32965 24052
rect 32824 24012 32830 24024
rect 32953 24021 32965 24024
rect 32999 24021 33011 24055
rect 33060 24052 33088 24080
rect 35268 24064 35296 24092
rect 36912 24074 36964 24080
rect 35069 24055 35127 24061
rect 35069 24052 35081 24055
rect 33060 24024 35081 24052
rect 32953 24015 33011 24021
rect 35069 24021 35081 24024
rect 35115 24021 35127 24055
rect 35069 24015 35127 24021
rect 35250 24012 35256 24064
rect 35308 24012 35314 24064
rect 1104 23962 38272 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 38272 23962
rect 1104 23888 38272 23910
rect 2314 23808 2320 23860
rect 2372 23808 2378 23860
rect 2777 23851 2835 23857
rect 2777 23817 2789 23851
rect 2823 23848 2835 23851
rect 3786 23848 3792 23860
rect 2823 23820 3792 23848
rect 2823 23817 2835 23820
rect 2777 23811 2835 23817
rect 3786 23808 3792 23820
rect 3844 23808 3850 23860
rect 9490 23848 9496 23860
rect 5460 23820 9496 23848
rect 2332 23780 2360 23808
rect 1964 23752 2360 23780
rect 2409 23783 2467 23789
rect 1964 23721 1992 23752
rect 2409 23749 2421 23783
rect 2455 23780 2467 23783
rect 3878 23780 3884 23792
rect 2455 23752 3884 23780
rect 2455 23749 2467 23752
rect 2409 23743 2467 23749
rect 3878 23740 3884 23752
rect 3936 23740 3942 23792
rect 4062 23740 4068 23792
rect 4120 23740 4126 23792
rect 5460 23724 5488 23820
rect 9490 23808 9496 23820
rect 9548 23808 9554 23860
rect 9582 23808 9588 23860
rect 9640 23808 9646 23860
rect 11422 23808 11428 23860
rect 11480 23848 11486 23860
rect 11974 23848 11980 23860
rect 11480 23820 11980 23848
rect 11480 23808 11486 23820
rect 11974 23808 11980 23820
rect 12032 23848 12038 23860
rect 13081 23851 13139 23857
rect 13081 23848 13093 23851
rect 12032 23820 13093 23848
rect 12032 23808 12038 23820
rect 13081 23817 13093 23820
rect 13127 23817 13139 23851
rect 13081 23811 13139 23817
rect 13449 23851 13507 23857
rect 13449 23817 13461 23851
rect 13495 23848 13507 23851
rect 13998 23848 14004 23860
rect 13495 23820 14004 23848
rect 13495 23817 13507 23820
rect 13449 23811 13507 23817
rect 13998 23808 14004 23820
rect 14056 23808 14062 23860
rect 16390 23808 16396 23860
rect 16448 23848 16454 23860
rect 16669 23851 16727 23857
rect 16669 23848 16681 23851
rect 16448 23820 16681 23848
rect 16448 23808 16454 23820
rect 16669 23817 16681 23820
rect 16715 23817 16727 23851
rect 24026 23848 24032 23860
rect 16669 23811 16727 23817
rect 16776 23820 24032 23848
rect 6822 23780 6828 23792
rect 6656 23752 6828 23780
rect 1949 23715 2007 23721
rect 1949 23681 1961 23715
rect 1995 23681 2007 23715
rect 1949 23675 2007 23681
rect 2225 23715 2283 23721
rect 2225 23681 2237 23715
rect 2271 23681 2283 23715
rect 2225 23675 2283 23681
rect 2501 23715 2559 23721
rect 2501 23681 2513 23715
rect 2547 23681 2559 23715
rect 2501 23675 2559 23681
rect 2593 23715 2651 23721
rect 2593 23681 2605 23715
rect 2639 23712 2651 23715
rect 2639 23684 4384 23712
rect 2639 23681 2651 23684
rect 2593 23675 2651 23681
rect 1762 23468 1768 23520
rect 1820 23468 1826 23520
rect 2240 23508 2268 23675
rect 2516 23576 2544 23675
rect 3510 23604 3516 23656
rect 3568 23644 3574 23656
rect 3970 23644 3976 23656
rect 3568 23616 3976 23644
rect 3568 23604 3574 23616
rect 3970 23604 3976 23616
rect 4028 23604 4034 23656
rect 4356 23644 4384 23684
rect 5442 23672 5448 23724
rect 5500 23672 5506 23724
rect 6656 23721 6684 23752
rect 6822 23740 6828 23752
rect 6880 23740 6886 23792
rect 7374 23740 7380 23792
rect 7432 23740 7438 23792
rect 9398 23740 9404 23792
rect 9456 23780 9462 23792
rect 9600 23780 9628 23808
rect 9456 23752 9628 23780
rect 9456 23740 9462 23752
rect 11330 23740 11336 23792
rect 11388 23780 11394 23792
rect 12342 23780 12348 23792
rect 11388 23752 12348 23780
rect 11388 23740 11394 23752
rect 12342 23740 12348 23752
rect 12400 23780 12406 23792
rect 13173 23783 13231 23789
rect 13173 23780 13185 23783
rect 12400 23752 13185 23780
rect 12400 23740 12406 23752
rect 13173 23749 13185 23752
rect 13219 23749 13231 23783
rect 13173 23743 13231 23749
rect 13630 23740 13636 23792
rect 13688 23780 13694 23792
rect 16776 23780 16804 23820
rect 24026 23808 24032 23820
rect 24084 23808 24090 23860
rect 27246 23848 27252 23860
rect 25332 23820 27252 23848
rect 13688 23752 16804 23780
rect 20901 23783 20959 23789
rect 13688 23740 13694 23752
rect 20901 23749 20913 23783
rect 20947 23780 20959 23783
rect 21174 23780 21180 23792
rect 20947 23752 21180 23780
rect 20947 23749 20959 23752
rect 20901 23743 20959 23749
rect 21174 23740 21180 23752
rect 21232 23740 21238 23792
rect 21358 23740 21364 23792
rect 21416 23780 21422 23792
rect 23842 23780 23848 23792
rect 21416 23752 23848 23780
rect 21416 23740 21422 23752
rect 23842 23740 23848 23752
rect 23900 23740 23906 23792
rect 23937 23783 23995 23789
rect 23937 23749 23949 23783
rect 23983 23780 23995 23783
rect 24210 23780 24216 23792
rect 23983 23752 24216 23780
rect 23983 23749 23995 23752
rect 23937 23743 23995 23749
rect 24210 23740 24216 23752
rect 24268 23780 24274 23792
rect 25332 23780 25360 23820
rect 27246 23808 27252 23820
rect 27304 23808 27310 23860
rect 27338 23808 27344 23860
rect 27396 23848 27402 23860
rect 28994 23848 29000 23860
rect 27396 23820 29000 23848
rect 27396 23808 27402 23820
rect 28994 23808 29000 23820
rect 29052 23808 29058 23860
rect 31021 23851 31079 23857
rect 31021 23817 31033 23851
rect 31067 23848 31079 23851
rect 31938 23848 31944 23860
rect 31067 23820 31944 23848
rect 31067 23817 31079 23820
rect 31021 23811 31079 23817
rect 31938 23808 31944 23820
rect 31996 23808 32002 23860
rect 32398 23808 32404 23860
rect 32456 23848 32462 23860
rect 32456 23820 32904 23848
rect 32456 23808 32462 23820
rect 24268 23752 25360 23780
rect 25501 23783 25559 23789
rect 24268 23740 24274 23752
rect 25501 23749 25513 23783
rect 25547 23780 25559 23783
rect 29270 23780 29276 23792
rect 25547 23752 29276 23780
rect 25547 23749 25559 23752
rect 25501 23743 25559 23749
rect 29270 23740 29276 23752
rect 29328 23780 29334 23792
rect 29454 23780 29460 23792
rect 29328 23752 29460 23780
rect 29328 23740 29334 23752
rect 29454 23740 29460 23752
rect 29512 23740 29518 23792
rect 32766 23780 32772 23792
rect 31726 23752 32772 23780
rect 6641 23715 6699 23721
rect 6641 23681 6653 23715
rect 6687 23681 6699 23715
rect 6641 23675 6699 23681
rect 9309 23715 9367 23721
rect 9309 23681 9321 23715
rect 9355 23681 9367 23715
rect 9309 23675 9367 23681
rect 4614 23644 4620 23656
rect 4356 23616 4620 23644
rect 4614 23604 4620 23616
rect 4672 23604 4678 23656
rect 4798 23604 4804 23656
rect 4856 23644 4862 23656
rect 5077 23647 5135 23653
rect 5077 23644 5089 23647
rect 4856 23616 5089 23644
rect 4856 23604 4862 23616
rect 5077 23613 5089 23616
rect 5123 23613 5135 23647
rect 5077 23607 5135 23613
rect 6914 23604 6920 23656
rect 6972 23604 6978 23656
rect 9030 23604 9036 23656
rect 9088 23644 9094 23656
rect 9324 23644 9352 23675
rect 11514 23672 11520 23724
rect 11572 23672 11578 23724
rect 12897 23715 12955 23721
rect 12897 23712 12909 23715
rect 11624 23684 12909 23712
rect 11624 23644 11652 23684
rect 12897 23681 12909 23684
rect 12943 23712 12955 23715
rect 12943 23684 13216 23712
rect 12943 23681 12955 23684
rect 12897 23675 12955 23681
rect 9088 23616 11652 23644
rect 9088 23604 9094 23616
rect 11882 23604 11888 23656
rect 11940 23604 11946 23656
rect 13188 23644 13216 23684
rect 13262 23672 13268 23724
rect 13320 23712 13326 23724
rect 13725 23715 13783 23721
rect 13725 23712 13737 23715
rect 13320 23684 13737 23712
rect 13320 23672 13326 23684
rect 13725 23681 13737 23684
rect 13771 23681 13783 23715
rect 13725 23675 13783 23681
rect 14093 23715 14151 23721
rect 14093 23681 14105 23715
rect 14139 23712 14151 23715
rect 14182 23712 14188 23724
rect 14139 23684 14188 23712
rect 14139 23681 14151 23684
rect 14093 23675 14151 23681
rect 14182 23672 14188 23684
rect 14240 23672 14246 23724
rect 14461 23715 14519 23721
rect 14461 23681 14473 23715
rect 14507 23712 14519 23715
rect 14642 23712 14648 23724
rect 14507 23684 14648 23712
rect 14507 23681 14519 23684
rect 14461 23675 14519 23681
rect 14476 23644 14504 23675
rect 14642 23672 14648 23684
rect 14700 23672 14706 23724
rect 17034 23672 17040 23724
rect 17092 23672 17098 23724
rect 17586 23672 17592 23724
rect 17644 23712 17650 23724
rect 18417 23715 18475 23721
rect 18417 23712 18429 23715
rect 17644 23684 18429 23712
rect 17644 23672 17650 23684
rect 18417 23681 18429 23684
rect 18463 23681 18475 23715
rect 18417 23675 18475 23681
rect 18601 23715 18659 23721
rect 18601 23681 18613 23715
rect 18647 23681 18659 23715
rect 18601 23675 18659 23681
rect 13188 23616 14504 23644
rect 14568 23616 15700 23644
rect 3651 23579 3709 23585
rect 3651 23576 3663 23579
rect 2516 23548 3663 23576
rect 3651 23545 3663 23548
rect 3697 23576 3709 23579
rect 3697 23548 4384 23576
rect 3697 23545 3709 23548
rect 3651 23539 3709 23545
rect 2869 23511 2927 23517
rect 2869 23508 2881 23511
rect 2240 23480 2881 23508
rect 2869 23477 2881 23480
rect 2915 23477 2927 23511
rect 2869 23471 2927 23477
rect 2958 23468 2964 23520
rect 3016 23508 3022 23520
rect 3786 23508 3792 23520
rect 3016 23480 3792 23508
rect 3016 23468 3022 23480
rect 3786 23468 3792 23480
rect 3844 23508 3850 23520
rect 4062 23508 4068 23520
rect 3844 23480 4068 23508
rect 3844 23468 3850 23480
rect 4062 23468 4068 23480
rect 4120 23468 4126 23520
rect 4356 23508 4384 23548
rect 8386 23536 8392 23588
rect 8444 23576 8450 23588
rect 14568 23576 14596 23616
rect 8444 23548 14596 23576
rect 15672 23576 15700 23616
rect 15930 23604 15936 23656
rect 15988 23644 15994 23656
rect 17129 23647 17187 23653
rect 17129 23644 17141 23647
rect 15988 23616 17141 23644
rect 15988 23604 15994 23616
rect 17129 23613 17141 23616
rect 17175 23613 17187 23647
rect 17129 23607 17187 23613
rect 17313 23647 17371 23653
rect 17313 23613 17325 23647
rect 17359 23644 17371 23647
rect 17678 23644 17684 23656
rect 17359 23616 17684 23644
rect 17359 23613 17371 23616
rect 17313 23607 17371 23613
rect 17678 23604 17684 23616
rect 17736 23604 17742 23656
rect 18616 23644 18644 23675
rect 20622 23672 20628 23724
rect 20680 23672 20686 23724
rect 20809 23715 20867 23721
rect 20809 23712 20821 23715
rect 20732 23684 20821 23712
rect 20530 23644 20536 23656
rect 18616 23616 20536 23644
rect 20530 23604 20536 23616
rect 20588 23604 20594 23656
rect 20732 23644 20760 23684
rect 20809 23681 20821 23684
rect 20855 23681 20867 23715
rect 20809 23675 20867 23681
rect 20990 23672 20996 23724
rect 21048 23712 21054 23724
rect 23566 23712 23572 23724
rect 21048 23684 23572 23712
rect 21048 23672 21054 23684
rect 23566 23672 23572 23684
rect 23624 23672 23630 23724
rect 23661 23715 23719 23721
rect 23661 23681 23673 23715
rect 23707 23712 23719 23715
rect 23750 23712 23756 23724
rect 23707 23684 23756 23712
rect 23707 23681 23719 23684
rect 23661 23675 23719 23681
rect 23750 23672 23756 23684
rect 23808 23672 23814 23724
rect 24034 23715 24092 23721
rect 24034 23681 24046 23715
rect 24080 23681 24092 23715
rect 24034 23675 24092 23681
rect 21358 23644 21364 23656
rect 20732 23616 21364 23644
rect 21358 23604 21364 23616
rect 21416 23604 21422 23656
rect 23590 23644 23618 23672
rect 24049 23644 24077 23675
rect 25590 23672 25596 23724
rect 25648 23712 25654 23724
rect 28166 23712 28172 23724
rect 25648 23684 28172 23712
rect 25648 23672 25654 23684
rect 28166 23672 28172 23684
rect 28224 23672 28230 23724
rect 28810 23672 28816 23724
rect 28868 23712 28874 23724
rect 29549 23715 29607 23721
rect 29549 23712 29561 23715
rect 28868 23684 29561 23712
rect 28868 23672 28874 23684
rect 29549 23681 29561 23684
rect 29595 23681 29607 23715
rect 29549 23675 29607 23681
rect 30834 23672 30840 23724
rect 30892 23712 30898 23724
rect 30929 23715 30987 23721
rect 30929 23712 30941 23715
rect 30892 23684 30941 23712
rect 30892 23672 30898 23684
rect 30929 23681 30941 23684
rect 30975 23681 30987 23715
rect 30929 23675 30987 23681
rect 31113 23715 31171 23721
rect 31113 23681 31125 23715
rect 31159 23712 31171 23715
rect 31726 23712 31754 23752
rect 32766 23740 32772 23752
rect 32824 23740 32830 23792
rect 32876 23789 32904 23820
rect 33226 23808 33232 23860
rect 33284 23808 33290 23860
rect 34882 23808 34888 23860
rect 34940 23848 34946 23860
rect 34977 23851 35035 23857
rect 34977 23848 34989 23851
rect 34940 23820 34989 23848
rect 34940 23808 34946 23820
rect 34977 23817 34989 23820
rect 35023 23817 35035 23851
rect 34977 23811 35035 23817
rect 35805 23851 35863 23857
rect 35805 23817 35817 23851
rect 35851 23848 35863 23851
rect 35986 23848 35992 23860
rect 35851 23820 35992 23848
rect 35851 23817 35863 23820
rect 35805 23811 35863 23817
rect 32861 23783 32919 23789
rect 32861 23749 32873 23783
rect 32907 23749 32919 23783
rect 32861 23743 32919 23749
rect 31159 23684 31754 23712
rect 31159 23681 31171 23684
rect 31113 23675 31171 23681
rect 23590 23616 24077 23644
rect 25406 23604 25412 23656
rect 25464 23604 25470 23656
rect 25958 23604 25964 23656
rect 26016 23604 26022 23656
rect 27706 23604 27712 23656
rect 27764 23644 27770 23656
rect 28074 23644 28080 23656
rect 27764 23616 28080 23644
rect 27764 23604 27770 23616
rect 28074 23604 28080 23616
rect 28132 23604 28138 23656
rect 29270 23604 29276 23656
rect 29328 23644 29334 23656
rect 29365 23647 29423 23653
rect 29365 23644 29377 23647
rect 29328 23616 29377 23644
rect 29328 23604 29334 23616
rect 29365 23613 29377 23616
rect 29411 23644 29423 23647
rect 29638 23644 29644 23656
rect 29411 23616 29644 23644
rect 29411 23613 29423 23616
rect 29365 23607 29423 23613
rect 29638 23604 29644 23616
rect 29696 23604 29702 23656
rect 29733 23647 29791 23653
rect 29733 23613 29745 23647
rect 29779 23644 29791 23647
rect 30006 23644 30012 23656
rect 29779 23616 30012 23644
rect 29779 23613 29791 23616
rect 29733 23607 29791 23613
rect 30006 23604 30012 23616
rect 30064 23644 30070 23656
rect 31128 23644 31156 23675
rect 32122 23672 32128 23724
rect 32180 23672 32186 23724
rect 32306 23721 32312 23724
rect 32273 23715 32312 23721
rect 32273 23681 32285 23715
rect 32273 23675 32312 23681
rect 32306 23672 32312 23675
rect 32364 23672 32370 23724
rect 32398 23672 32404 23724
rect 32456 23672 32462 23724
rect 32493 23715 32551 23721
rect 32493 23681 32505 23715
rect 32539 23681 32551 23715
rect 32493 23675 32551 23681
rect 30064 23616 31156 23644
rect 30064 23604 30070 23616
rect 20070 23576 20076 23588
rect 15672 23548 20076 23576
rect 8444 23536 8450 23548
rect 20070 23536 20076 23548
rect 20128 23536 20134 23588
rect 21177 23579 21235 23585
rect 21177 23545 21189 23579
rect 21223 23576 21235 23579
rect 21634 23576 21640 23588
rect 21223 23548 21640 23576
rect 21223 23545 21235 23548
rect 21177 23539 21235 23545
rect 21634 23536 21640 23548
rect 21692 23536 21698 23588
rect 5258 23508 5264 23520
rect 4356 23480 5264 23508
rect 5258 23468 5264 23480
rect 5316 23468 5322 23520
rect 6638 23468 6644 23520
rect 6696 23508 6702 23520
rect 11606 23508 11612 23520
rect 6696 23480 11612 23508
rect 6696 23468 6702 23480
rect 11606 23468 11612 23480
rect 11664 23468 11670 23520
rect 16666 23468 16672 23520
rect 16724 23508 16730 23520
rect 17586 23508 17592 23520
rect 16724 23480 17592 23508
rect 16724 23468 16730 23480
rect 17586 23468 17592 23480
rect 17644 23468 17650 23520
rect 18322 23468 18328 23520
rect 18380 23508 18386 23520
rect 18509 23511 18567 23517
rect 18509 23508 18521 23511
rect 18380 23480 18521 23508
rect 18380 23468 18386 23480
rect 18509 23477 18521 23480
rect 18555 23477 18567 23511
rect 18509 23471 18567 23477
rect 24210 23468 24216 23520
rect 24268 23468 24274 23520
rect 25976 23517 26004 23604
rect 26142 23536 26148 23588
rect 26200 23576 26206 23588
rect 29914 23576 29920 23588
rect 26200 23548 29920 23576
rect 26200 23536 26206 23548
rect 29914 23536 29920 23548
rect 29972 23536 29978 23588
rect 30466 23536 30472 23588
rect 30524 23576 30530 23588
rect 32508 23576 32536 23675
rect 32582 23672 32588 23724
rect 32640 23721 32646 23724
rect 32640 23712 32648 23721
rect 32640 23684 32685 23712
rect 32640 23675 32648 23684
rect 32640 23672 32646 23675
rect 33134 23672 33140 23724
rect 33192 23672 33198 23724
rect 33244 23712 33272 23808
rect 34606 23740 34612 23792
rect 34664 23780 34670 23792
rect 35820 23780 35848 23811
rect 35986 23808 35992 23820
rect 36044 23808 36050 23860
rect 36262 23808 36268 23860
rect 36320 23808 36326 23860
rect 36630 23808 36636 23860
rect 36688 23848 36694 23860
rect 36725 23851 36783 23857
rect 36725 23848 36737 23851
rect 36688 23820 36737 23848
rect 36688 23808 36694 23820
rect 36725 23817 36737 23820
rect 36771 23817 36783 23851
rect 36725 23811 36783 23817
rect 36814 23808 36820 23860
rect 36872 23808 36878 23860
rect 36832 23780 36860 23808
rect 34664 23752 35848 23780
rect 36464 23752 36860 23780
rect 34664 23740 34670 23752
rect 33321 23715 33379 23721
rect 33321 23712 33333 23715
rect 33244 23684 33333 23712
rect 33321 23681 33333 23684
rect 33367 23681 33379 23715
rect 33321 23675 33379 23681
rect 35250 23672 35256 23724
rect 35308 23712 35314 23724
rect 35434 23712 35440 23724
rect 35308 23684 35440 23712
rect 35308 23672 35314 23684
rect 35434 23672 35440 23684
rect 35492 23712 35498 23724
rect 36464 23721 36492 23752
rect 36906 23740 36912 23792
rect 36964 23740 36970 23792
rect 35713 23715 35771 23721
rect 35713 23712 35725 23715
rect 35492 23684 35725 23712
rect 35492 23672 35498 23684
rect 35713 23681 35725 23684
rect 35759 23681 35771 23715
rect 35713 23675 35771 23681
rect 35897 23715 35955 23721
rect 35897 23681 35909 23715
rect 35943 23681 35955 23715
rect 35897 23675 35955 23681
rect 36449 23715 36507 23721
rect 36449 23681 36461 23715
rect 36495 23681 36507 23715
rect 36449 23675 36507 23681
rect 36541 23715 36599 23721
rect 36541 23681 36553 23715
rect 36587 23681 36599 23715
rect 36541 23675 36599 23681
rect 36633 23715 36691 23721
rect 36633 23681 36645 23715
rect 36679 23681 36691 23715
rect 36633 23675 36691 23681
rect 34790 23604 34796 23656
rect 34848 23644 34854 23656
rect 35161 23647 35219 23653
rect 35161 23644 35173 23647
rect 34848 23616 35173 23644
rect 34848 23604 34854 23616
rect 35161 23613 35173 23616
rect 35207 23613 35219 23647
rect 35161 23607 35219 23613
rect 30524 23548 32536 23576
rect 35176 23576 35204 23607
rect 35342 23604 35348 23656
rect 35400 23644 35406 23656
rect 35621 23647 35679 23653
rect 35621 23644 35633 23647
rect 35400 23616 35633 23644
rect 35400 23604 35406 23616
rect 35621 23613 35633 23616
rect 35667 23613 35679 23647
rect 35621 23607 35679 23613
rect 35912 23576 35940 23675
rect 36262 23604 36268 23656
rect 36320 23604 36326 23656
rect 35176 23548 35940 23576
rect 36556 23576 36584 23675
rect 36648 23644 36676 23675
rect 36722 23644 36728 23656
rect 36648 23616 36728 23644
rect 36722 23604 36728 23616
rect 36780 23644 36786 23656
rect 36780 23616 37044 23644
rect 36780 23604 36786 23616
rect 36909 23579 36967 23585
rect 36909 23576 36921 23579
rect 36556 23548 36921 23576
rect 30524 23536 30530 23548
rect 36909 23545 36921 23548
rect 36955 23545 36967 23579
rect 36909 23539 36967 23545
rect 25961 23511 26019 23517
rect 25961 23477 25973 23511
rect 26007 23477 26019 23511
rect 25961 23471 26019 23477
rect 26234 23468 26240 23520
rect 26292 23508 26298 23520
rect 31202 23508 31208 23520
rect 26292 23480 31208 23508
rect 26292 23468 26298 23480
rect 31202 23468 31208 23480
rect 31260 23468 31266 23520
rect 32769 23511 32827 23517
rect 32769 23477 32781 23511
rect 32815 23508 32827 23511
rect 32953 23511 33011 23517
rect 32953 23508 32965 23511
rect 32815 23480 32965 23508
rect 32815 23477 32827 23480
rect 32769 23471 32827 23477
rect 32953 23477 32965 23480
rect 32999 23477 33011 23511
rect 32953 23471 33011 23477
rect 33505 23511 33563 23517
rect 33505 23477 33517 23511
rect 33551 23508 33563 23511
rect 34514 23508 34520 23520
rect 33551 23480 34520 23508
rect 33551 23477 33563 23480
rect 33505 23471 33563 23477
rect 34514 23468 34520 23480
rect 34572 23468 34578 23520
rect 36078 23468 36084 23520
rect 36136 23508 36142 23520
rect 37016 23508 37044 23616
rect 36136 23480 37044 23508
rect 36136 23468 36142 23480
rect 1104 23418 38272 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38272 23418
rect 1104 23344 38272 23366
rect 2866 23264 2872 23316
rect 2924 23264 2930 23316
rect 3145 23307 3203 23313
rect 3145 23273 3157 23307
rect 3191 23304 3203 23307
rect 3510 23304 3516 23316
rect 3191 23276 3516 23304
rect 3191 23273 3203 23276
rect 3145 23267 3203 23273
rect 3510 23264 3516 23276
rect 3568 23264 3574 23316
rect 3878 23264 3884 23316
rect 3936 23264 3942 23316
rect 4249 23307 4307 23313
rect 4249 23273 4261 23307
rect 4295 23304 4307 23307
rect 4614 23304 4620 23316
rect 4295 23276 4620 23304
rect 4295 23273 4307 23276
rect 4249 23267 4307 23273
rect 4614 23264 4620 23276
rect 4672 23264 4678 23316
rect 6914 23264 6920 23316
rect 6972 23304 6978 23316
rect 7009 23307 7067 23313
rect 7009 23304 7021 23307
rect 6972 23276 7021 23304
rect 6972 23264 6978 23276
rect 7009 23273 7021 23276
rect 7055 23273 7067 23307
rect 9585 23307 9643 23313
rect 9585 23304 9597 23307
rect 7009 23267 7067 23273
rect 7116 23276 9597 23304
rect 1673 23171 1731 23177
rect 1673 23137 1685 23171
rect 1719 23168 1731 23171
rect 1762 23168 1768 23180
rect 1719 23140 1768 23168
rect 1719 23137 1731 23140
rect 1673 23131 1731 23137
rect 1762 23128 1768 23140
rect 1820 23128 1826 23180
rect 1394 23060 1400 23112
rect 1452 23060 1458 23112
rect 2884 23100 2912 23264
rect 3694 23196 3700 23248
rect 3752 23236 3758 23248
rect 7116 23236 7144 23276
rect 9585 23273 9597 23276
rect 9631 23273 9643 23307
rect 9585 23267 9643 23273
rect 9769 23307 9827 23313
rect 9769 23273 9781 23307
rect 9815 23273 9827 23307
rect 9769 23267 9827 23273
rect 3752 23208 7144 23236
rect 7285 23239 7343 23245
rect 3752 23196 3758 23208
rect 3988 23109 4016 23208
rect 7285 23205 7297 23239
rect 7331 23205 7343 23239
rect 7285 23199 7343 23205
rect 7300 23168 7328 23199
rect 7742 23196 7748 23248
rect 7800 23236 7806 23248
rect 9784 23236 9812 23267
rect 10226 23264 10232 23316
rect 10284 23304 10290 23316
rect 15746 23304 15752 23316
rect 10284 23276 15752 23304
rect 10284 23264 10290 23276
rect 15746 23264 15752 23276
rect 15804 23264 15810 23316
rect 15841 23307 15899 23313
rect 15841 23273 15853 23307
rect 15887 23304 15899 23307
rect 16666 23304 16672 23316
rect 15887 23276 16672 23304
rect 15887 23273 15899 23276
rect 15841 23267 15899 23273
rect 16666 23264 16672 23276
rect 16724 23264 16730 23316
rect 16758 23264 16764 23316
rect 16816 23264 16822 23316
rect 16945 23307 17003 23313
rect 16945 23273 16957 23307
rect 16991 23304 17003 23307
rect 17034 23304 17040 23316
rect 16991 23276 17040 23304
rect 16991 23273 17003 23276
rect 16945 23267 17003 23273
rect 17034 23264 17040 23276
rect 17092 23264 17098 23316
rect 17144 23276 17954 23304
rect 7800 23208 9812 23236
rect 7800 23196 7806 23208
rect 7208 23140 7328 23168
rect 7929 23171 7987 23177
rect 7208 23109 7236 23140
rect 7929 23137 7941 23171
rect 7975 23168 7987 23171
rect 8110 23168 8116 23180
rect 7975 23140 8116 23168
rect 7975 23137 7987 23140
rect 7929 23131 7987 23137
rect 8110 23128 8116 23140
rect 8168 23128 8174 23180
rect 8386 23128 8392 23180
rect 8444 23128 8450 23180
rect 9784 23168 9812 23208
rect 10318 23196 10324 23248
rect 10376 23196 10382 23248
rect 13262 23236 13268 23248
rect 10428 23208 13268 23236
rect 10336 23168 10364 23196
rect 9784 23140 10364 23168
rect 2806 23072 2912 23100
rect 3973 23103 4031 23109
rect 3973 23069 3985 23103
rect 4019 23069 4031 23103
rect 3973 23063 4031 23069
rect 4341 23103 4399 23109
rect 4341 23069 4353 23103
rect 4387 23069 4399 23103
rect 4341 23063 4399 23069
rect 7193 23103 7251 23109
rect 7193 23069 7205 23103
rect 7239 23069 7251 23103
rect 7193 23063 7251 23069
rect 4356 22964 4384 23063
rect 7282 23060 7288 23112
rect 7340 23100 7346 23112
rect 7653 23103 7711 23109
rect 7653 23100 7665 23103
rect 7340 23072 7665 23100
rect 7340 23060 7346 23072
rect 7653 23069 7665 23072
rect 7699 23069 7711 23103
rect 7653 23063 7711 23069
rect 7745 23035 7803 23041
rect 7745 23001 7757 23035
rect 7791 23032 7803 23035
rect 8404 23032 8432 23128
rect 10428 23100 10456 23208
rect 13262 23196 13268 23208
rect 13320 23236 13326 23248
rect 13449 23239 13507 23245
rect 13449 23236 13461 23239
rect 13320 23208 13461 23236
rect 13320 23196 13326 23208
rect 13449 23205 13461 23208
rect 13495 23205 13507 23239
rect 13449 23199 13507 23205
rect 14366 23196 14372 23248
rect 14424 23236 14430 23248
rect 17144 23236 17172 23276
rect 14424 23208 17172 23236
rect 17681 23239 17739 23245
rect 14424 23196 14430 23208
rect 17681 23205 17693 23239
rect 17727 23205 17739 23239
rect 17926 23236 17954 23276
rect 18874 23264 18880 23316
rect 18932 23304 18938 23316
rect 19245 23307 19303 23313
rect 19245 23304 19257 23307
rect 18932 23276 19257 23304
rect 18932 23264 18938 23276
rect 19245 23273 19257 23276
rect 19291 23273 19303 23307
rect 19245 23267 19303 23273
rect 20162 23264 20168 23316
rect 20220 23264 20226 23316
rect 20898 23264 20904 23316
rect 20956 23304 20962 23316
rect 21358 23304 21364 23316
rect 20956 23276 21364 23304
rect 20956 23264 20962 23276
rect 21358 23264 21364 23276
rect 21416 23264 21422 23316
rect 22094 23264 22100 23316
rect 22152 23304 22158 23316
rect 22373 23307 22431 23313
rect 22373 23304 22385 23307
rect 22152 23276 22385 23304
rect 22152 23264 22158 23276
rect 22373 23273 22385 23276
rect 22419 23273 22431 23307
rect 22373 23267 22431 23273
rect 24578 23264 24584 23316
rect 24636 23304 24642 23316
rect 24949 23307 25007 23313
rect 24949 23304 24961 23307
rect 24636 23276 24961 23304
rect 24636 23264 24642 23276
rect 24949 23273 24961 23276
rect 24995 23273 25007 23307
rect 24949 23267 25007 23273
rect 27614 23264 27620 23316
rect 27672 23264 27678 23316
rect 28810 23304 28816 23316
rect 28000 23276 28816 23304
rect 17926 23208 21220 23236
rect 17681 23199 17739 23205
rect 12621 23171 12679 23177
rect 12621 23168 12633 23171
rect 10888 23140 12633 23168
rect 10888 23109 10916 23140
rect 12621 23137 12633 23140
rect 12667 23137 12679 23171
rect 17696 23168 17724 23199
rect 12621 23131 12679 23137
rect 13556 23140 15240 23168
rect 13556 23112 13584 23140
rect 15212 23112 15240 23140
rect 16500 23140 17724 23168
rect 7791 23004 8432 23032
rect 8496 23072 10456 23100
rect 10873 23103 10931 23109
rect 7791 23001 7803 23004
rect 7745 22995 7803 23001
rect 4706 22964 4712 22976
rect 4356 22936 4712 22964
rect 4706 22924 4712 22936
rect 4764 22964 4770 22976
rect 8496 22964 8524 23072
rect 10873 23069 10885 23103
rect 10919 23069 10931 23103
rect 10873 23063 10931 23069
rect 11054 23060 11060 23112
rect 11112 23060 11118 23112
rect 11606 23060 11612 23112
rect 11664 23100 11670 23112
rect 11977 23103 12035 23109
rect 11977 23100 11989 23103
rect 11664 23072 11989 23100
rect 11664 23060 11670 23072
rect 11977 23069 11989 23072
rect 12023 23100 12035 23103
rect 12069 23103 12127 23109
rect 12069 23100 12081 23103
rect 12023 23072 12081 23100
rect 12023 23069 12035 23072
rect 11977 23063 12035 23069
rect 12069 23069 12081 23072
rect 12115 23069 12127 23103
rect 12069 23063 12127 23069
rect 8662 22992 8668 23044
rect 8720 23032 8726 23044
rect 9953 23035 10011 23041
rect 8720 23004 9904 23032
rect 8720 22992 8726 23004
rect 4764 22936 8524 22964
rect 4764 22924 4770 22936
rect 9766 22924 9772 22976
rect 9824 22924 9830 22976
rect 9876 22964 9904 23004
rect 9953 23001 9965 23035
rect 9999 23032 10011 23035
rect 10778 23032 10784 23044
rect 9999 23004 10784 23032
rect 9999 23001 10011 23004
rect 9953 22995 10011 23001
rect 10778 22992 10784 23004
rect 10836 22992 10842 23044
rect 11514 22992 11520 23044
rect 11572 22992 11578 23044
rect 12084 23032 12112 23063
rect 12158 23060 12164 23112
rect 12216 23100 12222 23112
rect 12253 23103 12311 23109
rect 12253 23100 12265 23103
rect 12216 23072 12265 23100
rect 12216 23060 12222 23072
rect 12253 23069 12265 23072
rect 12299 23100 12311 23103
rect 12299 23072 13032 23100
rect 12299 23069 12311 23072
rect 12253 23063 12311 23069
rect 13004 23041 13032 23072
rect 13538 23060 13544 23112
rect 13596 23060 13602 23112
rect 13722 23060 13728 23112
rect 13780 23060 13786 23112
rect 14458 23060 14464 23112
rect 14516 23100 14522 23112
rect 14553 23103 14611 23109
rect 14553 23100 14565 23103
rect 14516 23072 14565 23100
rect 14516 23060 14522 23072
rect 14553 23069 14565 23072
rect 14599 23069 14611 23103
rect 14553 23063 14611 23069
rect 14918 23060 14924 23112
rect 14976 23060 14982 23112
rect 15102 23060 15108 23112
rect 15160 23060 15166 23112
rect 15194 23060 15200 23112
rect 15252 23060 15258 23112
rect 15654 23060 15660 23112
rect 15712 23060 15718 23112
rect 15838 23060 15844 23112
rect 15896 23060 15902 23112
rect 16500 23109 16528 23140
rect 18322 23128 18328 23180
rect 18380 23128 18386 23180
rect 18616 23140 18828 23168
rect 18616 23112 18644 23140
rect 16485 23103 16543 23109
rect 16485 23069 16497 23103
rect 16531 23069 16543 23103
rect 16485 23063 16543 23069
rect 16669 23103 16727 23109
rect 16669 23069 16681 23103
rect 16715 23100 16727 23103
rect 16715 23072 16988 23100
rect 16715 23069 16727 23072
rect 16669 23063 16727 23069
rect 12805 23035 12863 23041
rect 12805 23032 12817 23035
rect 12084 23004 12817 23032
rect 12805 23001 12817 23004
rect 12851 23001 12863 23035
rect 12805 22995 12863 23001
rect 12989 23035 13047 23041
rect 12989 23001 13001 23035
rect 13035 23032 13047 23035
rect 14476 23032 14504 23060
rect 13035 23004 14504 23032
rect 15856 23032 15884 23060
rect 16960 23044 16988 23072
rect 17034 23060 17040 23112
rect 17092 23100 17098 23112
rect 17221 23103 17279 23109
rect 17221 23100 17233 23103
rect 17092 23072 17233 23100
rect 17092 23060 17098 23072
rect 17221 23069 17233 23072
rect 17267 23069 17279 23103
rect 17221 23063 17279 23069
rect 17310 23060 17316 23112
rect 17368 23060 17374 23112
rect 17402 23060 17408 23112
rect 17460 23060 17466 23112
rect 17589 23103 17647 23109
rect 17589 23069 17601 23103
rect 17635 23069 17647 23103
rect 17589 23063 17647 23069
rect 17972 23072 18368 23100
rect 15856 23004 16804 23032
rect 13035 23001 13047 23004
rect 12989 22995 13047 23001
rect 10226 22964 10232 22976
rect 9876 22936 10232 22964
rect 10226 22924 10232 22936
rect 10284 22924 10290 22976
rect 10502 22924 10508 22976
rect 10560 22964 10566 22976
rect 10597 22967 10655 22973
rect 10597 22964 10609 22967
rect 10560 22936 10609 22964
rect 10560 22924 10566 22936
rect 10597 22933 10609 22936
rect 10643 22964 10655 22967
rect 11606 22964 11612 22976
rect 10643 22936 11612 22964
rect 10643 22933 10655 22936
rect 10597 22927 10655 22933
rect 11606 22924 11612 22936
rect 11664 22924 11670 22976
rect 12434 22924 12440 22976
rect 12492 22924 12498 22976
rect 16022 22924 16028 22976
rect 16080 22924 16086 22976
rect 16776 22964 16804 23004
rect 16850 22992 16856 23044
rect 16908 22992 16914 23044
rect 16942 22992 16948 23044
rect 17000 23032 17006 23044
rect 17604 23032 17632 23063
rect 17000 23004 17632 23032
rect 17000 22992 17006 23004
rect 17972 22964 18000 23072
rect 18049 23035 18107 23041
rect 18049 23001 18061 23035
rect 18095 23032 18107 23035
rect 18095 23004 18276 23032
rect 18095 23001 18107 23004
rect 18049 22995 18107 23001
rect 18248 22976 18276 23004
rect 18340 22976 18368 23072
rect 18414 23060 18420 23112
rect 18472 23100 18478 23112
rect 18509 23103 18567 23109
rect 18509 23100 18521 23103
rect 18472 23072 18521 23100
rect 18472 23060 18478 23072
rect 18509 23069 18521 23072
rect 18555 23069 18567 23103
rect 18509 23063 18567 23069
rect 18598 23060 18604 23112
rect 18656 23060 18662 23112
rect 18690 23060 18696 23112
rect 18748 23060 18754 23112
rect 18800 23032 18828 23140
rect 19702 23128 19708 23180
rect 19760 23128 19766 23180
rect 19889 23171 19947 23177
rect 19889 23137 19901 23171
rect 19935 23168 19947 23171
rect 20806 23168 20812 23180
rect 19935 23140 20812 23168
rect 19935 23137 19947 23140
rect 19889 23131 19947 23137
rect 20272 23109 20300 23140
rect 20806 23128 20812 23140
rect 20864 23128 20870 23180
rect 21192 23168 21220 23208
rect 24854 23196 24860 23248
rect 24912 23196 24918 23248
rect 28000 23236 28028 23276
rect 28810 23264 28816 23276
rect 28868 23264 28874 23316
rect 30285 23307 30343 23313
rect 30285 23273 30297 23307
rect 30331 23304 30343 23307
rect 31294 23304 31300 23316
rect 30331 23276 31300 23304
rect 30331 23273 30343 23276
rect 30285 23267 30343 23273
rect 31294 23264 31300 23276
rect 31352 23264 31358 23316
rect 32674 23264 32680 23316
rect 32732 23264 32738 23316
rect 36262 23264 36268 23316
rect 36320 23304 36326 23316
rect 36449 23307 36507 23313
rect 36449 23304 36461 23307
rect 36320 23276 36461 23304
rect 36320 23264 36326 23276
rect 36449 23273 36461 23276
rect 36495 23273 36507 23307
rect 36449 23267 36507 23273
rect 30742 23236 30748 23248
rect 25332 23208 28028 23236
rect 28092 23208 30748 23236
rect 22557 23171 22615 23177
rect 22557 23168 22569 23171
rect 21192 23140 22569 23168
rect 22557 23137 22569 23140
rect 22603 23168 22615 23171
rect 23382 23168 23388 23180
rect 22603 23140 23388 23168
rect 22603 23137 22615 23140
rect 22557 23131 22615 23137
rect 23382 23128 23388 23140
rect 23440 23128 23446 23180
rect 25041 23171 25099 23177
rect 25041 23168 25053 23171
rect 23860 23140 25053 23168
rect 23860 23112 23888 23140
rect 25041 23137 25053 23140
rect 25087 23168 25099 23171
rect 25332 23168 25360 23208
rect 28092 23177 28120 23208
rect 30742 23196 30748 23208
rect 30800 23236 30806 23248
rect 32122 23236 32128 23248
rect 30800 23208 32128 23236
rect 30800 23196 30806 23208
rect 32122 23196 32128 23208
rect 32180 23196 32186 23248
rect 32217 23239 32275 23245
rect 32217 23205 32229 23239
rect 32263 23236 32275 23239
rect 32692 23236 32720 23264
rect 32263 23208 32720 23236
rect 32263 23205 32275 23208
rect 32217 23199 32275 23205
rect 27985 23171 28043 23177
rect 27985 23168 27997 23171
rect 25087 23140 25360 23168
rect 25424 23140 27997 23168
rect 25087 23137 25099 23140
rect 25041 23131 25099 23137
rect 25424 23112 25452 23140
rect 27985 23137 27997 23140
rect 28031 23137 28043 23171
rect 27985 23131 28043 23137
rect 28077 23171 28135 23177
rect 28077 23137 28089 23171
rect 28123 23137 28135 23171
rect 28077 23131 28135 23137
rect 20257 23103 20315 23109
rect 20257 23069 20269 23103
rect 20303 23069 20315 23103
rect 20257 23063 20315 23069
rect 20441 23103 20499 23109
rect 20441 23069 20453 23103
rect 20487 23100 20499 23103
rect 20993 23103 21051 23109
rect 20993 23100 21005 23103
rect 20487 23072 21005 23100
rect 20487 23069 20499 23072
rect 20441 23063 20499 23069
rect 20993 23069 21005 23072
rect 21039 23069 21051 23103
rect 20993 23063 21051 23069
rect 21177 23103 21235 23109
rect 21177 23069 21189 23103
rect 21223 23069 21235 23103
rect 21177 23063 21235 23069
rect 20456 23032 20484 23063
rect 18800 23004 20484 23032
rect 20717 23035 20775 23041
rect 20717 23001 20729 23035
rect 20763 23032 20775 23035
rect 21192 23032 21220 23063
rect 21358 23060 21364 23112
rect 21416 23060 21422 23112
rect 22925 23103 22983 23109
rect 22925 23069 22937 23103
rect 22971 23100 22983 23103
rect 23290 23100 23296 23112
rect 22971 23072 23296 23100
rect 22971 23069 22983 23072
rect 22925 23063 22983 23069
rect 23290 23060 23296 23072
rect 23348 23060 23354 23112
rect 23842 23060 23848 23112
rect 23900 23060 23906 23112
rect 24765 23103 24823 23109
rect 24765 23069 24777 23103
rect 24811 23100 24823 23103
rect 25406 23100 25412 23112
rect 24811 23072 25412 23100
rect 24811 23069 24823 23072
rect 24765 23063 24823 23069
rect 25406 23060 25412 23072
rect 25464 23060 25470 23112
rect 25774 23060 25780 23112
rect 25832 23100 25838 23112
rect 26510 23100 26516 23112
rect 25832 23072 26516 23100
rect 25832 23060 25838 23072
rect 26510 23060 26516 23072
rect 26568 23060 26574 23112
rect 26697 23103 26755 23109
rect 26697 23069 26709 23103
rect 26743 23069 26755 23103
rect 26697 23063 26755 23069
rect 26881 23103 26939 23109
rect 26881 23069 26893 23103
rect 26927 23100 26939 23103
rect 27430 23100 27436 23112
rect 26927 23072 27436 23100
rect 26927 23069 26939 23072
rect 26881 23063 26939 23069
rect 21266 23032 21272 23044
rect 20763 23004 21128 23032
rect 21192 23004 21272 23032
rect 20763 23001 20775 23004
rect 20717 22995 20775 23001
rect 18141 22967 18199 22973
rect 18141 22964 18153 22967
rect 16776 22936 18153 22964
rect 18141 22933 18153 22936
rect 18187 22933 18199 22967
rect 18141 22927 18199 22933
rect 18230 22924 18236 22976
rect 18288 22924 18294 22976
rect 18322 22924 18328 22976
rect 18380 22964 18386 22976
rect 18601 22967 18659 22973
rect 18601 22964 18613 22967
rect 18380 22936 18613 22964
rect 18380 22924 18386 22936
rect 18601 22933 18613 22936
rect 18647 22933 18659 22967
rect 18601 22927 18659 22933
rect 19610 22924 19616 22976
rect 19668 22924 19674 22976
rect 21100 22964 21128 23004
rect 21266 22992 21272 23004
rect 21324 22992 21330 23044
rect 24394 23032 24400 23044
rect 22664 23004 24400 23032
rect 22664 22964 22692 23004
rect 24394 22992 24400 23004
rect 24452 23032 24458 23044
rect 26234 23032 26240 23044
rect 24452 23004 26240 23032
rect 24452 22992 24458 23004
rect 26234 22992 26240 23004
rect 26292 22992 26298 23044
rect 26712 23032 26740 23063
rect 27430 23060 27436 23072
rect 27488 23100 27494 23112
rect 27614 23100 27620 23112
rect 27488 23072 27620 23100
rect 27488 23060 27494 23072
rect 27614 23060 27620 23072
rect 27672 23060 27678 23112
rect 27798 23060 27804 23112
rect 27856 23060 27862 23112
rect 27893 23103 27951 23109
rect 27893 23069 27905 23103
rect 27939 23069 27951 23103
rect 27893 23063 27951 23069
rect 27908 23032 27936 23063
rect 26344 23004 26740 23032
rect 27264 23004 27936 23032
rect 28000 23032 28028 23131
rect 28718 23128 28724 23180
rect 28776 23168 28782 23180
rect 28776 23140 29040 23168
rect 28776 23128 28782 23140
rect 28810 23060 28816 23112
rect 28868 23060 28874 23112
rect 29012 23109 29040 23140
rect 29178 23128 29184 23180
rect 29236 23128 29242 23180
rect 29917 23171 29975 23177
rect 29917 23137 29929 23171
rect 29963 23168 29975 23171
rect 30466 23168 30472 23180
rect 29963 23140 30472 23168
rect 29963 23137 29975 23140
rect 29917 23131 29975 23137
rect 30466 23128 30472 23140
rect 30524 23128 30530 23180
rect 31662 23168 31668 23180
rect 31623 23140 31668 23168
rect 31662 23128 31668 23140
rect 31720 23168 31726 23180
rect 33870 23168 33876 23180
rect 31720 23140 33876 23168
rect 31720 23128 31726 23140
rect 33870 23128 33876 23140
rect 33928 23128 33934 23180
rect 34514 23128 34520 23180
rect 34572 23128 34578 23180
rect 28997 23103 29055 23109
rect 28997 23069 29009 23103
rect 29043 23069 29055 23103
rect 28997 23063 29055 23069
rect 30098 23060 30104 23112
rect 30156 23060 30162 23112
rect 30282 23060 30288 23112
rect 30340 23060 30346 23112
rect 34532 23100 34560 23128
rect 36633 23103 36691 23109
rect 36633 23100 36645 23103
rect 34532 23072 36645 23100
rect 36633 23069 36645 23072
rect 36679 23069 36691 23103
rect 36633 23063 36691 23069
rect 36814 23060 36820 23112
rect 36872 23100 36878 23112
rect 36909 23103 36967 23109
rect 36909 23100 36921 23103
rect 36872 23072 36921 23100
rect 36872 23060 36878 23072
rect 36909 23069 36921 23072
rect 36955 23069 36967 23103
rect 36909 23063 36967 23069
rect 37093 23103 37151 23109
rect 37093 23069 37105 23103
rect 37139 23069 37151 23103
rect 37093 23063 37151 23069
rect 29178 23032 29184 23044
rect 28000 23004 29184 23032
rect 26344 22976 26372 23004
rect 27264 22976 27292 23004
rect 21100 22936 22692 22964
rect 22738 22924 22744 22976
rect 22796 22924 22802 22976
rect 24854 22924 24860 22976
rect 24912 22964 24918 22976
rect 25590 22964 25596 22976
rect 24912 22936 25596 22964
rect 24912 22924 24918 22936
rect 25590 22924 25596 22936
rect 25648 22924 25654 22976
rect 26326 22924 26332 22976
rect 26384 22924 26390 22976
rect 27246 22924 27252 22976
rect 27304 22924 27310 22976
rect 27908 22964 27936 23004
rect 29178 22992 29184 23004
rect 29236 22992 29242 23044
rect 29270 22992 29276 23044
rect 29328 22992 29334 23044
rect 29638 22992 29644 23044
rect 29696 22992 29702 23044
rect 31478 23032 31484 23044
rect 29748 23004 31484 23032
rect 29288 22964 29316 22992
rect 29748 22976 29776 23004
rect 31478 22992 31484 23004
rect 31536 23032 31542 23044
rect 31849 23035 31907 23041
rect 31849 23032 31861 23035
rect 31536 23004 31861 23032
rect 31536 22992 31542 23004
rect 31849 23001 31861 23004
rect 31895 23032 31907 23035
rect 32214 23032 32220 23044
rect 31895 23004 32220 23032
rect 31895 23001 31907 23004
rect 31849 22995 31907 23001
rect 32214 22992 32220 23004
rect 32272 22992 32278 23044
rect 32674 22992 32680 23044
rect 32732 23032 32738 23044
rect 37108 23032 37136 23063
rect 32732 23004 37136 23032
rect 32732 22992 32738 23004
rect 27908 22936 29316 22964
rect 29730 22924 29736 22976
rect 29788 22924 29794 22976
rect 30466 22924 30472 22976
rect 30524 22924 30530 22976
rect 31018 22924 31024 22976
rect 31076 22964 31082 22976
rect 31757 22967 31815 22973
rect 31757 22964 31769 22967
rect 31076 22936 31769 22964
rect 31076 22924 31082 22936
rect 31757 22933 31769 22936
rect 31803 22933 31815 22967
rect 31757 22927 31815 22933
rect 33870 22924 33876 22976
rect 33928 22964 33934 22976
rect 36722 22964 36728 22976
rect 33928 22936 36728 22964
rect 33928 22924 33934 22936
rect 36722 22924 36728 22936
rect 36780 22924 36786 22976
rect 1104 22874 38272 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 38272 22874
rect 1104 22800 38272 22822
rect 5534 22720 5540 22772
rect 5592 22720 5598 22772
rect 6825 22763 6883 22769
rect 6825 22729 6837 22763
rect 6871 22760 6883 22763
rect 7098 22760 7104 22772
rect 6871 22732 7104 22760
rect 6871 22729 6883 22732
rect 6825 22723 6883 22729
rect 7098 22720 7104 22732
rect 7156 22720 7162 22772
rect 9217 22763 9275 22769
rect 9217 22729 9229 22763
rect 9263 22760 9275 22763
rect 9398 22760 9404 22772
rect 9263 22732 9404 22760
rect 9263 22729 9275 22732
rect 9217 22723 9275 22729
rect 9398 22720 9404 22732
rect 9456 22720 9462 22772
rect 9766 22720 9772 22772
rect 9824 22720 9830 22772
rect 10594 22720 10600 22772
rect 10652 22720 10658 22772
rect 13538 22760 13544 22772
rect 12268 22732 13544 22760
rect 5350 22516 5356 22568
rect 5408 22556 5414 22568
rect 5552 22556 5580 22720
rect 6917 22695 6975 22701
rect 6917 22661 6929 22695
rect 6963 22692 6975 22695
rect 7742 22692 7748 22704
rect 6963 22664 7748 22692
rect 6963 22661 6975 22664
rect 6917 22655 6975 22661
rect 7742 22652 7748 22664
rect 7800 22652 7806 22704
rect 9585 22695 9643 22701
rect 9585 22661 9597 22695
rect 9631 22692 9643 22695
rect 9784 22692 9812 22720
rect 9631 22664 9812 22692
rect 9631 22661 9643 22664
rect 9585 22655 9643 22661
rect 9306 22584 9312 22636
rect 9364 22584 9370 22636
rect 9398 22584 9404 22636
rect 9456 22584 9462 22636
rect 9674 22584 9680 22636
rect 9732 22584 9738 22636
rect 9784 22633 9812 22664
rect 9769 22627 9827 22633
rect 9769 22593 9781 22627
rect 9815 22593 9827 22627
rect 9769 22587 9827 22593
rect 9858 22584 9864 22636
rect 9916 22624 9922 22636
rect 9953 22627 10011 22633
rect 9953 22624 9965 22627
rect 9916 22596 9965 22624
rect 9916 22584 9922 22596
rect 9953 22593 9965 22596
rect 9999 22593 10011 22627
rect 10612 22624 10640 22720
rect 12268 22701 12296 22732
rect 13538 22720 13544 22732
rect 13596 22720 13602 22772
rect 13722 22720 13728 22772
rect 13780 22760 13786 22772
rect 14553 22763 14611 22769
rect 13780 22732 14228 22760
rect 13780 22720 13786 22732
rect 12253 22695 12311 22701
rect 12253 22661 12265 22695
rect 12299 22661 12311 22695
rect 12253 22655 12311 22661
rect 12434 22652 12440 22704
rect 12492 22692 12498 22704
rect 12492 22664 14136 22692
rect 12492 22652 12498 22664
rect 11517 22627 11575 22633
rect 11517 22624 11529 22627
rect 10612 22596 11529 22624
rect 9953 22587 10011 22593
rect 11517 22593 11529 22596
rect 11563 22593 11575 22627
rect 11517 22587 11575 22593
rect 7009 22559 7067 22565
rect 7009 22556 7021 22559
rect 5408 22528 7021 22556
rect 5408 22516 5414 22528
rect 7009 22525 7021 22528
rect 7055 22525 7067 22559
rect 7009 22519 7067 22525
rect 7190 22516 7196 22568
rect 7248 22556 7254 22568
rect 9692 22556 9720 22584
rect 7248 22528 9720 22556
rect 9968 22556 9996 22587
rect 11606 22584 11612 22636
rect 11664 22584 11670 22636
rect 11793 22627 11851 22633
rect 11793 22593 11805 22627
rect 11839 22624 11851 22627
rect 11839 22596 12296 22624
rect 11839 22593 11851 22596
rect 11793 22587 11851 22593
rect 11882 22556 11888 22568
rect 9968 22528 11888 22556
rect 7248 22516 7254 22528
rect 11882 22516 11888 22528
rect 11940 22516 11946 22568
rect 5534 22448 5540 22500
rect 5592 22488 5598 22500
rect 5902 22488 5908 22500
rect 5592 22460 5908 22488
rect 5592 22448 5598 22460
rect 5902 22448 5908 22460
rect 5960 22448 5966 22500
rect 8294 22448 8300 22500
rect 8352 22488 8358 22500
rect 9033 22491 9091 22497
rect 9033 22488 9045 22491
rect 8352 22460 9045 22488
rect 8352 22448 8358 22460
rect 9033 22457 9045 22460
rect 9079 22488 9091 22491
rect 12158 22488 12164 22500
rect 9079 22460 10456 22488
rect 9079 22457 9091 22460
rect 9033 22451 9091 22457
rect 6454 22380 6460 22432
rect 6512 22380 6518 22432
rect 9766 22380 9772 22432
rect 9824 22380 9830 22432
rect 10428 22420 10456 22460
rect 11716 22460 12164 22488
rect 11716 22432 11744 22460
rect 12158 22448 12164 22460
rect 12216 22448 12222 22500
rect 12268 22432 12296 22596
rect 12894 22584 12900 22636
rect 12952 22624 12958 22636
rect 14108 22633 14136 22664
rect 14200 22633 14228 22732
rect 14553 22729 14565 22763
rect 14599 22760 14611 22763
rect 15654 22760 15660 22772
rect 14599 22732 15660 22760
rect 14599 22729 14611 22732
rect 14553 22723 14611 22729
rect 15654 22720 15660 22732
rect 15712 22720 15718 22772
rect 15930 22720 15936 22772
rect 15988 22720 15994 22772
rect 16761 22763 16819 22769
rect 16761 22729 16773 22763
rect 16807 22760 16819 22763
rect 16942 22760 16948 22772
rect 16807 22732 16948 22760
rect 16807 22729 16819 22732
rect 16761 22723 16819 22729
rect 16942 22720 16948 22732
rect 17000 22720 17006 22772
rect 17218 22720 17224 22772
rect 17276 22760 17282 22772
rect 17402 22760 17408 22772
rect 17276 22732 17408 22760
rect 17276 22720 17282 22732
rect 17402 22720 17408 22732
rect 17460 22720 17466 22772
rect 17586 22720 17592 22772
rect 17644 22720 17650 22772
rect 19426 22720 19432 22772
rect 19484 22760 19490 22772
rect 19889 22763 19947 22769
rect 19889 22760 19901 22763
rect 19484 22732 19901 22760
rect 19484 22720 19490 22732
rect 19889 22729 19901 22732
rect 19935 22729 19947 22763
rect 19889 22723 19947 22729
rect 20162 22720 20168 22772
rect 20220 22720 20226 22772
rect 23677 22763 23735 22769
rect 23677 22760 23689 22763
rect 22066 22732 22416 22760
rect 15746 22652 15752 22704
rect 15804 22652 15810 22704
rect 17034 22692 17040 22704
rect 16684 22664 17040 22692
rect 13909 22627 13967 22633
rect 13909 22624 13921 22627
rect 12952 22596 13921 22624
rect 12952 22584 12958 22596
rect 13909 22593 13921 22596
rect 13955 22593 13967 22627
rect 13909 22587 13967 22593
rect 14093 22627 14151 22633
rect 14093 22593 14105 22627
rect 14139 22593 14151 22627
rect 14093 22587 14151 22593
rect 14185 22627 14243 22633
rect 14185 22593 14197 22627
rect 14231 22593 14243 22627
rect 14185 22587 14243 22593
rect 14277 22627 14335 22633
rect 14277 22593 14289 22627
rect 14323 22624 14335 22627
rect 14366 22624 14372 22636
rect 14323 22596 14372 22624
rect 14323 22593 14335 22596
rect 14277 22587 14335 22593
rect 14108 22488 14136 22587
rect 14366 22584 14372 22596
rect 14424 22624 14430 22636
rect 14550 22624 14556 22636
rect 14424 22596 14556 22624
rect 14424 22584 14430 22596
rect 14550 22584 14556 22596
rect 14608 22584 14614 22636
rect 14918 22584 14924 22636
rect 14976 22624 14982 22636
rect 16022 22624 16028 22636
rect 14976 22596 16028 22624
rect 14976 22584 14982 22596
rect 16022 22584 16028 22596
rect 16080 22624 16086 22636
rect 16684 22633 16712 22664
rect 17034 22652 17040 22664
rect 17092 22652 17098 22704
rect 17144 22664 19840 22692
rect 16669 22627 16727 22633
rect 16669 22624 16681 22627
rect 16080 22596 16681 22624
rect 16080 22584 16086 22596
rect 16669 22593 16681 22596
rect 16715 22593 16727 22627
rect 16669 22587 16727 22593
rect 16853 22627 16911 22633
rect 16853 22593 16865 22627
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 15381 22559 15439 22565
rect 15381 22556 15393 22559
rect 14752 22528 15393 22556
rect 14752 22500 14780 22528
rect 15381 22525 15393 22528
rect 15427 22556 15439 22559
rect 16758 22556 16764 22568
rect 15427 22528 16764 22556
rect 15427 22525 15439 22528
rect 15381 22519 15439 22525
rect 16758 22516 16764 22528
rect 16816 22556 16822 22568
rect 16868 22556 16896 22587
rect 17144 22556 17172 22664
rect 17310 22584 17316 22636
rect 17368 22624 17374 22636
rect 17497 22627 17555 22633
rect 17497 22624 17509 22627
rect 17368 22596 17509 22624
rect 17368 22584 17374 22596
rect 17497 22593 17509 22596
rect 17543 22593 17555 22627
rect 17497 22587 17555 22593
rect 17681 22627 17739 22633
rect 17681 22593 17693 22627
rect 17727 22593 17739 22627
rect 18414 22624 18420 22636
rect 17681 22587 17739 22593
rect 18248 22596 18420 22624
rect 16816 22528 16896 22556
rect 16960 22528 17172 22556
rect 16816 22516 16822 22528
rect 14182 22488 14188 22500
rect 14108 22460 14188 22488
rect 14182 22448 14188 22460
rect 14240 22448 14246 22500
rect 14734 22448 14740 22500
rect 14792 22448 14798 22500
rect 14918 22448 14924 22500
rect 14976 22488 14982 22500
rect 15102 22488 15108 22500
rect 14976 22460 15108 22488
rect 14976 22448 14982 22460
rect 15102 22448 15108 22460
rect 15160 22488 15166 22500
rect 16960 22488 16988 22528
rect 15160 22460 16988 22488
rect 15160 22448 15166 22460
rect 17034 22448 17040 22500
rect 17092 22448 17098 22500
rect 17218 22448 17224 22500
rect 17276 22488 17282 22500
rect 17586 22488 17592 22500
rect 17276 22460 17592 22488
rect 17276 22448 17282 22460
rect 17586 22448 17592 22460
rect 17644 22448 17650 22500
rect 17696 22488 17724 22587
rect 17770 22516 17776 22568
rect 17828 22556 17834 22568
rect 18248 22556 18276 22596
rect 18414 22584 18420 22596
rect 18472 22584 18478 22636
rect 19705 22627 19763 22633
rect 19705 22593 19717 22627
rect 19751 22593 19763 22627
rect 19705 22587 19763 22593
rect 17828 22528 18276 22556
rect 17828 22516 17834 22528
rect 18322 22516 18328 22568
rect 18380 22516 18386 22568
rect 18690 22488 18696 22500
rect 17696 22460 18696 22488
rect 11054 22420 11060 22432
rect 10428 22392 11060 22420
rect 11054 22380 11060 22392
rect 11112 22420 11118 22432
rect 11698 22420 11704 22432
rect 11112 22392 11704 22420
rect 11112 22380 11118 22392
rect 11698 22380 11704 22392
rect 11756 22380 11762 22432
rect 12250 22380 12256 22432
rect 12308 22380 12314 22432
rect 15749 22423 15807 22429
rect 15749 22389 15761 22423
rect 15795 22420 15807 22423
rect 15838 22420 15844 22432
rect 15795 22392 15844 22420
rect 15795 22389 15807 22392
rect 15749 22383 15807 22389
rect 15838 22380 15844 22392
rect 15896 22380 15902 22432
rect 17052 22420 17080 22448
rect 17696 22420 17724 22460
rect 18690 22448 18696 22460
rect 18748 22448 18754 22500
rect 19720 22488 19748 22587
rect 19812 22556 19840 22664
rect 19981 22627 20039 22633
rect 19981 22593 19993 22627
rect 20027 22624 20039 22627
rect 20180 22624 20208 22720
rect 22066 22704 22094 22732
rect 22066 22692 22100 22704
rect 20732 22664 22100 22692
rect 20732 22633 20760 22664
rect 22094 22652 22100 22664
rect 22152 22652 22158 22704
rect 20027 22596 20208 22624
rect 20717 22627 20775 22633
rect 20027 22593 20039 22596
rect 19981 22587 20039 22593
rect 20717 22593 20729 22627
rect 20763 22593 20775 22627
rect 20717 22587 20775 22593
rect 20732 22556 20760 22587
rect 20806 22584 20812 22636
rect 20864 22624 20870 22636
rect 22002 22624 22008 22636
rect 20864 22596 22008 22624
rect 20864 22584 20870 22596
rect 22002 22584 22008 22596
rect 22060 22584 22066 22636
rect 22189 22627 22247 22633
rect 22189 22593 22201 22627
rect 22235 22593 22247 22627
rect 22189 22587 22247 22593
rect 19812 22528 20760 22556
rect 21082 22516 21088 22568
rect 21140 22516 21146 22568
rect 22204 22556 22232 22587
rect 22278 22584 22284 22636
rect 22336 22584 22342 22636
rect 22388 22633 22416 22732
rect 23308 22732 23689 22760
rect 22738 22652 22744 22704
rect 22796 22652 22802 22704
rect 23308 22692 23336 22732
rect 23677 22729 23689 22732
rect 23723 22729 23735 22763
rect 23677 22723 23735 22729
rect 23842 22720 23848 22772
rect 23900 22720 23906 22772
rect 24578 22720 24584 22772
rect 24636 22760 24642 22772
rect 25961 22763 26019 22769
rect 24636 22732 25176 22760
rect 24636 22720 24642 22732
rect 23124 22664 23336 22692
rect 22388 22627 22465 22633
rect 22388 22596 22419 22627
rect 22407 22593 22419 22596
rect 22453 22624 22465 22627
rect 23014 22624 23020 22636
rect 22453 22596 23020 22624
rect 22453 22593 22465 22596
rect 22407 22587 22465 22593
rect 23014 22584 23020 22596
rect 23072 22584 23078 22636
rect 23124 22633 23152 22664
rect 23308 22636 23336 22664
rect 23477 22695 23535 22701
rect 23477 22661 23489 22695
rect 23523 22661 23535 22695
rect 23477 22655 23535 22661
rect 23109 22627 23167 22633
rect 23109 22593 23121 22627
rect 23155 22593 23167 22627
rect 23109 22587 23167 22593
rect 23201 22627 23259 22633
rect 23201 22593 23213 22627
rect 23247 22593 23259 22627
rect 23201 22587 23259 22593
rect 23216 22556 23244 22587
rect 23290 22584 23296 22636
rect 23348 22584 23354 22636
rect 23382 22584 23388 22636
rect 23440 22624 23446 22636
rect 23492 22624 23520 22655
rect 23566 22624 23572 22636
rect 23440 22596 23572 22624
rect 23440 22584 23446 22596
rect 23566 22584 23572 22596
rect 23624 22584 23630 22636
rect 24118 22584 24124 22636
rect 24176 22584 24182 22636
rect 24854 22584 24860 22636
rect 24912 22584 24918 22636
rect 25148 22624 25176 22732
rect 25961 22729 25973 22763
rect 26007 22760 26019 22763
rect 26050 22760 26056 22772
rect 26007 22732 26056 22760
rect 26007 22729 26019 22732
rect 25961 22723 26019 22729
rect 26050 22720 26056 22732
rect 26108 22720 26114 22772
rect 26326 22720 26332 22772
rect 26384 22720 26390 22772
rect 26510 22720 26516 22772
rect 26568 22760 26574 22772
rect 26568 22732 27200 22760
rect 26568 22720 26574 22732
rect 25590 22652 25596 22704
rect 25648 22692 25654 22704
rect 26344 22692 26372 22720
rect 27172 22701 27200 22732
rect 29178 22720 29184 22772
rect 29236 22760 29242 22772
rect 29236 22732 30144 22760
rect 29236 22720 29242 22732
rect 26973 22695 27031 22701
rect 26973 22692 26985 22695
rect 25648 22664 25728 22692
rect 25648 22652 25654 22664
rect 25700 22633 25728 22664
rect 26344 22664 26985 22692
rect 25501 22627 25559 22633
rect 25501 22624 25513 22627
rect 25148 22596 25513 22624
rect 25501 22593 25513 22596
rect 25547 22593 25559 22627
rect 25501 22587 25559 22593
rect 25685 22627 25743 22633
rect 25685 22593 25697 22627
rect 25731 22593 25743 22627
rect 25685 22587 25743 22593
rect 25774 22584 25780 22636
rect 25832 22584 25838 22636
rect 26344 22633 26372 22664
rect 26973 22661 26985 22664
rect 27019 22661 27031 22695
rect 26973 22655 27031 22661
rect 27157 22695 27215 22701
rect 27157 22661 27169 22695
rect 27203 22661 27215 22695
rect 27157 22655 27215 22661
rect 27338 22652 27344 22704
rect 27396 22652 27402 22704
rect 27614 22652 27620 22704
rect 27672 22692 27678 22704
rect 28629 22695 28687 22701
rect 27672 22664 28580 22692
rect 27672 22652 27678 22664
rect 26145 22627 26203 22633
rect 26145 22624 26157 22627
rect 25884 22596 26157 22624
rect 22204 22528 23244 22556
rect 24581 22559 24639 22565
rect 22388 22500 22416 22528
rect 24581 22525 24593 22559
rect 24627 22556 24639 22559
rect 24762 22556 24768 22568
rect 24627 22528 24768 22556
rect 24627 22525 24639 22528
rect 24581 22519 24639 22525
rect 24762 22516 24768 22528
rect 24820 22516 24826 22568
rect 24872 22556 24900 22584
rect 24872 22528 25360 22556
rect 22278 22488 22284 22500
rect 19720 22460 22284 22488
rect 22278 22448 22284 22460
rect 22336 22448 22342 22500
rect 22370 22448 22376 22500
rect 22428 22448 22434 22500
rect 22649 22491 22707 22497
rect 22649 22457 22661 22491
rect 22695 22488 22707 22491
rect 25332 22488 25360 22528
rect 25406 22516 25412 22568
rect 25464 22556 25470 22568
rect 25593 22559 25651 22565
rect 25593 22556 25605 22559
rect 25464 22528 25605 22556
rect 25464 22516 25470 22528
rect 25593 22525 25605 22528
rect 25639 22525 25651 22559
rect 25593 22519 25651 22525
rect 25884 22488 25912 22596
rect 26145 22593 26157 22596
rect 26191 22593 26203 22627
rect 26145 22587 26203 22593
rect 26329 22627 26387 22633
rect 26329 22593 26341 22627
rect 26375 22593 26387 22627
rect 26329 22587 26387 22593
rect 27798 22584 27804 22636
rect 27856 22584 27862 22636
rect 27982 22584 27988 22636
rect 28040 22584 28046 22636
rect 28258 22584 28264 22636
rect 28316 22584 28322 22636
rect 28445 22627 28503 22633
rect 28445 22593 28457 22627
rect 28491 22593 28503 22627
rect 28552 22624 28580 22664
rect 28629 22661 28641 22695
rect 28675 22692 28687 22695
rect 29822 22692 29828 22704
rect 28675 22664 29828 22692
rect 28675 22661 28687 22664
rect 28629 22655 28687 22661
rect 29822 22652 29828 22664
rect 29880 22652 29886 22704
rect 30006 22701 30012 22704
rect 29983 22695 30012 22701
rect 29983 22661 29995 22695
rect 29983 22655 30012 22661
rect 30006 22652 30012 22655
rect 30064 22652 30070 22704
rect 30116 22701 30144 22732
rect 30282 22720 30288 22772
rect 30340 22720 30346 22772
rect 30466 22720 30472 22772
rect 30524 22720 30530 22772
rect 30742 22720 30748 22772
rect 30800 22720 30806 22772
rect 31113 22763 31171 22769
rect 31113 22729 31125 22763
rect 31159 22760 31171 22763
rect 31202 22760 31208 22772
rect 31159 22732 31208 22760
rect 31159 22729 31171 22732
rect 31113 22723 31171 22729
rect 31202 22720 31208 22732
rect 31260 22720 31266 22772
rect 31294 22720 31300 22772
rect 31352 22720 31358 22772
rect 31938 22720 31944 22772
rect 31996 22760 32002 22772
rect 32582 22760 32588 22772
rect 31996 22732 32588 22760
rect 31996 22720 32002 22732
rect 32582 22720 32588 22732
rect 32640 22720 32646 22772
rect 33962 22720 33968 22772
rect 34020 22760 34026 22772
rect 34020 22732 34560 22760
rect 34020 22720 34026 22732
rect 30101 22695 30159 22701
rect 30101 22661 30113 22695
rect 30147 22661 30159 22695
rect 30101 22655 30159 22661
rect 30190 22652 30196 22704
rect 30248 22652 30254 22704
rect 30300 22692 30328 22720
rect 30300 22664 30420 22692
rect 28552 22596 28994 22624
rect 28445 22587 28503 22593
rect 26513 22559 26571 22565
rect 26513 22525 26525 22559
rect 26559 22556 26571 22559
rect 27816 22556 27844 22584
rect 26559 22528 27844 22556
rect 28000 22556 28028 22584
rect 28460 22556 28488 22587
rect 28000 22528 28488 22556
rect 26559 22525 26571 22528
rect 26513 22519 26571 22525
rect 22695 22460 25268 22488
rect 25332 22460 25912 22488
rect 22695 22457 22707 22460
rect 22649 22451 22707 22457
rect 17052 22392 17724 22420
rect 17770 22380 17776 22432
rect 17828 22420 17834 22432
rect 18141 22423 18199 22429
rect 18141 22420 18153 22423
rect 17828 22392 18153 22420
rect 17828 22380 17834 22392
rect 18141 22389 18153 22392
rect 18187 22389 18199 22423
rect 18141 22383 18199 22389
rect 19521 22423 19579 22429
rect 19521 22389 19533 22423
rect 19567 22420 19579 22423
rect 20254 22420 20260 22432
rect 19567 22392 20260 22420
rect 19567 22389 19579 22392
rect 19521 22383 19579 22389
rect 20254 22380 20260 22392
rect 20312 22380 20318 22432
rect 23198 22380 23204 22432
rect 23256 22420 23262 22432
rect 23661 22423 23719 22429
rect 23661 22420 23673 22423
rect 23256 22392 23673 22420
rect 23256 22380 23262 22392
rect 23661 22389 23673 22392
rect 23707 22389 23719 22423
rect 25240 22420 25268 22460
rect 25774 22420 25780 22432
rect 25240 22392 25780 22420
rect 23661 22383 23719 22389
rect 25774 22380 25780 22392
rect 25832 22380 25838 22432
rect 28460 22420 28488 22528
rect 28966 22488 28994 22596
rect 29730 22584 29736 22636
rect 29788 22624 29794 22636
rect 30285 22627 30343 22633
rect 29788 22596 29868 22624
rect 29788 22584 29794 22596
rect 29840 22565 29868 22596
rect 30285 22593 30297 22627
rect 30331 22593 30343 22627
rect 30285 22587 30343 22593
rect 29825 22559 29883 22565
rect 29825 22525 29837 22559
rect 29871 22525 29883 22559
rect 29825 22519 29883 22525
rect 30300 22488 30328 22587
rect 30392 22556 30420 22664
rect 30484 22624 30512 22720
rect 30561 22627 30619 22633
rect 30561 22624 30573 22627
rect 30484 22596 30573 22624
rect 30561 22593 30573 22596
rect 30607 22593 30619 22627
rect 30561 22587 30619 22593
rect 30653 22627 30711 22633
rect 30653 22593 30665 22627
rect 30699 22593 30711 22627
rect 30760 22624 30788 22720
rect 31849 22695 31907 22701
rect 31849 22661 31861 22695
rect 31895 22692 31907 22695
rect 32306 22692 32312 22704
rect 31895 22664 32312 22692
rect 31895 22661 31907 22664
rect 31849 22655 31907 22661
rect 32306 22652 32312 22664
rect 32364 22692 32370 22704
rect 33781 22695 33839 22701
rect 32364 22664 32536 22692
rect 32364 22652 32370 22664
rect 32508 22636 32536 22664
rect 33781 22661 33793 22695
rect 33827 22692 33839 22695
rect 33827 22664 34192 22692
rect 33827 22661 33839 22664
rect 33781 22655 33839 22661
rect 30837 22627 30895 22633
rect 30837 22624 30849 22627
rect 30760 22596 30849 22624
rect 30653 22587 30711 22593
rect 30837 22593 30849 22596
rect 30883 22593 30895 22627
rect 30837 22587 30895 22593
rect 30929 22627 30987 22633
rect 30929 22593 30941 22627
rect 30975 22624 30987 22627
rect 31018 22624 31024 22636
rect 30975 22596 31024 22624
rect 30975 22593 30987 22596
rect 30929 22587 30987 22593
rect 30469 22559 30527 22565
rect 30469 22556 30481 22559
rect 30392 22528 30481 22556
rect 30469 22525 30481 22528
rect 30515 22525 30527 22559
rect 30469 22519 30527 22525
rect 30668 22500 30696 22587
rect 31018 22584 31024 22596
rect 31076 22584 31082 22636
rect 31202 22584 31208 22636
rect 31260 22624 31266 22636
rect 31478 22624 31484 22636
rect 31260 22596 31484 22624
rect 31260 22584 31266 22596
rect 31478 22584 31484 22596
rect 31536 22584 31542 22636
rect 31573 22627 31631 22633
rect 31573 22593 31585 22627
rect 31619 22624 31631 22627
rect 32030 22624 32036 22636
rect 31619 22596 32036 22624
rect 31619 22593 31631 22596
rect 31573 22587 31631 22593
rect 32030 22584 32036 22596
rect 32088 22584 32094 22636
rect 32122 22584 32128 22636
rect 32180 22584 32186 22636
rect 32214 22584 32220 22636
rect 32272 22624 32278 22636
rect 32272 22596 32317 22624
rect 32272 22584 32278 22596
rect 32398 22584 32404 22636
rect 32456 22584 32462 22636
rect 32490 22584 32496 22636
rect 32548 22584 32554 22636
rect 32631 22627 32689 22633
rect 32631 22593 32643 22627
rect 32677 22624 32689 22627
rect 32766 22624 32772 22636
rect 32677 22596 32772 22624
rect 32677 22593 32689 22596
rect 32631 22587 32689 22593
rect 32766 22584 32772 22596
rect 32824 22584 32830 22636
rect 33689 22627 33747 22633
rect 33689 22593 33701 22627
rect 33735 22593 33747 22627
rect 33689 22587 33747 22593
rect 31938 22516 31944 22568
rect 31996 22516 32002 22568
rect 30558 22488 30564 22500
rect 28966 22460 30564 22488
rect 30558 22448 30564 22460
rect 30616 22448 30622 22500
rect 30650 22448 30656 22500
rect 30708 22448 30714 22500
rect 28718 22420 28724 22432
rect 28460 22392 28724 22420
rect 28718 22380 28724 22392
rect 28776 22420 28782 22432
rect 29730 22420 29736 22432
rect 28776 22392 29736 22420
rect 28776 22380 28782 22392
rect 29730 22380 29736 22392
rect 29788 22380 29794 22432
rect 30576 22420 30604 22448
rect 32416 22420 32444 22584
rect 33704 22556 33732 22587
rect 33870 22584 33876 22636
rect 33928 22584 33934 22636
rect 34164 22633 34192 22664
rect 34149 22627 34207 22633
rect 34149 22593 34161 22627
rect 34195 22593 34207 22627
rect 34149 22587 34207 22593
rect 34330 22584 34336 22636
rect 34388 22584 34394 22636
rect 34532 22633 34560 22732
rect 34606 22720 34612 22772
rect 34664 22760 34670 22772
rect 35069 22763 35127 22769
rect 35069 22760 35081 22763
rect 34664 22732 35081 22760
rect 34664 22720 34670 22732
rect 35069 22729 35081 22732
rect 35115 22729 35127 22763
rect 35069 22723 35127 22729
rect 35253 22763 35311 22769
rect 35253 22729 35265 22763
rect 35299 22760 35311 22763
rect 35342 22760 35348 22772
rect 35299 22732 35348 22760
rect 35299 22729 35311 22732
rect 35253 22723 35311 22729
rect 35342 22720 35348 22732
rect 35400 22720 35406 22772
rect 35894 22760 35900 22772
rect 35820 22732 35900 22760
rect 35161 22695 35219 22701
rect 35161 22661 35173 22695
rect 35207 22692 35219 22695
rect 35820 22692 35848 22732
rect 35894 22720 35900 22732
rect 35952 22720 35958 22772
rect 35986 22720 35992 22772
rect 36044 22720 36050 22772
rect 36173 22763 36231 22769
rect 36173 22729 36185 22763
rect 36219 22760 36231 22763
rect 36639 22763 36697 22769
rect 36219 22732 36584 22760
rect 36219 22729 36231 22732
rect 36173 22723 36231 22729
rect 36004 22692 36032 22720
rect 36556 22701 36584 22732
rect 36639 22729 36651 22763
rect 36685 22760 36697 22763
rect 36685 22732 37688 22760
rect 36685 22729 36697 22732
rect 36639 22723 36697 22729
rect 35207 22664 35848 22692
rect 35912 22664 36032 22692
rect 36541 22695 36599 22701
rect 35207 22661 35219 22664
rect 35161 22655 35219 22661
rect 34517 22627 34575 22633
rect 34517 22593 34529 22627
rect 34563 22593 34575 22627
rect 34517 22587 34575 22593
rect 34701 22627 34759 22633
rect 34701 22593 34713 22627
rect 34747 22593 34759 22627
rect 34701 22587 34759 22593
rect 34054 22556 34060 22568
rect 33704 22528 34060 22556
rect 34054 22516 34060 22528
rect 34112 22516 34118 22568
rect 34422 22516 34428 22568
rect 34480 22516 34486 22568
rect 34716 22500 34744 22587
rect 34790 22584 34796 22636
rect 34848 22624 34854 22636
rect 35385 22627 35443 22633
rect 35385 22624 35397 22627
rect 34848 22596 35397 22624
rect 34848 22584 34854 22596
rect 35385 22593 35397 22596
rect 35431 22593 35443 22627
rect 35385 22587 35443 22593
rect 35526 22584 35532 22636
rect 35584 22584 35590 22636
rect 35618 22584 35624 22636
rect 35676 22584 35682 22636
rect 35710 22584 35716 22636
rect 35768 22624 35774 22636
rect 35912 22633 35940 22664
rect 36541 22661 36553 22695
rect 36587 22661 36599 22695
rect 36541 22655 36599 22661
rect 36722 22652 36728 22704
rect 36780 22652 36786 22704
rect 35805 22627 35863 22633
rect 35805 22624 35817 22627
rect 35768 22596 35817 22624
rect 35768 22584 35774 22596
rect 35805 22593 35817 22596
rect 35851 22593 35863 22627
rect 35805 22587 35863 22593
rect 35897 22627 35955 22633
rect 35897 22593 35909 22627
rect 35943 22593 35955 22627
rect 35897 22587 35955 22593
rect 35989 22627 36047 22633
rect 35989 22593 36001 22627
rect 36035 22624 36047 22627
rect 36262 22624 36268 22636
rect 36035 22596 36268 22624
rect 36035 22593 36047 22596
rect 35989 22587 36047 22593
rect 36262 22584 36268 22596
rect 36320 22584 36326 22636
rect 36814 22584 36820 22636
rect 36872 22584 36878 22636
rect 37660 22633 37688 22732
rect 37645 22627 37703 22633
rect 37645 22593 37657 22627
rect 37691 22593 37703 22627
rect 37645 22587 37703 22593
rect 34882 22516 34888 22568
rect 34940 22516 34946 22568
rect 37553 22559 37611 22565
rect 37553 22556 37565 22559
rect 36280 22528 37565 22556
rect 36280 22500 36308 22528
rect 37553 22525 37565 22528
rect 37599 22525 37611 22559
rect 37553 22519 37611 22525
rect 33594 22448 33600 22500
rect 33652 22448 33658 22500
rect 34698 22448 34704 22500
rect 34756 22448 34762 22500
rect 36262 22448 36268 22500
rect 36320 22448 36326 22500
rect 30576 22392 32444 22420
rect 32769 22423 32827 22429
rect 32769 22389 32781 22423
rect 32815 22420 32827 22423
rect 32950 22420 32956 22432
rect 32815 22392 32956 22420
rect 32815 22389 32827 22392
rect 32769 22383 32827 22389
rect 32950 22380 32956 22392
rect 33008 22380 33014 22432
rect 33612 22420 33640 22448
rect 35986 22420 35992 22432
rect 33612 22392 35992 22420
rect 35986 22380 35992 22392
rect 36044 22380 36050 22432
rect 37274 22380 37280 22432
rect 37332 22420 37338 22432
rect 37369 22423 37427 22429
rect 37369 22420 37381 22423
rect 37332 22392 37381 22420
rect 37332 22380 37338 22392
rect 37369 22389 37381 22392
rect 37415 22389 37427 22423
rect 37369 22383 37427 22389
rect 1104 22330 38272 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38272 22330
rect 1104 22256 38272 22278
rect 3786 22176 3792 22228
rect 3844 22216 3850 22228
rect 7098 22216 7104 22228
rect 3844 22188 7104 22216
rect 3844 22176 3850 22188
rect 7098 22176 7104 22188
rect 7156 22176 7162 22228
rect 10137 22219 10195 22225
rect 10137 22185 10149 22219
rect 10183 22216 10195 22219
rect 10962 22216 10968 22228
rect 10183 22188 10968 22216
rect 10183 22185 10195 22188
rect 10137 22179 10195 22185
rect 10962 22176 10968 22188
rect 11020 22176 11026 22228
rect 13449 22219 13507 22225
rect 13449 22185 13461 22219
rect 13495 22216 13507 22219
rect 13722 22216 13728 22228
rect 13495 22188 13728 22216
rect 13495 22185 13507 22188
rect 13449 22179 13507 22185
rect 13722 22176 13728 22188
rect 13780 22176 13786 22228
rect 16758 22176 16764 22228
rect 16816 22176 16822 22228
rect 16850 22176 16856 22228
rect 16908 22216 16914 22228
rect 17129 22219 17187 22225
rect 17129 22216 17141 22219
rect 16908 22188 17141 22216
rect 16908 22176 16914 22188
rect 17129 22185 17141 22188
rect 17175 22185 17187 22219
rect 17129 22179 17187 22185
rect 17497 22219 17555 22225
rect 17497 22185 17509 22219
rect 17543 22216 17555 22219
rect 17770 22216 17776 22228
rect 17543 22188 17776 22216
rect 17543 22185 17555 22188
rect 17497 22179 17555 22185
rect 17770 22176 17776 22188
rect 17828 22176 17834 22228
rect 17862 22176 17868 22228
rect 17920 22216 17926 22228
rect 18138 22216 18144 22228
rect 17920 22188 18144 22216
rect 17920 22176 17926 22188
rect 18138 22176 18144 22188
rect 18196 22176 18202 22228
rect 18414 22176 18420 22228
rect 18472 22216 18478 22228
rect 20622 22216 20628 22228
rect 18472 22188 20628 22216
rect 18472 22176 18478 22188
rect 20622 22176 20628 22188
rect 20680 22176 20686 22228
rect 23014 22176 23020 22228
rect 23072 22216 23078 22228
rect 23661 22219 23719 22225
rect 23661 22216 23673 22219
rect 23072 22188 23673 22216
rect 23072 22176 23078 22188
rect 23661 22185 23673 22188
rect 23707 22185 23719 22219
rect 23661 22179 23719 22185
rect 25038 22176 25044 22228
rect 25096 22216 25102 22228
rect 28442 22216 28448 22228
rect 25096 22188 25176 22216
rect 25096 22176 25102 22188
rect 5350 22148 5356 22160
rect 4356 22120 5356 22148
rect 3145 22083 3203 22089
rect 3145 22049 3157 22083
rect 3191 22080 3203 22083
rect 3326 22080 3332 22092
rect 3191 22052 3332 22080
rect 3191 22049 3203 22052
rect 3145 22043 3203 22049
rect 3326 22040 3332 22052
rect 3384 22040 3390 22092
rect 4356 22089 4384 22120
rect 5350 22108 5356 22120
rect 5408 22108 5414 22160
rect 9490 22108 9496 22160
rect 9548 22108 9554 22160
rect 9858 22108 9864 22160
rect 9916 22148 9922 22160
rect 9916 22120 10548 22148
rect 9916 22108 9922 22120
rect 10520 22092 10548 22120
rect 11882 22108 11888 22160
rect 11940 22148 11946 22160
rect 14918 22148 14924 22160
rect 11940 22120 14924 22148
rect 11940 22108 11946 22120
rect 14918 22108 14924 22120
rect 14976 22108 14982 22160
rect 15746 22148 15752 22160
rect 15304 22120 15752 22148
rect 4341 22083 4399 22089
rect 3436 22052 4200 22080
rect 2869 22015 2927 22021
rect 2869 21981 2881 22015
rect 2915 22012 2927 22015
rect 3436 22012 3464 22052
rect 4172 22021 4200 22052
rect 4341 22049 4353 22083
rect 4387 22080 4399 22083
rect 5166 22080 5172 22092
rect 4387 22052 4421 22080
rect 4540 22052 5172 22080
rect 4387 22049 4399 22052
rect 4341 22043 4399 22049
rect 2915 21984 3464 22012
rect 3513 22015 3571 22021
rect 2915 21981 2927 21984
rect 2869 21975 2927 21981
rect 3513 21981 3525 22015
rect 3559 21981 3571 22015
rect 3513 21975 3571 21981
rect 4157 22015 4215 22021
rect 4157 21981 4169 22015
rect 4203 22012 4215 22015
rect 4540 22012 4568 22052
rect 5166 22040 5172 22052
rect 5224 22040 5230 22092
rect 9306 22080 9312 22092
rect 8956 22052 9312 22080
rect 4203 21984 4568 22012
rect 4985 22015 5043 22021
rect 4203 21981 4215 21984
rect 4157 21975 4215 21981
rect 4985 21981 4997 22015
rect 5031 22012 5043 22015
rect 5258 22012 5264 22024
rect 5031 21984 5264 22012
rect 5031 21981 5043 21984
rect 4985 21975 5043 21981
rect 2961 21947 3019 21953
rect 2961 21913 2973 21947
rect 3007 21944 3019 21947
rect 3142 21944 3148 21956
rect 3007 21916 3148 21944
rect 3007 21913 3019 21916
rect 2961 21907 3019 21913
rect 3142 21904 3148 21916
rect 3200 21904 3206 21956
rect 2498 21836 2504 21888
rect 2556 21836 2562 21888
rect 3050 21836 3056 21888
rect 3108 21876 3114 21888
rect 3329 21879 3387 21885
rect 3329 21876 3341 21879
rect 3108 21848 3341 21876
rect 3108 21836 3114 21848
rect 3329 21845 3341 21848
rect 3375 21845 3387 21879
rect 3528 21876 3556 21975
rect 5258 21972 5264 21984
rect 5316 21972 5322 22024
rect 5442 21972 5448 22024
rect 5500 22012 5506 22024
rect 5721 22015 5779 22021
rect 5721 22012 5733 22015
rect 5500 21984 5733 22012
rect 5500 21972 5506 21984
rect 5721 21981 5733 21984
rect 5767 21981 5779 22015
rect 5721 21975 5779 21981
rect 3789 21879 3847 21885
rect 3789 21876 3801 21879
rect 3528 21848 3801 21876
rect 3329 21839 3387 21845
rect 3789 21845 3801 21848
rect 3835 21845 3847 21879
rect 3789 21839 3847 21845
rect 4249 21879 4307 21885
rect 4249 21845 4261 21879
rect 4295 21876 4307 21879
rect 4522 21876 4528 21888
rect 4295 21848 4528 21876
rect 4295 21845 4307 21848
rect 4249 21839 4307 21845
rect 4522 21836 4528 21848
rect 4580 21836 4586 21888
rect 4614 21836 4620 21888
rect 4672 21876 4678 21888
rect 4801 21879 4859 21885
rect 4801 21876 4813 21879
rect 4672 21848 4813 21876
rect 4672 21836 4678 21848
rect 4801 21845 4813 21848
rect 4847 21845 4859 21879
rect 5736 21876 5764 21975
rect 7098 21972 7104 22024
rect 7156 21972 7162 22024
rect 8956 22021 8984 22052
rect 9306 22040 9312 22052
rect 9364 22080 9370 22092
rect 9364 22052 10088 22080
rect 9364 22040 9370 22052
rect 8389 22015 8447 22021
rect 8389 21981 8401 22015
rect 8435 21981 8447 22015
rect 8389 21975 8447 21981
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 21981 8631 22015
rect 8573 21975 8631 21981
rect 8757 22015 8815 22021
rect 8757 21981 8769 22015
rect 8803 22012 8815 22015
rect 8941 22015 8999 22021
rect 8941 22012 8953 22015
rect 8803 21984 8953 22012
rect 8803 21981 8815 21984
rect 8757 21975 8815 21981
rect 8941 21981 8953 21984
rect 8987 21981 8999 22015
rect 8941 21975 8999 21981
rect 5994 21904 6000 21956
rect 6052 21904 6058 21956
rect 7742 21904 7748 21956
rect 7800 21944 7806 21956
rect 8404 21944 8432 21975
rect 7800 21916 8432 21944
rect 8588 21944 8616 21975
rect 9030 21972 9036 22024
rect 9088 22012 9094 22024
rect 9125 22015 9183 22021
rect 9125 22012 9137 22015
rect 9088 21984 9137 22012
rect 9088 21972 9094 21984
rect 9125 21981 9137 21984
rect 9171 21981 9183 22015
rect 9125 21975 9183 21981
rect 9217 22015 9275 22021
rect 9217 21981 9229 22015
rect 9263 22012 9275 22015
rect 9263 21984 9444 22012
rect 9263 21981 9275 21984
rect 9217 21975 9275 21981
rect 8846 21944 8852 21956
rect 8588 21916 8852 21944
rect 7800 21904 7806 21916
rect 8846 21904 8852 21916
rect 8904 21904 8910 21956
rect 6178 21876 6184 21888
rect 5736 21848 6184 21876
rect 4801 21839 4859 21845
rect 6178 21836 6184 21848
rect 6236 21836 6242 21888
rect 9125 21879 9183 21885
rect 9125 21845 9137 21879
rect 9171 21876 9183 21879
rect 9214 21876 9220 21888
rect 9171 21848 9220 21876
rect 9171 21845 9183 21848
rect 9125 21839 9183 21845
rect 9214 21836 9220 21848
rect 9272 21836 9278 21888
rect 9306 21836 9312 21888
rect 9364 21836 9370 21888
rect 9416 21876 9444 21984
rect 9766 21972 9772 22024
rect 9824 22012 9830 22024
rect 9953 22015 10011 22021
rect 9953 22012 9965 22015
rect 9824 21984 9965 22012
rect 9824 21972 9830 21984
rect 9953 21981 9965 21984
rect 9999 21981 10011 22015
rect 10060 22012 10088 22052
rect 10502 22040 10508 22092
rect 10560 22080 10566 22092
rect 10870 22080 10876 22092
rect 10560 22052 10876 22080
rect 10560 22040 10566 22052
rect 10870 22040 10876 22052
rect 10928 22040 10934 22092
rect 14369 22083 14427 22089
rect 14369 22049 14381 22083
rect 14415 22080 14427 22083
rect 15304 22080 15332 22120
rect 15746 22108 15752 22120
rect 15804 22148 15810 22160
rect 16206 22148 16212 22160
rect 15804 22120 16212 22148
rect 15804 22108 15810 22120
rect 16206 22108 16212 22120
rect 16264 22108 16270 22160
rect 16776 22148 16804 22176
rect 17681 22151 17739 22157
rect 17681 22148 17693 22151
rect 16776 22120 17693 22148
rect 17681 22117 17693 22120
rect 17727 22148 17739 22151
rect 17727 22120 18644 22148
rect 17727 22117 17739 22120
rect 17681 22111 17739 22117
rect 14415 22052 15332 22080
rect 14415 22049 14427 22052
rect 14369 22043 14427 22049
rect 16022 22040 16028 22092
rect 16080 22040 16086 22092
rect 17034 22040 17040 22092
rect 17092 22040 17098 22092
rect 17310 22040 17316 22092
rect 17368 22080 17374 22092
rect 17589 22083 17647 22089
rect 17589 22080 17601 22083
rect 17368 22052 17601 22080
rect 17368 22040 17374 22052
rect 17589 22049 17601 22052
rect 17635 22049 17647 22083
rect 18233 22083 18291 22089
rect 18233 22080 18245 22083
rect 17589 22043 17647 22049
rect 17788 22052 18245 22080
rect 10229 22015 10287 22021
rect 10229 22012 10241 22015
rect 10060 21984 10241 22012
rect 9953 21975 10011 21981
rect 10229 21981 10241 21984
rect 10275 21981 10287 22015
rect 12345 22015 12403 22021
rect 12345 22012 12357 22015
rect 10229 21975 10287 21981
rect 12268 21984 12357 22012
rect 12268 21956 12296 21984
rect 12345 21981 12357 21984
rect 12391 22012 12403 22015
rect 12805 22015 12863 22021
rect 12805 22012 12817 22015
rect 12391 21984 12817 22012
rect 12391 21981 12403 21984
rect 12345 21975 12403 21981
rect 12805 21981 12817 21984
rect 12851 21981 12863 22015
rect 12805 21975 12863 21981
rect 13541 22015 13599 22021
rect 13541 21981 13553 22015
rect 13587 22012 13599 22015
rect 14277 22015 14335 22021
rect 13587 21984 13860 22012
rect 13587 21981 13599 21984
rect 13541 21975 13599 21981
rect 9493 21947 9551 21953
rect 9493 21913 9505 21947
rect 9539 21944 9551 21947
rect 9858 21944 9864 21956
rect 9539 21916 9864 21944
rect 9539 21913 9551 21916
rect 9493 21907 9551 21913
rect 9858 21904 9864 21916
rect 9916 21904 9922 21956
rect 10962 21904 10968 21956
rect 11020 21944 11026 21956
rect 11885 21947 11943 21953
rect 11885 21944 11897 21947
rect 11020 21916 11897 21944
rect 11020 21904 11026 21916
rect 11885 21913 11897 21916
rect 11931 21913 11943 21947
rect 11885 21907 11943 21913
rect 11974 21904 11980 21956
rect 12032 21904 12038 21956
rect 12250 21904 12256 21956
rect 12308 21904 12314 21956
rect 12434 21904 12440 21956
rect 12492 21904 12498 21956
rect 13725 21947 13783 21953
rect 13725 21913 13737 21947
rect 13771 21913 13783 21947
rect 13832 21944 13860 21984
rect 14277 21981 14289 22015
rect 14323 22012 14335 22015
rect 15841 22015 15899 22021
rect 14323 21984 14872 22012
rect 14323 21981 14335 21984
rect 14277 21975 14335 21981
rect 14366 21944 14372 21956
rect 13832 21916 14372 21944
rect 13725 21907 13783 21913
rect 9677 21879 9735 21885
rect 9677 21876 9689 21879
rect 9416 21848 9689 21876
rect 9677 21845 9689 21848
rect 9723 21845 9735 21879
rect 9677 21839 9735 21845
rect 9766 21836 9772 21888
rect 9824 21876 9830 21888
rect 10042 21876 10048 21888
rect 9824 21848 10048 21876
rect 9824 21836 9830 21848
rect 10042 21836 10048 21848
rect 10100 21876 10106 21888
rect 12894 21876 12900 21888
rect 10100 21848 12900 21876
rect 10100 21836 10106 21848
rect 12894 21836 12900 21848
rect 12952 21836 12958 21888
rect 13538 21836 13544 21888
rect 13596 21876 13602 21888
rect 13740 21876 13768 21907
rect 14366 21904 14372 21916
rect 14424 21904 14430 21956
rect 14844 21888 14872 21984
rect 15841 21981 15853 22015
rect 15887 22012 15899 22015
rect 16040 22012 16068 22040
rect 15887 21984 16068 22012
rect 17052 22012 17080 22040
rect 17405 22015 17463 22021
rect 17405 22012 17417 22015
rect 17052 21984 17417 22012
rect 15887 21981 15899 21984
rect 15841 21975 15899 21981
rect 17405 21981 17417 21984
rect 17451 21981 17463 22015
rect 17405 21975 17463 21981
rect 17494 21972 17500 22024
rect 17552 22012 17558 22024
rect 17788 22012 17816 22052
rect 18233 22049 18245 22052
rect 18279 22049 18291 22083
rect 18233 22043 18291 22049
rect 17552 21984 17816 22012
rect 17552 21972 17558 21984
rect 17862 21972 17868 22024
rect 17920 21972 17926 22024
rect 18046 21972 18052 22024
rect 18104 22012 18110 22024
rect 18616 22021 18644 22120
rect 19702 22108 19708 22160
rect 19760 22148 19766 22160
rect 20070 22148 20076 22160
rect 19760 22120 20076 22148
rect 19760 22108 19766 22120
rect 20070 22108 20076 22120
rect 20128 22108 20134 22160
rect 22186 22108 22192 22160
rect 22244 22148 22250 22160
rect 23290 22148 23296 22160
rect 22244 22120 23296 22148
rect 22244 22108 22250 22120
rect 23290 22108 23296 22120
rect 23348 22108 23354 22160
rect 20533 22083 20591 22089
rect 20533 22049 20545 22083
rect 20579 22080 20591 22083
rect 20990 22080 20996 22092
rect 20579 22052 20996 22080
rect 20579 22049 20591 22052
rect 20533 22043 20591 22049
rect 20990 22040 20996 22052
rect 21048 22040 21054 22092
rect 22002 22040 22008 22092
rect 22060 22080 22066 22092
rect 22060 22052 23060 22080
rect 22060 22040 22066 22052
rect 18141 22015 18199 22021
rect 18141 22012 18153 22015
rect 18104 21984 18153 22012
rect 18104 21972 18110 21984
rect 18141 21981 18153 21984
rect 18187 21981 18199 22015
rect 18141 21975 18199 21981
rect 18601 22015 18659 22021
rect 18601 21981 18613 22015
rect 18647 21981 18659 22015
rect 18601 21975 18659 21981
rect 20625 22015 20683 22021
rect 20625 21981 20637 22015
rect 20671 22012 20683 22015
rect 20898 22012 20904 22024
rect 20671 21984 20904 22012
rect 20671 21981 20683 21984
rect 20625 21975 20683 21981
rect 20898 21972 20904 21984
rect 20956 21972 20962 22024
rect 22094 21972 22100 22024
rect 22152 21972 22158 22024
rect 22186 21972 22192 22024
rect 22244 22012 22250 22024
rect 23032 22021 23060 22052
rect 23382 22040 23388 22092
rect 23440 22040 23446 22092
rect 25148 22089 25176 22188
rect 25976 22188 28448 22216
rect 25976 22157 26004 22188
rect 28442 22176 28448 22188
rect 28500 22176 28506 22228
rect 28534 22176 28540 22228
rect 28592 22216 28598 22228
rect 28592 22188 31754 22216
rect 28592 22176 28598 22188
rect 25961 22151 26019 22157
rect 25961 22117 25973 22151
rect 26007 22117 26019 22151
rect 25961 22111 26019 22117
rect 26786 22108 26792 22160
rect 26844 22148 26850 22160
rect 27341 22151 27399 22157
rect 27341 22148 27353 22151
rect 26844 22120 27353 22148
rect 26844 22108 26850 22120
rect 27341 22117 27353 22120
rect 27387 22148 27399 22151
rect 28994 22148 29000 22160
rect 27387 22120 29000 22148
rect 27387 22117 27399 22120
rect 27341 22111 27399 22117
rect 28994 22108 29000 22120
rect 29052 22108 29058 22160
rect 29730 22148 29736 22160
rect 29656 22120 29736 22148
rect 29656 22094 29684 22120
rect 29730 22108 29736 22120
rect 29788 22108 29794 22160
rect 30098 22108 30104 22160
rect 30156 22108 30162 22160
rect 31726 22148 31754 22188
rect 32122 22176 32128 22228
rect 32180 22216 32186 22228
rect 32309 22219 32367 22225
rect 32309 22216 32321 22219
rect 32180 22188 32321 22216
rect 32180 22176 32186 22188
rect 32309 22185 32321 22188
rect 32355 22185 32367 22219
rect 32309 22179 32367 22185
rect 32674 22176 32680 22228
rect 32732 22176 32738 22228
rect 33502 22176 33508 22228
rect 33560 22176 33566 22228
rect 35250 22176 35256 22228
rect 35308 22176 35314 22228
rect 35437 22219 35495 22225
rect 35437 22185 35449 22219
rect 35483 22216 35495 22219
rect 35526 22216 35532 22228
rect 35483 22188 35532 22216
rect 35483 22185 35495 22188
rect 35437 22179 35495 22185
rect 35526 22176 35532 22188
rect 35584 22176 35590 22228
rect 35894 22176 35900 22228
rect 35952 22176 35958 22228
rect 32692 22148 32720 22176
rect 31726 22120 32720 22148
rect 25133 22083 25191 22089
rect 25133 22049 25145 22083
rect 25179 22080 25191 22083
rect 26881 22083 26939 22089
rect 25179 22052 26832 22080
rect 25179 22049 25191 22052
rect 25133 22043 25191 22049
rect 22281 22015 22339 22021
rect 22281 22012 22293 22015
rect 22244 21984 22293 22012
rect 22244 21972 22250 21984
rect 22281 21981 22293 21984
rect 22327 21981 22339 22015
rect 22281 21975 22339 21981
rect 22833 22015 22891 22021
rect 22833 21981 22845 22015
rect 22879 21981 22891 22015
rect 22833 21975 22891 21981
rect 23017 22015 23075 22021
rect 23017 21981 23029 22015
rect 23063 21981 23075 22015
rect 23017 21975 23075 21981
rect 23124 21984 23704 22012
rect 15378 21904 15384 21956
rect 15436 21944 15442 21956
rect 15565 21947 15623 21953
rect 15565 21944 15577 21947
rect 15436 21916 15577 21944
rect 15436 21904 15442 21916
rect 15565 21913 15577 21916
rect 15611 21913 15623 21947
rect 15565 21907 15623 21913
rect 16025 21947 16083 21953
rect 16025 21913 16037 21947
rect 16071 21944 16083 21947
rect 17034 21944 17040 21956
rect 16071 21916 17040 21944
rect 16071 21913 16083 21916
rect 16025 21907 16083 21913
rect 17034 21904 17040 21916
rect 17092 21904 17098 21956
rect 17678 21904 17684 21956
rect 17736 21944 17742 21956
rect 22370 21944 22376 21956
rect 17736 21916 22376 21944
rect 17736 21904 17742 21916
rect 22370 21904 22376 21916
rect 22428 21944 22434 21956
rect 22848 21944 22876 21975
rect 23124 21944 23152 21984
rect 22428 21916 23152 21944
rect 23477 21947 23535 21953
rect 22428 21904 22434 21916
rect 23477 21913 23489 21947
rect 23523 21944 23535 21947
rect 23566 21944 23572 21956
rect 23523 21916 23572 21944
rect 23523 21913 23535 21916
rect 23477 21907 23535 21913
rect 23566 21904 23572 21916
rect 23624 21904 23630 21956
rect 23676 21953 23704 21984
rect 24118 21972 24124 22024
rect 24176 21972 24182 22024
rect 24578 21972 24584 22024
rect 24636 21972 24642 22024
rect 25317 22015 25375 22021
rect 25317 22012 25329 22015
rect 24688 21984 25329 22012
rect 23676 21947 23735 21953
rect 23676 21916 23689 21947
rect 23677 21913 23689 21916
rect 23723 21913 23735 21947
rect 24136 21944 24164 21972
rect 24688 21944 24716 21984
rect 25317 21981 25329 21984
rect 25363 21981 25375 22015
rect 25317 21975 25375 21981
rect 25774 21972 25780 22024
rect 25832 22012 25838 22024
rect 26234 22012 26240 22024
rect 25832 21984 26240 22012
rect 25832 21972 25838 21984
rect 26234 21972 26240 21984
rect 26292 22012 26298 22024
rect 26513 22015 26571 22021
rect 26513 22012 26525 22015
rect 26292 21984 26525 22012
rect 26292 21972 26298 21984
rect 26513 21981 26525 21984
rect 26559 21981 26571 22015
rect 26513 21975 26571 21981
rect 26697 22015 26755 22021
rect 26697 21981 26709 22015
rect 26743 21981 26755 22015
rect 26697 21975 26755 21981
rect 26712 21944 26740 21975
rect 24136 21916 24716 21944
rect 25792 21916 26740 21944
rect 26804 21944 26832 22052
rect 26881 22049 26893 22083
rect 26927 22080 26939 22083
rect 27709 22083 27767 22089
rect 27709 22080 27721 22083
rect 26927 22052 27721 22080
rect 26927 22049 26939 22052
rect 26881 22043 26939 22049
rect 27709 22049 27721 22052
rect 27755 22080 27767 22083
rect 27755 22052 28304 22080
rect 27755 22049 27767 22052
rect 27709 22043 27767 22049
rect 28276 22024 28304 22052
rect 28534 22040 28540 22092
rect 28592 22080 28598 22092
rect 28813 22083 28871 22089
rect 28813 22080 28825 22083
rect 28592 22052 28825 22080
rect 28592 22040 28598 22052
rect 28813 22049 28825 22052
rect 28859 22049 28871 22083
rect 28813 22043 28871 22049
rect 28902 22040 28908 22092
rect 28960 22080 28966 22092
rect 28960 22052 29408 22080
rect 28960 22040 28966 22052
rect 27246 21972 27252 22024
rect 27304 22012 27310 22024
rect 27525 22015 27583 22021
rect 27525 22012 27537 22015
rect 27304 21984 27537 22012
rect 27304 21972 27310 21984
rect 27525 21981 27537 21984
rect 27571 21981 27583 22015
rect 27525 21975 27583 21981
rect 27801 22015 27859 22021
rect 27801 21981 27813 22015
rect 27847 22012 27859 22015
rect 28077 22015 28135 22021
rect 28077 22012 28089 22015
rect 27847 21984 28089 22012
rect 27847 21981 27859 21984
rect 27801 21975 27859 21981
rect 28077 21981 28089 21984
rect 28123 21981 28135 22015
rect 28077 21975 28135 21981
rect 27816 21944 27844 21975
rect 26804 21916 27844 21944
rect 28092 21944 28120 21975
rect 28258 21972 28264 22024
rect 28316 21972 28322 22024
rect 28721 22015 28779 22021
rect 28721 21981 28733 22015
rect 28767 22012 28779 22015
rect 29270 22012 29276 22024
rect 28767 21984 29276 22012
rect 28767 21981 28779 21984
rect 28721 21975 28779 21981
rect 29270 21972 29276 21984
rect 29328 21972 29334 22024
rect 29380 21944 29408 22052
rect 29564 22066 29684 22094
rect 31662 22080 31668 22092
rect 29564 22021 29592 22066
rect 30024 22052 31668 22080
rect 29549 22015 29607 22021
rect 29549 21981 29561 22015
rect 29595 21981 29607 22015
rect 29549 21975 29607 21981
rect 29914 21972 29920 22024
rect 29972 21972 29978 22024
rect 29733 21947 29791 21953
rect 29733 21944 29745 21947
rect 28092 21916 28994 21944
rect 29380 21916 29745 21944
rect 23677 21907 23735 21913
rect 25792 21888 25820 21916
rect 13596 21848 13768 21876
rect 13596 21836 13602 21848
rect 14826 21836 14832 21888
rect 14884 21836 14890 21888
rect 15102 21836 15108 21888
rect 15160 21876 15166 21888
rect 15657 21879 15715 21885
rect 15657 21876 15669 21879
rect 15160 21848 15669 21876
rect 15160 21836 15166 21848
rect 15657 21845 15669 21848
rect 15703 21845 15715 21879
rect 15657 21839 15715 21845
rect 17770 21836 17776 21888
rect 17828 21876 17834 21888
rect 17957 21879 18015 21885
rect 17957 21876 17969 21879
rect 17828 21848 17969 21876
rect 17828 21836 17834 21848
rect 17957 21845 17969 21848
rect 18003 21845 18015 21879
rect 17957 21839 18015 21845
rect 20346 21836 20352 21888
rect 20404 21876 20410 21888
rect 20717 21879 20775 21885
rect 20717 21876 20729 21879
rect 20404 21848 20729 21876
rect 20404 21836 20410 21848
rect 20717 21845 20729 21848
rect 20763 21845 20775 21879
rect 20717 21839 20775 21845
rect 21082 21836 21088 21888
rect 21140 21836 21146 21888
rect 23845 21879 23903 21885
rect 23845 21845 23857 21879
rect 23891 21876 23903 21879
rect 25774 21876 25780 21888
rect 23891 21848 25780 21876
rect 23891 21845 23903 21848
rect 23845 21839 23903 21845
rect 25774 21836 25780 21848
rect 25832 21836 25838 21888
rect 27522 21836 27528 21888
rect 27580 21876 27586 21888
rect 27706 21876 27712 21888
rect 27580 21848 27712 21876
rect 27580 21836 27586 21848
rect 27706 21836 27712 21848
rect 27764 21836 27770 21888
rect 28966 21876 28994 21916
rect 29733 21913 29745 21916
rect 29779 21913 29791 21947
rect 29733 21907 29791 21913
rect 29822 21904 29828 21956
rect 29880 21904 29886 21956
rect 30024 21876 30052 22052
rect 31662 22040 31668 22052
rect 31720 22040 31726 22092
rect 32030 21972 32036 22024
rect 32088 21972 32094 22024
rect 32692 22021 32720 22120
rect 33873 22151 33931 22157
rect 33873 22117 33885 22151
rect 33919 22148 33931 22151
rect 35268 22148 35296 22176
rect 35710 22148 35716 22160
rect 33919 22120 34560 22148
rect 35268 22120 35716 22148
rect 33919 22117 33931 22120
rect 33873 22111 33931 22117
rect 33321 22083 33379 22089
rect 33321 22049 33333 22083
rect 33367 22080 33379 22083
rect 33781 22083 33839 22089
rect 33781 22080 33793 22083
rect 33367 22052 33793 22080
rect 33367 22049 33379 22052
rect 33321 22043 33379 22049
rect 33781 22049 33793 22052
rect 33827 22049 33839 22083
rect 33781 22043 33839 22049
rect 32125 22015 32183 22021
rect 32125 21981 32137 22015
rect 32171 22012 32183 22015
rect 32677 22015 32735 22021
rect 32171 21984 32536 22012
rect 32171 21981 32183 21984
rect 32125 21975 32183 21981
rect 31294 21944 31300 21956
rect 30116 21916 31300 21944
rect 30116 21888 30144 21916
rect 31294 21904 31300 21916
rect 31352 21944 31358 21956
rect 31665 21947 31723 21953
rect 31665 21944 31677 21947
rect 31352 21916 31677 21944
rect 31352 21904 31358 21916
rect 31665 21913 31677 21916
rect 31711 21913 31723 21947
rect 31665 21907 31723 21913
rect 31757 21947 31815 21953
rect 31757 21913 31769 21947
rect 31803 21944 31815 21947
rect 32398 21944 32404 21956
rect 31803 21916 32404 21944
rect 31803 21913 31815 21916
rect 31757 21907 31815 21913
rect 32398 21904 32404 21916
rect 32456 21904 32462 21956
rect 32508 21888 32536 21984
rect 32677 21981 32689 22015
rect 32723 21981 32735 22015
rect 32677 21975 32735 21981
rect 32861 22015 32919 22021
rect 32861 21981 32873 22015
rect 32907 21981 32919 22015
rect 32861 21975 32919 21981
rect 32876 21944 32904 21975
rect 32950 21972 32956 22024
rect 33008 22012 33014 22024
rect 33137 22015 33195 22021
rect 33137 22012 33149 22015
rect 33008 21984 33149 22012
rect 33008 21972 33014 21984
rect 33137 21981 33149 21984
rect 33183 21981 33195 22015
rect 33137 21975 33195 21981
rect 33413 22015 33471 22021
rect 33413 21981 33425 22015
rect 33459 22012 33471 22015
rect 33502 22012 33508 22024
rect 33459 21984 33508 22012
rect 33459 21981 33471 21984
rect 33413 21975 33471 21981
rect 33502 21972 33508 21984
rect 33560 21972 33566 22024
rect 33686 21972 33692 22024
rect 33744 21972 33750 22024
rect 34054 21972 34060 22024
rect 34112 21972 34118 22024
rect 34422 21972 34428 22024
rect 34480 21972 34486 22024
rect 34532 22012 34560 22120
rect 35710 22108 35716 22120
rect 35768 22108 35774 22160
rect 34606 22040 34612 22092
rect 34664 22080 34670 22092
rect 34664 22052 34928 22080
rect 34664 22040 34670 22052
rect 34900 22021 34928 22052
rect 34992 22052 35572 22080
rect 34793 22015 34851 22021
rect 34793 22012 34805 22015
rect 34532 21984 34805 22012
rect 34793 21981 34805 21984
rect 34839 21981 34851 22015
rect 34793 21975 34851 21981
rect 34886 22015 34944 22021
rect 34886 21981 34898 22015
rect 34932 21981 34944 22015
rect 34886 21975 34944 21981
rect 34072 21944 34100 21972
rect 32876 21916 34100 21944
rect 34440 21944 34468 21972
rect 34992 21944 35020 22052
rect 35158 21972 35164 22024
rect 35216 21972 35222 22024
rect 35268 22021 35296 22052
rect 35544 22021 35572 22052
rect 35258 22015 35316 22021
rect 35258 21981 35270 22015
rect 35304 21981 35316 22015
rect 35258 21975 35316 21981
rect 35529 22015 35587 22021
rect 35529 21981 35541 22015
rect 35575 21981 35587 22015
rect 35529 21975 35587 21981
rect 34440 21916 35020 21944
rect 35069 21947 35127 21953
rect 35069 21913 35081 21947
rect 35115 21913 35127 21947
rect 35069 21907 35127 21913
rect 35713 21947 35771 21953
rect 35713 21913 35725 21947
rect 35759 21913 35771 21947
rect 35713 21907 35771 21913
rect 28966 21848 30052 21876
rect 30098 21836 30104 21888
rect 30156 21836 30162 21888
rect 32490 21836 32496 21888
rect 32548 21876 32554 21888
rect 34698 21876 34704 21888
rect 32548 21848 34704 21876
rect 32548 21836 32554 21848
rect 34698 21836 34704 21848
rect 34756 21836 34762 21888
rect 34790 21836 34796 21888
rect 34848 21876 34854 21888
rect 35084 21876 35112 21907
rect 34848 21848 35112 21876
rect 34848 21836 34854 21848
rect 35158 21836 35164 21888
rect 35216 21876 35222 21888
rect 35728 21876 35756 21907
rect 35216 21848 35756 21876
rect 35216 21836 35222 21848
rect 1104 21786 38272 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 38272 21786
rect 1104 21712 38272 21734
rect 2498 21632 2504 21684
rect 2556 21632 2562 21684
rect 5169 21675 5227 21681
rect 5169 21641 5181 21675
rect 5215 21672 5227 21675
rect 5258 21672 5264 21684
rect 5215 21644 5264 21672
rect 5215 21641 5227 21644
rect 5169 21635 5227 21641
rect 5258 21632 5264 21644
rect 5316 21632 5322 21684
rect 5994 21632 6000 21684
rect 6052 21672 6058 21684
rect 6365 21675 6423 21681
rect 6365 21672 6377 21675
rect 6052 21644 6377 21672
rect 6052 21632 6058 21644
rect 6365 21641 6377 21644
rect 6411 21641 6423 21675
rect 6365 21635 6423 21641
rect 9125 21675 9183 21681
rect 9125 21641 9137 21675
rect 9171 21672 9183 21675
rect 9306 21672 9312 21684
rect 9171 21644 9312 21672
rect 9171 21641 9183 21644
rect 9125 21635 9183 21641
rect 9306 21632 9312 21644
rect 9364 21632 9370 21684
rect 9493 21675 9551 21681
rect 9493 21641 9505 21675
rect 9539 21672 9551 21675
rect 10686 21672 10692 21684
rect 9539 21644 10692 21672
rect 9539 21641 9551 21644
rect 9493 21635 9551 21641
rect 10686 21632 10692 21644
rect 10744 21632 10750 21684
rect 11514 21672 11520 21684
rect 10796 21644 11520 21672
rect 1762 21496 1768 21548
rect 1820 21496 1826 21548
rect 2133 21539 2191 21545
rect 2133 21505 2145 21539
rect 2179 21536 2191 21539
rect 2516 21536 2544 21632
rect 3050 21564 3056 21616
rect 3108 21564 3114 21616
rect 3786 21564 3792 21616
rect 3844 21564 3850 21616
rect 4522 21564 4528 21616
rect 4580 21604 4586 21616
rect 4801 21607 4859 21613
rect 4801 21604 4813 21607
rect 4580 21576 4813 21604
rect 4580 21564 4586 21576
rect 4801 21573 4813 21576
rect 4847 21604 4859 21607
rect 4847 21576 8984 21604
rect 4847 21573 4859 21576
rect 4801 21567 4859 21573
rect 2179 21508 2544 21536
rect 2179 21505 2191 21508
rect 2133 21499 2191 21505
rect 2774 21496 2780 21548
rect 2832 21496 2838 21548
rect 5534 21496 5540 21548
rect 5592 21496 5598 21548
rect 5629 21539 5687 21545
rect 5629 21505 5641 21539
rect 5675 21536 5687 21539
rect 6086 21536 6092 21548
rect 5675 21508 6092 21536
rect 5675 21505 5687 21508
rect 5629 21499 5687 21505
rect 6086 21496 6092 21508
rect 6144 21496 6150 21548
rect 6546 21496 6552 21548
rect 6604 21496 6610 21548
rect 8956 21545 8984 21576
rect 9214 21564 9220 21616
rect 9272 21604 9278 21616
rect 10796 21604 10824 21644
rect 11514 21632 11520 21644
rect 11572 21632 11578 21684
rect 14826 21672 14832 21684
rect 13464 21644 14688 21672
rect 13464 21616 13492 21644
rect 9272 21576 9720 21604
rect 9272 21564 9278 21576
rect 8573 21539 8631 21545
rect 8573 21536 8585 21539
rect 8220 21508 8585 21536
rect 5813 21471 5871 21477
rect 5813 21437 5825 21471
rect 5859 21468 5871 21471
rect 8110 21468 8116 21480
rect 5859 21440 8116 21468
rect 5859 21437 5871 21440
rect 5813 21431 5871 21437
rect 8110 21428 8116 21440
rect 8168 21428 8174 21480
rect 8220 21412 8248 21508
rect 8573 21505 8585 21508
rect 8619 21505 8631 21539
rect 8573 21499 8631 21505
rect 8665 21539 8723 21545
rect 8665 21505 8677 21539
rect 8711 21505 8723 21539
rect 8665 21499 8723 21505
rect 8849 21539 8907 21545
rect 8849 21505 8861 21539
rect 8895 21505 8907 21539
rect 8849 21499 8907 21505
rect 8941 21539 8999 21545
rect 8941 21505 8953 21539
rect 8987 21536 8999 21539
rect 8987 21508 9076 21536
rect 8987 21505 8999 21508
rect 8941 21499 8999 21505
rect 8680 21468 8708 21499
rect 8496 21440 8708 21468
rect 8496 21412 8524 21440
rect 8202 21360 8208 21412
rect 8260 21360 8266 21412
rect 8478 21360 8484 21412
rect 8536 21360 8542 21412
rect 8570 21360 8576 21412
rect 8628 21400 8634 21412
rect 8864 21400 8892 21499
rect 9048 21412 9076 21508
rect 9490 21496 9496 21548
rect 9548 21496 9554 21548
rect 9692 21545 9720 21576
rect 9876 21576 10824 21604
rect 9876 21545 9904 21576
rect 10962 21564 10968 21616
rect 11020 21604 11026 21616
rect 11698 21604 11704 21616
rect 11020 21576 11192 21604
rect 11020 21564 11026 21576
rect 9677 21539 9735 21545
rect 9677 21505 9689 21539
rect 9723 21505 9735 21539
rect 9677 21499 9735 21505
rect 9861 21539 9919 21545
rect 9861 21505 9873 21539
rect 9907 21505 9919 21539
rect 9861 21499 9919 21505
rect 10686 21496 10692 21548
rect 10744 21496 10750 21548
rect 11164 21545 11192 21576
rect 11348 21576 11704 21604
rect 11348 21545 11376 21576
rect 11698 21564 11704 21576
rect 11756 21564 11762 21616
rect 13446 21564 13452 21616
rect 13504 21564 13510 21616
rect 13722 21564 13728 21616
rect 13780 21604 13786 21616
rect 14660 21613 14688 21644
rect 14752 21644 14832 21672
rect 14752 21613 14780 21644
rect 14826 21632 14832 21644
rect 14884 21632 14890 21684
rect 15013 21675 15071 21681
rect 15013 21641 15025 21675
rect 15059 21641 15071 21675
rect 15013 21635 15071 21641
rect 14645 21607 14703 21613
rect 13780 21576 14228 21604
rect 13780 21564 13786 21576
rect 14200 21548 14228 21576
rect 14645 21573 14657 21607
rect 14691 21573 14703 21607
rect 14645 21567 14703 21573
rect 14737 21607 14795 21613
rect 14737 21573 14749 21607
rect 14783 21573 14795 21607
rect 15028 21604 15056 21635
rect 16022 21632 16028 21684
rect 16080 21672 16086 21684
rect 16080 21644 16988 21672
rect 16080 21632 16086 21644
rect 16960 21604 16988 21644
rect 17310 21632 17316 21684
rect 17368 21632 17374 21684
rect 17494 21632 17500 21684
rect 17552 21672 17558 21684
rect 17681 21675 17739 21681
rect 17681 21672 17693 21675
rect 17552 21644 17693 21672
rect 17552 21632 17558 21644
rect 17681 21641 17693 21644
rect 17727 21641 17739 21675
rect 17681 21635 17739 21641
rect 18230 21632 18236 21684
rect 18288 21632 18294 21684
rect 20806 21672 20812 21684
rect 18340 21644 20812 21672
rect 17862 21604 17868 21616
rect 15028 21576 16160 21604
rect 14737 21567 14795 21573
rect 10873 21539 10931 21545
rect 10873 21505 10885 21539
rect 10919 21505 10931 21539
rect 10873 21499 10931 21505
rect 11057 21539 11115 21545
rect 11057 21505 11069 21539
rect 11103 21505 11115 21539
rect 11057 21499 11115 21505
rect 11149 21539 11207 21545
rect 11149 21505 11161 21539
rect 11195 21505 11207 21539
rect 11149 21499 11207 21505
rect 11333 21539 11391 21545
rect 11333 21505 11345 21539
rect 11379 21505 11391 21539
rect 11333 21499 11391 21505
rect 8628 21372 8892 21400
rect 8628 21360 8634 21372
rect 9030 21360 9036 21412
rect 9088 21360 9094 21412
rect 9508 21400 9536 21496
rect 9766 21428 9772 21480
rect 9824 21428 9830 21480
rect 9950 21428 9956 21480
rect 10008 21468 10014 21480
rect 10318 21468 10324 21480
rect 10008 21440 10324 21468
rect 10008 21428 10014 21440
rect 10318 21428 10324 21440
rect 10376 21428 10382 21480
rect 10413 21471 10471 21477
rect 10413 21437 10425 21471
rect 10459 21437 10471 21471
rect 10888 21468 10916 21499
rect 10413 21431 10471 21437
rect 10704 21440 10916 21468
rect 10428 21400 10456 21431
rect 10704 21412 10732 21440
rect 9508 21372 10456 21400
rect 10686 21360 10692 21412
rect 10744 21360 10750 21412
rect 11072 21400 11100 21499
rect 11606 21496 11612 21548
rect 11664 21496 11670 21548
rect 11974 21496 11980 21548
rect 12032 21496 12038 21548
rect 12250 21496 12256 21548
rect 12308 21536 12314 21548
rect 12308 21508 13400 21536
rect 12308 21496 12314 21508
rect 13372 21468 13400 21508
rect 13630 21496 13636 21548
rect 13688 21496 13694 21548
rect 13814 21496 13820 21548
rect 13872 21496 13878 21548
rect 13909 21539 13967 21545
rect 13909 21505 13921 21539
rect 13955 21505 13967 21539
rect 13909 21499 13967 21505
rect 14001 21539 14059 21545
rect 14001 21505 14013 21539
rect 14047 21505 14059 21539
rect 14001 21499 14059 21505
rect 13924 21468 13952 21499
rect 13372 21440 13952 21468
rect 11974 21400 11980 21412
rect 11072 21372 11980 21400
rect 11974 21360 11980 21372
rect 12032 21400 12038 21412
rect 13814 21400 13820 21412
rect 12032 21372 13820 21400
rect 12032 21360 12038 21372
rect 13814 21360 13820 21372
rect 13872 21400 13878 21412
rect 14016 21400 14044 21499
rect 14182 21496 14188 21548
rect 14240 21536 14246 21548
rect 14918 21545 14924 21548
rect 14369 21539 14427 21545
rect 14369 21536 14381 21539
rect 14240 21508 14381 21536
rect 14240 21496 14246 21508
rect 14369 21505 14381 21508
rect 14415 21505 14427 21539
rect 14369 21499 14427 21505
rect 14462 21539 14520 21545
rect 14462 21505 14474 21539
rect 14508 21505 14520 21539
rect 14462 21499 14520 21505
rect 14875 21539 14924 21545
rect 14875 21505 14887 21539
rect 14921 21505 14924 21539
rect 14875 21499 14924 21505
rect 14277 21471 14335 21477
rect 14277 21437 14289 21471
rect 14323 21468 14335 21471
rect 14476 21468 14504 21499
rect 14918 21496 14924 21499
rect 14976 21496 14982 21548
rect 15286 21496 15292 21548
rect 15344 21536 15350 21548
rect 16132 21545 16160 21576
rect 16960 21576 17868 21604
rect 15749 21539 15807 21545
rect 16117 21539 16175 21545
rect 15749 21536 15761 21539
rect 15344 21508 15761 21536
rect 15344 21496 15350 21508
rect 15749 21505 15761 21508
rect 15795 21536 15807 21539
rect 15851 21536 15947 21539
rect 15795 21511 15947 21536
rect 15795 21508 15879 21511
rect 15795 21505 15807 21508
rect 15749 21499 15807 21505
rect 14323 21440 14504 21468
rect 15473 21471 15531 21477
rect 14323 21437 14335 21440
rect 14277 21431 14335 21437
rect 15473 21437 15485 21471
rect 15519 21437 15531 21471
rect 15919 21468 15947 21511
rect 16117 21505 16129 21539
rect 16163 21536 16175 21539
rect 16853 21539 16911 21545
rect 16853 21536 16865 21539
rect 16163 21508 16865 21536
rect 16163 21505 16175 21508
rect 16117 21499 16175 21505
rect 16853 21505 16865 21508
rect 16899 21505 16911 21539
rect 16960 21536 16988 21576
rect 17862 21564 17868 21576
rect 17920 21564 17926 21616
rect 18049 21607 18107 21613
rect 18049 21573 18061 21607
rect 18095 21604 18107 21607
rect 18248 21604 18276 21632
rect 18095 21576 18276 21604
rect 18095 21573 18107 21576
rect 18049 21567 18107 21573
rect 17129 21539 17187 21545
rect 17129 21536 17141 21539
rect 16960 21508 17141 21536
rect 16853 21499 16911 21505
rect 17129 21505 17141 21508
rect 17175 21505 17187 21539
rect 17129 21499 17187 21505
rect 17221 21539 17279 21545
rect 17221 21505 17233 21539
rect 17267 21536 17279 21539
rect 17405 21539 17463 21545
rect 17267 21508 17356 21536
rect 17267 21505 17279 21508
rect 17221 21499 17279 21505
rect 17328 21480 17356 21508
rect 17405 21505 17417 21539
rect 17451 21536 17463 21539
rect 17494 21536 17500 21548
rect 17451 21508 17500 21536
rect 17451 21505 17463 21508
rect 17405 21499 17463 21505
rect 17494 21496 17500 21508
rect 17552 21496 17558 21548
rect 18340 21545 18368 21644
rect 20806 21632 20812 21644
rect 20864 21632 20870 21684
rect 20916 21644 21037 21672
rect 20916 21604 20944 21644
rect 20364 21576 20944 21604
rect 20364 21548 20392 21576
rect 21009 21551 21037 21644
rect 21174 21632 21180 21684
rect 21232 21672 21238 21684
rect 23198 21672 23204 21684
rect 21232 21644 23204 21672
rect 21232 21632 21238 21644
rect 23198 21632 23204 21644
rect 23256 21632 23262 21684
rect 23382 21632 23388 21684
rect 23440 21632 23446 21684
rect 24489 21675 24547 21681
rect 24489 21641 24501 21675
rect 24535 21672 24547 21675
rect 24578 21672 24584 21684
rect 24535 21644 24584 21672
rect 24535 21641 24547 21644
rect 24489 21635 24547 21641
rect 24578 21632 24584 21644
rect 24636 21632 24642 21684
rect 25774 21632 25780 21684
rect 25832 21681 25838 21684
rect 25832 21675 25851 21681
rect 25839 21641 25851 21675
rect 25832 21635 25851 21641
rect 25961 21675 26019 21681
rect 25961 21641 25973 21675
rect 26007 21672 26019 21675
rect 26510 21672 26516 21684
rect 26007 21644 26516 21672
rect 26007 21641 26019 21644
rect 25961 21635 26019 21641
rect 25832 21632 25838 21635
rect 26510 21632 26516 21644
rect 26568 21632 26574 21684
rect 26602 21632 26608 21684
rect 26660 21632 26666 21684
rect 27154 21632 27160 21684
rect 27212 21672 27218 21684
rect 27614 21672 27620 21684
rect 27212 21644 27620 21672
rect 27212 21632 27218 21644
rect 27614 21632 27620 21644
rect 27672 21632 27678 21684
rect 28258 21632 28264 21684
rect 28316 21632 28322 21684
rect 28905 21675 28963 21681
rect 28905 21641 28917 21675
rect 28951 21672 28963 21675
rect 29638 21672 29644 21684
rect 28951 21644 29644 21672
rect 28951 21641 28963 21644
rect 28905 21635 28963 21641
rect 29638 21632 29644 21644
rect 29696 21632 29702 21684
rect 29914 21632 29920 21684
rect 29972 21672 29978 21684
rect 30009 21675 30067 21681
rect 30009 21672 30021 21675
rect 29972 21644 30021 21672
rect 29972 21632 29978 21644
rect 30009 21641 30021 21644
rect 30055 21641 30067 21675
rect 30009 21635 30067 21641
rect 34882 21632 34888 21684
rect 34940 21672 34946 21684
rect 34977 21675 35035 21681
rect 34977 21672 34989 21675
rect 34940 21644 34989 21672
rect 34940 21632 34946 21644
rect 34977 21641 34989 21644
rect 35023 21641 35035 21675
rect 35158 21672 35164 21684
rect 34977 21635 35035 21641
rect 35084 21644 35164 21672
rect 21269 21607 21327 21613
rect 21269 21573 21281 21607
rect 21315 21604 21327 21607
rect 21910 21604 21916 21616
rect 21315 21576 21916 21604
rect 21315 21573 21327 21576
rect 21269 21567 21327 21573
rect 21910 21564 21916 21576
rect 21968 21564 21974 21616
rect 18141 21539 18199 21545
rect 18141 21505 18153 21539
rect 18187 21505 18199 21539
rect 18141 21499 18199 21505
rect 18325 21539 18383 21545
rect 18325 21505 18337 21539
rect 18371 21505 18383 21539
rect 18325 21499 18383 21505
rect 17037 21471 17095 21477
rect 17037 21468 17049 21471
rect 15919 21440 17049 21468
rect 15473 21431 15531 21437
rect 17037 21437 17049 21440
rect 17083 21437 17095 21471
rect 17037 21431 17095 21437
rect 15102 21400 15108 21412
rect 13872 21372 15108 21400
rect 13872 21360 13878 21372
rect 15102 21360 15108 21372
rect 15160 21360 15166 21412
rect 15488 21400 15516 21431
rect 17310 21428 17316 21480
rect 17368 21468 17374 21480
rect 18156 21468 18184 21499
rect 17368 21440 18184 21468
rect 17368 21428 17374 21440
rect 16022 21400 16028 21412
rect 15488 21372 16028 21400
rect 16022 21360 16028 21372
rect 16080 21360 16086 21412
rect 16114 21360 16120 21412
rect 16172 21360 16178 21412
rect 18340 21400 18368 21499
rect 19426 21496 19432 21548
rect 19484 21496 19490 21548
rect 19702 21496 19708 21548
rect 19760 21536 19766 21548
rect 19797 21539 19855 21545
rect 19797 21536 19809 21539
rect 19760 21508 19809 21536
rect 19760 21496 19766 21508
rect 19797 21505 19809 21508
rect 19843 21505 19855 21539
rect 19797 21499 19855 21505
rect 20257 21539 20315 21545
rect 20257 21505 20269 21539
rect 20303 21505 20315 21539
rect 20257 21499 20315 21505
rect 20272 21468 20300 21499
rect 20346 21496 20352 21548
rect 20404 21496 20410 21548
rect 20622 21496 20628 21548
rect 20680 21496 20686 21548
rect 20806 21496 20812 21548
rect 20864 21496 20870 21548
rect 20994 21545 21052 21551
rect 20901 21539 20959 21545
rect 20901 21505 20913 21539
rect 20947 21505 20959 21539
rect 20994 21511 21006 21545
rect 21040 21511 21052 21545
rect 20994 21505 21052 21511
rect 22649 21539 22707 21545
rect 22649 21505 22661 21539
rect 22695 21536 22707 21539
rect 22738 21536 22744 21548
rect 22695 21508 22744 21536
rect 22695 21505 22707 21508
rect 20901 21499 20959 21505
rect 22649 21499 22707 21505
rect 16224 21372 18368 21400
rect 19812 21440 20300 21468
rect 20916 21468 20944 21499
rect 22738 21496 22744 21508
rect 22796 21496 22802 21548
rect 23216 21545 23244 21632
rect 23201 21539 23259 21545
rect 23201 21505 23213 21539
rect 23247 21505 23259 21539
rect 23201 21499 23259 21505
rect 23290 21496 23296 21548
rect 23348 21496 23354 21548
rect 23400 21536 23428 21632
rect 25130 21564 25136 21616
rect 25188 21604 25194 21616
rect 25590 21604 25596 21616
rect 25188 21576 25596 21604
rect 25188 21564 25194 21576
rect 25590 21564 25596 21576
rect 25648 21604 25654 21616
rect 28276 21604 28304 21632
rect 30834 21604 30840 21616
rect 25648 21576 27108 21604
rect 25648 21564 25654 21576
rect 24305 21539 24363 21545
rect 24305 21536 24317 21539
rect 23400 21508 24317 21536
rect 24305 21505 24317 21508
rect 24351 21536 24363 21539
rect 24854 21536 24860 21548
rect 24351 21508 24860 21536
rect 24351 21505 24363 21508
rect 24305 21499 24363 21505
rect 24854 21496 24860 21508
rect 24912 21496 24918 21548
rect 25866 21496 25872 21548
rect 25924 21536 25930 21548
rect 26789 21539 26847 21545
rect 26789 21536 26801 21539
rect 25924 21508 26801 21536
rect 25924 21496 25930 21508
rect 26789 21505 26801 21508
rect 26835 21536 26847 21539
rect 26973 21539 27031 21545
rect 26973 21536 26985 21539
rect 26835 21508 26985 21536
rect 26835 21505 26847 21508
rect 26789 21499 26847 21505
rect 26973 21505 26985 21508
rect 27019 21505 27031 21539
rect 27080 21536 27108 21576
rect 27816 21576 28304 21604
rect 28368 21576 30840 21604
rect 27246 21536 27252 21548
rect 27080 21508 27252 21536
rect 26973 21499 27031 21505
rect 27246 21496 27252 21508
rect 27304 21496 27310 21548
rect 27816 21545 27844 21576
rect 27801 21539 27859 21545
rect 27801 21505 27813 21539
rect 27847 21505 27859 21539
rect 27801 21499 27859 21505
rect 27982 21496 27988 21548
rect 28040 21496 28046 21548
rect 24118 21468 24124 21480
rect 20916 21440 21128 21468
rect 934 21292 940 21344
rect 992 21332 998 21344
rect 1489 21335 1547 21341
rect 1489 21332 1501 21335
rect 992 21304 1501 21332
rect 992 21292 998 21304
rect 1489 21301 1501 21304
rect 1535 21301 1547 21335
rect 1489 21295 1547 21301
rect 1854 21292 1860 21344
rect 1912 21332 1918 21344
rect 1949 21335 2007 21341
rect 1949 21332 1961 21335
rect 1912 21304 1961 21332
rect 1912 21292 1918 21304
rect 1949 21301 1961 21304
rect 1995 21301 2007 21335
rect 1949 21295 2007 21301
rect 7742 21292 7748 21344
rect 7800 21332 7806 21344
rect 9950 21332 9956 21344
rect 7800 21304 9956 21332
rect 7800 21292 7806 21304
rect 9950 21292 9956 21304
rect 10008 21292 10014 21344
rect 10134 21292 10140 21344
rect 10192 21292 10198 21344
rect 10594 21292 10600 21344
rect 10652 21292 10658 21344
rect 11146 21292 11152 21344
rect 11204 21292 11210 21344
rect 13630 21292 13636 21344
rect 13688 21332 13694 21344
rect 13998 21332 14004 21344
rect 13688 21304 14004 21332
rect 13688 21292 13694 21304
rect 13998 21292 14004 21304
rect 14056 21292 14062 21344
rect 14642 21292 14648 21344
rect 14700 21332 14706 21344
rect 16224 21332 16252 21372
rect 19812 21344 19840 21440
rect 21100 21412 21128 21440
rect 22756 21440 24124 21468
rect 20349 21403 20407 21409
rect 20349 21369 20361 21403
rect 20395 21369 20407 21403
rect 20349 21363 20407 21369
rect 14700 21304 16252 21332
rect 14700 21292 14706 21304
rect 16666 21292 16672 21344
rect 16724 21292 16730 21344
rect 17494 21292 17500 21344
rect 17552 21332 17558 21344
rect 18046 21332 18052 21344
rect 17552 21304 18052 21332
rect 17552 21292 17558 21304
rect 18046 21292 18052 21304
rect 18104 21292 18110 21344
rect 19794 21292 19800 21344
rect 19852 21292 19858 21344
rect 20364 21332 20392 21363
rect 21082 21360 21088 21412
rect 21140 21360 21146 21412
rect 22756 21409 22784 21440
rect 24118 21428 24124 21440
rect 24176 21428 24182 21480
rect 22741 21403 22799 21409
rect 22741 21369 22753 21403
rect 22787 21369 22799 21403
rect 24872 21400 24900 21496
rect 26234 21428 26240 21480
rect 26292 21428 26298 21480
rect 26326 21428 26332 21480
rect 26384 21428 26390 21480
rect 26510 21428 26516 21480
rect 26568 21468 26574 21480
rect 28368 21468 28396 21576
rect 28718 21496 28724 21548
rect 28776 21496 28782 21548
rect 28994 21496 29000 21548
rect 29052 21536 29058 21548
rect 29549 21539 29607 21545
rect 29549 21536 29561 21539
rect 29052 21508 29561 21536
rect 29052 21496 29058 21508
rect 29549 21505 29561 21508
rect 29595 21505 29607 21539
rect 29549 21499 29607 21505
rect 29638 21496 29644 21548
rect 29696 21496 29702 21548
rect 29840 21545 29868 21576
rect 30834 21564 30840 21576
rect 30892 21564 30898 21616
rect 35084 21604 35112 21644
rect 35158 21632 35164 21644
rect 35216 21632 35222 21684
rect 36725 21675 36783 21681
rect 36725 21641 36737 21675
rect 36771 21672 36783 21675
rect 36814 21672 36820 21684
rect 36771 21644 36820 21672
rect 36771 21641 36783 21644
rect 36725 21635 36783 21641
rect 36814 21632 36820 21644
rect 36872 21632 36878 21684
rect 31496 21576 35112 21604
rect 31496 21548 31524 21576
rect 29825 21539 29883 21545
rect 29825 21505 29837 21539
rect 29871 21505 29883 21539
rect 29825 21499 29883 21505
rect 31478 21496 31484 21548
rect 31536 21496 31542 21548
rect 34514 21496 34520 21548
rect 34572 21536 34578 21548
rect 34977 21539 35035 21545
rect 34977 21536 34989 21539
rect 34572 21508 34989 21536
rect 34572 21496 34578 21508
rect 34977 21505 34989 21508
rect 35023 21505 35035 21539
rect 35084 21536 35112 21576
rect 35154 21539 35212 21545
rect 35154 21536 35166 21539
rect 35084 21508 35166 21536
rect 34977 21499 35035 21505
rect 35154 21505 35166 21508
rect 35200 21505 35212 21539
rect 35154 21499 35212 21505
rect 36906 21496 36912 21548
rect 36964 21496 36970 21548
rect 37090 21496 37096 21548
rect 37148 21496 37154 21548
rect 37642 21496 37648 21548
rect 37700 21496 37706 21548
rect 26568 21440 28396 21468
rect 28537 21471 28595 21477
rect 26568 21428 26574 21440
rect 28537 21437 28549 21471
rect 28583 21468 28595 21471
rect 28626 21468 28632 21480
rect 28583 21440 28632 21468
rect 28583 21437 28595 21440
rect 28537 21431 28595 21437
rect 28626 21428 28632 21440
rect 28684 21428 28690 21480
rect 28810 21428 28816 21480
rect 28868 21468 28874 21480
rect 28868 21440 31754 21468
rect 28868 21428 28874 21440
rect 26252 21400 26280 21428
rect 24872 21372 25820 21400
rect 26252 21372 27108 21400
rect 22741 21363 22799 21369
rect 25590 21332 25596 21344
rect 20364 21304 25596 21332
rect 25590 21292 25596 21304
rect 25648 21292 25654 21344
rect 25792 21341 25820 21372
rect 27080 21341 27108 21372
rect 27614 21360 27620 21412
rect 27672 21400 27678 21412
rect 30098 21400 30104 21412
rect 27672 21372 30104 21400
rect 27672 21360 27678 21372
rect 30098 21360 30104 21372
rect 30156 21360 30162 21412
rect 25777 21335 25835 21341
rect 25777 21301 25789 21335
rect 25823 21301 25835 21335
rect 25777 21295 25835 21301
rect 27065 21335 27123 21341
rect 27065 21301 27077 21335
rect 27111 21301 27123 21335
rect 27065 21295 27123 21301
rect 27338 21292 27344 21344
rect 27396 21332 27402 21344
rect 27525 21335 27583 21341
rect 27525 21332 27537 21335
rect 27396 21304 27537 21332
rect 27396 21292 27402 21304
rect 27525 21301 27537 21304
rect 27571 21301 27583 21335
rect 27525 21295 27583 21301
rect 28442 21292 28448 21344
rect 28500 21332 28506 21344
rect 31570 21332 31576 21344
rect 28500 21304 31576 21332
rect 28500 21292 28506 21304
rect 31570 21292 31576 21304
rect 31628 21292 31634 21344
rect 31726 21332 31754 21440
rect 34146 21332 34152 21344
rect 31726 21304 34152 21332
rect 34146 21292 34152 21304
rect 34204 21292 34210 21344
rect 37826 21292 37832 21344
rect 37884 21292 37890 21344
rect 1104 21242 38272 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38272 21242
rect 1104 21168 38272 21190
rect 1660 21131 1718 21137
rect 1660 21097 1672 21131
rect 1706 21128 1718 21131
rect 1854 21128 1860 21140
rect 1706 21100 1860 21128
rect 1706 21097 1718 21100
rect 1660 21091 1718 21097
rect 1854 21088 1860 21100
rect 1912 21088 1918 21140
rect 6086 21088 6092 21140
rect 6144 21088 6150 21140
rect 8202 21088 8208 21140
rect 8260 21128 8266 21140
rect 10686 21128 10692 21140
rect 8260 21100 10692 21128
rect 8260 21088 8266 21100
rect 10686 21088 10692 21100
rect 10744 21088 10750 21140
rect 11146 21088 11152 21140
rect 11204 21088 11210 21140
rect 12894 21088 12900 21140
rect 12952 21088 12958 21140
rect 13725 21131 13783 21137
rect 13725 21097 13737 21131
rect 13771 21128 13783 21131
rect 13814 21128 13820 21140
rect 13771 21100 13820 21128
rect 13771 21097 13783 21100
rect 13725 21091 13783 21097
rect 13814 21088 13820 21100
rect 13872 21088 13878 21140
rect 13909 21131 13967 21137
rect 13909 21097 13921 21131
rect 13955 21128 13967 21131
rect 13955 21100 14780 21128
rect 13955 21097 13967 21100
rect 13909 21091 13967 21097
rect 2774 21020 2780 21072
rect 2832 21020 2838 21072
rect 10134 21020 10140 21072
rect 10192 21020 10198 21072
rect 1394 20952 1400 21004
rect 1452 20992 1458 21004
rect 2792 20992 2820 21020
rect 4062 20992 4068 21004
rect 1452 20964 4068 20992
rect 1452 20952 1458 20964
rect 4062 20952 4068 20964
rect 4120 20992 4126 21004
rect 4341 20995 4399 21001
rect 4341 20992 4353 20995
rect 4120 20964 4353 20992
rect 4120 20952 4126 20964
rect 4341 20961 4353 20964
rect 4387 20992 4399 20995
rect 4387 20964 6224 20992
rect 4387 20961 4399 20964
rect 4341 20955 4399 20961
rect 2898 20828 3832 20856
rect 3804 20800 3832 20828
rect 4614 20816 4620 20868
rect 4672 20816 4678 20868
rect 6196 20856 6224 20964
rect 8018 20884 8024 20936
rect 8076 20884 8082 20936
rect 9953 20927 10011 20933
rect 9953 20893 9965 20927
rect 9999 20924 10011 20927
rect 10152 20924 10180 21020
rect 10594 20924 10600 20936
rect 9999 20896 10180 20924
rect 10244 20896 10600 20924
rect 9999 20893 10011 20896
rect 9953 20887 10011 20893
rect 6273 20859 6331 20865
rect 6273 20856 6285 20859
rect 4724 20828 5106 20856
rect 6196 20828 6285 20856
rect 3142 20748 3148 20800
rect 3200 20748 3206 20800
rect 3786 20748 3792 20800
rect 3844 20788 3850 20800
rect 4724 20788 4752 20828
rect 6196 20800 6224 20828
rect 6273 20825 6285 20828
rect 6319 20825 6331 20859
rect 6273 20819 6331 20825
rect 9030 20816 9036 20868
rect 9088 20856 9094 20868
rect 10244 20856 10272 20896
rect 10594 20884 10600 20896
rect 10652 20884 10658 20936
rect 10870 20884 10876 20936
rect 10928 20924 10934 20936
rect 11164 20933 11192 21088
rect 12912 21060 12940 21088
rect 12912 21032 13952 21060
rect 11698 20992 11704 21004
rect 11532 20964 11704 20992
rect 11532 20933 11560 20964
rect 11698 20952 11704 20964
rect 11756 20952 11762 21004
rect 13538 20952 13544 21004
rect 13596 20952 13602 21004
rect 13924 20992 13952 21032
rect 13998 21020 14004 21072
rect 14056 21060 14062 21072
rect 14093 21063 14151 21069
rect 14093 21060 14105 21063
rect 14056 21032 14105 21060
rect 14056 21020 14062 21032
rect 14093 21029 14105 21032
rect 14139 21029 14151 21063
rect 14093 21023 14151 21029
rect 13924 20964 14504 20992
rect 10965 20927 11023 20933
rect 10965 20924 10977 20927
rect 10928 20896 10977 20924
rect 10928 20884 10934 20896
rect 10965 20893 10977 20896
rect 11011 20893 11023 20927
rect 10965 20887 11023 20893
rect 11149 20927 11207 20933
rect 11149 20893 11161 20927
rect 11195 20893 11207 20927
rect 11149 20887 11207 20893
rect 11517 20927 11575 20933
rect 11517 20893 11529 20927
rect 11563 20893 11575 20927
rect 11517 20887 11575 20893
rect 11606 20884 11612 20936
rect 11664 20884 11670 20936
rect 11885 20927 11943 20933
rect 11885 20893 11897 20927
rect 11931 20893 11943 20927
rect 13556 20924 13584 20952
rect 14231 20927 14289 20933
rect 14231 20924 14243 20927
rect 13556 20896 14243 20924
rect 11885 20887 11943 20893
rect 14231 20893 14243 20896
rect 14277 20893 14289 20927
rect 14231 20887 14289 20893
rect 9088 20828 10272 20856
rect 9088 20816 9094 20828
rect 10318 20816 10324 20868
rect 10376 20856 10382 20868
rect 11900 20856 11928 20887
rect 14366 20884 14372 20936
rect 14424 20884 14430 20936
rect 14476 20933 14504 20964
rect 14461 20927 14519 20933
rect 14461 20893 14473 20927
rect 14507 20893 14519 20927
rect 14642 20924 14648 20936
rect 14603 20896 14648 20924
rect 14461 20887 14519 20893
rect 14642 20884 14648 20896
rect 14700 20884 14706 20936
rect 14752 20933 14780 21100
rect 16666 21088 16672 21140
rect 16724 21088 16730 21140
rect 19521 21131 19579 21137
rect 19521 21097 19533 21131
rect 19567 21128 19579 21131
rect 20622 21128 20628 21140
rect 19567 21100 20628 21128
rect 19567 21097 19579 21100
rect 19521 21091 19579 21097
rect 20622 21088 20628 21100
rect 20680 21088 20686 21140
rect 21266 21128 21272 21140
rect 20824 21100 21272 21128
rect 14737 20927 14795 20933
rect 14737 20893 14749 20927
rect 14783 20924 14795 20927
rect 15286 20924 15292 20936
rect 14783 20896 15292 20924
rect 14783 20893 14795 20896
rect 14737 20887 14795 20893
rect 15286 20884 15292 20896
rect 15344 20884 15350 20936
rect 16485 20927 16543 20933
rect 16485 20893 16497 20927
rect 16531 20924 16543 20927
rect 16684 20924 16712 21088
rect 20824 21069 20852 21100
rect 21266 21088 21272 21100
rect 21324 21128 21330 21140
rect 22554 21128 22560 21140
rect 21324 21100 22560 21128
rect 21324 21088 21330 21100
rect 22554 21088 22560 21100
rect 22612 21088 22618 21140
rect 25406 21088 25412 21140
rect 25464 21088 25470 21140
rect 28718 21128 28724 21140
rect 25516 21100 28724 21128
rect 20809 21063 20867 21069
rect 16531 20896 16712 20924
rect 17696 21032 20760 21060
rect 16531 20893 16543 20896
rect 16485 20887 16543 20893
rect 10376 20828 11928 20856
rect 10376 20816 10382 20828
rect 12342 20816 12348 20868
rect 12400 20816 12406 20868
rect 13541 20859 13599 20865
rect 13541 20825 13553 20859
rect 13587 20856 13599 20859
rect 14826 20856 14832 20868
rect 13587 20828 14832 20856
rect 13587 20825 13599 20828
rect 13541 20819 13599 20825
rect 14826 20816 14832 20828
rect 14884 20816 14890 20868
rect 15470 20816 15476 20868
rect 15528 20856 15534 20868
rect 15749 20859 15807 20865
rect 15749 20856 15761 20859
rect 15528 20828 15761 20856
rect 15528 20816 15534 20828
rect 15749 20825 15761 20828
rect 15795 20856 15807 20859
rect 17696 20856 17724 21032
rect 20732 20992 20760 21032
rect 20809 21029 20821 21063
rect 20855 21029 20867 21063
rect 20809 21023 20867 21029
rect 20898 21020 20904 21072
rect 20956 21060 20962 21072
rect 25516 21060 25544 21100
rect 28718 21088 28724 21100
rect 28776 21088 28782 21140
rect 30650 21088 30656 21140
rect 30708 21128 30714 21140
rect 30745 21131 30803 21137
rect 30745 21128 30757 21131
rect 30708 21100 30757 21128
rect 30708 21088 30714 21100
rect 30745 21097 30757 21100
rect 30791 21097 30803 21131
rect 31846 21128 31852 21140
rect 30745 21091 30803 21097
rect 31036 21100 31852 21128
rect 20956 21032 25544 21060
rect 20956 21020 20962 21032
rect 25590 21020 25596 21072
rect 25648 21020 25654 21072
rect 27338 21020 27344 21072
rect 27396 21020 27402 21072
rect 27614 21020 27620 21072
rect 27672 21060 27678 21072
rect 28810 21060 28816 21072
rect 27672 21032 28816 21060
rect 27672 21020 27678 21032
rect 28810 21020 28816 21032
rect 28868 21020 28874 21072
rect 30282 21060 30288 21072
rect 28966 21032 30288 21060
rect 25130 20992 25136 21004
rect 19352 20964 20484 20992
rect 20732 20964 25136 20992
rect 19352 20936 19380 20964
rect 19334 20884 19340 20936
rect 19392 20884 19398 20936
rect 19429 20927 19487 20933
rect 19429 20893 19441 20927
rect 19475 20924 19487 20927
rect 19702 20924 19708 20936
rect 19475 20896 19708 20924
rect 19475 20893 19487 20896
rect 19429 20887 19487 20893
rect 15795 20828 17724 20856
rect 15795 20825 15807 20828
rect 15749 20819 15807 20825
rect 3844 20760 4752 20788
rect 3844 20748 3850 20760
rect 6178 20748 6184 20800
rect 6236 20748 6242 20800
rect 9861 20791 9919 20797
rect 9861 20757 9873 20791
rect 9907 20788 9919 20791
rect 10410 20788 10416 20800
rect 9907 20760 10416 20788
rect 9907 20757 9919 20760
rect 9861 20751 9919 20757
rect 10410 20748 10416 20760
rect 10468 20748 10474 20800
rect 11146 20748 11152 20800
rect 11204 20788 11210 20800
rect 12250 20788 12256 20800
rect 11204 20760 12256 20788
rect 11204 20748 11210 20760
rect 12250 20748 12256 20760
rect 12308 20788 12314 20800
rect 13741 20791 13799 20797
rect 13741 20788 13753 20791
rect 12308 20760 13753 20788
rect 12308 20748 12314 20760
rect 13741 20757 13753 20760
rect 13787 20757 13799 20791
rect 14844 20788 14872 20816
rect 19444 20800 19472 20887
rect 19702 20884 19708 20896
rect 19760 20924 19766 20936
rect 20456 20933 20484 20964
rect 25130 20952 25136 20964
rect 25188 20952 25194 21004
rect 25222 20952 25228 21004
rect 25280 20952 25286 21004
rect 25608 20992 25636 21020
rect 25608 20964 27200 20992
rect 19797 20927 19855 20933
rect 19797 20924 19809 20927
rect 19760 20896 19809 20924
rect 19760 20884 19766 20896
rect 19797 20893 19809 20896
rect 19843 20924 19855 20927
rect 20441 20927 20499 20933
rect 19843 20896 20392 20924
rect 19843 20893 19855 20896
rect 19797 20887 19855 20893
rect 20364 20856 20392 20896
rect 20441 20893 20453 20927
rect 20487 20924 20499 20927
rect 21082 20924 21088 20936
rect 20487 20896 21088 20924
rect 20487 20893 20499 20896
rect 20441 20887 20499 20893
rect 21082 20884 21088 20896
rect 21140 20924 21146 20936
rect 21177 20927 21235 20933
rect 21177 20924 21189 20927
rect 21140 20896 21189 20924
rect 21140 20884 21146 20896
rect 21177 20893 21189 20896
rect 21223 20893 21235 20927
rect 21177 20887 21235 20893
rect 21634 20884 21640 20936
rect 21692 20924 21698 20936
rect 24026 20924 24032 20936
rect 21692 20896 24032 20924
rect 21692 20884 21698 20896
rect 24026 20884 24032 20896
rect 24084 20884 24090 20936
rect 25685 20927 25743 20933
rect 25685 20893 25697 20927
rect 25731 20924 25743 20927
rect 25731 20896 25820 20924
rect 25731 20893 25743 20896
rect 25685 20887 25743 20893
rect 25792 20868 25820 20896
rect 21361 20859 21419 20865
rect 21361 20856 21373 20859
rect 20364 20828 21373 20856
rect 21361 20825 21373 20828
rect 21407 20825 21419 20859
rect 21361 20819 21419 20825
rect 21545 20859 21603 20865
rect 21545 20825 21557 20859
rect 21591 20856 21603 20859
rect 24397 20859 24455 20865
rect 24397 20856 24409 20859
rect 21591 20828 24409 20856
rect 21591 20825 21603 20828
rect 21545 20819 21603 20825
rect 24397 20825 24409 20828
rect 24443 20825 24455 20859
rect 24397 20819 24455 20825
rect 24762 20816 24768 20868
rect 24820 20856 24826 20868
rect 25409 20859 25467 20865
rect 25409 20856 25421 20859
rect 24820 20828 25421 20856
rect 24820 20816 24826 20828
rect 25409 20825 25421 20828
rect 25455 20825 25467 20859
rect 25409 20819 25467 20825
rect 25774 20816 25780 20868
rect 25832 20816 25838 20868
rect 27172 20856 27200 20964
rect 27249 20927 27307 20933
rect 27249 20893 27261 20927
rect 27295 20924 27307 20927
rect 27356 20924 27384 21020
rect 28966 20992 28994 21032
rect 30282 21020 30288 21032
rect 30340 21020 30346 21072
rect 31036 21069 31064 21100
rect 31846 21088 31852 21100
rect 31904 21088 31910 21140
rect 32398 21088 32404 21140
rect 32456 21088 32462 21140
rect 32861 21131 32919 21137
rect 32861 21097 32873 21131
rect 32907 21128 32919 21131
rect 33686 21128 33692 21140
rect 32907 21100 33692 21128
rect 32907 21097 32919 21100
rect 32861 21091 32919 21097
rect 33686 21088 33692 21100
rect 33744 21088 33750 21140
rect 34256 21100 34652 21128
rect 31021 21063 31079 21069
rect 31021 21029 31033 21063
rect 31067 21029 31079 21063
rect 31021 21023 31079 21029
rect 31481 21063 31539 21069
rect 31481 21029 31493 21063
rect 31527 21029 31539 21063
rect 31481 21023 31539 21029
rect 27295 20896 27384 20924
rect 27632 20964 28994 20992
rect 27295 20893 27307 20896
rect 27249 20887 27307 20893
rect 27632 20856 27660 20964
rect 29822 20952 29828 21004
rect 29880 20992 29886 21004
rect 30190 20992 30196 21004
rect 29880 20964 30196 20992
rect 29880 20952 29886 20964
rect 30190 20952 30196 20964
rect 30248 20992 30254 21004
rect 31205 20995 31263 21001
rect 30248 20964 30328 20992
rect 30248 20952 30254 20964
rect 27706 20884 27712 20936
rect 27764 20884 27770 20936
rect 29638 20884 29644 20936
rect 29696 20924 29702 20936
rect 30300 20933 30328 20964
rect 31205 20961 31217 20995
rect 31251 20992 31263 20995
rect 31496 20992 31524 21023
rect 31570 21020 31576 21072
rect 31628 21060 31634 21072
rect 31754 21060 31760 21072
rect 31628 21032 31760 21060
rect 31628 21020 31634 21032
rect 31754 21020 31760 21032
rect 31812 21020 31818 21072
rect 32416 21060 32444 21088
rect 34256 21072 34284 21100
rect 32416 21032 34100 21060
rect 31251 20964 31524 20992
rect 31251 20961 31263 20964
rect 31205 20955 31263 20961
rect 30101 20927 30159 20933
rect 30101 20924 30113 20927
rect 29696 20896 30113 20924
rect 29696 20884 29702 20896
rect 30101 20893 30113 20896
rect 30147 20893 30159 20927
rect 30101 20887 30159 20893
rect 30285 20927 30343 20933
rect 30285 20893 30297 20927
rect 30331 20893 30343 20927
rect 30285 20887 30343 20893
rect 30469 20927 30527 20933
rect 30469 20893 30481 20927
rect 30515 20924 30527 20927
rect 30929 20927 30987 20933
rect 30929 20924 30941 20927
rect 30515 20896 30941 20924
rect 30515 20893 30527 20896
rect 30469 20887 30527 20893
rect 30929 20893 30941 20896
rect 30975 20924 30987 20927
rect 31018 20924 31024 20936
rect 30975 20896 31024 20924
rect 30975 20893 30987 20896
rect 30929 20887 30987 20893
rect 27172 20828 27660 20856
rect 15562 20788 15568 20800
rect 14844 20760 15568 20788
rect 13741 20751 13799 20757
rect 15562 20748 15568 20760
rect 15620 20748 15626 20800
rect 16298 20748 16304 20800
rect 16356 20788 16362 20800
rect 17310 20788 17316 20800
rect 16356 20760 17316 20788
rect 16356 20748 16362 20760
rect 17310 20748 17316 20760
rect 17368 20748 17374 20800
rect 19426 20748 19432 20800
rect 19484 20748 19490 20800
rect 20714 20748 20720 20800
rect 20772 20788 20778 20800
rect 21450 20788 21456 20800
rect 20772 20760 21456 20788
rect 20772 20748 20778 20760
rect 21450 20748 21456 20760
rect 21508 20748 21514 20800
rect 22554 20748 22560 20800
rect 22612 20788 22618 20800
rect 23474 20788 23480 20800
rect 22612 20760 23480 20788
rect 22612 20748 22618 20760
rect 23474 20748 23480 20760
rect 23532 20748 23538 20800
rect 24210 20748 24216 20800
rect 24268 20788 24274 20800
rect 25498 20788 25504 20800
rect 24268 20760 25504 20788
rect 24268 20748 24274 20760
rect 25498 20748 25504 20760
rect 25556 20748 25562 20800
rect 25593 20791 25651 20797
rect 25593 20757 25605 20791
rect 25639 20788 25651 20791
rect 26786 20788 26792 20800
rect 25639 20760 26792 20788
rect 25639 20757 25651 20760
rect 25593 20751 25651 20757
rect 26786 20748 26792 20760
rect 26844 20748 26850 20800
rect 27065 20791 27123 20797
rect 27065 20757 27077 20791
rect 27111 20788 27123 20791
rect 27724 20788 27752 20884
rect 30116 20856 30144 20887
rect 31018 20884 31024 20896
rect 31076 20884 31082 20936
rect 31110 20884 31116 20936
rect 31168 20884 31174 20936
rect 31294 20884 31300 20936
rect 31352 20924 31358 20936
rect 31772 20933 31800 21020
rect 33318 20952 33324 21004
rect 33376 20952 33382 21004
rect 33870 20952 33876 21004
rect 33928 20992 33934 21004
rect 33965 20995 34023 21001
rect 33965 20992 33977 20995
rect 33928 20964 33977 20992
rect 33928 20952 33934 20964
rect 33965 20961 33977 20964
rect 34011 20961 34023 20995
rect 33965 20955 34023 20961
rect 34072 20992 34100 21032
rect 34238 21020 34244 21072
rect 34296 21020 34302 21072
rect 34422 21020 34428 21072
rect 34480 21020 34486 21072
rect 34624 21060 34652 21100
rect 34698 21088 34704 21140
rect 34756 21088 34762 21140
rect 37182 21128 37188 21140
rect 36280 21100 37188 21128
rect 36280 21060 36308 21100
rect 37182 21088 37188 21100
rect 37240 21088 37246 21140
rect 34624 21032 36308 21060
rect 34514 20992 34520 21004
rect 34072 20964 34520 20992
rect 31389 20927 31447 20933
rect 31389 20924 31401 20927
rect 31352 20896 31401 20924
rect 31352 20884 31358 20896
rect 31389 20893 31401 20896
rect 31435 20893 31447 20927
rect 31389 20887 31447 20893
rect 31757 20927 31815 20933
rect 31757 20893 31769 20927
rect 31803 20893 31815 20927
rect 31757 20887 31815 20893
rect 32858 20884 32864 20936
rect 32916 20924 32922 20936
rect 33045 20927 33103 20933
rect 33045 20924 33057 20927
rect 32916 20896 33057 20924
rect 32916 20884 32922 20896
rect 33045 20893 33057 20896
rect 33091 20893 33103 20927
rect 33045 20887 33103 20893
rect 33137 20927 33195 20933
rect 33137 20893 33149 20927
rect 33183 20924 33195 20927
rect 33226 20924 33232 20936
rect 33183 20896 33232 20924
rect 33183 20893 33195 20896
rect 33137 20887 33195 20893
rect 33226 20884 33232 20896
rect 33284 20884 33290 20936
rect 33410 20884 33416 20936
rect 33468 20884 33474 20936
rect 30116 20828 30420 20856
rect 30392 20800 30420 20828
rect 30558 20816 30564 20868
rect 30616 20856 30622 20868
rect 31478 20856 31484 20868
rect 30616 20828 31484 20856
rect 30616 20816 30622 20828
rect 31478 20816 31484 20828
rect 31536 20816 31542 20868
rect 31570 20816 31576 20868
rect 31628 20856 31634 20868
rect 31665 20859 31723 20865
rect 31665 20856 31677 20859
rect 31628 20828 31677 20856
rect 31628 20816 31634 20828
rect 31665 20825 31677 20828
rect 31711 20856 31723 20859
rect 33888 20856 33916 20952
rect 34072 20933 34100 20964
rect 34514 20952 34520 20964
rect 34572 20952 34578 21004
rect 36280 21001 36308 21032
rect 36725 21063 36783 21069
rect 36725 21029 36737 21063
rect 36771 21060 36783 21063
rect 36771 21032 36860 21060
rect 36771 21029 36783 21032
rect 36725 21023 36783 21029
rect 36832 21004 36860 21032
rect 36906 21020 36912 21072
rect 36964 21020 36970 21072
rect 36265 20995 36323 21001
rect 36265 20961 36277 20995
rect 36311 20961 36323 20995
rect 36265 20955 36323 20961
rect 36814 20952 36820 21004
rect 36872 20952 36878 21004
rect 34057 20927 34115 20933
rect 34057 20893 34069 20927
rect 34103 20893 34115 20927
rect 34057 20887 34115 20893
rect 34146 20884 34152 20936
rect 34204 20924 34210 20936
rect 34422 20924 34428 20936
rect 34204 20896 34428 20924
rect 34204 20884 34210 20896
rect 34422 20884 34428 20896
rect 34480 20924 34486 20936
rect 34701 20927 34759 20933
rect 34701 20924 34713 20927
rect 34480 20896 34713 20924
rect 34480 20884 34486 20896
rect 34701 20893 34713 20896
rect 34747 20893 34759 20927
rect 34701 20887 34759 20893
rect 34885 20927 34943 20933
rect 34885 20893 34897 20927
rect 34931 20893 34943 20927
rect 34885 20887 34943 20893
rect 31711 20828 33916 20856
rect 31711 20825 31723 20828
rect 31665 20819 31723 20825
rect 34606 20816 34612 20868
rect 34664 20856 34670 20868
rect 34900 20856 34928 20887
rect 35986 20884 35992 20936
rect 36044 20924 36050 20936
rect 36357 20927 36415 20933
rect 36357 20924 36369 20927
rect 36044 20896 36369 20924
rect 36044 20884 36050 20896
rect 36357 20893 36369 20896
rect 36403 20893 36415 20927
rect 36357 20887 36415 20893
rect 36906 20884 36912 20936
rect 36964 20924 36970 20936
rect 37047 20927 37105 20933
rect 37047 20924 37059 20927
rect 36964 20896 37059 20924
rect 36964 20884 36970 20896
rect 37047 20893 37059 20896
rect 37093 20893 37105 20927
rect 37047 20887 37105 20893
rect 37182 20884 37188 20936
rect 37240 20884 37246 20936
rect 34664 20828 34928 20856
rect 34664 20816 34670 20828
rect 27111 20760 27752 20788
rect 27111 20757 27123 20760
rect 27065 20751 27123 20757
rect 30374 20748 30380 20800
rect 30432 20788 30438 20800
rect 31588 20788 31616 20816
rect 30432 20760 31616 20788
rect 30432 20748 30438 20760
rect 1104 20698 38272 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 38272 20698
rect 1104 20624 38272 20646
rect 6733 20587 6791 20593
rect 6733 20553 6745 20587
rect 6779 20553 6791 20587
rect 6733 20547 6791 20553
rect 9401 20587 9459 20593
rect 9401 20553 9413 20587
rect 9447 20584 9459 20587
rect 9674 20584 9680 20596
rect 9447 20556 9680 20584
rect 9447 20553 9459 20556
rect 9401 20547 9459 20553
rect 6641 20451 6699 20457
rect 6641 20417 6653 20451
rect 6687 20448 6699 20451
rect 6748 20448 6776 20547
rect 9674 20544 9680 20556
rect 9732 20544 9738 20596
rect 9766 20544 9772 20596
rect 9824 20544 9830 20596
rect 10226 20544 10232 20596
rect 10284 20584 10290 20596
rect 11606 20584 11612 20596
rect 10284 20556 11612 20584
rect 10284 20544 10290 20556
rect 11606 20544 11612 20556
rect 11664 20544 11670 20596
rect 17037 20587 17095 20593
rect 17037 20553 17049 20587
rect 17083 20584 17095 20587
rect 17218 20584 17224 20596
rect 17083 20556 17224 20584
rect 17083 20553 17095 20556
rect 17037 20547 17095 20553
rect 17218 20544 17224 20556
rect 17276 20544 17282 20596
rect 19429 20587 19487 20593
rect 19429 20553 19441 20587
rect 19475 20584 19487 20587
rect 19518 20584 19524 20596
rect 19475 20556 19524 20584
rect 19475 20553 19487 20556
rect 19429 20547 19487 20553
rect 19518 20544 19524 20556
rect 19576 20544 19582 20596
rect 20530 20544 20536 20596
rect 20588 20584 20594 20596
rect 21266 20584 21272 20596
rect 20588 20556 21272 20584
rect 20588 20544 20594 20556
rect 21266 20544 21272 20556
rect 21324 20544 21330 20596
rect 21450 20544 21456 20596
rect 21508 20584 21514 20596
rect 22649 20587 22707 20593
rect 22649 20584 22661 20587
rect 21508 20556 22661 20584
rect 21508 20544 21514 20556
rect 22649 20553 22661 20556
rect 22695 20553 22707 20587
rect 22649 20547 22707 20553
rect 23934 20544 23940 20596
rect 23992 20544 23998 20596
rect 24026 20544 24032 20596
rect 24084 20544 24090 20596
rect 24394 20544 24400 20596
rect 24452 20544 24458 20596
rect 24673 20587 24731 20593
rect 24673 20553 24685 20587
rect 24719 20584 24731 20587
rect 24762 20584 24768 20596
rect 24719 20556 24768 20584
rect 24719 20553 24731 20556
rect 24673 20547 24731 20553
rect 24762 20544 24768 20556
rect 24820 20544 24826 20596
rect 27798 20544 27804 20596
rect 27856 20584 27862 20596
rect 28626 20584 28632 20596
rect 27856 20556 28632 20584
rect 27856 20544 27862 20556
rect 28626 20544 28632 20556
rect 28684 20584 28690 20596
rect 30006 20584 30012 20596
rect 28684 20556 30012 20584
rect 28684 20544 28690 20556
rect 6822 20476 6828 20528
rect 6880 20516 6886 20528
rect 7101 20519 7159 20525
rect 7101 20516 7113 20519
rect 6880 20488 7113 20516
rect 6880 20476 6886 20488
rect 7101 20485 7113 20488
rect 7147 20485 7159 20519
rect 7101 20479 7159 20485
rect 7193 20519 7251 20525
rect 7193 20485 7205 20519
rect 7239 20516 7251 20519
rect 7926 20516 7932 20528
rect 7239 20488 7932 20516
rect 7239 20485 7251 20488
rect 7193 20479 7251 20485
rect 7926 20476 7932 20488
rect 7984 20476 7990 20528
rect 8294 20476 8300 20528
rect 8352 20476 8358 20528
rect 8478 20476 8484 20528
rect 8536 20476 8542 20528
rect 10428 20488 12434 20516
rect 6687 20420 6776 20448
rect 8113 20451 8171 20457
rect 6687 20417 6699 20420
rect 6641 20411 6699 20417
rect 8113 20417 8125 20451
rect 8159 20448 8171 20451
rect 8202 20448 8208 20460
rect 8159 20420 8208 20448
rect 8159 20417 8171 20420
rect 8113 20411 8171 20417
rect 8202 20408 8208 20420
rect 8260 20408 8266 20460
rect 8312 20448 8340 20476
rect 10428 20460 10456 20488
rect 9033 20451 9091 20457
rect 9033 20448 9045 20451
rect 8312 20420 9045 20448
rect 9033 20417 9045 20420
rect 9079 20417 9091 20451
rect 9033 20411 9091 20417
rect 9309 20451 9367 20457
rect 9309 20417 9321 20451
rect 9355 20417 9367 20451
rect 9309 20411 9367 20417
rect 7285 20383 7343 20389
rect 7285 20349 7297 20383
rect 7331 20349 7343 20383
rect 7285 20343 7343 20349
rect 7300 20312 7328 20343
rect 9122 20340 9128 20392
rect 9180 20380 9186 20392
rect 9324 20380 9352 20411
rect 9398 20408 9404 20460
rect 9456 20448 9462 20460
rect 9585 20451 9643 20457
rect 9585 20448 9597 20451
rect 9456 20420 9597 20448
rect 9456 20408 9462 20420
rect 9585 20417 9597 20420
rect 9631 20417 9643 20451
rect 9585 20411 9643 20417
rect 10410 20408 10416 20460
rect 10468 20408 10474 20460
rect 10689 20451 10747 20457
rect 10689 20417 10701 20451
rect 10735 20448 10747 20451
rect 10870 20448 10876 20460
rect 10735 20420 10876 20448
rect 10735 20417 10747 20420
rect 10689 20411 10747 20417
rect 10870 20408 10876 20420
rect 10928 20408 10934 20460
rect 10962 20408 10968 20460
rect 11020 20408 11026 20460
rect 12406 20448 12434 20488
rect 15194 20476 15200 20528
rect 15252 20516 15258 20528
rect 15473 20519 15531 20525
rect 15473 20516 15485 20519
rect 15252 20488 15485 20516
rect 15252 20476 15258 20488
rect 15473 20485 15485 20488
rect 15519 20516 15531 20519
rect 19334 20516 19340 20528
rect 15519 20488 16160 20516
rect 15519 20485 15531 20488
rect 15473 20479 15531 20485
rect 16132 20460 16160 20488
rect 16776 20488 19340 20516
rect 12526 20448 12532 20460
rect 12406 20420 12532 20448
rect 12526 20408 12532 20420
rect 12584 20408 12590 20460
rect 13078 20408 13084 20460
rect 13136 20408 13142 20460
rect 13449 20451 13507 20457
rect 13449 20417 13461 20451
rect 13495 20417 13507 20451
rect 13449 20411 13507 20417
rect 9180 20352 9352 20380
rect 9180 20340 9186 20352
rect 8110 20312 8116 20324
rect 7300 20284 8116 20312
rect 8110 20272 8116 20284
rect 8168 20272 8174 20324
rect 8665 20315 8723 20321
rect 8665 20281 8677 20315
rect 8711 20312 8723 20315
rect 9416 20312 9444 20408
rect 10778 20340 10784 20392
rect 10836 20340 10842 20392
rect 10980 20380 11008 20408
rect 13170 20380 13176 20392
rect 10980 20352 13176 20380
rect 13170 20340 13176 20352
rect 13228 20380 13234 20392
rect 13464 20380 13492 20411
rect 13906 20408 13912 20460
rect 13964 20408 13970 20460
rect 15654 20408 15660 20460
rect 15712 20408 15718 20460
rect 16114 20408 16120 20460
rect 16172 20408 16178 20460
rect 13228 20352 13492 20380
rect 14185 20383 14243 20389
rect 13228 20340 13234 20352
rect 14185 20349 14197 20383
rect 14231 20380 14243 20383
rect 16776 20380 16804 20488
rect 19334 20476 19340 20488
rect 19392 20476 19398 20528
rect 19720 20488 22876 20516
rect 17126 20408 17132 20460
rect 17184 20408 17190 20460
rect 17770 20408 17776 20460
rect 17828 20408 17834 20460
rect 18138 20408 18144 20460
rect 18196 20448 18202 20460
rect 18509 20451 18567 20457
rect 18509 20448 18521 20451
rect 18196 20420 18521 20448
rect 18196 20408 18202 20420
rect 18509 20417 18521 20420
rect 18555 20417 18567 20451
rect 18509 20411 18567 20417
rect 18693 20451 18751 20457
rect 18693 20417 18705 20451
rect 18739 20417 18751 20451
rect 18693 20411 18751 20417
rect 14231 20352 16804 20380
rect 16853 20383 16911 20389
rect 14231 20349 14243 20352
rect 14185 20343 14243 20349
rect 16853 20349 16865 20383
rect 16899 20380 16911 20383
rect 18598 20380 18604 20392
rect 16899 20352 18604 20380
rect 16899 20349 16911 20352
rect 16853 20343 16911 20349
rect 8711 20284 9444 20312
rect 8711 20281 8723 20284
rect 8665 20275 8723 20281
rect 6454 20204 6460 20256
rect 6512 20204 6518 20256
rect 8018 20204 8024 20256
rect 8076 20244 8082 20256
rect 8481 20247 8539 20253
rect 8481 20244 8493 20247
rect 8076 20216 8493 20244
rect 8076 20204 8082 20216
rect 8481 20213 8493 20216
rect 8527 20244 8539 20247
rect 8570 20244 8576 20256
rect 8527 20216 8576 20244
rect 8527 20213 8539 20216
rect 8481 20207 8539 20213
rect 8570 20204 8576 20216
rect 8628 20204 8634 20256
rect 9122 20204 9128 20256
rect 9180 20204 9186 20256
rect 9416 20244 9444 20284
rect 12158 20272 12164 20324
rect 12216 20312 12222 20324
rect 12434 20312 12440 20324
rect 12216 20284 12440 20312
rect 12216 20272 12222 20284
rect 12434 20272 12440 20284
rect 12492 20272 12498 20324
rect 12526 20272 12532 20324
rect 12584 20312 12590 20324
rect 16868 20312 16896 20343
rect 18598 20340 18604 20352
rect 18656 20380 18662 20392
rect 18708 20380 18736 20411
rect 19426 20408 19432 20460
rect 19484 20448 19490 20460
rect 19610 20448 19616 20460
rect 19484 20420 19616 20448
rect 19484 20408 19490 20420
rect 19610 20408 19616 20420
rect 19668 20408 19674 20460
rect 19720 20380 19748 20488
rect 19794 20408 19800 20460
rect 19852 20448 19858 20460
rect 19889 20451 19947 20457
rect 19889 20448 19901 20451
rect 19852 20420 19901 20448
rect 19852 20408 19858 20420
rect 19889 20417 19901 20420
rect 19935 20417 19947 20451
rect 20993 20451 21051 20457
rect 20993 20448 21005 20451
rect 19889 20411 19947 20417
rect 19996 20420 21005 20448
rect 18656 20352 19748 20380
rect 18656 20340 18662 20352
rect 12584 20284 16896 20312
rect 12584 20272 12590 20284
rect 19996 20256 20024 20420
rect 20993 20417 21005 20420
rect 21039 20417 21051 20451
rect 20993 20411 21051 20417
rect 22554 20408 22560 20460
rect 22612 20408 22618 20460
rect 20714 20340 20720 20392
rect 20772 20340 20778 20392
rect 20898 20340 20904 20392
rect 20956 20340 20962 20392
rect 22848 20389 22876 20488
rect 22833 20383 22891 20389
rect 22833 20349 22845 20383
rect 22879 20380 22891 20383
rect 23753 20383 23811 20389
rect 23753 20380 23765 20383
rect 22879 20352 23765 20380
rect 22879 20349 22891 20352
rect 22833 20343 22891 20349
rect 23753 20349 23765 20352
rect 23799 20349 23811 20383
rect 23753 20343 23811 20349
rect 24044 20312 24072 20544
rect 25774 20516 25780 20528
rect 24872 20488 25780 20516
rect 24872 20460 24900 20488
rect 25774 20476 25780 20488
rect 25832 20525 25838 20528
rect 25832 20519 25895 20525
rect 25832 20485 25849 20519
rect 25883 20485 25895 20519
rect 25832 20479 25895 20485
rect 25832 20476 25838 20479
rect 26050 20476 26056 20528
rect 26108 20476 26114 20528
rect 24581 20451 24639 20457
rect 24581 20417 24593 20451
rect 24627 20448 24639 20451
rect 24670 20448 24676 20460
rect 24627 20420 24676 20448
rect 24627 20417 24639 20420
rect 24581 20411 24639 20417
rect 24670 20408 24676 20420
rect 24728 20408 24734 20460
rect 24765 20451 24823 20457
rect 24765 20417 24777 20451
rect 24811 20448 24823 20451
rect 24854 20448 24860 20460
rect 24811 20420 24860 20448
rect 24811 20417 24823 20420
rect 24765 20411 24823 20417
rect 24854 20408 24860 20420
rect 24912 20408 24918 20460
rect 26970 20408 26976 20460
rect 27028 20448 27034 20460
rect 29012 20457 29040 20556
rect 30006 20544 30012 20556
rect 30064 20544 30070 20596
rect 30190 20544 30196 20596
rect 30248 20544 30254 20596
rect 31021 20587 31079 20593
rect 31021 20553 31033 20587
rect 31067 20584 31079 20587
rect 31570 20584 31576 20596
rect 31067 20556 31576 20584
rect 31067 20553 31079 20556
rect 31021 20547 31079 20553
rect 31570 20544 31576 20556
rect 31628 20544 31634 20596
rect 33502 20584 33508 20596
rect 31864 20556 33508 20584
rect 31386 20516 31392 20528
rect 29104 20488 31392 20516
rect 29104 20457 29132 20488
rect 31386 20476 31392 20488
rect 31444 20516 31450 20528
rect 31864 20516 31892 20556
rect 33502 20544 33508 20556
rect 33560 20544 33566 20596
rect 33778 20544 33784 20596
rect 33836 20584 33842 20596
rect 33873 20587 33931 20593
rect 33873 20584 33885 20587
rect 33836 20556 33885 20584
rect 33836 20544 33842 20556
rect 33873 20553 33885 20556
rect 33919 20553 33931 20587
rect 33873 20547 33931 20553
rect 34054 20544 34060 20596
rect 34112 20544 34118 20596
rect 37090 20544 37096 20596
rect 37148 20544 37154 20596
rect 31444 20488 31892 20516
rect 31941 20519 31999 20525
rect 31444 20476 31450 20488
rect 31941 20485 31953 20519
rect 31987 20516 31999 20519
rect 33318 20516 33324 20528
rect 31987 20488 33324 20516
rect 31987 20485 31999 20488
rect 31941 20479 31999 20485
rect 33318 20476 33324 20488
rect 33376 20476 33382 20528
rect 33410 20476 33416 20528
rect 33468 20476 33474 20528
rect 36725 20519 36783 20525
rect 36725 20485 36737 20519
rect 36771 20516 36783 20519
rect 36814 20516 36820 20528
rect 36771 20488 36820 20516
rect 36771 20485 36783 20488
rect 36725 20479 36783 20485
rect 36814 20476 36820 20488
rect 36872 20476 36878 20528
rect 36906 20476 36912 20528
rect 36964 20525 36970 20528
rect 36964 20519 36983 20525
rect 36971 20485 36983 20519
rect 36964 20479 36983 20485
rect 36964 20476 36970 20479
rect 27157 20451 27215 20457
rect 27157 20448 27169 20451
rect 27028 20420 27169 20448
rect 27028 20408 27034 20420
rect 27157 20417 27169 20420
rect 27203 20417 27215 20451
rect 27157 20411 27215 20417
rect 27893 20451 27951 20457
rect 27893 20417 27905 20451
rect 27939 20417 27951 20451
rect 27893 20411 27951 20417
rect 28997 20451 29055 20457
rect 28997 20417 29009 20451
rect 29043 20417 29055 20451
rect 28997 20411 29055 20417
rect 29089 20451 29147 20457
rect 29089 20417 29101 20451
rect 29135 20417 29147 20451
rect 29089 20411 29147 20417
rect 29365 20451 29423 20457
rect 29365 20417 29377 20451
rect 29411 20448 29423 20451
rect 29454 20448 29460 20460
rect 29411 20420 29460 20448
rect 29411 20417 29423 20420
rect 29365 20411 29423 20417
rect 24210 20340 24216 20392
rect 24268 20380 24274 20392
rect 27908 20380 27936 20411
rect 29454 20408 29460 20420
rect 29512 20408 29518 20460
rect 29549 20451 29607 20457
rect 29549 20417 29561 20451
rect 29595 20417 29607 20451
rect 29549 20411 29607 20417
rect 24268 20352 27936 20380
rect 29564 20380 29592 20411
rect 29638 20408 29644 20460
rect 29696 20448 29702 20460
rect 29733 20451 29791 20457
rect 29733 20448 29745 20451
rect 29696 20420 29745 20448
rect 29696 20408 29702 20420
rect 29733 20417 29745 20420
rect 29779 20417 29791 20451
rect 30006 20448 30012 20460
rect 29733 20411 29791 20417
rect 29840 20420 30012 20448
rect 29840 20380 29868 20420
rect 30006 20408 30012 20420
rect 30064 20408 30070 20460
rect 30098 20408 30104 20460
rect 30156 20408 30162 20460
rect 30282 20408 30288 20460
rect 30340 20448 30346 20460
rect 30377 20451 30435 20457
rect 30377 20448 30389 20451
rect 30340 20420 30389 20448
rect 30340 20408 30346 20420
rect 30377 20417 30389 20420
rect 30423 20417 30435 20451
rect 30377 20411 30435 20417
rect 30466 20408 30472 20460
rect 30524 20408 30530 20460
rect 30561 20451 30619 20457
rect 30561 20417 30573 20451
rect 30607 20448 30619 20451
rect 30650 20448 30656 20460
rect 30607 20420 30656 20448
rect 30607 20417 30619 20420
rect 30561 20411 30619 20417
rect 30650 20408 30656 20420
rect 30708 20448 30714 20460
rect 31114 20451 31172 20457
rect 31114 20448 31126 20451
rect 30708 20420 31126 20448
rect 30708 20408 30714 20420
rect 31114 20417 31126 20420
rect 31160 20448 31172 20451
rect 31202 20448 31208 20460
rect 31160 20420 31208 20448
rect 31160 20417 31172 20420
rect 31114 20411 31172 20417
rect 31202 20408 31208 20420
rect 31260 20408 31266 20460
rect 31554 20454 31612 20457
rect 31665 20454 31723 20457
rect 31554 20451 31723 20454
rect 31554 20448 31566 20451
rect 31312 20420 31566 20448
rect 31312 20392 31340 20420
rect 31554 20417 31566 20420
rect 31600 20426 31677 20451
rect 31600 20420 31616 20426
rect 31600 20417 31612 20420
rect 31554 20411 31612 20417
rect 31665 20417 31677 20426
rect 31711 20417 31723 20451
rect 31665 20411 31723 20417
rect 31757 20451 31815 20457
rect 31757 20417 31769 20451
rect 31803 20417 31815 20451
rect 33428 20448 33456 20476
rect 33689 20451 33747 20457
rect 33689 20448 33701 20451
rect 33428 20420 33701 20448
rect 31757 20411 31815 20417
rect 33689 20417 33701 20420
rect 33735 20417 33747 20451
rect 33689 20411 33747 20417
rect 29564 20352 29868 20380
rect 29917 20383 29975 20389
rect 24268 20340 24274 20352
rect 29917 20349 29929 20383
rect 29963 20380 29975 20383
rect 30926 20380 30932 20392
rect 29963 20352 30932 20380
rect 29963 20349 29975 20352
rect 29917 20343 29975 20349
rect 30926 20340 30932 20352
rect 30984 20340 30990 20392
rect 31294 20340 31300 20392
rect 31352 20340 31358 20392
rect 31461 20383 31519 20389
rect 31461 20349 31473 20383
rect 31507 20380 31519 20383
rect 31772 20380 31800 20411
rect 33962 20408 33968 20460
rect 34020 20408 34026 20460
rect 34149 20451 34207 20457
rect 34149 20417 34161 20451
rect 34195 20448 34207 20451
rect 36924 20448 36952 20476
rect 34195 20420 36952 20448
rect 34195 20417 34207 20420
rect 34149 20411 34207 20417
rect 31507 20352 31800 20380
rect 31507 20349 31519 20352
rect 31461 20343 31519 20349
rect 24044 20284 31156 20312
rect 10689 20247 10747 20253
rect 10689 20244 10701 20247
rect 9416 20216 10701 20244
rect 10689 20213 10701 20216
rect 10735 20213 10747 20247
rect 10689 20207 10747 20213
rect 11054 20204 11060 20256
rect 11112 20204 11118 20256
rect 15838 20204 15844 20256
rect 15896 20204 15902 20256
rect 17494 20204 17500 20256
rect 17552 20204 17558 20256
rect 17586 20204 17592 20256
rect 17644 20244 17650 20256
rect 17681 20247 17739 20253
rect 17681 20244 17693 20247
rect 17644 20216 17693 20244
rect 17644 20204 17650 20216
rect 17681 20213 17693 20216
rect 17727 20213 17739 20247
rect 17681 20207 17739 20213
rect 18601 20247 18659 20253
rect 18601 20213 18613 20247
rect 18647 20244 18659 20247
rect 19426 20244 19432 20256
rect 18647 20216 19432 20244
rect 18647 20213 18659 20216
rect 18601 20207 18659 20213
rect 19426 20204 19432 20216
rect 19484 20204 19490 20256
rect 19978 20204 19984 20256
rect 20036 20204 20042 20256
rect 21361 20247 21419 20253
rect 21361 20213 21373 20247
rect 21407 20244 21419 20247
rect 21542 20244 21548 20256
rect 21407 20216 21548 20244
rect 21407 20213 21419 20216
rect 21361 20207 21419 20213
rect 21542 20204 21548 20216
rect 21600 20204 21606 20256
rect 22186 20204 22192 20256
rect 22244 20204 22250 20256
rect 22278 20204 22284 20256
rect 22336 20244 22342 20256
rect 25685 20247 25743 20253
rect 25685 20244 25697 20247
rect 22336 20216 25697 20244
rect 22336 20204 22342 20216
rect 25685 20213 25697 20216
rect 25731 20213 25743 20247
rect 25685 20207 25743 20213
rect 25869 20247 25927 20253
rect 25869 20213 25881 20247
rect 25915 20244 25927 20247
rect 27062 20244 27068 20256
rect 25915 20216 27068 20244
rect 25915 20213 25927 20216
rect 25869 20207 25927 20213
rect 27062 20204 27068 20216
rect 27120 20204 27126 20256
rect 27341 20247 27399 20253
rect 27341 20213 27353 20247
rect 27387 20244 27399 20247
rect 30650 20244 30656 20256
rect 27387 20216 30656 20244
rect 27387 20213 27399 20216
rect 27341 20207 27399 20213
rect 30650 20204 30656 20216
rect 30708 20244 30714 20256
rect 30926 20244 30932 20256
rect 30708 20216 30932 20244
rect 30708 20204 30714 20216
rect 30926 20204 30932 20216
rect 30984 20204 30990 20256
rect 31128 20244 31156 20284
rect 31202 20272 31208 20324
rect 31260 20312 31266 20324
rect 31680 20312 31708 20352
rect 31846 20340 31852 20392
rect 31904 20340 31910 20392
rect 33226 20340 33232 20392
rect 33284 20380 33290 20392
rect 33413 20383 33471 20389
rect 33413 20380 33425 20383
rect 33284 20352 33425 20380
rect 33284 20340 33290 20352
rect 33413 20349 33425 20352
rect 33459 20380 33471 20383
rect 33778 20380 33784 20392
rect 33459 20352 33784 20380
rect 33459 20349 33471 20352
rect 33413 20343 33471 20349
rect 33778 20340 33784 20352
rect 33836 20340 33842 20392
rect 33870 20340 33876 20392
rect 33928 20340 33934 20392
rect 31260 20284 31708 20312
rect 31864 20312 31892 20340
rect 31941 20315 31999 20321
rect 31941 20312 31953 20315
rect 31864 20284 31953 20312
rect 31260 20272 31266 20284
rect 31941 20281 31953 20284
rect 31987 20281 31999 20315
rect 31941 20275 31999 20281
rect 33505 20315 33563 20321
rect 33505 20281 33517 20315
rect 33551 20312 33563 20315
rect 33888 20312 33916 20340
rect 33551 20284 33916 20312
rect 33551 20281 33563 20284
rect 33505 20275 33563 20281
rect 33134 20244 33140 20256
rect 31128 20216 33140 20244
rect 33134 20204 33140 20216
rect 33192 20204 33198 20256
rect 33226 20204 33232 20256
rect 33284 20244 33290 20256
rect 34164 20244 34192 20411
rect 33284 20216 34192 20244
rect 33284 20204 33290 20216
rect 36538 20204 36544 20256
rect 36596 20244 36602 20256
rect 36909 20247 36967 20253
rect 36909 20244 36921 20247
rect 36596 20216 36921 20244
rect 36596 20204 36602 20216
rect 36909 20213 36921 20216
rect 36955 20244 36967 20247
rect 37182 20244 37188 20256
rect 36955 20216 37188 20244
rect 36955 20213 36967 20216
rect 36909 20207 36967 20213
rect 37182 20204 37188 20216
rect 37240 20204 37246 20256
rect 1104 20154 38272 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38272 20154
rect 1104 20080 38272 20102
rect 2976 20012 5488 20040
rect 2593 19975 2651 19981
rect 2593 19941 2605 19975
rect 2639 19941 2651 19975
rect 2593 19935 2651 19941
rect 2133 19839 2191 19845
rect 2133 19805 2145 19839
rect 2179 19836 2191 19839
rect 2608 19836 2636 19935
rect 2976 19845 3004 20012
rect 5460 19984 5488 20012
rect 7926 20000 7932 20052
rect 7984 20000 7990 20052
rect 9766 20000 9772 20052
rect 9824 20000 9830 20052
rect 13906 20000 13912 20052
rect 13964 20000 13970 20052
rect 14274 20000 14280 20052
rect 14332 20040 14338 20052
rect 14553 20043 14611 20049
rect 14553 20040 14565 20043
rect 14332 20012 14565 20040
rect 14332 20000 14338 20012
rect 14553 20009 14565 20012
rect 14599 20009 14611 20043
rect 19794 20040 19800 20052
rect 14553 20003 14611 20009
rect 17052 20012 19800 20040
rect 5442 19932 5448 19984
rect 5500 19932 5506 19984
rect 3237 19907 3295 19913
rect 3237 19873 3249 19907
rect 3283 19904 3295 19907
rect 3326 19904 3332 19916
rect 3283 19876 3332 19904
rect 3283 19873 3295 19876
rect 3237 19867 3295 19873
rect 3326 19864 3332 19876
rect 3384 19864 3390 19916
rect 3789 19907 3847 19913
rect 3789 19873 3801 19907
rect 3835 19904 3847 19907
rect 4062 19904 4068 19916
rect 3835 19876 4068 19904
rect 3835 19873 3847 19876
rect 3789 19867 3847 19873
rect 4062 19864 4068 19876
rect 4120 19864 4126 19916
rect 6178 19864 6184 19916
rect 6236 19864 6242 19916
rect 6454 19864 6460 19916
rect 6512 19864 6518 19916
rect 9493 19907 9551 19913
rect 9493 19873 9505 19907
rect 9539 19904 9551 19907
rect 9784 19904 9812 20000
rect 13446 19972 13452 19984
rect 9539 19876 9812 19904
rect 12360 19944 13452 19972
rect 9539 19873 9551 19876
rect 9493 19867 9551 19873
rect 2179 19808 2636 19836
rect 2961 19839 3019 19845
rect 2179 19805 2191 19808
rect 2133 19799 2191 19805
rect 2961 19805 2973 19839
rect 3007 19805 3019 19839
rect 2961 19799 3019 19805
rect 9401 19839 9459 19845
rect 9401 19805 9413 19839
rect 9447 19836 9459 19839
rect 9674 19836 9680 19848
rect 9447 19808 9680 19836
rect 9447 19805 9459 19808
rect 9401 19799 9459 19805
rect 9674 19796 9680 19808
rect 9732 19796 9738 19848
rect 9766 19796 9772 19848
rect 9824 19796 9830 19848
rect 9858 19796 9864 19848
rect 9916 19796 9922 19848
rect 11054 19796 11060 19848
rect 11112 19796 11118 19848
rect 11606 19796 11612 19848
rect 11664 19836 11670 19848
rect 11882 19836 11888 19848
rect 11664 19808 11888 19836
rect 11664 19796 11670 19808
rect 11882 19796 11888 19808
rect 11940 19836 11946 19848
rect 12360 19845 12388 19944
rect 13446 19932 13452 19944
rect 13504 19932 13510 19984
rect 12805 19907 12863 19913
rect 12805 19873 12817 19907
rect 12851 19904 12863 19907
rect 13357 19907 13415 19913
rect 13357 19904 13369 19907
rect 12851 19876 13369 19904
rect 12851 19873 12863 19876
rect 12805 19867 12863 19873
rect 13357 19873 13369 19876
rect 13403 19904 13415 19907
rect 13924 19904 13952 20000
rect 17052 19972 17080 20012
rect 19794 20000 19800 20012
rect 19852 20000 19858 20052
rect 20898 20000 20904 20052
rect 20956 20040 20962 20052
rect 24210 20040 24216 20052
rect 20956 20012 24216 20040
rect 20956 20000 20962 20012
rect 24210 20000 24216 20012
rect 24268 20000 24274 20052
rect 24394 20000 24400 20052
rect 24452 20000 24458 20052
rect 27246 20040 27252 20052
rect 25148 20012 27252 20040
rect 13403 19876 13952 19904
rect 14016 19944 17080 19972
rect 13403 19873 13415 19876
rect 13357 19867 13415 19873
rect 12161 19839 12219 19845
rect 12161 19836 12173 19839
rect 11940 19808 12173 19836
rect 11940 19796 11946 19808
rect 12161 19805 12173 19808
rect 12207 19805 12219 19839
rect 12161 19799 12219 19805
rect 12345 19839 12403 19845
rect 12345 19805 12357 19839
rect 12391 19805 12403 19839
rect 12345 19799 12403 19805
rect 12437 19839 12495 19845
rect 12437 19805 12449 19839
rect 12483 19805 12495 19839
rect 12437 19799 12495 19805
rect 3326 19728 3332 19780
rect 3384 19728 3390 19780
rect 4062 19728 4068 19780
rect 4120 19728 4126 19780
rect 4448 19740 4554 19768
rect 1946 19660 1952 19712
rect 2004 19660 2010 19712
rect 3053 19703 3111 19709
rect 3053 19669 3065 19703
rect 3099 19700 3111 19703
rect 3142 19700 3148 19712
rect 3099 19672 3148 19700
rect 3099 19669 3111 19672
rect 3053 19663 3111 19669
rect 3142 19660 3148 19672
rect 3200 19660 3206 19712
rect 3344 19700 3372 19728
rect 4448 19700 4476 19740
rect 5994 19728 6000 19780
rect 6052 19768 6058 19780
rect 8294 19768 8300 19780
rect 6052 19740 6946 19768
rect 7760 19740 8300 19768
rect 6052 19728 6058 19740
rect 3344 19672 4476 19700
rect 4798 19660 4804 19712
rect 4856 19700 4862 19712
rect 5537 19703 5595 19709
rect 5537 19700 5549 19703
rect 4856 19672 5549 19700
rect 4856 19660 4862 19672
rect 5537 19669 5549 19672
rect 5583 19700 5595 19703
rect 7760 19700 7788 19740
rect 8294 19728 8300 19740
rect 8352 19728 8358 19780
rect 9306 19728 9312 19780
rect 9364 19768 9370 19780
rect 10137 19771 10195 19777
rect 10137 19768 10149 19771
rect 9364 19740 10149 19768
rect 9364 19728 9370 19740
rect 10137 19737 10149 19740
rect 10183 19737 10195 19771
rect 10505 19771 10563 19777
rect 10505 19768 10517 19771
rect 10137 19731 10195 19737
rect 10244 19740 10517 19768
rect 5583 19672 7788 19700
rect 10045 19703 10103 19709
rect 5583 19669 5595 19672
rect 5537 19663 5595 19669
rect 10045 19669 10057 19703
rect 10091 19700 10103 19703
rect 10244 19700 10272 19740
rect 10505 19737 10517 19740
rect 10551 19737 10563 19771
rect 11072 19768 11100 19796
rect 12452 19768 12480 19799
rect 12526 19796 12532 19848
rect 12584 19796 12590 19848
rect 13078 19796 13084 19848
rect 13136 19796 13142 19848
rect 13170 19796 13176 19848
rect 13228 19796 13234 19848
rect 13541 19839 13599 19845
rect 13541 19805 13553 19839
rect 13587 19836 13599 19839
rect 14016 19836 14044 19944
rect 17494 19932 17500 19984
rect 17552 19932 17558 19984
rect 17589 19975 17647 19981
rect 17589 19941 17601 19975
rect 17635 19972 17647 19975
rect 17862 19972 17868 19984
rect 17635 19944 17868 19972
rect 17635 19941 17647 19944
rect 17589 19935 17647 19941
rect 17862 19932 17868 19944
rect 17920 19932 17926 19984
rect 19150 19932 19156 19984
rect 19208 19972 19214 19984
rect 19208 19944 20484 19972
rect 19208 19932 19214 19944
rect 16942 19904 16948 19916
rect 14292 19876 16948 19904
rect 13587 19808 14044 19836
rect 14185 19839 14243 19845
rect 13587 19805 13599 19808
rect 13541 19799 13599 19805
rect 14185 19805 14197 19839
rect 14231 19805 14243 19839
rect 14185 19799 14243 19805
rect 11072 19740 12480 19768
rect 13188 19768 13216 19796
rect 14200 19768 14228 19799
rect 13188 19740 14228 19768
rect 10505 19731 10563 19737
rect 10091 19672 10272 19700
rect 10091 19669 10103 19672
rect 10045 19663 10103 19669
rect 10318 19660 10324 19712
rect 10376 19660 10382 19712
rect 10410 19660 10416 19712
rect 10468 19660 10474 19712
rect 10597 19703 10655 19709
rect 10597 19669 10609 19703
rect 10643 19700 10655 19703
rect 14292 19700 14320 19876
rect 16942 19864 16948 19876
rect 17000 19864 17006 19916
rect 17129 19907 17187 19913
rect 17129 19873 17141 19907
rect 17175 19904 17187 19907
rect 17512 19904 17540 19932
rect 19978 19904 19984 19916
rect 17175 19876 17540 19904
rect 17788 19876 19984 19904
rect 17175 19873 17187 19876
rect 17129 19867 17187 19873
rect 14366 19796 14372 19848
rect 14424 19836 14430 19848
rect 14921 19839 14979 19845
rect 14921 19836 14933 19839
rect 14424 19808 14933 19836
rect 14424 19796 14430 19808
rect 14921 19805 14933 19808
rect 14967 19805 14979 19839
rect 14921 19799 14979 19805
rect 15102 19796 15108 19848
rect 15160 19796 15166 19848
rect 15654 19836 15660 19848
rect 15212 19808 15660 19836
rect 10643 19672 14320 19700
rect 14553 19703 14611 19709
rect 10643 19669 10655 19672
rect 10597 19663 10655 19669
rect 14553 19669 14565 19703
rect 14599 19700 14611 19703
rect 14642 19700 14648 19712
rect 14599 19672 14648 19700
rect 14599 19669 14611 19672
rect 14553 19663 14611 19669
rect 14642 19660 14648 19672
rect 14700 19660 14706 19712
rect 14737 19703 14795 19709
rect 14737 19669 14749 19703
rect 14783 19700 14795 19703
rect 14826 19700 14832 19712
rect 14783 19672 14832 19700
rect 14783 19669 14795 19672
rect 14737 19663 14795 19669
rect 14826 19660 14832 19672
rect 14884 19660 14890 19712
rect 15212 19709 15240 19808
rect 15654 19796 15660 19808
rect 15712 19796 15718 19848
rect 16114 19796 16120 19848
rect 16172 19796 16178 19848
rect 16482 19796 16488 19848
rect 16540 19836 16546 19848
rect 17788 19836 17816 19876
rect 19978 19864 19984 19876
rect 20036 19864 20042 19916
rect 20456 19913 20484 19944
rect 20714 19932 20720 19984
rect 20772 19972 20778 19984
rect 20990 19972 20996 19984
rect 20772 19944 20996 19972
rect 20772 19932 20778 19944
rect 20990 19932 20996 19944
rect 21048 19972 21054 19984
rect 24412 19972 24440 20000
rect 21048 19944 22232 19972
rect 24412 19944 24716 19972
rect 21048 19932 21054 19944
rect 20441 19907 20499 19913
rect 20441 19873 20453 19907
rect 20487 19873 20499 19907
rect 20441 19867 20499 19873
rect 21637 19907 21695 19913
rect 21637 19873 21649 19907
rect 21683 19904 21695 19907
rect 22097 19907 22155 19913
rect 22097 19904 22109 19907
rect 21683 19876 22109 19904
rect 21683 19873 21695 19876
rect 21637 19867 21695 19873
rect 22097 19873 22109 19876
rect 22143 19873 22155 19907
rect 22204 19904 22232 19944
rect 22204 19876 24532 19904
rect 22097 19867 22155 19873
rect 16540 19808 17816 19836
rect 16540 19796 16546 19808
rect 17862 19796 17868 19848
rect 17920 19796 17926 19848
rect 19058 19796 19064 19848
rect 19116 19796 19122 19848
rect 19334 19796 19340 19848
rect 19392 19836 19398 19848
rect 20165 19839 20223 19845
rect 20165 19836 20177 19839
rect 19392 19808 20177 19836
rect 19392 19796 19398 19808
rect 20165 19805 20177 19808
rect 20211 19805 20223 19839
rect 20165 19799 20223 19805
rect 20533 19839 20591 19845
rect 20533 19805 20545 19839
rect 20579 19836 20591 19839
rect 20622 19836 20628 19848
rect 20579 19808 20628 19836
rect 20579 19805 20591 19808
rect 20533 19799 20591 19805
rect 20622 19796 20628 19808
rect 20680 19796 20686 19848
rect 21545 19839 21603 19845
rect 21545 19805 21557 19839
rect 21591 19805 21603 19839
rect 21545 19799 21603 19805
rect 17770 19768 17776 19780
rect 15764 19740 17776 19768
rect 15764 19712 15792 19740
rect 17770 19728 17776 19740
rect 17828 19768 17834 19780
rect 18233 19771 18291 19777
rect 17828 19740 18184 19768
rect 17828 19728 17834 19740
rect 15197 19703 15255 19709
rect 15197 19669 15209 19703
rect 15243 19669 15255 19703
rect 15197 19663 15255 19669
rect 15470 19660 15476 19712
rect 15528 19660 15534 19712
rect 15746 19660 15752 19712
rect 15804 19660 15810 19712
rect 17218 19660 17224 19712
rect 17276 19660 17282 19712
rect 17402 19660 17408 19712
rect 17460 19700 17466 19712
rect 17681 19703 17739 19709
rect 17681 19700 17693 19703
rect 17460 19672 17693 19700
rect 17460 19660 17466 19672
rect 17681 19669 17693 19672
rect 17727 19669 17739 19703
rect 18156 19700 18184 19740
rect 18233 19737 18245 19771
rect 18279 19768 18291 19771
rect 18322 19768 18328 19780
rect 18279 19740 18328 19768
rect 18279 19737 18291 19740
rect 18233 19731 18291 19737
rect 18322 19728 18328 19740
rect 18380 19728 18386 19780
rect 19242 19728 19248 19780
rect 19300 19768 19306 19780
rect 19521 19771 19579 19777
rect 19521 19768 19533 19771
rect 19300 19740 19533 19768
rect 19300 19728 19306 19740
rect 19521 19737 19533 19740
rect 19567 19737 19579 19771
rect 19521 19731 19579 19737
rect 19610 19728 19616 19780
rect 19668 19768 19674 19780
rect 19705 19771 19763 19777
rect 19705 19768 19717 19771
rect 19668 19740 19717 19768
rect 19668 19728 19674 19740
rect 19705 19737 19717 19740
rect 19751 19737 19763 19771
rect 19705 19731 19763 19737
rect 19794 19728 19800 19780
rect 19852 19768 19858 19780
rect 19889 19771 19947 19777
rect 19889 19768 19901 19771
rect 19852 19740 19901 19768
rect 19852 19728 19858 19740
rect 19889 19737 19901 19740
rect 19935 19737 19947 19771
rect 19889 19731 19947 19737
rect 21174 19728 21180 19780
rect 21232 19728 21238 19780
rect 19334 19700 19340 19712
rect 18156 19672 19340 19700
rect 17681 19663 17739 19669
rect 19334 19660 19340 19672
rect 19392 19700 19398 19712
rect 21560 19700 21588 19799
rect 21818 19796 21824 19848
rect 21876 19796 21882 19848
rect 24504 19836 24532 19876
rect 24578 19864 24584 19916
rect 24636 19864 24642 19916
rect 24688 19913 24716 19944
rect 24673 19907 24731 19913
rect 24673 19873 24685 19907
rect 24719 19873 24731 19907
rect 24673 19867 24731 19873
rect 24854 19836 24860 19848
rect 24504 19808 24860 19836
rect 24854 19796 24860 19808
rect 24912 19796 24918 19848
rect 25148 19836 25176 20012
rect 27246 20000 27252 20012
rect 27304 20040 27310 20052
rect 29178 20040 29184 20052
rect 27304 20012 29184 20040
rect 27304 20000 27310 20012
rect 29178 20000 29184 20012
rect 29236 20040 29242 20052
rect 30282 20040 30288 20052
rect 29236 20012 30288 20040
rect 29236 20000 29242 20012
rect 30282 20000 30288 20012
rect 30340 20000 30346 20052
rect 30374 20000 30380 20052
rect 30432 20000 30438 20052
rect 30558 20000 30564 20052
rect 30616 20000 30622 20052
rect 30837 20043 30895 20049
rect 30837 20009 30849 20043
rect 30883 20040 30895 20043
rect 31110 20040 31116 20052
rect 30883 20012 31116 20040
rect 30883 20009 30895 20012
rect 30837 20003 30895 20009
rect 31110 20000 31116 20012
rect 31168 20000 31174 20052
rect 31481 20043 31539 20049
rect 31481 20009 31493 20043
rect 31527 20040 31539 20043
rect 33873 20043 33931 20049
rect 31527 20012 33825 20040
rect 31527 20009 31539 20012
rect 31481 20003 31539 20009
rect 26510 19932 26516 19984
rect 26568 19972 26574 19984
rect 28077 19975 28135 19981
rect 26568 19944 28028 19972
rect 26568 19932 26574 19944
rect 26234 19864 26240 19916
rect 26292 19904 26298 19916
rect 26292 19876 27384 19904
rect 26292 19864 26298 19876
rect 27356 19848 27384 19876
rect 24964 19808 25176 19836
rect 24964 19780 24992 19808
rect 25222 19796 25228 19848
rect 25280 19796 25286 19848
rect 27246 19796 27252 19848
rect 27304 19796 27310 19848
rect 27338 19796 27344 19848
rect 27396 19796 27402 19848
rect 27709 19839 27767 19845
rect 27709 19805 27721 19839
rect 27755 19836 27767 19839
rect 27798 19836 27804 19848
rect 27755 19808 27804 19836
rect 27755 19805 27767 19808
rect 27709 19799 27767 19805
rect 27798 19796 27804 19808
rect 27856 19796 27862 19848
rect 27893 19839 27951 19845
rect 27893 19805 27905 19839
rect 27939 19805 27951 19839
rect 28000 19836 28028 19944
rect 28077 19941 28089 19975
rect 28123 19972 28135 19975
rect 29086 19972 29092 19984
rect 28123 19944 29092 19972
rect 28123 19941 28135 19944
rect 28077 19935 28135 19941
rect 29086 19932 29092 19944
rect 29144 19932 29150 19984
rect 30101 19975 30159 19981
rect 30101 19941 30113 19975
rect 30147 19972 30159 19975
rect 30742 19972 30748 19984
rect 30147 19944 30748 19972
rect 30147 19941 30159 19944
rect 30101 19935 30159 19941
rect 30742 19932 30748 19944
rect 30800 19932 30806 19984
rect 31754 19972 31760 19984
rect 30852 19944 31760 19972
rect 28166 19864 28172 19916
rect 28224 19904 28230 19916
rect 28224 19876 29868 19904
rect 28224 19864 28230 19876
rect 28261 19839 28319 19845
rect 28261 19836 28273 19839
rect 28000 19808 28273 19836
rect 27893 19799 27951 19805
rect 28261 19805 28273 19808
rect 28307 19805 28319 19839
rect 28261 19799 28319 19805
rect 22373 19771 22431 19777
rect 22373 19768 22385 19771
rect 22020 19740 22385 19768
rect 22020 19709 22048 19740
rect 22373 19737 22385 19740
rect 22419 19737 22431 19771
rect 24026 19768 24032 19780
rect 23598 19740 24032 19768
rect 22373 19731 22431 19737
rect 24026 19728 24032 19740
rect 24084 19728 24090 19780
rect 24765 19771 24823 19777
rect 24765 19737 24777 19771
rect 24811 19768 24823 19771
rect 24946 19768 24952 19780
rect 24811 19740 24952 19768
rect 24811 19737 24823 19740
rect 24765 19731 24823 19737
rect 24946 19728 24952 19740
rect 25004 19728 25010 19780
rect 25038 19728 25044 19780
rect 25096 19768 25102 19780
rect 25501 19771 25559 19777
rect 25501 19768 25513 19771
rect 25096 19740 25513 19768
rect 25096 19728 25102 19740
rect 25501 19737 25513 19740
rect 25547 19737 25559 19771
rect 27356 19768 27384 19796
rect 27908 19768 27936 19799
rect 28626 19796 28632 19848
rect 28684 19796 28690 19848
rect 29454 19796 29460 19848
rect 29512 19836 29518 19848
rect 29840 19845 29868 19876
rect 30190 19864 30196 19916
rect 30248 19904 30254 19916
rect 30248 19876 30436 19904
rect 30248 19864 30254 19876
rect 29549 19839 29607 19845
rect 29549 19836 29561 19839
rect 29512 19808 29561 19836
rect 29512 19796 29518 19808
rect 29549 19805 29561 19808
rect 29595 19805 29607 19839
rect 29549 19799 29607 19805
rect 29825 19839 29883 19845
rect 29825 19805 29837 19839
rect 29871 19805 29883 19839
rect 29825 19799 29883 19805
rect 29917 19839 29975 19845
rect 29917 19805 29929 19839
rect 29963 19836 29975 19839
rect 30098 19836 30104 19848
rect 29963 19808 30104 19836
rect 29963 19805 29975 19808
rect 29917 19799 29975 19805
rect 30098 19796 30104 19808
rect 30156 19796 30162 19848
rect 30408 19811 30436 19876
rect 30852 19845 30880 19944
rect 31754 19932 31760 19944
rect 31812 19932 31818 19984
rect 32033 19975 32091 19981
rect 32033 19941 32045 19975
rect 32079 19941 32091 19975
rect 32033 19935 32091 19941
rect 30926 19864 30932 19916
rect 30984 19904 30990 19916
rect 31113 19907 31171 19913
rect 31113 19904 31125 19907
rect 30984 19876 31125 19904
rect 30984 19864 30990 19876
rect 31113 19873 31125 19876
rect 31159 19873 31171 19907
rect 31113 19867 31171 19873
rect 30653 19839 30711 19845
rect 30408 19805 30481 19811
rect 26726 19740 27292 19768
rect 27356 19740 27936 19768
rect 29733 19771 29791 19777
rect 25501 19731 25559 19737
rect 19392 19672 21588 19700
rect 22005 19703 22063 19709
rect 19392 19660 19398 19672
rect 22005 19669 22017 19703
rect 22051 19669 22063 19703
rect 22005 19663 22063 19669
rect 23658 19660 23664 19712
rect 23716 19700 23722 19712
rect 23845 19703 23903 19709
rect 23845 19700 23857 19703
rect 23716 19672 23857 19700
rect 23716 19660 23722 19672
rect 23845 19669 23857 19672
rect 23891 19669 23903 19703
rect 23845 19663 23903 19669
rect 25130 19660 25136 19712
rect 25188 19660 25194 19712
rect 26326 19660 26332 19712
rect 26384 19700 26390 19712
rect 26804 19700 26832 19740
rect 27264 19712 27292 19740
rect 29733 19737 29745 19771
rect 29779 19737 29791 19771
rect 29733 19731 29791 19737
rect 26384 19672 26832 19700
rect 26384 19660 26390 19672
rect 27246 19660 27252 19712
rect 27304 19660 27310 19712
rect 29748 19700 29776 19731
rect 30006 19728 30012 19780
rect 30064 19728 30070 19780
rect 30193 19771 30251 19777
rect 30193 19737 30205 19771
rect 30239 19768 30251 19771
rect 30282 19768 30288 19780
rect 30239 19740 30288 19768
rect 30239 19737 30251 19740
rect 30193 19731 30251 19737
rect 30282 19728 30288 19740
rect 30340 19728 30346 19780
rect 30408 19774 30435 19805
rect 30423 19771 30435 19774
rect 30469 19771 30481 19805
rect 30653 19805 30665 19839
rect 30699 19805 30711 19839
rect 30653 19799 30711 19805
rect 30837 19839 30895 19845
rect 30837 19805 30849 19839
rect 30883 19805 30895 19839
rect 30837 19799 30895 19805
rect 31021 19839 31079 19845
rect 31021 19805 31033 19839
rect 31067 19805 31079 19839
rect 31021 19799 31079 19805
rect 30423 19765 30481 19771
rect 30668 19768 30696 19799
rect 31036 19768 31064 19799
rect 30668 19740 31064 19768
rect 31128 19768 31156 19867
rect 31202 19864 31208 19916
rect 31260 19904 31266 19916
rect 31260 19876 31892 19904
rect 31260 19864 31266 19876
rect 31294 19796 31300 19848
rect 31352 19836 31358 19848
rect 31864 19845 31892 19876
rect 31757 19839 31815 19845
rect 31757 19836 31769 19839
rect 31352 19808 31769 19836
rect 31352 19796 31358 19808
rect 31757 19805 31769 19808
rect 31803 19805 31815 19839
rect 31757 19799 31815 19805
rect 31849 19839 31907 19845
rect 31849 19805 31861 19839
rect 31895 19805 31907 19839
rect 32048 19836 32076 19935
rect 33226 19932 33232 19984
rect 33284 19932 33290 19984
rect 33797 19972 33825 20012
rect 33873 20009 33885 20043
rect 33919 20040 33931 20043
rect 33962 20040 33968 20052
rect 33919 20012 33968 20040
rect 33919 20009 33931 20012
rect 33873 20003 33931 20009
rect 33962 20000 33968 20012
rect 34020 20000 34026 20052
rect 34790 20000 34796 20052
rect 34848 20000 34854 20052
rect 35342 20000 35348 20052
rect 35400 20040 35406 20052
rect 35400 20012 35848 20040
rect 35400 20000 35406 20012
rect 35158 19972 35164 19984
rect 33797 19944 35164 19972
rect 35158 19932 35164 19944
rect 35216 19972 35222 19984
rect 35216 19944 35572 19972
rect 35216 19932 35222 19944
rect 33870 19904 33876 19916
rect 33704 19876 33876 19904
rect 33704 19845 33732 19876
rect 33870 19864 33876 19876
rect 33928 19864 33934 19916
rect 34514 19864 34520 19916
rect 34572 19864 34578 19916
rect 35250 19864 35256 19916
rect 35308 19864 35314 19916
rect 35544 19913 35572 19944
rect 35529 19907 35587 19913
rect 35529 19873 35541 19907
rect 35575 19873 35587 19907
rect 35529 19867 35587 19873
rect 33413 19839 33471 19845
rect 33413 19836 33425 19839
rect 32048 19808 33425 19836
rect 31849 19799 31907 19805
rect 33413 19805 33425 19808
rect 33459 19805 33471 19839
rect 33413 19799 33471 19805
rect 33689 19839 33747 19845
rect 33689 19805 33701 19839
rect 33735 19805 33747 19839
rect 33689 19799 33747 19805
rect 33781 19839 33839 19845
rect 33781 19805 33793 19839
rect 33827 19805 33839 19839
rect 33781 19799 33839 19805
rect 33965 19839 34023 19845
rect 33965 19805 33977 19839
rect 34011 19836 34023 19839
rect 34532 19836 34560 19864
rect 35066 19836 35072 19848
rect 34011 19808 35072 19836
rect 34011 19805 34023 19808
rect 33965 19799 34023 19805
rect 31662 19768 31668 19780
rect 31128 19740 31668 19768
rect 30024 19700 30052 19728
rect 30668 19712 30696 19740
rect 31662 19728 31668 19740
rect 31720 19768 31726 19780
rect 32033 19771 32091 19777
rect 32033 19768 32045 19771
rect 31720 19740 32045 19768
rect 31720 19728 31726 19740
rect 32033 19737 32045 19740
rect 32079 19737 32091 19771
rect 33428 19768 33456 19799
rect 33796 19768 33824 19799
rect 35066 19796 35072 19808
rect 35124 19836 35130 19848
rect 35820 19845 35848 20012
rect 36078 20000 36084 20052
rect 36136 20000 36142 20052
rect 36538 20000 36544 20052
rect 36596 20000 36602 20052
rect 36630 20000 36636 20052
rect 36688 20040 36694 20052
rect 36725 20043 36783 20049
rect 36725 20040 36737 20043
rect 36688 20012 36737 20040
rect 36688 20000 36694 20012
rect 36725 20009 36737 20012
rect 36771 20009 36783 20043
rect 36725 20003 36783 20009
rect 35161 19839 35219 19845
rect 35161 19836 35173 19839
rect 35124 19808 35173 19836
rect 35124 19796 35130 19808
rect 35161 19805 35173 19808
rect 35207 19805 35219 19839
rect 35161 19799 35219 19805
rect 35437 19839 35495 19845
rect 35437 19805 35449 19839
rect 35483 19805 35495 19839
rect 35437 19799 35495 19805
rect 35805 19839 35863 19845
rect 35805 19805 35817 19839
rect 35851 19805 35863 19839
rect 35805 19799 35863 19805
rect 35897 19839 35955 19845
rect 35897 19805 35909 19839
rect 35943 19836 35955 19839
rect 35986 19836 35992 19848
rect 35943 19808 35992 19836
rect 35943 19805 35955 19808
rect 35897 19799 35955 19805
rect 33428 19740 33824 19768
rect 32033 19731 32091 19737
rect 35452 19712 35480 19799
rect 35820 19768 35848 19799
rect 35986 19796 35992 19808
rect 36044 19836 36050 19848
rect 36357 19839 36415 19845
rect 36357 19836 36369 19839
rect 36044 19808 36369 19836
rect 36044 19796 36050 19808
rect 36357 19805 36369 19808
rect 36403 19836 36415 19839
rect 36633 19839 36691 19845
rect 36633 19836 36645 19839
rect 36403 19808 36645 19836
rect 36403 19805 36415 19808
rect 36357 19799 36415 19805
rect 36633 19805 36645 19808
rect 36679 19805 36691 19839
rect 36633 19799 36691 19805
rect 36817 19839 36875 19845
rect 36817 19805 36829 19839
rect 36863 19805 36875 19839
rect 36817 19799 36875 19805
rect 36173 19771 36231 19777
rect 36173 19768 36185 19771
rect 35820 19740 36185 19768
rect 36173 19737 36185 19740
rect 36219 19768 36231 19771
rect 36832 19768 36860 19799
rect 36219 19740 36860 19768
rect 36219 19737 36231 19740
rect 36173 19731 36231 19737
rect 29748 19672 30052 19700
rect 30650 19660 30656 19712
rect 30708 19660 30714 19712
rect 33410 19660 33416 19712
rect 33468 19700 33474 19712
rect 33597 19703 33655 19709
rect 33597 19700 33609 19703
rect 33468 19672 33609 19700
rect 33468 19660 33474 19672
rect 33597 19669 33609 19672
rect 33643 19669 33655 19703
rect 33597 19663 33655 19669
rect 35434 19660 35440 19712
rect 35492 19660 35498 19712
rect 1104 19610 38272 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 38272 19610
rect 1104 19536 38272 19558
rect 4062 19456 4068 19508
rect 4120 19456 4126 19508
rect 4341 19499 4399 19505
rect 4341 19465 4353 19499
rect 4387 19465 4399 19499
rect 4341 19459 4399 19465
rect 1673 19431 1731 19437
rect 1673 19397 1685 19431
rect 1719 19428 1731 19431
rect 1946 19428 1952 19440
rect 1719 19400 1952 19428
rect 1719 19397 1731 19400
rect 1673 19391 1731 19397
rect 1946 19388 1952 19400
rect 2004 19388 2010 19440
rect 3142 19388 3148 19440
rect 3200 19388 3206 19440
rect 1394 19320 1400 19372
rect 1452 19320 1458 19372
rect 2792 19156 2820 19346
rect 3160 19301 3188 19388
rect 4249 19363 4307 19369
rect 4249 19329 4261 19363
rect 4295 19360 4307 19363
rect 4356 19360 4384 19459
rect 4798 19456 4804 19508
rect 4856 19456 4862 19508
rect 5810 19456 5816 19508
rect 5868 19456 5874 19508
rect 6733 19499 6791 19505
rect 6733 19465 6745 19499
rect 6779 19496 6791 19499
rect 6822 19496 6828 19508
rect 6779 19468 6828 19496
rect 6779 19465 6791 19468
rect 6733 19459 6791 19465
rect 6822 19456 6828 19468
rect 6880 19456 6886 19508
rect 11882 19456 11888 19508
rect 11940 19496 11946 19508
rect 12647 19499 12705 19505
rect 11940 19468 12296 19496
rect 11940 19456 11946 19468
rect 4706 19388 4712 19440
rect 4764 19428 4770 19440
rect 5828 19428 5856 19456
rect 4764 19400 5856 19428
rect 4764 19388 4770 19400
rect 9490 19388 9496 19440
rect 9548 19428 9554 19440
rect 10229 19431 10287 19437
rect 10229 19428 10241 19431
rect 9548 19400 10241 19428
rect 9548 19388 9554 19400
rect 10229 19397 10241 19400
rect 10275 19428 10287 19431
rect 10686 19428 10692 19440
rect 10275 19400 10692 19428
rect 10275 19397 10287 19400
rect 10229 19391 10287 19397
rect 10686 19388 10692 19400
rect 10744 19428 10750 19440
rect 11606 19428 11612 19440
rect 10744 19400 11612 19428
rect 10744 19388 10750 19400
rect 11606 19388 11612 19400
rect 11664 19388 11670 19440
rect 12268 19428 12296 19468
rect 12647 19465 12659 19499
rect 12693 19496 12705 19499
rect 12693 19468 13768 19496
rect 12693 19465 12705 19468
rect 12647 19459 12705 19465
rect 13740 19440 13768 19468
rect 14550 19456 14556 19508
rect 14608 19456 14614 19508
rect 15102 19456 15108 19508
rect 15160 19496 15166 19508
rect 15160 19468 15608 19496
rect 15160 19456 15166 19468
rect 12437 19431 12495 19437
rect 12437 19428 12449 19431
rect 12268 19400 12449 19428
rect 12437 19397 12449 19400
rect 12483 19397 12495 19431
rect 13633 19431 13691 19437
rect 13633 19428 13645 19431
rect 12437 19391 12495 19397
rect 13280 19400 13645 19428
rect 4295 19332 4384 19360
rect 6825 19363 6883 19369
rect 4295 19329 4307 19332
rect 4249 19323 4307 19329
rect 6825 19329 6837 19363
rect 6871 19360 6883 19363
rect 8018 19360 8024 19372
rect 6871 19332 8024 19360
rect 6871 19329 6883 19332
rect 6825 19323 6883 19329
rect 8018 19320 8024 19332
rect 8076 19320 8082 19372
rect 9674 19320 9680 19372
rect 9732 19320 9738 19372
rect 9766 19320 9772 19372
rect 9824 19360 9830 19372
rect 10045 19363 10103 19369
rect 10045 19360 10057 19363
rect 9824 19332 10057 19360
rect 9824 19320 9830 19332
rect 10045 19329 10057 19332
rect 10091 19360 10103 19363
rect 10321 19363 10379 19369
rect 10091 19332 10272 19360
rect 10091 19329 10103 19332
rect 10045 19323 10103 19329
rect 3145 19295 3203 19301
rect 3145 19261 3157 19295
rect 3191 19261 3203 19295
rect 3145 19255 3203 19261
rect 3234 19252 3240 19304
rect 3292 19252 3298 19304
rect 4893 19295 4951 19301
rect 4893 19261 4905 19295
rect 4939 19261 4951 19295
rect 4893 19255 4951 19261
rect 3252 19224 3280 19252
rect 4908 19224 4936 19255
rect 5350 19252 5356 19304
rect 5408 19252 5414 19304
rect 6917 19295 6975 19301
rect 6917 19261 6929 19295
rect 6963 19261 6975 19295
rect 6917 19255 6975 19261
rect 9493 19295 9551 19301
rect 9493 19261 9505 19295
rect 9539 19292 9551 19295
rect 9858 19292 9864 19304
rect 9539 19264 9864 19292
rect 9539 19261 9551 19264
rect 9493 19255 9551 19261
rect 3252 19196 4936 19224
rect 5368 19224 5396 19252
rect 6932 19224 6960 19255
rect 9858 19252 9864 19264
rect 9916 19252 9922 19304
rect 9953 19295 10011 19301
rect 9953 19261 9965 19295
rect 9999 19292 10011 19295
rect 10134 19292 10140 19304
rect 9999 19264 10140 19292
rect 9999 19261 10011 19264
rect 9953 19255 10011 19261
rect 10134 19252 10140 19264
rect 10192 19252 10198 19304
rect 5368 19196 6960 19224
rect 10244 19224 10272 19332
rect 10321 19329 10333 19363
rect 10367 19329 10379 19363
rect 11624 19360 11652 19388
rect 11701 19363 11759 19369
rect 11701 19360 11713 19363
rect 11624 19332 11713 19360
rect 10321 19323 10379 19329
rect 11701 19329 11713 19332
rect 11747 19360 11759 19363
rect 11882 19360 11888 19372
rect 11747 19332 11888 19360
rect 11747 19329 11759 19332
rect 11701 19323 11759 19329
rect 10336 19292 10364 19323
rect 11882 19320 11888 19332
rect 11940 19320 11946 19372
rect 11974 19320 11980 19372
rect 12032 19360 12038 19372
rect 12069 19363 12127 19369
rect 12069 19360 12081 19363
rect 12032 19332 12081 19360
rect 12032 19320 12038 19332
rect 12069 19329 12081 19332
rect 12115 19329 12127 19363
rect 12069 19323 12127 19329
rect 12268 19358 12848 19360
rect 12894 19358 12900 19372
rect 12268 19332 12900 19358
rect 10502 19292 10508 19304
rect 10336 19264 10508 19292
rect 10502 19252 10508 19264
rect 10560 19252 10566 19304
rect 10594 19252 10600 19304
rect 10652 19292 10658 19304
rect 11609 19295 11667 19301
rect 11609 19292 11621 19295
rect 10652 19264 11621 19292
rect 10652 19252 10658 19264
rect 11609 19261 11621 19264
rect 11655 19261 11667 19295
rect 11609 19255 11667 19261
rect 11054 19224 11060 19236
rect 10244 19196 11060 19224
rect 11054 19184 11060 19196
rect 11112 19184 11118 19236
rect 3326 19156 3332 19168
rect 2792 19128 3332 19156
rect 3326 19116 3332 19128
rect 3384 19116 3390 19168
rect 6362 19116 6368 19168
rect 6420 19116 6426 19168
rect 7742 19116 7748 19168
rect 7800 19156 7806 19168
rect 8478 19156 8484 19168
rect 7800 19128 8484 19156
rect 7800 19116 7806 19128
rect 8478 19116 8484 19128
rect 8536 19116 8542 19168
rect 9861 19159 9919 19165
rect 9861 19125 9873 19159
rect 9907 19156 9919 19159
rect 10045 19159 10103 19165
rect 10045 19156 10057 19159
rect 9907 19128 10057 19156
rect 9907 19125 9919 19128
rect 9861 19119 9919 19125
rect 10045 19125 10057 19128
rect 10091 19125 10103 19159
rect 10045 19119 10103 19125
rect 11974 19116 11980 19168
rect 12032 19116 12038 19168
rect 12084 19156 12112 19323
rect 12268 19233 12296 19332
rect 12820 19330 12900 19332
rect 12894 19320 12900 19330
rect 12952 19320 12958 19372
rect 13081 19363 13139 19369
rect 13081 19329 13093 19363
rect 13127 19360 13139 19363
rect 13170 19360 13176 19372
rect 13127 19332 13176 19360
rect 13127 19329 13139 19332
rect 13081 19323 13139 19329
rect 13170 19320 13176 19332
rect 13228 19320 13234 19372
rect 13280 19292 13308 19400
rect 13633 19397 13645 19400
rect 13679 19397 13691 19431
rect 13633 19391 13691 19397
rect 13722 19388 13728 19440
rect 13780 19388 13786 19440
rect 14568 19428 14596 19456
rect 14568 19400 15424 19428
rect 13446 19320 13452 19372
rect 13504 19360 13510 19372
rect 14568 19360 14596 19400
rect 14737 19363 14795 19369
rect 14737 19360 14749 19363
rect 13504 19332 13768 19360
rect 14568 19332 14749 19360
rect 13504 19320 13510 19332
rect 12820 19264 13308 19292
rect 13740 19292 13768 19332
rect 14737 19329 14749 19332
rect 14783 19329 14795 19363
rect 14737 19323 14795 19329
rect 15286 19320 15292 19372
rect 15344 19320 15350 19372
rect 15396 19369 15424 19400
rect 15580 19369 15608 19468
rect 17218 19456 17224 19508
rect 17276 19496 17282 19508
rect 18785 19499 18843 19505
rect 18785 19496 18797 19499
rect 17276 19468 18797 19496
rect 17276 19456 17282 19468
rect 18785 19465 18797 19468
rect 18831 19465 18843 19499
rect 18785 19459 18843 19465
rect 15654 19388 15660 19440
rect 15712 19428 15718 19440
rect 15933 19431 15991 19437
rect 15933 19428 15945 19431
rect 15712 19400 15945 19428
rect 15712 19388 15718 19400
rect 15933 19397 15945 19400
rect 15979 19397 15991 19431
rect 17586 19428 17592 19440
rect 15933 19391 15991 19397
rect 17052 19400 17592 19428
rect 17052 19369 17080 19400
rect 17586 19388 17592 19400
rect 17644 19388 17650 19440
rect 18322 19388 18328 19440
rect 18380 19388 18386 19440
rect 18800 19372 18828 19459
rect 21818 19456 21824 19508
rect 21876 19496 21882 19508
rect 22005 19499 22063 19505
rect 22005 19496 22017 19499
rect 21876 19468 22017 19496
rect 21876 19456 21882 19468
rect 22005 19465 22017 19468
rect 22051 19465 22063 19499
rect 22005 19459 22063 19465
rect 22186 19456 22192 19508
rect 22244 19496 22250 19508
rect 22465 19499 22523 19505
rect 22465 19496 22477 19499
rect 22244 19468 22477 19496
rect 22244 19456 22250 19468
rect 22465 19465 22477 19468
rect 22511 19465 22523 19499
rect 22465 19459 22523 19465
rect 25038 19456 25044 19508
rect 25096 19456 25102 19508
rect 25222 19456 25228 19508
rect 25280 19496 25286 19508
rect 25409 19499 25467 19505
rect 25409 19496 25421 19499
rect 25280 19468 25421 19496
rect 25280 19456 25286 19468
rect 25409 19465 25421 19468
rect 25455 19465 25467 19499
rect 25409 19459 25467 19465
rect 25516 19468 26924 19496
rect 19058 19388 19064 19440
rect 19116 19428 19122 19440
rect 25516 19428 25544 19468
rect 26896 19428 26924 19468
rect 26970 19456 26976 19508
rect 27028 19456 27034 19508
rect 30374 19496 30380 19508
rect 27080 19468 30380 19496
rect 27080 19428 27108 19468
rect 30374 19456 30380 19468
rect 30432 19456 30438 19508
rect 30561 19499 30619 19505
rect 30561 19465 30573 19499
rect 30607 19496 30619 19499
rect 30650 19496 30656 19508
rect 30607 19468 30656 19496
rect 30607 19465 30619 19468
rect 30561 19459 30619 19465
rect 30650 19456 30656 19468
rect 30708 19456 30714 19508
rect 31202 19456 31208 19508
rect 31260 19496 31266 19508
rect 31481 19499 31539 19505
rect 31481 19496 31493 19499
rect 31260 19468 31493 19496
rect 31260 19456 31266 19468
rect 31481 19465 31493 19468
rect 31527 19465 31539 19499
rect 31481 19459 31539 19465
rect 35066 19456 35072 19508
rect 35124 19456 35130 19508
rect 35158 19456 35164 19508
rect 35216 19456 35222 19508
rect 35250 19456 35256 19508
rect 35308 19496 35314 19508
rect 35437 19499 35495 19505
rect 35437 19496 35449 19499
rect 35308 19468 35449 19496
rect 35308 19456 35314 19468
rect 35437 19465 35449 19468
rect 35483 19465 35495 19499
rect 35437 19459 35495 19465
rect 27154 19437 27160 19440
rect 19116 19400 25544 19428
rect 26068 19400 26280 19428
rect 26896 19400 27108 19428
rect 27141 19431 27160 19437
rect 19116 19388 19122 19400
rect 15381 19363 15439 19369
rect 15381 19329 15393 19363
rect 15427 19329 15439 19363
rect 15381 19323 15439 19329
rect 15565 19363 15623 19369
rect 15565 19329 15577 19363
rect 15611 19329 15623 19363
rect 15565 19323 15623 19329
rect 17037 19363 17095 19369
rect 17037 19329 17049 19363
rect 17083 19329 17095 19363
rect 17037 19323 17095 19329
rect 18782 19320 18788 19372
rect 18840 19320 18846 19372
rect 19518 19320 19524 19372
rect 19576 19360 19582 19372
rect 22094 19360 22100 19372
rect 19576 19332 22100 19360
rect 19576 19320 19582 19332
rect 22094 19320 22100 19332
rect 22152 19320 22158 19372
rect 22373 19363 22431 19369
rect 22373 19329 22385 19363
rect 22419 19360 22431 19363
rect 23658 19360 23664 19372
rect 22419 19332 23664 19360
rect 22419 19329 22431 19332
rect 22373 19323 22431 19329
rect 23658 19320 23664 19332
rect 23716 19320 23722 19372
rect 24857 19363 24915 19369
rect 24857 19329 24869 19363
rect 24903 19360 24915 19363
rect 25130 19360 25136 19372
rect 24903 19332 25136 19360
rect 24903 19329 24915 19332
rect 24857 19323 24915 19329
rect 25130 19320 25136 19332
rect 25188 19320 25194 19372
rect 25501 19363 25559 19369
rect 25501 19329 25513 19363
rect 25547 19360 25559 19363
rect 26068 19360 26096 19400
rect 25547 19332 26096 19360
rect 25547 19329 25559 19332
rect 25501 19323 25559 19329
rect 26142 19320 26148 19372
rect 26200 19320 26206 19372
rect 26252 19360 26280 19400
rect 27141 19397 27153 19431
rect 27141 19391 27160 19397
rect 27154 19388 27160 19391
rect 27212 19388 27218 19440
rect 27341 19431 27399 19437
rect 27341 19397 27353 19431
rect 27387 19428 27399 19431
rect 27798 19428 27804 19440
rect 27387 19400 27804 19428
rect 27387 19397 27399 19400
rect 27341 19391 27399 19397
rect 27798 19388 27804 19400
rect 27856 19388 27862 19440
rect 30190 19388 30196 19440
rect 30248 19428 30254 19440
rect 34149 19431 34207 19437
rect 30248 19400 30512 19428
rect 30248 19388 30254 19400
rect 27430 19360 27436 19372
rect 26252 19332 27436 19360
rect 27430 19320 27436 19332
rect 27488 19320 27494 19372
rect 28353 19363 28411 19369
rect 28353 19329 28365 19363
rect 28399 19360 28411 19363
rect 28626 19360 28632 19372
rect 28399 19332 28632 19360
rect 28399 19329 28411 19332
rect 28353 19323 28411 19329
rect 28626 19320 28632 19332
rect 28684 19320 28690 19372
rect 30484 19369 30512 19400
rect 34149 19397 34161 19431
rect 34195 19428 34207 19431
rect 34977 19431 35035 19437
rect 34977 19428 34989 19431
rect 34195 19400 34989 19428
rect 34195 19397 34207 19400
rect 34149 19391 34207 19397
rect 34977 19397 34989 19400
rect 35023 19397 35035 19431
rect 35176 19428 35204 19456
rect 35176 19400 35664 19428
rect 34977 19391 35035 19397
rect 30469 19363 30527 19369
rect 30469 19329 30481 19363
rect 30515 19329 30527 19363
rect 30469 19323 30527 19329
rect 30742 19320 30748 19372
rect 30800 19360 30806 19372
rect 31294 19360 31300 19372
rect 30800 19332 31300 19360
rect 30800 19320 30806 19332
rect 31294 19320 31300 19332
rect 31352 19360 31358 19372
rect 31389 19363 31447 19369
rect 31389 19360 31401 19363
rect 31352 19332 31401 19360
rect 31352 19320 31358 19332
rect 31389 19329 31401 19332
rect 31435 19329 31447 19363
rect 31389 19323 31447 19329
rect 31662 19320 31668 19372
rect 31720 19320 31726 19372
rect 33410 19320 33416 19372
rect 33468 19360 33474 19372
rect 33781 19363 33839 19369
rect 33781 19360 33793 19363
rect 33468 19332 33793 19360
rect 33468 19320 33474 19332
rect 33781 19329 33793 19332
rect 33827 19329 33839 19363
rect 33781 19323 33839 19329
rect 33870 19320 33876 19372
rect 33928 19360 33934 19372
rect 33965 19363 34023 19369
rect 33965 19360 33977 19363
rect 33928 19332 33977 19360
rect 33928 19320 33934 19332
rect 33965 19329 33977 19332
rect 34011 19329 34023 19363
rect 33965 19323 34023 19329
rect 34422 19320 34428 19372
rect 34480 19320 34486 19372
rect 34606 19320 34612 19372
rect 34664 19320 34670 19372
rect 35434 19360 35440 19372
rect 34716 19332 35440 19360
rect 14550 19292 14556 19304
rect 13740 19264 14556 19292
rect 12820 19233 12848 19264
rect 14550 19252 14556 19264
rect 14608 19252 14614 19304
rect 17313 19295 17371 19301
rect 17313 19261 17325 19295
rect 17359 19292 17371 19295
rect 17402 19292 17408 19304
rect 17359 19264 17408 19292
rect 17359 19261 17371 19264
rect 17313 19255 17371 19261
rect 17402 19252 17408 19264
rect 17460 19252 17466 19304
rect 22649 19295 22707 19301
rect 22649 19292 22661 19295
rect 18432 19264 22661 19292
rect 18432 19236 18460 19264
rect 22649 19261 22661 19264
rect 22695 19292 22707 19295
rect 24578 19292 24584 19304
rect 22695 19264 24584 19292
rect 22695 19261 22707 19264
rect 22649 19255 22707 19261
rect 24578 19252 24584 19264
rect 24636 19252 24642 19304
rect 26326 19292 26332 19304
rect 24688 19264 26332 19292
rect 12253 19227 12311 19233
rect 12253 19193 12265 19227
rect 12299 19193 12311 19227
rect 12253 19187 12311 19193
rect 12805 19227 12863 19233
rect 12805 19193 12817 19227
rect 12851 19193 12863 19227
rect 12805 19187 12863 19193
rect 15010 19184 15016 19236
rect 15068 19224 15074 19236
rect 16666 19224 16672 19236
rect 15068 19196 16672 19224
rect 15068 19184 15074 19196
rect 16666 19184 16672 19196
rect 16724 19184 16730 19236
rect 18414 19184 18420 19236
rect 18472 19184 18478 19236
rect 22278 19184 22284 19236
rect 22336 19224 22342 19236
rect 24688 19224 24716 19264
rect 26326 19252 26332 19264
rect 26384 19252 26390 19304
rect 26418 19252 26424 19304
rect 26476 19292 26482 19304
rect 26694 19292 26700 19304
rect 26476 19264 26700 19292
rect 26476 19252 26482 19264
rect 26694 19252 26700 19264
rect 26752 19292 26758 19304
rect 28537 19295 28595 19301
rect 28537 19292 28549 19295
rect 26752 19264 28549 19292
rect 26752 19252 26758 19264
rect 28537 19261 28549 19264
rect 28583 19261 28595 19295
rect 28537 19255 28595 19261
rect 31849 19295 31907 19301
rect 31849 19261 31861 19295
rect 31895 19292 31907 19295
rect 34716 19292 34744 19332
rect 35434 19320 35440 19332
rect 35492 19320 35498 19372
rect 35636 19369 35664 19400
rect 35621 19363 35679 19369
rect 35621 19329 35633 19363
rect 35667 19329 35679 19363
rect 35621 19323 35679 19329
rect 37921 19363 37979 19369
rect 37921 19329 37933 19363
rect 37967 19360 37979 19363
rect 38286 19360 38292 19372
rect 37967 19332 38292 19360
rect 37967 19329 37979 19332
rect 37921 19323 37979 19329
rect 38286 19320 38292 19332
rect 38344 19320 38350 19372
rect 31895 19264 34744 19292
rect 34793 19295 34851 19301
rect 31895 19261 31907 19264
rect 31849 19255 31907 19261
rect 34793 19261 34805 19295
rect 34839 19292 34851 19295
rect 35986 19292 35992 19304
rect 34839 19264 35992 19292
rect 34839 19261 34851 19264
rect 34793 19255 34851 19261
rect 35986 19252 35992 19264
rect 36044 19252 36050 19304
rect 22336 19196 24716 19224
rect 26068 19196 27200 19224
rect 22336 19184 22342 19196
rect 26068 19168 26096 19196
rect 12342 19156 12348 19168
rect 12084 19128 12348 19156
rect 12342 19116 12348 19128
rect 12400 19116 12406 19168
rect 12526 19116 12532 19168
rect 12584 19156 12590 19168
rect 12621 19159 12679 19165
rect 12621 19156 12633 19159
rect 12584 19128 12633 19156
rect 12584 19116 12590 19128
rect 12621 19125 12633 19128
rect 12667 19156 12679 19159
rect 13081 19159 13139 19165
rect 13081 19156 13093 19159
rect 12667 19128 13093 19156
rect 12667 19125 12679 19128
rect 12621 19119 12679 19125
rect 13081 19125 13093 19128
rect 13127 19125 13139 19159
rect 13081 19119 13139 19125
rect 13906 19116 13912 19168
rect 13964 19116 13970 19168
rect 14366 19116 14372 19168
rect 14424 19156 14430 19168
rect 14645 19159 14703 19165
rect 14645 19156 14657 19159
rect 14424 19128 14657 19156
rect 14424 19116 14430 19128
rect 14645 19125 14657 19128
rect 14691 19125 14703 19159
rect 14645 19119 14703 19125
rect 14734 19116 14740 19168
rect 14792 19156 14798 19168
rect 18966 19156 18972 19168
rect 14792 19128 18972 19156
rect 14792 19116 14798 19128
rect 18966 19116 18972 19128
rect 19024 19116 19030 19168
rect 19242 19116 19248 19168
rect 19300 19156 19306 19168
rect 20898 19156 20904 19168
rect 19300 19128 20904 19156
rect 19300 19116 19306 19128
rect 20898 19116 20904 19128
rect 20956 19116 20962 19168
rect 24578 19116 24584 19168
rect 24636 19156 24642 19168
rect 25314 19156 25320 19168
rect 24636 19128 25320 19156
rect 24636 19116 24642 19128
rect 25314 19116 25320 19128
rect 25372 19116 25378 19168
rect 25682 19116 25688 19168
rect 25740 19156 25746 19168
rect 25961 19159 26019 19165
rect 25961 19156 25973 19159
rect 25740 19128 25973 19156
rect 25740 19116 25746 19128
rect 25961 19125 25973 19128
rect 26007 19125 26019 19159
rect 25961 19119 26019 19125
rect 26050 19116 26056 19168
rect 26108 19116 26114 19168
rect 26234 19116 26240 19168
rect 26292 19156 26298 19168
rect 27172 19165 27200 19196
rect 26329 19159 26387 19165
rect 26329 19156 26341 19159
rect 26292 19128 26341 19156
rect 26292 19116 26298 19128
rect 26329 19125 26341 19128
rect 26375 19125 26387 19159
rect 26329 19119 26387 19125
rect 27157 19159 27215 19165
rect 27157 19125 27169 19159
rect 27203 19125 27215 19159
rect 27157 19119 27215 19125
rect 37734 19116 37740 19168
rect 37792 19116 37798 19168
rect 1104 19066 38272 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38272 19066
rect 1104 18992 38272 19014
rect 5902 18952 5908 18964
rect 1688 18924 5908 18952
rect 1688 18825 1716 18924
rect 5902 18912 5908 18924
rect 5960 18912 5966 18964
rect 8386 18952 8392 18964
rect 6012 18924 8392 18952
rect 6012 18884 6040 18924
rect 8386 18912 8392 18924
rect 8444 18912 8450 18964
rect 9585 18955 9643 18961
rect 9585 18921 9597 18955
rect 9631 18952 9643 18955
rect 9674 18952 9680 18964
rect 9631 18924 9680 18952
rect 9631 18921 9643 18924
rect 9585 18915 9643 18921
rect 9674 18912 9680 18924
rect 9732 18912 9738 18964
rect 9766 18912 9772 18964
rect 9824 18912 9830 18964
rect 11146 18912 11152 18964
rect 11204 18952 11210 18964
rect 11606 18952 11612 18964
rect 11204 18924 11612 18952
rect 11204 18912 11210 18924
rect 11606 18912 11612 18924
rect 11664 18952 11670 18964
rect 11974 18952 11980 18964
rect 11664 18924 11980 18952
rect 11664 18912 11670 18924
rect 11974 18912 11980 18924
rect 12032 18952 12038 18964
rect 12713 18955 12771 18961
rect 12713 18952 12725 18955
rect 12032 18924 12725 18952
rect 12032 18912 12038 18924
rect 12713 18921 12725 18924
rect 12759 18952 12771 18955
rect 12759 18924 13676 18952
rect 12759 18921 12771 18924
rect 12713 18915 12771 18921
rect 4264 18856 6040 18884
rect 1673 18819 1731 18825
rect 1673 18785 1685 18819
rect 1719 18785 1731 18819
rect 1673 18779 1731 18785
rect 3602 18776 3608 18828
rect 3660 18816 3666 18828
rect 4264 18825 4292 18856
rect 8202 18844 8208 18896
rect 8260 18884 8266 18896
rect 8260 18856 8432 18884
rect 8260 18844 8266 18856
rect 4249 18819 4307 18825
rect 4249 18816 4261 18819
rect 3660 18788 4261 18816
rect 3660 18776 3666 18788
rect 4249 18785 4261 18788
rect 4295 18785 4307 18819
rect 4249 18779 4307 18785
rect 4433 18819 4491 18825
rect 4433 18785 4445 18819
rect 4479 18816 4491 18819
rect 5350 18816 5356 18828
rect 4479 18788 5356 18816
rect 4479 18785 4491 18788
rect 4433 18779 4491 18785
rect 5350 18776 5356 18788
rect 5408 18776 5414 18828
rect 934 18708 940 18760
rect 992 18748 998 18760
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 992 18720 1409 18748
rect 992 18708 998 18720
rect 1397 18717 1409 18720
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 2501 18751 2559 18757
rect 2501 18717 2513 18751
rect 2547 18748 2559 18751
rect 4157 18751 4215 18757
rect 2547 18720 2774 18748
rect 2547 18717 2559 18720
rect 2501 18711 2559 18717
rect 2038 18572 2044 18624
rect 2096 18612 2102 18624
rect 2317 18615 2375 18621
rect 2317 18612 2329 18615
rect 2096 18584 2329 18612
rect 2096 18572 2102 18584
rect 2317 18581 2329 18584
rect 2363 18581 2375 18615
rect 2746 18612 2774 18720
rect 4157 18717 4169 18751
rect 4203 18748 4215 18751
rect 5442 18748 5448 18760
rect 4203 18720 5448 18748
rect 4203 18717 4215 18720
rect 4157 18711 4215 18717
rect 5442 18708 5448 18720
rect 5500 18708 5506 18760
rect 5813 18751 5871 18757
rect 5813 18717 5825 18751
rect 5859 18748 5871 18751
rect 6362 18748 6368 18760
rect 5859 18720 6368 18748
rect 5859 18717 5871 18720
rect 5813 18711 5871 18717
rect 6362 18708 6368 18720
rect 6420 18708 6426 18760
rect 8404 18757 8432 18856
rect 8481 18819 8539 18825
rect 8481 18785 8493 18819
rect 8527 18816 8539 18819
rect 9784 18816 9812 18912
rect 10870 18884 10876 18896
rect 8527 18788 9812 18816
rect 9968 18856 10876 18884
rect 8527 18785 8539 18788
rect 8481 18779 8539 18785
rect 9324 18757 9352 18788
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18717 8447 18751
rect 8389 18711 8447 18717
rect 9309 18751 9367 18757
rect 9309 18717 9321 18751
rect 9355 18717 9367 18751
rect 9309 18711 9367 18717
rect 9490 18708 9496 18760
rect 9548 18708 9554 18760
rect 9582 18708 9588 18760
rect 9640 18748 9646 18760
rect 9769 18751 9827 18757
rect 9769 18748 9781 18751
rect 9640 18720 9781 18748
rect 9640 18708 9646 18720
rect 9769 18717 9781 18720
rect 9815 18717 9827 18751
rect 9769 18711 9827 18717
rect 7742 18640 7748 18692
rect 7800 18680 7806 18692
rect 7837 18683 7895 18689
rect 7837 18680 7849 18683
rect 7800 18652 7849 18680
rect 7800 18640 7806 18652
rect 7837 18649 7849 18652
rect 7883 18649 7895 18683
rect 9968 18680 9996 18856
rect 10870 18844 10876 18856
rect 10928 18844 10934 18896
rect 11054 18844 11060 18896
rect 11112 18884 11118 18896
rect 13538 18884 13544 18896
rect 11112 18856 13544 18884
rect 11112 18844 11118 18856
rect 13538 18844 13544 18856
rect 13596 18844 13602 18896
rect 13648 18884 13676 18924
rect 13722 18912 13728 18964
rect 13780 18912 13786 18964
rect 13906 18912 13912 18964
rect 13964 18952 13970 18964
rect 20714 18952 20720 18964
rect 13964 18924 20720 18952
rect 13964 18912 13970 18924
rect 20714 18912 20720 18924
rect 20772 18912 20778 18964
rect 22094 18912 22100 18964
rect 22152 18952 22158 18964
rect 24397 18955 24455 18961
rect 22152 18924 24348 18952
rect 22152 18912 22158 18924
rect 15378 18884 15384 18896
rect 13648 18856 15384 18884
rect 15378 18844 15384 18856
rect 15436 18844 15442 18896
rect 16206 18844 16212 18896
rect 16264 18844 16270 18896
rect 18414 18844 18420 18896
rect 18472 18884 18478 18896
rect 18472 18856 18920 18884
rect 18472 18844 18478 18856
rect 12342 18816 12348 18828
rect 10060 18788 11836 18816
rect 10060 18757 10088 18788
rect 10045 18751 10103 18757
rect 10045 18717 10057 18751
rect 10091 18717 10103 18751
rect 10045 18711 10103 18717
rect 10144 18751 10202 18757
rect 10144 18717 10156 18751
rect 10190 18717 10202 18751
rect 10144 18711 10202 18717
rect 10291 18751 10349 18757
rect 10291 18717 10303 18751
rect 10337 18748 10349 18751
rect 10410 18748 10416 18760
rect 10337 18720 10416 18748
rect 10337 18717 10349 18720
rect 10291 18711 10349 18717
rect 7837 18643 7895 18649
rect 8312 18652 9996 18680
rect 3789 18615 3847 18621
rect 3789 18612 3801 18615
rect 2746 18584 3801 18612
rect 2317 18575 2375 18581
rect 3789 18581 3801 18584
rect 3835 18581 3847 18615
rect 3789 18575 3847 18581
rect 5626 18572 5632 18624
rect 5684 18572 5690 18624
rect 8312 18621 8340 18652
rect 8297 18615 8355 18621
rect 8297 18581 8309 18615
rect 8343 18581 8355 18615
rect 8297 18575 8355 18581
rect 9493 18615 9551 18621
rect 9493 18581 9505 18615
rect 9539 18612 9551 18615
rect 9953 18615 10011 18621
rect 9953 18612 9965 18615
rect 9539 18584 9965 18612
rect 9539 18581 9551 18584
rect 9493 18575 9551 18581
rect 9953 18581 9965 18584
rect 9999 18581 10011 18615
rect 9953 18575 10011 18581
rect 10042 18572 10048 18624
rect 10100 18612 10106 18624
rect 10152 18612 10180 18711
rect 10410 18708 10416 18720
rect 10468 18708 10474 18760
rect 10520 18680 10548 18788
rect 10336 18652 10548 18680
rect 10336 18624 10364 18652
rect 10100 18584 10180 18612
rect 10100 18572 10106 18584
rect 10318 18572 10324 18624
rect 10376 18572 10382 18624
rect 10502 18572 10508 18624
rect 10560 18572 10566 18624
rect 11808 18612 11836 18788
rect 12176 18788 12348 18816
rect 11882 18708 11888 18760
rect 11940 18708 11946 18760
rect 12176 18757 12204 18788
rect 12342 18776 12348 18788
rect 12400 18816 12406 18828
rect 12400 18788 12664 18816
rect 12400 18776 12406 18788
rect 12636 18760 12664 18788
rect 12894 18776 12900 18828
rect 12952 18776 12958 18828
rect 12161 18751 12219 18757
rect 12161 18717 12173 18751
rect 12207 18717 12219 18751
rect 12161 18711 12219 18717
rect 12529 18751 12587 18757
rect 12529 18717 12541 18751
rect 12575 18717 12587 18751
rect 12529 18711 12587 18717
rect 11900 18680 11928 18708
rect 12544 18680 12572 18711
rect 12618 18708 12624 18760
rect 12676 18708 12682 18760
rect 12802 18708 12808 18760
rect 12860 18708 12866 18760
rect 13081 18751 13139 18757
rect 13081 18717 13093 18751
rect 13127 18717 13139 18751
rect 13081 18711 13139 18717
rect 11900 18652 12572 18680
rect 13096 18680 13124 18711
rect 13170 18708 13176 18760
rect 13228 18708 13234 18760
rect 13556 18689 13584 18844
rect 14829 18819 14887 18825
rect 13832 18788 14596 18816
rect 13630 18708 13636 18760
rect 13688 18708 13694 18760
rect 13541 18683 13599 18689
rect 13096 18652 13492 18680
rect 12345 18615 12403 18621
rect 12345 18612 12357 18615
rect 11808 18584 12357 18612
rect 12345 18581 12357 18584
rect 12391 18612 12403 18615
rect 13096 18612 13124 18652
rect 12391 18584 13124 18612
rect 12391 18581 12403 18584
rect 12345 18575 12403 18581
rect 13354 18572 13360 18624
rect 13412 18572 13418 18624
rect 13464 18612 13492 18652
rect 13541 18649 13553 18683
rect 13587 18649 13599 18683
rect 13648 18680 13676 18708
rect 13741 18683 13799 18689
rect 13741 18680 13753 18683
rect 13648 18652 13753 18680
rect 13541 18643 13599 18649
rect 13741 18649 13753 18652
rect 13787 18649 13799 18683
rect 13741 18643 13799 18649
rect 13832 18612 13860 18788
rect 14366 18708 14372 18760
rect 14424 18708 14430 18760
rect 14568 18757 14596 18788
rect 14829 18785 14841 18819
rect 14875 18785 14887 18819
rect 16224 18816 16252 18844
rect 14829 18779 14887 18785
rect 15764 18788 16252 18816
rect 14553 18751 14611 18757
rect 14553 18717 14565 18751
rect 14599 18717 14611 18751
rect 14553 18711 14611 18717
rect 14182 18640 14188 18692
rect 14240 18680 14246 18692
rect 14844 18680 14872 18779
rect 14921 18751 14979 18757
rect 14921 18717 14933 18751
rect 14967 18717 14979 18751
rect 14921 18711 14979 18717
rect 14240 18652 14872 18680
rect 14240 18640 14246 18652
rect 13464 18584 13860 18612
rect 13906 18572 13912 18624
rect 13964 18572 13970 18624
rect 14550 18572 14556 18624
rect 14608 18612 14614 18624
rect 14936 18612 14964 18711
rect 15286 18708 15292 18760
rect 15344 18708 15350 18760
rect 15764 18757 15792 18788
rect 16666 18776 16672 18828
rect 16724 18816 16730 18828
rect 18693 18819 18751 18825
rect 18693 18816 18705 18819
rect 16724 18788 18705 18816
rect 16724 18776 16730 18788
rect 18693 18785 18705 18788
rect 18739 18785 18751 18819
rect 18693 18779 18751 18785
rect 15749 18751 15807 18757
rect 15749 18717 15761 18751
rect 15795 18717 15807 18751
rect 15749 18711 15807 18717
rect 15838 18708 15844 18760
rect 15896 18748 15902 18760
rect 16301 18751 16359 18757
rect 16301 18748 16313 18751
rect 15896 18720 16313 18748
rect 15896 18708 15902 18720
rect 16301 18717 16313 18720
rect 16347 18717 16359 18751
rect 16301 18711 16359 18717
rect 18598 18708 18604 18760
rect 18656 18708 18662 18760
rect 18892 18757 18920 18856
rect 21082 18844 21088 18896
rect 21140 18884 21146 18896
rect 24320 18884 24348 18924
rect 24397 18921 24409 18955
rect 24443 18952 24455 18955
rect 24486 18952 24492 18964
rect 24443 18924 24492 18952
rect 24443 18921 24455 18924
rect 24397 18915 24455 18921
rect 24486 18912 24492 18924
rect 24544 18912 24550 18964
rect 24670 18912 24676 18964
rect 24728 18952 24734 18964
rect 29730 18952 29736 18964
rect 24728 18924 29736 18952
rect 24728 18912 24734 18924
rect 29730 18912 29736 18924
rect 29788 18912 29794 18964
rect 33410 18912 33416 18964
rect 33468 18952 33474 18964
rect 33873 18955 33931 18961
rect 33873 18952 33885 18955
rect 33468 18924 33885 18952
rect 33468 18912 33474 18924
rect 33873 18921 33885 18924
rect 33919 18921 33931 18955
rect 33873 18915 33931 18921
rect 34241 18955 34299 18961
rect 34241 18921 34253 18955
rect 34287 18952 34299 18955
rect 34330 18952 34336 18964
rect 34287 18924 34336 18952
rect 34287 18921 34299 18924
rect 34241 18915 34299 18921
rect 34330 18912 34336 18924
rect 34388 18912 34394 18964
rect 34425 18955 34483 18961
rect 34425 18921 34437 18955
rect 34471 18952 34483 18955
rect 35342 18952 35348 18964
rect 34471 18924 35348 18952
rect 34471 18921 34483 18924
rect 34425 18915 34483 18921
rect 35342 18912 35348 18924
rect 35400 18912 35406 18964
rect 37553 18955 37611 18961
rect 37553 18921 37565 18955
rect 37599 18952 37611 18955
rect 37642 18952 37648 18964
rect 37599 18924 37648 18952
rect 37599 18921 37611 18924
rect 37553 18915 37611 18921
rect 37642 18912 37648 18924
rect 37700 18912 37706 18964
rect 30650 18884 30656 18896
rect 21140 18856 23152 18884
rect 24320 18856 30656 18884
rect 21140 18844 21146 18856
rect 19334 18776 19340 18828
rect 19392 18776 19398 18828
rect 20530 18776 20536 18828
rect 20588 18816 20594 18828
rect 21913 18819 21971 18825
rect 21913 18816 21925 18819
rect 20588 18788 21925 18816
rect 20588 18776 20594 18788
rect 21913 18785 21925 18788
rect 21959 18816 21971 18819
rect 21959 18788 22600 18816
rect 21959 18785 21971 18788
rect 21913 18779 21971 18785
rect 18877 18751 18935 18757
rect 18877 18717 18889 18751
rect 18923 18717 18935 18751
rect 19352 18748 19380 18776
rect 19429 18751 19487 18757
rect 19429 18748 19441 18751
rect 19352 18720 19441 18748
rect 18877 18711 18935 18717
rect 19429 18717 19441 18720
rect 19475 18717 19487 18751
rect 19429 18711 19487 18717
rect 19521 18751 19579 18757
rect 19521 18717 19533 18751
rect 19567 18748 19579 18751
rect 19705 18751 19763 18757
rect 19705 18748 19717 18751
rect 19567 18720 19717 18748
rect 19567 18717 19579 18720
rect 19521 18711 19579 18717
rect 19705 18717 19717 18720
rect 19751 18717 19763 18751
rect 19705 18711 19763 18717
rect 21542 18708 21548 18760
rect 21600 18708 21606 18760
rect 22094 18708 22100 18760
rect 22152 18708 22158 18760
rect 22278 18708 22284 18760
rect 22336 18708 22342 18760
rect 22370 18708 22376 18760
rect 22428 18708 22434 18760
rect 22462 18708 22468 18760
rect 22520 18708 22526 18760
rect 22572 18748 22600 18788
rect 22646 18776 22652 18828
rect 22704 18816 22710 18828
rect 23017 18819 23075 18825
rect 23017 18816 23029 18819
rect 22704 18788 23029 18816
rect 22704 18776 22710 18788
rect 23017 18785 23029 18788
rect 23063 18785 23075 18819
rect 23124 18816 23152 18856
rect 30650 18844 30656 18856
rect 30708 18844 30714 18896
rect 33502 18884 33508 18896
rect 32600 18856 33508 18884
rect 23124 18788 24808 18816
rect 23017 18779 23075 18785
rect 23842 18748 23848 18760
rect 22572 18720 23848 18748
rect 23842 18708 23848 18720
rect 23900 18708 23906 18760
rect 24670 18708 24676 18760
rect 24728 18708 24734 18760
rect 24780 18757 24808 18788
rect 25130 18776 25136 18828
rect 25188 18816 25194 18828
rect 30098 18816 30104 18828
rect 25188 18788 30104 18816
rect 25188 18776 25194 18788
rect 30098 18776 30104 18788
rect 30156 18816 30162 18828
rect 32600 18816 32628 18856
rect 33502 18844 33508 18856
rect 33560 18844 33566 18896
rect 33778 18844 33784 18896
rect 33836 18844 33842 18896
rect 34054 18844 34060 18896
rect 34112 18884 34118 18896
rect 34606 18884 34612 18896
rect 34112 18856 34612 18884
rect 34112 18844 34118 18856
rect 34606 18844 34612 18856
rect 34664 18844 34670 18896
rect 33686 18816 33692 18828
rect 30156 18788 32628 18816
rect 30156 18776 30162 18788
rect 24765 18751 24823 18757
rect 24765 18717 24777 18751
rect 24811 18717 24823 18751
rect 24765 18711 24823 18717
rect 24857 18751 24915 18757
rect 24857 18717 24869 18751
rect 24903 18717 24915 18751
rect 24857 18711 24915 18717
rect 17129 18683 17187 18689
rect 17129 18649 17141 18683
rect 17175 18680 17187 18683
rect 17586 18680 17592 18692
rect 17175 18652 17592 18680
rect 17175 18649 17187 18652
rect 17129 18643 17187 18649
rect 17586 18640 17592 18652
rect 17644 18640 17650 18692
rect 19978 18640 19984 18692
rect 20036 18640 20042 18692
rect 22296 18680 22324 18708
rect 21206 18652 22324 18680
rect 14608 18584 14964 18612
rect 14608 18572 14614 18584
rect 16114 18572 16120 18624
rect 16172 18612 16178 18624
rect 18322 18612 18328 18624
rect 16172 18584 18328 18612
rect 16172 18572 16178 18584
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 19058 18572 19064 18624
rect 19116 18572 19122 18624
rect 21266 18572 21272 18624
rect 21324 18612 21330 18624
rect 21453 18615 21511 18621
rect 21453 18612 21465 18615
rect 21324 18584 21465 18612
rect 21324 18572 21330 18584
rect 21453 18581 21465 18584
rect 21499 18581 21511 18615
rect 21453 18575 21511 18581
rect 23014 18572 23020 18624
rect 23072 18612 23078 18624
rect 24872 18612 24900 18711
rect 25038 18708 25044 18760
rect 25096 18708 25102 18760
rect 25314 18708 25320 18760
rect 25372 18748 25378 18760
rect 28721 18751 28779 18757
rect 28721 18748 28733 18751
rect 25372 18720 28733 18748
rect 25372 18708 25378 18720
rect 28721 18717 28733 18720
rect 28767 18748 28779 18751
rect 28810 18748 28816 18760
rect 28767 18720 28816 18748
rect 28767 18717 28779 18720
rect 28721 18711 28779 18717
rect 28810 18708 28816 18720
rect 28868 18708 28874 18760
rect 28997 18751 29055 18757
rect 28997 18717 29009 18751
rect 29043 18717 29055 18751
rect 28997 18711 29055 18717
rect 29365 18751 29423 18757
rect 29365 18717 29377 18751
rect 29411 18748 29423 18751
rect 29914 18748 29920 18760
rect 29411 18720 29920 18748
rect 29411 18717 29423 18720
rect 29365 18711 29423 18717
rect 29012 18680 29040 18711
rect 29914 18708 29920 18720
rect 29972 18708 29978 18760
rect 32398 18708 32404 18760
rect 32456 18708 32462 18760
rect 32600 18757 32628 18788
rect 33152 18788 33692 18816
rect 33152 18757 33180 18788
rect 33686 18776 33692 18788
rect 33744 18816 33750 18828
rect 33744 18788 34192 18816
rect 33744 18776 33750 18788
rect 32585 18751 32643 18757
rect 32585 18717 32597 18751
rect 32631 18717 32643 18751
rect 32585 18711 32643 18717
rect 33137 18751 33195 18757
rect 33137 18717 33149 18751
rect 33183 18717 33195 18751
rect 33321 18751 33379 18757
rect 33321 18748 33333 18751
rect 33137 18711 33195 18717
rect 33244 18720 33333 18748
rect 33244 18692 33272 18720
rect 33321 18717 33333 18720
rect 33367 18717 33379 18751
rect 33321 18711 33379 18717
rect 33410 18708 33416 18760
rect 33468 18708 33474 18760
rect 33502 18708 33508 18760
rect 33560 18748 33566 18760
rect 34054 18748 34060 18760
rect 33560 18720 34060 18748
rect 33560 18708 33566 18720
rect 34054 18708 34060 18720
rect 34112 18708 34118 18760
rect 34164 18745 34192 18788
rect 34241 18751 34299 18757
rect 34241 18745 34253 18751
rect 34164 18717 34253 18745
rect 34287 18745 34299 18751
rect 34333 18751 34391 18757
rect 34333 18745 34345 18751
rect 34287 18717 34345 18745
rect 34379 18717 34391 18751
rect 34241 18711 34299 18717
rect 34333 18711 34391 18717
rect 34517 18751 34575 18757
rect 34517 18717 34529 18751
rect 34563 18717 34575 18751
rect 34517 18711 34575 18717
rect 27448 18652 29040 18680
rect 32493 18683 32551 18689
rect 27448 18624 27476 18652
rect 32493 18649 32505 18683
rect 32539 18680 32551 18683
rect 33226 18680 33232 18692
rect 32539 18652 33232 18680
rect 32539 18649 32551 18652
rect 32493 18643 32551 18649
rect 33226 18640 33232 18652
rect 33284 18680 33290 18692
rect 34532 18680 34560 18711
rect 37366 18708 37372 18760
rect 37424 18708 37430 18760
rect 33284 18652 34560 18680
rect 33284 18640 33290 18652
rect 23072 18584 24900 18612
rect 23072 18572 23078 18584
rect 27430 18572 27436 18624
rect 27488 18572 27494 18624
rect 28629 18615 28687 18621
rect 28629 18581 28641 18615
rect 28675 18612 28687 18615
rect 28718 18612 28724 18624
rect 28675 18584 28724 18612
rect 28675 18581 28687 18584
rect 28629 18575 28687 18581
rect 28718 18572 28724 18584
rect 28776 18572 28782 18624
rect 28902 18572 28908 18624
rect 28960 18572 28966 18624
rect 29270 18572 29276 18624
rect 29328 18572 29334 18624
rect 1104 18522 38272 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 38272 18522
rect 1104 18448 38272 18470
rect 2038 18408 2044 18420
rect 1872 18380 2044 18408
rect 1872 18349 1900 18380
rect 2038 18368 2044 18380
rect 2096 18368 2102 18420
rect 3602 18368 3608 18420
rect 3660 18368 3666 18420
rect 4065 18411 4123 18417
rect 4065 18377 4077 18411
rect 4111 18408 4123 18411
rect 4706 18408 4712 18420
rect 4111 18380 4712 18408
rect 4111 18377 4123 18380
rect 4065 18371 4123 18377
rect 4706 18368 4712 18380
rect 4764 18368 4770 18420
rect 5445 18411 5503 18417
rect 5445 18377 5457 18411
rect 5491 18408 5503 18411
rect 5534 18408 5540 18420
rect 5491 18380 5540 18408
rect 5491 18377 5503 18380
rect 5445 18371 5503 18377
rect 5534 18368 5540 18380
rect 5592 18368 5598 18420
rect 10502 18408 10508 18420
rect 10428 18380 10508 18408
rect 1857 18343 1915 18349
rect 1857 18309 1869 18343
rect 1903 18309 1915 18343
rect 1857 18303 1915 18309
rect 1394 18232 1400 18284
rect 1452 18272 1458 18284
rect 1581 18275 1639 18281
rect 1581 18272 1593 18275
rect 1452 18244 1593 18272
rect 1452 18232 1458 18244
rect 1581 18241 1593 18244
rect 1627 18241 1639 18275
rect 3234 18272 3240 18284
rect 2990 18244 3240 18272
rect 1581 18235 1639 18241
rect 3234 18232 3240 18244
rect 3292 18232 3298 18284
rect 3620 18281 3648 18368
rect 8846 18340 8852 18352
rect 8786 18312 8852 18340
rect 8846 18300 8852 18312
rect 8904 18340 8910 18352
rect 8904 18312 9674 18340
rect 8904 18300 8910 18312
rect 3605 18275 3663 18281
rect 3605 18241 3617 18275
rect 3651 18241 3663 18275
rect 3605 18235 3663 18241
rect 5368 18244 5672 18272
rect 5368 18216 5396 18244
rect 4157 18207 4215 18213
rect 4157 18173 4169 18207
rect 4203 18173 4215 18207
rect 4157 18167 4215 18173
rect 4341 18207 4399 18213
rect 4341 18173 4353 18207
rect 4387 18204 4399 18207
rect 5350 18204 5356 18216
rect 4387 18176 5356 18204
rect 4387 18173 4399 18176
rect 4341 18167 4399 18173
rect 4172 18136 4200 18167
rect 5350 18164 5356 18176
rect 5408 18164 5414 18216
rect 5644 18213 5672 18244
rect 7742 18232 7748 18284
rect 7800 18272 7806 18284
rect 7837 18275 7895 18281
rect 7837 18272 7849 18275
rect 7800 18244 7849 18272
rect 7800 18232 7806 18244
rect 7837 18241 7849 18244
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 8294 18232 8300 18284
rect 8352 18272 8358 18284
rect 8389 18275 8447 18281
rect 8389 18272 8401 18275
rect 8352 18244 8401 18272
rect 8352 18232 8358 18244
rect 8389 18241 8401 18244
rect 8435 18241 8447 18275
rect 8389 18235 8447 18241
rect 5537 18207 5595 18213
rect 5537 18173 5549 18207
rect 5583 18173 5595 18207
rect 5537 18167 5595 18173
rect 5629 18207 5687 18213
rect 5629 18173 5641 18207
rect 5675 18173 5687 18207
rect 9646 18204 9674 18312
rect 10229 18275 10287 18281
rect 10229 18241 10241 18275
rect 10275 18272 10287 18275
rect 10318 18272 10324 18284
rect 10275 18244 10324 18272
rect 10275 18241 10287 18244
rect 10229 18235 10287 18241
rect 10318 18232 10324 18244
rect 10376 18232 10382 18284
rect 10428 18281 10456 18380
rect 10502 18368 10508 18380
rect 10560 18408 10566 18420
rect 13170 18408 13176 18420
rect 10560 18380 13176 18408
rect 10560 18368 10566 18380
rect 13170 18368 13176 18380
rect 13228 18368 13234 18420
rect 13906 18368 13912 18420
rect 13964 18368 13970 18420
rect 14645 18411 14703 18417
rect 14645 18377 14657 18411
rect 14691 18408 14703 18411
rect 17770 18408 17776 18420
rect 14691 18380 17776 18408
rect 14691 18377 14703 18380
rect 14645 18371 14703 18377
rect 17770 18368 17776 18380
rect 17828 18368 17834 18420
rect 19058 18368 19064 18420
rect 19116 18368 19122 18420
rect 19705 18411 19763 18417
rect 19705 18377 19717 18411
rect 19751 18408 19763 18411
rect 19978 18408 19984 18420
rect 19751 18380 19984 18408
rect 19751 18377 19763 18380
rect 19705 18371 19763 18377
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 22189 18411 22247 18417
rect 22189 18377 22201 18411
rect 22235 18408 22247 18411
rect 22462 18408 22468 18420
rect 22235 18380 22468 18408
rect 22235 18377 22247 18380
rect 22189 18371 22247 18377
rect 22462 18368 22468 18380
rect 22520 18368 22526 18420
rect 24670 18368 24676 18420
rect 24728 18408 24734 18420
rect 25409 18411 25467 18417
rect 25409 18408 25421 18411
rect 24728 18380 25421 18408
rect 24728 18368 24734 18380
rect 25409 18377 25421 18380
rect 25455 18408 25467 18411
rect 25455 18380 26012 18408
rect 25455 18377 25467 18380
rect 25409 18371 25467 18377
rect 11514 18300 11520 18352
rect 11572 18340 11578 18352
rect 13924 18340 13952 18368
rect 18601 18343 18659 18349
rect 18601 18340 18613 18343
rect 11572 18312 13860 18340
rect 13924 18312 18613 18340
rect 11572 18300 11578 18312
rect 10413 18275 10471 18281
rect 10413 18241 10425 18275
rect 10459 18241 10471 18275
rect 10413 18235 10471 18241
rect 11698 18204 11704 18216
rect 9646 18176 11704 18204
rect 5629 18167 5687 18173
rect 4798 18136 4804 18148
rect 4172 18108 4804 18136
rect 4798 18096 4804 18108
rect 4856 18096 4862 18148
rect 3694 18028 3700 18080
rect 3752 18028 3758 18080
rect 4890 18028 4896 18080
rect 4948 18068 4954 18080
rect 5077 18071 5135 18077
rect 5077 18068 5089 18071
rect 4948 18040 5089 18068
rect 4948 18028 4954 18040
rect 5077 18037 5089 18040
rect 5123 18037 5135 18071
rect 5552 18068 5580 18167
rect 11698 18164 11704 18176
rect 11756 18164 11762 18216
rect 13832 18204 13860 18312
rect 18601 18309 18613 18312
rect 18647 18309 18659 18343
rect 18601 18303 18659 18309
rect 14274 18232 14280 18284
rect 14332 18232 14338 18284
rect 14458 18232 14464 18284
rect 14516 18232 14522 18284
rect 15562 18232 15568 18284
rect 15620 18272 15626 18284
rect 15620 18244 16252 18272
rect 15620 18232 15626 18244
rect 15654 18204 15660 18216
rect 13832 18176 15660 18204
rect 15654 18164 15660 18176
rect 15712 18204 15718 18216
rect 16224 18213 16252 18244
rect 16298 18232 16304 18284
rect 16356 18232 16362 18284
rect 16574 18232 16580 18284
rect 16632 18272 16638 18284
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 16632 18244 16865 18272
rect 16632 18232 16638 18244
rect 16853 18241 16865 18244
rect 16899 18241 16911 18275
rect 16853 18235 16911 18241
rect 17221 18275 17279 18281
rect 17221 18241 17233 18275
rect 17267 18241 17279 18275
rect 17221 18235 17279 18241
rect 15841 18207 15899 18213
rect 15841 18204 15853 18207
rect 15712 18176 15853 18204
rect 15712 18164 15718 18176
rect 15841 18173 15853 18176
rect 15887 18173 15899 18207
rect 15841 18167 15899 18173
rect 16209 18207 16267 18213
rect 16209 18173 16221 18207
rect 16255 18173 16267 18207
rect 16945 18207 17003 18213
rect 16945 18204 16957 18207
rect 16209 18167 16267 18173
rect 16500 18176 16957 18204
rect 6454 18096 6460 18148
rect 6512 18136 6518 18148
rect 14734 18136 14740 18148
rect 6512 18108 14740 18136
rect 6512 18096 6518 18108
rect 14734 18096 14740 18108
rect 14792 18096 14798 18148
rect 16500 18080 16528 18176
rect 16945 18173 16957 18176
rect 16991 18173 17003 18207
rect 16945 18167 17003 18173
rect 17034 18164 17040 18216
rect 17092 18204 17098 18216
rect 17129 18207 17187 18213
rect 17129 18204 17141 18207
rect 17092 18176 17141 18204
rect 17092 18164 17098 18176
rect 17129 18173 17141 18176
rect 17175 18173 17187 18207
rect 17129 18167 17187 18173
rect 7834 18068 7840 18080
rect 5552 18040 7840 18068
rect 5077 18031 5135 18037
rect 7834 18028 7840 18040
rect 7892 18028 7898 18080
rect 10226 18028 10232 18080
rect 10284 18028 10290 18080
rect 11698 18028 11704 18080
rect 11756 18068 11762 18080
rect 14277 18071 14335 18077
rect 14277 18068 14289 18071
rect 11756 18040 14289 18068
rect 11756 18028 11762 18040
rect 14277 18037 14289 18040
rect 14323 18068 14335 18071
rect 14642 18068 14648 18080
rect 14323 18040 14648 18068
rect 14323 18037 14335 18040
rect 14277 18031 14335 18037
rect 14642 18028 14648 18040
rect 14700 18068 14706 18080
rect 15286 18068 15292 18080
rect 14700 18040 15292 18068
rect 14700 18028 14706 18040
rect 15286 18028 15292 18040
rect 15344 18028 15350 18080
rect 16482 18028 16488 18080
rect 16540 18028 16546 18080
rect 16850 18028 16856 18080
rect 16908 18068 16914 18080
rect 17236 18068 17264 18235
rect 18414 18232 18420 18284
rect 18472 18232 18478 18284
rect 19076 18272 19104 18368
rect 19334 18300 19340 18352
rect 19392 18300 19398 18352
rect 19429 18343 19487 18349
rect 19429 18309 19441 18343
rect 19475 18340 19487 18343
rect 20533 18343 20591 18349
rect 20533 18340 20545 18343
rect 19475 18312 20545 18340
rect 19475 18309 19487 18312
rect 19429 18303 19487 18309
rect 20533 18309 20545 18312
rect 20579 18309 20591 18343
rect 25984 18340 26012 18380
rect 26050 18368 26056 18420
rect 26108 18368 26114 18420
rect 28902 18368 28908 18420
rect 28960 18368 28966 18420
rect 33226 18368 33232 18420
rect 33284 18368 33290 18420
rect 33781 18411 33839 18417
rect 33781 18377 33793 18411
rect 33827 18408 33839 18411
rect 33870 18408 33876 18420
rect 33827 18380 33876 18408
rect 33827 18377 33839 18380
rect 33781 18371 33839 18377
rect 33870 18368 33876 18380
rect 33928 18368 33934 18420
rect 26602 18340 26608 18352
rect 25984 18312 26608 18340
rect 20533 18303 20591 18309
rect 26602 18300 26608 18312
rect 26660 18300 26666 18352
rect 28920 18340 28948 18368
rect 28736 18312 28948 18340
rect 33244 18340 33272 18368
rect 33244 18312 33640 18340
rect 19153 18275 19211 18281
rect 19153 18272 19165 18275
rect 19076 18244 19165 18272
rect 19153 18241 19165 18244
rect 19199 18241 19211 18275
rect 19521 18275 19579 18281
rect 19521 18272 19533 18275
rect 19153 18235 19211 18241
rect 19260 18244 19533 18272
rect 17862 18164 17868 18216
rect 17920 18164 17926 18216
rect 18432 18204 18460 18232
rect 19260 18204 19288 18244
rect 19521 18241 19533 18244
rect 19567 18241 19579 18275
rect 19521 18235 19579 18241
rect 18432 18176 19288 18204
rect 19536 18204 19564 18235
rect 20438 18232 20444 18284
rect 20496 18272 20502 18284
rect 21269 18275 21327 18281
rect 21269 18272 21281 18275
rect 20496 18244 21281 18272
rect 20496 18232 20502 18244
rect 21269 18241 21281 18244
rect 21315 18241 21327 18275
rect 21269 18235 21327 18241
rect 21358 18232 21364 18284
rect 21416 18232 21422 18284
rect 21818 18232 21824 18284
rect 21876 18232 21882 18284
rect 22005 18275 22063 18281
rect 22005 18241 22017 18275
rect 22051 18272 22063 18275
rect 23017 18275 23075 18281
rect 23017 18272 23029 18275
rect 22051 18244 23029 18272
rect 22051 18241 22063 18244
rect 22005 18235 22063 18241
rect 23017 18241 23029 18244
rect 23063 18241 23075 18275
rect 23017 18235 23075 18241
rect 20898 18204 20904 18216
rect 19536 18176 20904 18204
rect 20898 18164 20904 18176
rect 20956 18164 20962 18216
rect 21177 18207 21235 18213
rect 21177 18173 21189 18207
rect 21223 18204 21235 18207
rect 21376 18204 21404 18232
rect 22020 18204 22048 18235
rect 23842 18232 23848 18284
rect 23900 18272 23906 18284
rect 25130 18272 25136 18284
rect 23900 18244 25136 18272
rect 23900 18232 23906 18244
rect 25130 18232 25136 18244
rect 25188 18232 25194 18284
rect 25222 18232 25228 18284
rect 25280 18272 25286 18284
rect 25317 18275 25375 18281
rect 25317 18272 25329 18275
rect 25280 18244 25329 18272
rect 25280 18232 25286 18244
rect 25317 18241 25329 18244
rect 25363 18241 25375 18275
rect 25317 18235 25375 18241
rect 26970 18232 26976 18284
rect 27028 18232 27034 18284
rect 28736 18281 28764 18312
rect 28721 18275 28779 18281
rect 28721 18241 28733 18275
rect 28767 18241 28779 18275
rect 28721 18235 28779 18241
rect 21223 18176 21312 18204
rect 21376 18176 22048 18204
rect 21223 18173 21235 18176
rect 21177 18167 21235 18173
rect 18524 18108 19334 18136
rect 18524 18080 18552 18108
rect 16908 18040 17264 18068
rect 16908 18028 16914 18040
rect 18506 18028 18512 18080
rect 18564 18028 18570 18080
rect 18874 18028 18880 18080
rect 18932 18028 18938 18080
rect 19306 18068 19334 18108
rect 21284 18080 21312 18176
rect 22922 18164 22928 18216
rect 22980 18204 22986 18216
rect 23474 18204 23480 18216
rect 22980 18176 23480 18204
rect 22980 18164 22986 18176
rect 23474 18164 23480 18176
rect 23532 18204 23538 18216
rect 23532 18176 24348 18204
rect 23532 18164 23538 18176
rect 24320 18145 24348 18176
rect 24412 18176 25820 18204
rect 24305 18139 24363 18145
rect 24305 18105 24317 18139
rect 24351 18105 24363 18139
rect 24305 18099 24363 18105
rect 21082 18068 21088 18080
rect 19306 18040 21088 18068
rect 21082 18028 21088 18040
rect 21140 18028 21146 18080
rect 21266 18028 21272 18080
rect 21324 18028 21330 18080
rect 21453 18071 21511 18077
rect 21453 18037 21465 18071
rect 21499 18068 21511 18071
rect 22186 18068 22192 18080
rect 21499 18040 22192 18068
rect 21499 18037 21511 18040
rect 21453 18031 21511 18037
rect 22186 18028 22192 18040
rect 22244 18028 22250 18080
rect 23750 18028 23756 18080
rect 23808 18068 23814 18080
rect 24412 18068 24440 18176
rect 24670 18096 24676 18148
rect 24728 18136 24734 18148
rect 25792 18145 25820 18176
rect 28994 18164 29000 18216
rect 29052 18164 29058 18216
rect 30116 18204 30144 18258
rect 30374 18232 30380 18284
rect 30432 18272 30438 18284
rect 30653 18275 30711 18281
rect 30653 18272 30665 18275
rect 30432 18244 30665 18272
rect 30432 18232 30438 18244
rect 30653 18241 30665 18244
rect 30699 18272 30711 18275
rect 30699 18244 31754 18272
rect 30699 18241 30711 18244
rect 30653 18235 30711 18241
rect 31018 18204 31024 18216
rect 30116 18176 31024 18204
rect 25685 18139 25743 18145
rect 25685 18136 25697 18139
rect 24728 18108 25697 18136
rect 24728 18096 24734 18108
rect 25685 18105 25697 18108
rect 25731 18105 25743 18139
rect 25685 18099 25743 18105
rect 25777 18139 25835 18145
rect 25777 18105 25789 18139
rect 25823 18136 25835 18139
rect 28626 18136 28632 18148
rect 25823 18108 28632 18136
rect 25823 18105 25835 18108
rect 25777 18099 25835 18105
rect 28626 18096 28632 18108
rect 28684 18096 28690 18148
rect 23808 18040 24440 18068
rect 25593 18071 25651 18077
rect 23808 18028 23814 18040
rect 25593 18037 25605 18071
rect 25639 18068 25651 18071
rect 26050 18068 26056 18080
rect 25639 18040 26056 18068
rect 25639 18037 25651 18040
rect 25593 18031 25651 18037
rect 26050 18028 26056 18040
rect 26108 18028 26114 18080
rect 27154 18028 27160 18080
rect 27212 18028 27218 18080
rect 27246 18028 27252 18080
rect 27304 18068 27310 18080
rect 30116 18068 30144 18176
rect 31018 18164 31024 18176
rect 31076 18164 31082 18216
rect 31726 18136 31754 18244
rect 32214 18232 32220 18284
rect 32272 18232 32278 18284
rect 32306 18232 32312 18284
rect 32364 18232 32370 18284
rect 33321 18275 33379 18281
rect 33321 18241 33333 18275
rect 33367 18272 33379 18275
rect 33502 18272 33508 18284
rect 33367 18244 33508 18272
rect 33367 18241 33379 18244
rect 33321 18235 33379 18241
rect 33502 18232 33508 18244
rect 33560 18232 33566 18284
rect 33612 18281 33640 18312
rect 33597 18275 33655 18281
rect 33597 18241 33609 18275
rect 33643 18241 33655 18275
rect 33597 18235 33655 18241
rect 33686 18164 33692 18216
rect 33744 18164 33750 18216
rect 34330 18164 34336 18216
rect 34388 18164 34394 18216
rect 37274 18164 37280 18216
rect 37332 18164 37338 18216
rect 33134 18136 33140 18148
rect 31726 18108 33140 18136
rect 33134 18096 33140 18108
rect 33192 18096 33198 18148
rect 33410 18096 33416 18148
rect 33468 18136 33474 18148
rect 34348 18136 34376 18164
rect 33468 18108 34376 18136
rect 33468 18096 33474 18108
rect 27304 18040 30144 18068
rect 27304 18028 27310 18040
rect 30466 18028 30472 18080
rect 30524 18028 30530 18080
rect 32493 18071 32551 18077
rect 32493 18037 32505 18071
rect 32539 18068 32551 18071
rect 37292 18068 37320 18164
rect 32539 18040 37320 18068
rect 32539 18037 32551 18040
rect 32493 18031 32551 18037
rect 1104 17978 38272 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38272 17978
rect 1104 17904 38272 17926
rect 4798 17824 4804 17876
rect 4856 17864 4862 17876
rect 7742 17864 7748 17876
rect 4856 17836 7748 17864
rect 4856 17824 4862 17836
rect 7742 17824 7748 17836
rect 7800 17824 7806 17876
rect 7834 17824 7840 17876
rect 7892 17864 7898 17876
rect 9490 17864 9496 17876
rect 7892 17836 9496 17864
rect 7892 17824 7898 17836
rect 9490 17824 9496 17836
rect 9548 17864 9554 17876
rect 10042 17864 10048 17876
rect 9548 17836 10048 17864
rect 9548 17824 9554 17836
rect 10042 17824 10048 17836
rect 10100 17824 10106 17876
rect 10686 17824 10692 17876
rect 10744 17864 10750 17876
rect 10873 17867 10931 17873
rect 10873 17864 10885 17867
rect 10744 17836 10885 17864
rect 10744 17824 10750 17836
rect 10873 17833 10885 17836
rect 10919 17833 10931 17867
rect 10873 17827 10931 17833
rect 13722 17824 13728 17876
rect 13780 17864 13786 17876
rect 14090 17864 14096 17876
rect 13780 17836 14096 17864
rect 13780 17824 13786 17836
rect 14090 17824 14096 17836
rect 14148 17824 14154 17876
rect 17494 17824 17500 17876
rect 17552 17864 17558 17876
rect 17589 17867 17647 17873
rect 17589 17864 17601 17867
rect 17552 17836 17601 17864
rect 17552 17824 17558 17836
rect 17589 17833 17601 17836
rect 17635 17833 17647 17867
rect 17589 17827 17647 17833
rect 17770 17824 17776 17876
rect 17828 17864 17834 17876
rect 18690 17864 18696 17876
rect 17828 17836 18696 17864
rect 17828 17824 17834 17836
rect 18690 17824 18696 17836
rect 18748 17864 18754 17876
rect 19061 17867 19119 17873
rect 18748 17836 18920 17864
rect 18748 17824 18754 17836
rect 12621 17799 12679 17805
rect 8404 17768 12572 17796
rect 1394 17688 1400 17740
rect 1452 17728 1458 17740
rect 1854 17728 1860 17740
rect 1452 17700 1860 17728
rect 1452 17688 1458 17700
rect 1854 17688 1860 17700
rect 1912 17728 1918 17740
rect 3970 17728 3976 17740
rect 1912 17700 3976 17728
rect 1912 17688 1918 17700
rect 3970 17688 3976 17700
rect 4028 17728 4034 17740
rect 5077 17731 5135 17737
rect 5077 17728 5089 17731
rect 4028 17700 5089 17728
rect 4028 17688 4034 17700
rect 5077 17697 5089 17700
rect 5123 17697 5135 17731
rect 5077 17691 5135 17697
rect 4801 17663 4859 17669
rect 4801 17629 4813 17663
rect 4847 17660 4859 17663
rect 4890 17660 4896 17672
rect 4847 17632 4896 17660
rect 4847 17629 4859 17632
rect 4801 17623 4859 17629
rect 4890 17620 4896 17632
rect 4948 17620 4954 17672
rect 7101 17663 7159 17669
rect 5353 17595 5411 17601
rect 5353 17561 5365 17595
rect 5399 17592 5411 17595
rect 5626 17592 5632 17604
rect 5399 17564 5632 17592
rect 5399 17561 5411 17564
rect 5353 17555 5411 17561
rect 5626 17552 5632 17564
rect 5684 17552 5690 17604
rect 4614 17484 4620 17536
rect 4672 17484 4678 17536
rect 6178 17484 6184 17536
rect 6236 17524 6242 17536
rect 6472 17524 6500 17646
rect 7101 17629 7113 17663
rect 7147 17660 7159 17663
rect 7193 17663 7251 17669
rect 7193 17660 7205 17663
rect 7147 17632 7205 17660
rect 7147 17629 7159 17632
rect 7101 17623 7159 17629
rect 7193 17629 7205 17632
rect 7239 17660 7251 17663
rect 7282 17660 7288 17672
rect 7239 17632 7288 17660
rect 7239 17629 7251 17632
rect 7193 17623 7251 17629
rect 7282 17620 7288 17632
rect 7340 17660 7346 17672
rect 8110 17660 8116 17672
rect 7340 17632 8116 17660
rect 7340 17620 7346 17632
rect 8110 17620 8116 17632
rect 8168 17620 8174 17672
rect 8404 17604 8432 17768
rect 9692 17700 10548 17728
rect 9692 17672 9720 17700
rect 9674 17620 9680 17672
rect 9732 17620 9738 17672
rect 10042 17620 10048 17672
rect 10100 17660 10106 17672
rect 10520 17669 10548 17700
rect 10612 17669 10640 17768
rect 12544 17740 12572 17768
rect 12621 17765 12633 17799
rect 12667 17796 12679 17799
rect 12667 17768 18828 17796
rect 12667 17765 12679 17768
rect 12621 17759 12679 17765
rect 11808 17700 12480 17728
rect 10229 17663 10287 17669
rect 10229 17660 10241 17663
rect 10100 17632 10241 17660
rect 10100 17620 10106 17632
rect 10229 17629 10241 17632
rect 10275 17629 10287 17663
rect 10229 17623 10287 17629
rect 10413 17663 10471 17669
rect 10413 17629 10425 17663
rect 10459 17629 10471 17663
rect 10413 17623 10471 17629
rect 10505 17663 10563 17669
rect 10505 17629 10517 17663
rect 10551 17629 10563 17663
rect 10505 17623 10563 17629
rect 10597 17663 10655 17669
rect 10597 17629 10609 17663
rect 10643 17629 10655 17663
rect 11808 17660 11836 17700
rect 10597 17623 10655 17629
rect 10704 17632 11836 17660
rect 8018 17552 8024 17604
rect 8076 17592 8082 17604
rect 8386 17592 8392 17604
rect 8076 17564 8392 17592
rect 8076 17552 8082 17564
rect 8386 17552 8392 17564
rect 8444 17552 8450 17604
rect 10134 17552 10140 17604
rect 10192 17592 10198 17604
rect 10428 17592 10456 17623
rect 10704 17592 10732 17632
rect 12158 17620 12164 17672
rect 12216 17620 12222 17672
rect 12250 17620 12256 17672
rect 12308 17620 12314 17672
rect 12452 17669 12480 17700
rect 12526 17688 12532 17740
rect 12584 17688 12590 17740
rect 16669 17731 16727 17737
rect 16669 17728 16681 17731
rect 15856 17700 16681 17728
rect 12437 17663 12495 17669
rect 12437 17629 12449 17663
rect 12483 17660 12495 17663
rect 13722 17660 13728 17672
rect 12483 17632 13728 17660
rect 12483 17629 12495 17632
rect 12437 17623 12495 17629
rect 13722 17620 13728 17632
rect 13780 17620 13786 17672
rect 14734 17660 14740 17672
rect 14384 17632 14740 17660
rect 10192 17564 10732 17592
rect 10192 17552 10198 17564
rect 10778 17552 10784 17604
rect 10836 17592 10842 17604
rect 13446 17592 13452 17604
rect 10836 17564 13452 17592
rect 10836 17552 10842 17564
rect 13446 17552 13452 17564
rect 13504 17552 13510 17604
rect 6236 17496 6500 17524
rect 6236 17484 6242 17496
rect 7742 17484 7748 17536
rect 7800 17524 7806 17536
rect 11606 17524 11612 17536
rect 7800 17496 11612 17524
rect 7800 17484 7806 17496
rect 11606 17484 11612 17496
rect 11664 17484 11670 17536
rect 11974 17484 11980 17536
rect 12032 17524 12038 17536
rect 12250 17524 12256 17536
rect 12032 17496 12256 17524
rect 12032 17484 12038 17496
rect 12250 17484 12256 17496
rect 12308 17484 12314 17536
rect 12342 17484 12348 17536
rect 12400 17524 12406 17536
rect 14384 17524 14412 17632
rect 14734 17620 14740 17632
rect 14792 17620 14798 17672
rect 14826 17620 14832 17672
rect 14884 17660 14890 17672
rect 14921 17663 14979 17669
rect 14921 17660 14933 17663
rect 14884 17632 14933 17660
rect 14884 17620 14890 17632
rect 14921 17629 14933 17632
rect 14967 17629 14979 17663
rect 14921 17623 14979 17629
rect 15378 17620 15384 17672
rect 15436 17620 15442 17672
rect 15473 17663 15531 17669
rect 15473 17629 15485 17663
rect 15519 17660 15531 17663
rect 15654 17660 15660 17672
rect 15519 17632 15660 17660
rect 15519 17629 15531 17632
rect 15473 17623 15531 17629
rect 15654 17620 15660 17632
rect 15712 17660 15718 17672
rect 15856 17660 15884 17700
rect 16669 17697 16681 17700
rect 16715 17728 16727 17731
rect 17034 17728 17040 17740
rect 16715 17700 17040 17728
rect 16715 17697 16727 17700
rect 16669 17691 16727 17697
rect 17034 17688 17040 17700
rect 17092 17688 17098 17740
rect 17972 17700 18552 17728
rect 15712 17632 15884 17660
rect 16301 17663 16359 17669
rect 15712 17620 15718 17632
rect 16301 17629 16313 17663
rect 16347 17629 16359 17663
rect 16301 17623 16359 17629
rect 16393 17663 16451 17669
rect 16393 17629 16405 17663
rect 16439 17660 16451 17663
rect 16574 17660 16580 17672
rect 16439 17632 16580 17660
rect 16439 17629 16451 17632
rect 16393 17623 16451 17629
rect 16025 17595 16083 17601
rect 16025 17561 16037 17595
rect 16071 17592 16083 17595
rect 16206 17592 16212 17604
rect 16071 17564 16212 17592
rect 16071 17561 16083 17564
rect 16025 17555 16083 17561
rect 16206 17552 16212 17564
rect 16264 17552 16270 17604
rect 16316 17592 16344 17623
rect 16574 17620 16580 17632
rect 16632 17620 16638 17672
rect 16761 17663 16819 17669
rect 16761 17629 16773 17663
rect 16807 17660 16819 17663
rect 16850 17660 16856 17672
rect 16807 17632 16856 17660
rect 16807 17629 16819 17632
rect 16761 17623 16819 17629
rect 16850 17620 16856 17632
rect 16908 17620 16914 17672
rect 17218 17620 17224 17672
rect 17276 17620 17282 17672
rect 17770 17620 17776 17672
rect 17828 17660 17834 17672
rect 17972 17669 18000 17700
rect 18524 17672 18552 17700
rect 17865 17663 17923 17669
rect 17865 17660 17877 17663
rect 17828 17632 17877 17660
rect 17828 17620 17834 17632
rect 17865 17629 17877 17632
rect 17911 17629 17923 17663
rect 17865 17623 17923 17629
rect 17957 17663 18015 17669
rect 17957 17629 17969 17663
rect 18003 17629 18015 17663
rect 17957 17623 18015 17629
rect 18046 17620 18052 17672
rect 18104 17620 18110 17672
rect 18230 17620 18236 17672
rect 18288 17620 18294 17672
rect 18506 17620 18512 17672
rect 18564 17620 18570 17672
rect 18800 17669 18828 17768
rect 18892 17728 18920 17836
rect 19061 17833 19073 17867
rect 19107 17864 19119 17867
rect 19150 17864 19156 17876
rect 19107 17836 19156 17864
rect 19107 17833 19119 17836
rect 19061 17827 19119 17833
rect 19150 17824 19156 17836
rect 19208 17824 19214 17876
rect 20714 17824 20720 17876
rect 20772 17864 20778 17876
rect 21729 17867 21787 17873
rect 21729 17864 21741 17867
rect 20772 17836 21741 17864
rect 20772 17824 20778 17836
rect 21729 17833 21741 17836
rect 21775 17833 21787 17867
rect 24854 17864 24860 17876
rect 21729 17827 21787 17833
rect 22066 17836 24860 17864
rect 18966 17756 18972 17808
rect 19024 17796 19030 17808
rect 21637 17799 21695 17805
rect 19024 17768 20392 17796
rect 19024 17756 19030 17768
rect 20364 17740 20392 17768
rect 21637 17765 21649 17799
rect 21683 17796 21695 17799
rect 22066 17796 22094 17836
rect 24854 17824 24860 17836
rect 24912 17864 24918 17876
rect 25222 17864 25228 17876
rect 24912 17836 25228 17864
rect 24912 17824 24918 17836
rect 25222 17824 25228 17836
rect 25280 17824 25286 17876
rect 28721 17867 28779 17873
rect 25516 17836 28396 17864
rect 25516 17808 25544 17836
rect 23842 17796 23848 17808
rect 21683 17768 22094 17796
rect 23124 17768 23848 17796
rect 21683 17765 21695 17768
rect 21637 17759 21695 17765
rect 18892 17700 19656 17728
rect 18892 17669 18920 17700
rect 18785 17663 18843 17669
rect 18785 17629 18797 17663
rect 18831 17629 18843 17663
rect 18785 17623 18843 17629
rect 18877 17663 18935 17669
rect 18877 17629 18889 17663
rect 18923 17629 18935 17663
rect 19245 17663 19303 17669
rect 19245 17660 19257 17663
rect 18877 17623 18935 17629
rect 19168 17632 19257 17660
rect 16482 17592 16488 17604
rect 16316 17564 16488 17592
rect 16482 17552 16488 17564
rect 16540 17552 16546 17604
rect 16592 17592 16620 17620
rect 17034 17592 17040 17604
rect 16592 17564 17040 17592
rect 17034 17552 17040 17564
rect 17092 17552 17098 17604
rect 18138 17552 18144 17604
rect 18196 17592 18202 17604
rect 18325 17595 18383 17601
rect 18325 17592 18337 17595
rect 18196 17564 18337 17592
rect 18196 17552 18202 17564
rect 18325 17561 18337 17564
rect 18371 17561 18383 17595
rect 18800 17592 18828 17623
rect 18966 17592 18972 17604
rect 18800 17564 18972 17592
rect 18325 17555 18383 17561
rect 18966 17552 18972 17564
rect 19024 17592 19030 17604
rect 19168 17592 19196 17632
rect 19245 17629 19257 17632
rect 19291 17629 19303 17663
rect 19245 17623 19303 17629
rect 19334 17620 19340 17672
rect 19392 17620 19398 17672
rect 19628 17669 19656 17700
rect 20346 17688 20352 17740
rect 20404 17688 20410 17740
rect 20625 17731 20683 17737
rect 20625 17697 20637 17731
rect 20671 17728 20683 17731
rect 20671 17700 23060 17728
rect 20671 17697 20683 17700
rect 20625 17691 20683 17697
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17629 19671 17663
rect 19613 17623 19671 17629
rect 19981 17663 20039 17669
rect 19981 17629 19993 17663
rect 20027 17629 20039 17663
rect 19981 17623 20039 17629
rect 19024 17564 19196 17592
rect 19352 17592 19380 17620
rect 19996 17592 20024 17623
rect 20806 17620 20812 17672
rect 20864 17620 20870 17672
rect 21082 17620 21088 17672
rect 21140 17620 21146 17672
rect 21174 17620 21180 17672
rect 21232 17620 21238 17672
rect 21913 17663 21971 17669
rect 21913 17629 21925 17663
rect 21959 17629 21971 17663
rect 21913 17623 21971 17629
rect 21192 17592 21220 17620
rect 19352 17564 21220 17592
rect 21453 17595 21511 17601
rect 19024 17552 19030 17564
rect 21453 17561 21465 17595
rect 21499 17592 21511 17595
rect 21928 17592 21956 17623
rect 22278 17620 22284 17672
rect 22336 17660 22342 17672
rect 22664 17669 22692 17700
rect 23032 17672 23060 17700
rect 22431 17663 22489 17669
rect 22431 17660 22443 17663
rect 22336 17632 22443 17660
rect 22336 17620 22342 17632
rect 22431 17629 22443 17632
rect 22477 17629 22489 17663
rect 22431 17623 22489 17629
rect 22557 17663 22615 17669
rect 22557 17629 22569 17663
rect 22603 17629 22615 17663
rect 22557 17623 22615 17629
rect 22649 17663 22707 17669
rect 22649 17629 22661 17663
rect 22695 17629 22707 17663
rect 22649 17623 22707 17629
rect 22756 17647 22876 17660
rect 22756 17641 22892 17647
rect 22756 17632 22846 17641
rect 21499 17564 21956 17592
rect 22189 17595 22247 17601
rect 21499 17561 21511 17564
rect 21453 17555 21511 17561
rect 22189 17561 22201 17595
rect 22235 17561 22247 17595
rect 22189 17555 22247 17561
rect 12400 17496 14412 17524
rect 17129 17527 17187 17533
rect 12400 17484 12406 17496
rect 17129 17493 17141 17527
rect 17175 17524 17187 17527
rect 20438 17524 20444 17536
rect 17175 17496 20444 17524
rect 17175 17493 17187 17496
rect 17129 17487 17187 17493
rect 20438 17484 20444 17496
rect 20496 17484 20502 17536
rect 21174 17484 21180 17536
rect 21232 17524 21238 17536
rect 21468 17524 21496 17555
rect 21232 17496 21496 17524
rect 22204 17524 22232 17555
rect 22572 17536 22600 17623
rect 22756 17604 22784 17632
rect 22834 17607 22846 17632
rect 22880 17607 22892 17641
rect 23014 17620 23020 17672
rect 23072 17620 23078 17672
rect 23124 17669 23152 17768
rect 23842 17756 23848 17768
rect 23900 17756 23906 17808
rect 24412 17768 25268 17796
rect 23934 17688 23940 17740
rect 23992 17728 23998 17740
rect 24412 17737 24440 17768
rect 24397 17731 24455 17737
rect 24397 17728 24409 17731
rect 23992 17700 24409 17728
rect 23992 17688 23998 17700
rect 24397 17697 24409 17700
rect 24443 17697 24455 17731
rect 24397 17691 24455 17697
rect 25130 17688 25136 17740
rect 25188 17688 25194 17740
rect 25240 17737 25268 17768
rect 25498 17756 25504 17808
rect 25556 17756 25562 17808
rect 26605 17799 26663 17805
rect 26605 17765 26617 17799
rect 26651 17796 26663 17799
rect 26651 17768 26832 17796
rect 26651 17765 26663 17768
rect 26605 17759 26663 17765
rect 25225 17731 25283 17737
rect 25225 17697 25237 17731
rect 25271 17697 25283 17731
rect 25225 17691 25283 17697
rect 23109 17663 23167 17669
rect 23109 17629 23121 17663
rect 23155 17629 23167 17663
rect 23109 17623 23167 17629
rect 23474 17620 23480 17672
rect 23532 17620 23538 17672
rect 24489 17663 24547 17669
rect 24489 17660 24501 17663
rect 23860 17632 24501 17660
rect 22738 17552 22744 17604
rect 22796 17552 22802 17604
rect 22834 17601 22892 17607
rect 22922 17552 22928 17604
rect 22980 17552 22986 17604
rect 23860 17536 23888 17632
rect 24489 17629 24501 17632
rect 24535 17660 24547 17663
rect 25317 17663 25375 17669
rect 25317 17660 25329 17663
rect 24535 17632 25329 17660
rect 24535 17629 24547 17632
rect 24489 17623 24547 17629
rect 25317 17629 25329 17632
rect 25363 17629 25375 17663
rect 25317 17623 25375 17629
rect 25498 17620 25504 17672
rect 25556 17660 25562 17672
rect 26804 17669 26832 17768
rect 27065 17731 27123 17737
rect 27065 17697 27077 17731
rect 27111 17728 27123 17731
rect 27154 17728 27160 17740
rect 27111 17700 27160 17728
rect 27111 17697 27123 17700
rect 27065 17691 27123 17697
rect 27154 17688 27160 17700
rect 27212 17688 27218 17740
rect 25593 17663 25651 17669
rect 25593 17660 25605 17663
rect 25556 17632 25605 17660
rect 25556 17620 25562 17632
rect 25593 17629 25605 17632
rect 25639 17629 25651 17663
rect 25593 17623 25651 17629
rect 25685 17663 25743 17669
rect 25685 17629 25697 17663
rect 25731 17660 25743 17663
rect 26513 17663 26571 17669
rect 25731 17632 26372 17660
rect 25731 17629 25743 17632
rect 25685 17623 25743 17629
rect 24118 17552 24124 17604
rect 24176 17592 24182 17604
rect 24765 17595 24823 17601
rect 24765 17592 24777 17595
rect 24176 17564 24777 17592
rect 24176 17552 24182 17564
rect 24765 17561 24777 17564
rect 24811 17561 24823 17595
rect 24765 17555 24823 17561
rect 24851 17595 24909 17601
rect 24851 17561 24863 17595
rect 24897 17592 24909 17595
rect 24946 17592 24952 17604
rect 24897 17564 24952 17592
rect 24897 17561 24909 17564
rect 24851 17555 24909 17561
rect 24946 17552 24952 17564
rect 25004 17552 25010 17604
rect 25222 17552 25228 17604
rect 25280 17592 25286 17604
rect 25700 17592 25728 17623
rect 25280 17564 25728 17592
rect 25280 17552 25286 17564
rect 26344 17536 26372 17632
rect 26513 17629 26525 17663
rect 26559 17629 26571 17663
rect 26513 17623 26571 17629
rect 26789 17663 26847 17669
rect 26789 17629 26801 17663
rect 26835 17629 26847 17663
rect 26789 17623 26847 17629
rect 22462 17524 22468 17536
rect 22204 17496 22468 17524
rect 21232 17484 21238 17496
rect 22462 17484 22468 17496
rect 22520 17484 22526 17536
rect 22554 17484 22560 17536
rect 22612 17524 22618 17536
rect 23842 17524 23848 17536
rect 22612 17496 23848 17524
rect 22612 17484 22618 17496
rect 23842 17484 23848 17496
rect 23900 17484 23906 17536
rect 24578 17484 24584 17536
rect 24636 17524 24642 17536
rect 24673 17527 24731 17533
rect 24673 17524 24685 17527
rect 24636 17496 24685 17524
rect 24636 17484 24642 17496
rect 24673 17493 24685 17496
rect 24719 17524 24731 17527
rect 25501 17527 25559 17533
rect 25501 17524 25513 17527
rect 24719 17496 25513 17524
rect 24719 17493 24731 17496
rect 24673 17487 24731 17493
rect 25501 17493 25513 17496
rect 25547 17493 25559 17527
rect 25501 17487 25559 17493
rect 25958 17484 25964 17536
rect 26016 17484 26022 17536
rect 26326 17484 26332 17536
rect 26384 17484 26390 17536
rect 26528 17524 26556 17623
rect 27522 17552 27528 17604
rect 27580 17552 27586 17604
rect 28368 17592 28396 17836
rect 28721 17833 28733 17867
rect 28767 17864 28779 17867
rect 28994 17864 29000 17876
rect 28767 17836 29000 17864
rect 28767 17833 28779 17836
rect 28721 17827 28779 17833
rect 28994 17824 29000 17836
rect 29052 17824 29058 17876
rect 29181 17867 29239 17873
rect 29181 17833 29193 17867
rect 29227 17864 29239 17867
rect 29270 17864 29276 17876
rect 29227 17836 29276 17864
rect 29227 17833 29239 17836
rect 29181 17827 29239 17833
rect 29270 17824 29276 17836
rect 29328 17824 29334 17876
rect 30929 17867 30987 17873
rect 30929 17833 30941 17867
rect 30975 17864 30987 17867
rect 37366 17864 37372 17876
rect 30975 17836 37372 17864
rect 30975 17833 30987 17836
rect 30929 17827 30987 17833
rect 37366 17824 37372 17836
rect 37424 17824 37430 17876
rect 29733 17731 29791 17737
rect 29733 17728 29745 17731
rect 29012 17700 29745 17728
rect 28810 17620 28816 17672
rect 28868 17660 28874 17672
rect 29012 17669 29040 17700
rect 29733 17697 29745 17700
rect 29779 17697 29791 17731
rect 29733 17691 29791 17697
rect 30377 17731 30435 17737
rect 30377 17697 30389 17731
rect 30423 17728 30435 17731
rect 30466 17728 30472 17740
rect 30423 17700 30472 17728
rect 30423 17697 30435 17700
rect 30377 17691 30435 17697
rect 30466 17688 30472 17700
rect 30524 17728 30530 17740
rect 30834 17728 30840 17740
rect 30524 17700 30840 17728
rect 30524 17688 30530 17700
rect 30834 17688 30840 17700
rect 30892 17688 30898 17740
rect 28905 17663 28963 17669
rect 28905 17660 28917 17663
rect 28868 17632 28917 17660
rect 28868 17620 28874 17632
rect 28905 17629 28917 17632
rect 28951 17629 28963 17663
rect 28905 17623 28963 17629
rect 28997 17663 29055 17669
rect 28997 17629 29009 17663
rect 29043 17629 29055 17663
rect 28997 17623 29055 17629
rect 29273 17663 29331 17669
rect 29273 17629 29285 17663
rect 29319 17629 29331 17663
rect 29273 17623 29331 17629
rect 29288 17592 29316 17623
rect 30558 17620 30564 17672
rect 30616 17620 30622 17672
rect 30745 17663 30803 17669
rect 30745 17629 30757 17663
rect 30791 17660 30803 17663
rect 31202 17660 31208 17672
rect 30791 17632 31208 17660
rect 30791 17629 30803 17632
rect 30745 17623 30803 17629
rect 31202 17620 31208 17632
rect 31260 17620 31266 17672
rect 31294 17592 31300 17604
rect 28368 17564 31300 17592
rect 31294 17552 31300 17564
rect 31352 17552 31358 17604
rect 27430 17524 27436 17536
rect 26528 17496 27436 17524
rect 27430 17484 27436 17496
rect 27488 17484 27494 17536
rect 28534 17484 28540 17536
rect 28592 17484 28598 17536
rect 1104 17434 38272 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 38272 17434
rect 1104 17360 38272 17382
rect 3694 17280 3700 17332
rect 3752 17280 3758 17332
rect 4614 17320 4620 17332
rect 4356 17292 4620 17320
rect 3145 17187 3203 17193
rect 3145 17153 3157 17187
rect 3191 17184 3203 17187
rect 3712 17184 3740 17280
rect 4356 17261 4384 17292
rect 4614 17280 4620 17292
rect 4672 17280 4678 17332
rect 8846 17280 8852 17332
rect 8904 17280 8910 17332
rect 10686 17280 10692 17332
rect 10744 17320 10750 17332
rect 10744 17292 11192 17320
rect 10744 17280 10750 17292
rect 4341 17255 4399 17261
rect 4341 17221 4353 17255
rect 4387 17221 4399 17255
rect 6178 17252 6184 17264
rect 5566 17224 6184 17252
rect 4341 17215 4399 17221
rect 6178 17212 6184 17224
rect 6236 17212 6242 17264
rect 7193 17255 7251 17261
rect 7193 17221 7205 17255
rect 7239 17252 7251 17255
rect 7834 17252 7840 17264
rect 7239 17224 7840 17252
rect 7239 17221 7251 17224
rect 7193 17215 7251 17221
rect 7834 17212 7840 17224
rect 7892 17212 7898 17264
rect 8864 17252 8892 17280
rect 11054 17252 11060 17264
rect 8772 17224 8892 17252
rect 9416 17224 11060 17252
rect 3191 17156 3740 17184
rect 3191 17153 3203 17156
rect 3145 17147 3203 17153
rect 3970 17144 3976 17196
rect 4028 17184 4034 17196
rect 4065 17187 4123 17193
rect 4065 17184 4077 17187
rect 4028 17156 4077 17184
rect 4028 17144 4034 17156
rect 4065 17153 4077 17156
rect 4111 17153 4123 17187
rect 6365 17187 6423 17193
rect 6365 17184 6377 17187
rect 4065 17147 4123 17153
rect 5828 17156 6377 17184
rect 5828 17125 5856 17156
rect 6365 17153 6377 17156
rect 6411 17153 6423 17187
rect 6365 17147 6423 17153
rect 7926 17144 7932 17196
rect 7984 17144 7990 17196
rect 8772 17193 8800 17224
rect 8757 17187 8815 17193
rect 8757 17153 8769 17187
rect 8803 17153 8815 17187
rect 8757 17147 8815 17153
rect 8849 17187 8907 17193
rect 8849 17153 8861 17187
rect 8895 17184 8907 17187
rect 8895 17156 9168 17184
rect 8895 17153 8907 17156
rect 8849 17147 8907 17153
rect 5813 17119 5871 17125
rect 5813 17085 5825 17119
rect 5859 17085 5871 17119
rect 5813 17079 5871 17085
rect 2498 16940 2504 16992
rect 2556 16980 2562 16992
rect 2961 16983 3019 16989
rect 2961 16980 2973 16983
rect 2556 16952 2973 16980
rect 2556 16940 2562 16952
rect 2961 16949 2973 16952
rect 3007 16949 3019 16983
rect 2961 16943 3019 16949
rect 8202 16940 8208 16992
rect 8260 16980 8266 16992
rect 9140 16980 9168 17156
rect 9214 17144 9220 17196
rect 9272 17144 9278 17196
rect 9416 17057 9444 17224
rect 11054 17212 11060 17224
rect 11112 17212 11118 17264
rect 11164 17252 11192 17292
rect 11882 17280 11888 17332
rect 11940 17280 11946 17332
rect 12158 17280 12164 17332
rect 12216 17320 12222 17332
rect 12529 17323 12587 17329
rect 12529 17320 12541 17323
rect 12216 17292 12541 17320
rect 12216 17280 12222 17292
rect 12529 17289 12541 17292
rect 12575 17289 12587 17323
rect 12529 17283 12587 17289
rect 12802 17280 12808 17332
rect 12860 17320 12866 17332
rect 13173 17323 13231 17329
rect 13173 17320 13185 17323
rect 12860 17292 13185 17320
rect 12860 17280 12866 17292
rect 13173 17289 13185 17292
rect 13219 17289 13231 17323
rect 14642 17320 14648 17332
rect 13173 17283 13231 17289
rect 13832 17292 14648 17320
rect 12069 17255 12127 17261
rect 12069 17252 12081 17255
rect 11164 17224 12081 17252
rect 12069 17221 12081 17224
rect 12115 17221 12127 17255
rect 12069 17215 12127 17221
rect 12250 17212 12256 17264
rect 12308 17212 12314 17264
rect 12434 17212 12440 17264
rect 12492 17252 12498 17264
rect 13078 17252 13084 17264
rect 12492 17224 13084 17252
rect 12492 17212 12498 17224
rect 13078 17212 13084 17224
rect 13136 17212 13142 17264
rect 9674 17144 9680 17196
rect 9732 17144 9738 17196
rect 10226 17144 10232 17196
rect 10284 17144 10290 17196
rect 10321 17187 10379 17193
rect 10321 17153 10333 17187
rect 10367 17184 10379 17187
rect 10781 17187 10839 17193
rect 10781 17184 10793 17187
rect 10367 17156 10793 17184
rect 10367 17153 10379 17156
rect 10321 17147 10379 17153
rect 10781 17153 10793 17156
rect 10827 17184 10839 17187
rect 10870 17184 10876 17196
rect 10827 17156 10876 17184
rect 10827 17153 10839 17156
rect 10781 17147 10839 17153
rect 10870 17144 10876 17156
rect 10928 17144 10934 17196
rect 10965 17187 11023 17193
rect 10965 17153 10977 17187
rect 11011 17184 11023 17187
rect 11698 17184 11704 17196
rect 11011 17156 11704 17184
rect 11011 17153 11023 17156
rect 10965 17147 11023 17153
rect 9766 17076 9772 17128
rect 9824 17116 9830 17128
rect 10502 17116 10508 17128
rect 9824 17088 10508 17116
rect 9824 17076 9830 17088
rect 10502 17076 10508 17088
rect 10560 17116 10566 17128
rect 10597 17119 10655 17125
rect 10597 17116 10609 17119
rect 10560 17088 10609 17116
rect 10560 17076 10566 17088
rect 10597 17085 10609 17088
rect 10643 17085 10655 17119
rect 10597 17079 10655 17085
rect 10686 17076 10692 17128
rect 10744 17076 10750 17128
rect 9401 17051 9459 17057
rect 9401 17017 9413 17051
rect 9447 17017 9459 17051
rect 10980 17048 11008 17147
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 11977 17187 12035 17193
rect 11977 17153 11989 17187
rect 12023 17184 12035 17187
rect 13725 17187 13783 17193
rect 12023 17156 12664 17184
rect 12023 17153 12035 17156
rect 11977 17147 12035 17153
rect 12636 17128 12664 17156
rect 13725 17153 13737 17187
rect 13771 17153 13783 17187
rect 13832 17184 13860 17292
rect 14642 17280 14648 17292
rect 14700 17280 14706 17332
rect 14734 17280 14740 17332
rect 14792 17320 14798 17332
rect 15565 17323 15623 17329
rect 15565 17320 15577 17323
rect 14792 17292 15577 17320
rect 14792 17280 14798 17292
rect 15565 17289 15577 17292
rect 15611 17289 15623 17323
rect 15565 17283 15623 17289
rect 16408 17292 17264 17320
rect 13998 17212 14004 17264
rect 14056 17252 14062 17264
rect 14918 17252 14924 17264
rect 14056 17224 14924 17252
rect 14056 17212 14062 17224
rect 14918 17212 14924 17224
rect 14976 17252 14982 17264
rect 16408 17252 16436 17292
rect 17236 17264 17264 17292
rect 18690 17280 18696 17332
rect 18748 17280 18754 17332
rect 19153 17323 19211 17329
rect 19153 17289 19165 17323
rect 19199 17320 19211 17323
rect 19199 17292 19334 17320
rect 19199 17289 19211 17292
rect 19153 17283 19211 17289
rect 14976 17224 16436 17252
rect 14976 17212 14982 17224
rect 13909 17187 13967 17193
rect 13909 17184 13921 17187
rect 13832 17156 13921 17184
rect 13725 17147 13783 17153
rect 13909 17153 13921 17156
rect 13955 17153 13967 17187
rect 13909 17147 13967 17153
rect 11517 17119 11575 17125
rect 11517 17085 11529 17119
rect 11563 17116 11575 17119
rect 11606 17116 11612 17128
rect 11563 17088 11612 17116
rect 11563 17085 11575 17088
rect 11517 17079 11575 17085
rect 11606 17076 11612 17088
rect 11664 17076 11670 17128
rect 12618 17076 12624 17128
rect 12676 17116 12682 17128
rect 12713 17119 12771 17125
rect 12713 17116 12725 17119
rect 12676 17088 12725 17116
rect 12676 17076 12682 17088
rect 12713 17085 12725 17088
rect 12759 17085 12771 17119
rect 12713 17079 12771 17085
rect 12805 17119 12863 17125
rect 12805 17085 12817 17119
rect 12851 17085 12863 17119
rect 13740 17116 13768 17147
rect 14090 17144 14096 17196
rect 14148 17193 14154 17196
rect 14148 17147 14156 17193
rect 14148 17144 14154 17147
rect 14458 17144 14464 17196
rect 14516 17144 14522 17196
rect 14826 17144 14832 17196
rect 14884 17184 14890 17196
rect 15567 17187 15625 17193
rect 15567 17184 15579 17187
rect 14884 17156 15579 17184
rect 14884 17144 14890 17156
rect 15567 17153 15579 17156
rect 15613 17153 15625 17187
rect 15567 17147 15625 17153
rect 15654 17144 15660 17196
rect 15712 17144 15718 17196
rect 16408 17184 16436 17224
rect 16482 17212 16488 17264
rect 16540 17252 16546 17264
rect 16540 17224 17177 17252
rect 16540 17212 16546 17224
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 16408 17156 16681 17184
rect 16669 17153 16681 17156
rect 16715 17153 16727 17187
rect 16669 17147 16727 17153
rect 16762 17187 16820 17193
rect 16762 17153 16774 17187
rect 16808 17153 16820 17187
rect 16762 17147 16820 17153
rect 14476 17116 14504 17144
rect 13740 17088 14504 17116
rect 15105 17119 15163 17125
rect 12805 17079 12863 17085
rect 15105 17085 15117 17119
rect 15151 17116 15163 17119
rect 15672 17116 15700 17144
rect 16777 17116 16805 17147
rect 16850 17144 16856 17196
rect 16908 17184 16914 17196
rect 16945 17187 17003 17193
rect 16945 17184 16957 17187
rect 16908 17156 16957 17184
rect 16908 17144 16914 17156
rect 16945 17153 16957 17156
rect 16991 17153 17003 17187
rect 16945 17147 17003 17153
rect 17034 17144 17040 17196
rect 17092 17144 17098 17196
rect 17149 17193 17177 17224
rect 17218 17212 17224 17264
rect 17276 17212 17282 17264
rect 18708 17252 18736 17280
rect 19306 17252 19334 17292
rect 20806 17280 20812 17332
rect 20864 17280 20870 17332
rect 21174 17280 21180 17332
rect 21232 17280 21238 17332
rect 24578 17320 24584 17332
rect 24136 17292 24584 17320
rect 22278 17252 22284 17264
rect 18708 17224 18828 17252
rect 19306 17224 22284 17252
rect 17134 17187 17192 17193
rect 17134 17153 17146 17187
rect 17180 17153 17192 17187
rect 18800 17185 18828 17224
rect 22278 17212 22284 17224
rect 22336 17252 22342 17264
rect 22336 17224 22968 17252
rect 22336 17212 22342 17224
rect 18877 17187 18935 17193
rect 18877 17185 18889 17187
rect 18800 17157 18889 17185
rect 17134 17147 17192 17153
rect 18877 17153 18889 17157
rect 18923 17153 18935 17187
rect 18877 17147 18935 17153
rect 18966 17144 18972 17196
rect 19024 17144 19030 17196
rect 20346 17144 20352 17196
rect 20404 17184 20410 17196
rect 20441 17187 20499 17193
rect 20441 17184 20453 17187
rect 20404 17156 20453 17184
rect 20404 17144 20410 17156
rect 20441 17153 20453 17156
rect 20487 17184 20499 17187
rect 21269 17187 21327 17193
rect 20487 17156 21128 17184
rect 20487 17153 20499 17156
rect 20441 17147 20499 17153
rect 15151 17088 16805 17116
rect 18693 17119 18751 17125
rect 15151 17085 15163 17088
rect 15105 17079 15163 17085
rect 18693 17085 18705 17119
rect 18739 17085 18751 17119
rect 18693 17079 18751 17085
rect 18785 17119 18843 17125
rect 18785 17085 18797 17119
rect 18831 17116 18843 17119
rect 19150 17116 19156 17128
rect 18831 17088 19156 17116
rect 18831 17085 18843 17088
rect 18785 17079 18843 17085
rect 9401 17011 9459 17017
rect 9508 17020 11008 17048
rect 9508 16980 9536 17020
rect 11698 17008 11704 17060
rect 11756 17008 11762 17060
rect 11882 17008 11888 17060
rect 11940 17048 11946 17060
rect 12820 17048 12848 17079
rect 13538 17048 13544 17060
rect 11940 17020 13544 17048
rect 11940 17008 11946 17020
rect 13538 17008 13544 17020
rect 13596 17008 13602 17060
rect 18708 17048 18736 17079
rect 19150 17076 19156 17088
rect 19208 17076 19214 17128
rect 21100 17125 21128 17156
rect 21269 17153 21281 17187
rect 21315 17184 21327 17187
rect 21542 17184 21548 17196
rect 21315 17156 21548 17184
rect 21315 17153 21327 17156
rect 21269 17147 21327 17153
rect 21542 17144 21548 17156
rect 21600 17144 21606 17196
rect 22465 17187 22523 17193
rect 22465 17184 22477 17187
rect 21928 17156 22477 17184
rect 20533 17119 20591 17125
rect 20533 17085 20545 17119
rect 20579 17116 20591 17119
rect 20901 17119 20959 17125
rect 20901 17116 20913 17119
rect 20579 17088 20913 17116
rect 20579 17085 20591 17088
rect 20533 17079 20591 17085
rect 20901 17085 20913 17088
rect 20947 17085 20959 17119
rect 20901 17079 20959 17085
rect 21085 17119 21143 17125
rect 21085 17085 21097 17119
rect 21131 17116 21143 17119
rect 21928 17116 21956 17156
rect 22465 17153 22477 17156
rect 22511 17184 22523 17187
rect 22554 17184 22560 17196
rect 22511 17156 22560 17184
rect 22511 17153 22523 17156
rect 22465 17147 22523 17153
rect 22554 17144 22560 17156
rect 22612 17144 22618 17196
rect 21131 17088 21956 17116
rect 21131 17085 21143 17088
rect 21085 17079 21143 17085
rect 18874 17048 18880 17060
rect 18708 17020 18880 17048
rect 18874 17008 18880 17020
rect 18932 17008 18938 17060
rect 20548 17048 20576 17079
rect 22186 17076 22192 17128
rect 22244 17116 22250 17128
rect 22756 17125 22784 17224
rect 22833 17187 22891 17193
rect 22833 17153 22845 17187
rect 22879 17153 22891 17187
rect 22940 17184 22968 17224
rect 23014 17212 23020 17264
rect 23072 17252 23078 17264
rect 24136 17252 24164 17292
rect 24578 17280 24584 17292
rect 24636 17280 24642 17332
rect 24670 17280 24676 17332
rect 24728 17280 24734 17332
rect 25130 17280 25136 17332
rect 25188 17280 25194 17332
rect 25317 17323 25375 17329
rect 25317 17289 25329 17323
rect 25363 17320 25375 17323
rect 25866 17320 25872 17332
rect 25363 17292 25872 17320
rect 25363 17289 25375 17292
rect 25317 17283 25375 17289
rect 25866 17280 25872 17292
rect 25924 17280 25930 17332
rect 25958 17280 25964 17332
rect 26016 17280 26022 17332
rect 26970 17280 26976 17332
rect 27028 17280 27034 17332
rect 27433 17323 27491 17329
rect 27433 17289 27445 17323
rect 27479 17320 27491 17323
rect 28166 17320 28172 17332
rect 27479 17292 28172 17320
rect 27479 17289 27491 17292
rect 27433 17283 27491 17289
rect 23072 17224 24164 17252
rect 23072 17212 23078 17224
rect 24121 17187 24179 17193
rect 24121 17184 24133 17187
rect 22940 17156 24133 17184
rect 22833 17147 22891 17153
rect 24121 17153 24133 17156
rect 24167 17153 24179 17187
rect 24121 17147 24179 17153
rect 24213 17187 24271 17193
rect 24213 17153 24225 17187
rect 24259 17153 24271 17187
rect 24213 17147 24271 17153
rect 24305 17187 24363 17193
rect 24305 17153 24317 17187
rect 24351 17184 24363 17187
rect 24394 17184 24400 17196
rect 24351 17156 24400 17184
rect 24351 17153 24363 17156
rect 24305 17147 24363 17153
rect 22281 17119 22339 17125
rect 22281 17116 22293 17119
rect 22244 17088 22293 17116
rect 22244 17076 22250 17088
rect 22281 17085 22293 17088
rect 22327 17085 22339 17119
rect 22281 17079 22339 17085
rect 22741 17119 22799 17125
rect 22741 17085 22753 17119
rect 22787 17085 22799 17119
rect 22848 17116 22876 17147
rect 23198 17116 23204 17128
rect 22848 17088 23204 17116
rect 22741 17079 22799 17085
rect 20364 17020 20576 17048
rect 8260 16952 9536 16980
rect 8260 16940 8266 16952
rect 9766 16940 9772 16992
rect 9824 16980 9830 16992
rect 10045 16983 10103 16989
rect 10045 16980 10057 16983
rect 9824 16952 10057 16980
rect 9824 16940 9830 16952
rect 10045 16949 10057 16952
rect 10091 16949 10103 16983
rect 10045 16943 10103 16949
rect 10778 16940 10784 16992
rect 10836 16940 10842 16992
rect 10870 16940 10876 16992
rect 10928 16980 10934 16992
rect 12434 16980 12440 16992
rect 10928 16952 12440 16980
rect 10928 16940 10934 16952
rect 12434 16940 12440 16952
rect 12492 16940 12498 16992
rect 14274 16940 14280 16992
rect 14332 16940 14338 16992
rect 15197 16983 15255 16989
rect 15197 16949 15209 16983
rect 15243 16980 15255 16983
rect 15378 16980 15384 16992
rect 15243 16952 15384 16980
rect 15243 16949 15255 16952
rect 15197 16943 15255 16949
rect 15378 16940 15384 16952
rect 15436 16980 15442 16992
rect 15654 16980 15660 16992
rect 15436 16952 15660 16980
rect 15436 16940 15442 16952
rect 15654 16940 15660 16952
rect 15712 16940 15718 16992
rect 15749 16983 15807 16989
rect 15749 16949 15761 16983
rect 15795 16980 15807 16983
rect 16942 16980 16948 16992
rect 15795 16952 16948 16980
rect 15795 16949 15807 16952
rect 15749 16943 15807 16949
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 17313 16983 17371 16989
rect 17313 16949 17325 16983
rect 17359 16980 17371 16983
rect 17494 16980 17500 16992
rect 17359 16952 17500 16980
rect 17359 16949 17371 16952
rect 17313 16943 17371 16949
rect 17494 16940 17500 16952
rect 17552 16940 17558 16992
rect 18598 16940 18604 16992
rect 18656 16980 18662 16992
rect 20364 16980 20392 17020
rect 18656 16952 20392 16980
rect 18656 16940 18662 16952
rect 20438 16940 20444 16992
rect 20496 16940 20502 16992
rect 20548 16980 20576 17020
rect 20993 17051 21051 17057
rect 20993 17017 21005 17051
rect 21039 17048 21051 17051
rect 22296 17048 22324 17079
rect 23198 17076 23204 17088
rect 23256 17076 23262 17128
rect 23477 17119 23535 17125
rect 23477 17085 23489 17119
rect 23523 17116 23535 17119
rect 23566 17116 23572 17128
rect 23523 17088 23572 17116
rect 23523 17085 23535 17088
rect 23477 17079 23535 17085
rect 23566 17076 23572 17088
rect 23624 17076 23630 17128
rect 23845 17119 23903 17125
rect 23845 17085 23857 17119
rect 23891 17116 23903 17119
rect 23934 17116 23940 17128
rect 23891 17088 23940 17116
rect 23891 17085 23903 17088
rect 23845 17079 23903 17085
rect 22830 17048 22836 17060
rect 21039 17020 22836 17048
rect 21039 17017 21051 17020
rect 20993 17011 21051 17017
rect 22830 17008 22836 17020
rect 22888 17048 22894 17060
rect 23860 17048 23888 17079
rect 23934 17076 23940 17088
rect 23992 17076 23998 17128
rect 24228 17116 24256 17147
rect 24394 17144 24400 17156
rect 24452 17144 24458 17196
rect 24949 17187 25007 17193
rect 24949 17153 24961 17187
rect 24995 17184 25007 17187
rect 25148 17184 25176 17280
rect 24995 17156 25176 17184
rect 24995 17153 25007 17156
rect 24949 17147 25007 17153
rect 25406 17144 25412 17196
rect 25464 17144 25470 17196
rect 24136 17088 24256 17116
rect 25133 17119 25191 17125
rect 24136 17060 24164 17088
rect 25133 17085 25145 17119
rect 25179 17116 25191 17119
rect 25976 17116 26004 17280
rect 26326 17212 26332 17264
rect 26384 17252 26390 17264
rect 27448 17252 27476 17283
rect 28166 17280 28172 17292
rect 28224 17320 28230 17332
rect 28534 17320 28540 17332
rect 28224 17292 28540 17320
rect 28224 17280 28230 17292
rect 28534 17280 28540 17292
rect 28592 17280 28598 17332
rect 30561 17323 30619 17329
rect 30561 17289 30573 17323
rect 30607 17289 30619 17323
rect 30561 17283 30619 17289
rect 30101 17255 30159 17261
rect 30101 17252 30113 17255
rect 26384 17224 27476 17252
rect 27540 17224 30113 17252
rect 26384 17212 26390 17224
rect 27341 17187 27399 17193
rect 27341 17184 27353 17187
rect 25179 17088 26004 17116
rect 26068 17156 27353 17184
rect 25179 17085 25191 17088
rect 25133 17079 25191 17085
rect 22888 17020 23888 17048
rect 22888 17008 22894 17020
rect 24118 17008 24124 17060
rect 24176 17008 24182 17060
rect 24581 17051 24639 17057
rect 24581 17017 24593 17051
rect 24627 17048 24639 17051
rect 25041 17051 25099 17057
rect 25041 17048 25053 17051
rect 24627 17020 25053 17048
rect 24627 17017 24639 17020
rect 24581 17011 24639 17017
rect 25041 17017 25053 17020
rect 25087 17017 25099 17051
rect 25041 17011 25099 17017
rect 23198 16980 23204 16992
rect 20548 16952 23204 16980
rect 23198 16940 23204 16952
rect 23256 16940 23262 16992
rect 23842 16940 23848 16992
rect 23900 16980 23906 16992
rect 23937 16983 23995 16989
rect 23937 16980 23949 16983
rect 23900 16952 23949 16980
rect 23900 16940 23906 16952
rect 23937 16949 23949 16952
rect 23983 16949 23995 16983
rect 23937 16943 23995 16949
rect 24762 16940 24768 16992
rect 24820 16980 24826 16992
rect 26068 16980 26096 17156
rect 27341 17153 27353 17156
rect 27387 17184 27399 17187
rect 27540 17184 27568 17224
rect 30101 17221 30113 17224
rect 30147 17252 30159 17255
rect 30466 17252 30472 17264
rect 30147 17224 30472 17252
rect 30147 17221 30159 17224
rect 30101 17215 30159 17221
rect 30466 17212 30472 17224
rect 30524 17212 30530 17264
rect 27387 17156 27568 17184
rect 27387 17153 27399 17156
rect 27341 17147 27399 17153
rect 27982 17144 27988 17196
rect 28040 17184 28046 17196
rect 30193 17187 30251 17193
rect 30193 17184 30205 17187
rect 28040 17156 30205 17184
rect 28040 17144 28046 17156
rect 30193 17153 30205 17156
rect 30239 17153 30251 17187
rect 30576 17184 30604 17283
rect 35161 17255 35219 17261
rect 35161 17221 35173 17255
rect 35207 17252 35219 17255
rect 37734 17252 37740 17264
rect 35207 17224 37740 17252
rect 35207 17221 35219 17224
rect 35161 17215 35219 17221
rect 37734 17212 37740 17224
rect 37792 17212 37798 17264
rect 30653 17187 30711 17193
rect 30653 17184 30665 17187
rect 30576 17156 30665 17184
rect 30193 17147 30251 17153
rect 30653 17153 30665 17156
rect 30699 17153 30711 17187
rect 30653 17147 30711 17153
rect 27522 17076 27528 17128
rect 27580 17076 27586 17128
rect 29917 17119 29975 17125
rect 29917 17085 29929 17119
rect 29963 17085 29975 17119
rect 30208 17116 30236 17147
rect 33134 17144 33140 17196
rect 33192 17144 33198 17196
rect 33226 17144 33232 17196
rect 33284 17184 33290 17196
rect 33413 17187 33471 17193
rect 33413 17184 33425 17187
rect 33284 17156 33425 17184
rect 33284 17144 33290 17156
rect 33413 17153 33425 17156
rect 33459 17153 33471 17187
rect 33413 17147 33471 17153
rect 33689 17187 33747 17193
rect 33689 17153 33701 17187
rect 33735 17184 33747 17187
rect 34333 17187 34391 17193
rect 34333 17184 34345 17187
rect 33735 17156 34345 17184
rect 33735 17153 33747 17156
rect 33689 17147 33747 17153
rect 34333 17153 34345 17156
rect 34379 17153 34391 17187
rect 34333 17147 34391 17153
rect 32214 17116 32220 17128
rect 30208 17088 32220 17116
rect 29917 17079 29975 17085
rect 26142 17008 26148 17060
rect 26200 17048 26206 17060
rect 29932 17048 29960 17079
rect 32214 17076 32220 17088
rect 32272 17076 32278 17128
rect 33152 17116 33180 17144
rect 33704 17116 33732 17147
rect 33152 17088 33732 17116
rect 33962 17076 33968 17128
rect 34020 17076 34026 17128
rect 26200 17020 29960 17048
rect 26200 17008 26206 17020
rect 24820 16952 26096 16980
rect 30837 16983 30895 16989
rect 24820 16940 24826 16952
rect 30837 16949 30849 16983
rect 30883 16980 30895 16983
rect 30926 16980 30932 16992
rect 30883 16952 30932 16980
rect 30883 16949 30895 16952
rect 30837 16943 30895 16949
rect 30926 16940 30932 16952
rect 30984 16940 30990 16992
rect 33042 16940 33048 16992
rect 33100 16980 33106 16992
rect 33229 16983 33287 16989
rect 33229 16980 33241 16983
rect 33100 16952 33241 16980
rect 33100 16940 33106 16952
rect 33229 16949 33241 16952
rect 33275 16949 33287 16983
rect 33229 16943 33287 16949
rect 1104 16890 38272 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38272 16890
rect 1104 16816 38272 16838
rect 10594 16776 10600 16788
rect 8956 16748 10600 16776
rect 8956 16708 8984 16748
rect 10594 16736 10600 16748
rect 10652 16776 10658 16788
rect 10652 16748 11008 16776
rect 10652 16736 10658 16748
rect 7760 16680 8340 16708
rect 7760 16652 7788 16680
rect 1854 16600 1860 16652
rect 1912 16600 1918 16652
rect 2133 16643 2191 16649
rect 2133 16609 2145 16643
rect 2179 16640 2191 16643
rect 2498 16640 2504 16652
rect 2179 16612 2504 16640
rect 2179 16609 2191 16612
rect 2133 16603 2191 16609
rect 2498 16600 2504 16612
rect 2556 16600 2562 16652
rect 4798 16600 4804 16652
rect 4856 16640 4862 16652
rect 4893 16643 4951 16649
rect 4893 16640 4905 16643
rect 4856 16612 4905 16640
rect 4856 16600 4862 16612
rect 4893 16609 4905 16612
rect 4939 16609 4951 16643
rect 4893 16603 4951 16609
rect 5534 16600 5540 16652
rect 5592 16640 5598 16652
rect 6917 16643 6975 16649
rect 6917 16640 6929 16643
rect 5592 16612 6929 16640
rect 5592 16600 5598 16612
rect 6917 16609 6929 16612
rect 6963 16609 6975 16643
rect 7098 16640 7104 16652
rect 6917 16603 6975 16609
rect 7024 16612 7104 16640
rect 3234 16532 3240 16584
rect 3292 16572 3298 16584
rect 6825 16575 6883 16581
rect 3292 16544 6224 16572
rect 3292 16532 3298 16544
rect 6196 16516 6224 16544
rect 6825 16541 6837 16575
rect 6871 16572 6883 16575
rect 7024 16572 7052 16612
rect 7098 16600 7104 16612
rect 7156 16600 7162 16652
rect 7282 16600 7288 16652
rect 7340 16600 7346 16652
rect 7742 16600 7748 16652
rect 7800 16600 7806 16652
rect 8202 16600 8208 16652
rect 8260 16600 8266 16652
rect 8312 16649 8340 16680
rect 8864 16680 8984 16708
rect 8297 16643 8355 16649
rect 8297 16609 8309 16643
rect 8343 16609 8355 16643
rect 8297 16603 8355 16609
rect 6871 16544 7052 16572
rect 6871 16541 6883 16544
rect 6825 16535 6883 16541
rect 7834 16532 7840 16584
rect 7892 16572 7898 16584
rect 8110 16572 8116 16584
rect 7892 16544 8116 16572
rect 7892 16532 7898 16544
rect 8110 16532 8116 16544
rect 8168 16532 8174 16584
rect 4157 16507 4215 16513
rect 4157 16504 4169 16507
rect 3620 16476 4169 16504
rect 3620 16445 3648 16476
rect 4157 16473 4169 16476
rect 4203 16473 4215 16507
rect 4157 16467 4215 16473
rect 6178 16464 6184 16516
rect 6236 16464 6242 16516
rect 7745 16507 7803 16513
rect 7745 16473 7757 16507
rect 7791 16504 7803 16507
rect 8864 16504 8892 16680
rect 9582 16668 9588 16720
rect 9640 16708 9646 16720
rect 9640 16680 10916 16708
rect 9640 16668 9646 16680
rect 9214 16640 9220 16652
rect 8956 16612 9220 16640
rect 8956 16581 8984 16612
rect 9214 16600 9220 16612
rect 9272 16600 9278 16652
rect 9876 16584 9904 16680
rect 10778 16640 10784 16652
rect 10428 16612 10784 16640
rect 10428 16584 10456 16612
rect 10778 16600 10784 16612
rect 10836 16600 10842 16652
rect 8941 16575 8999 16581
rect 8941 16541 8953 16575
rect 8987 16541 8999 16575
rect 8941 16535 8999 16541
rect 9122 16532 9128 16584
rect 9180 16572 9186 16584
rect 9398 16572 9404 16584
rect 9180 16544 9404 16572
rect 9180 16532 9186 16544
rect 9398 16532 9404 16544
rect 9456 16532 9462 16584
rect 9490 16532 9496 16584
rect 9548 16532 9554 16584
rect 9674 16581 9680 16584
rect 9641 16575 9680 16581
rect 9641 16562 9653 16575
rect 9600 16541 9653 16562
rect 9732 16572 9738 16584
rect 9732 16544 9741 16572
rect 9600 16534 9680 16541
rect 9600 16504 9628 16534
rect 9674 16532 9680 16534
rect 9732 16532 9738 16544
rect 9858 16532 9864 16584
rect 9916 16532 9922 16584
rect 9999 16575 10057 16581
rect 9999 16541 10011 16575
rect 10045 16572 10057 16575
rect 10410 16572 10416 16584
rect 10045 16544 10416 16572
rect 10045 16541 10057 16544
rect 9999 16535 10057 16541
rect 10410 16532 10416 16544
rect 10468 16532 10474 16584
rect 10594 16581 10600 16584
rect 10592 16535 10600 16581
rect 10594 16532 10600 16535
rect 10652 16532 10658 16584
rect 10689 16575 10747 16581
rect 10689 16541 10701 16575
rect 10735 16572 10747 16575
rect 10888 16572 10916 16680
rect 10980 16581 11008 16748
rect 12342 16736 12348 16788
rect 12400 16736 12406 16788
rect 15562 16736 15568 16788
rect 15620 16736 15626 16788
rect 17129 16779 17187 16785
rect 17129 16745 17141 16779
rect 17175 16776 17187 16779
rect 17494 16776 17500 16788
rect 17175 16748 17500 16776
rect 17175 16745 17187 16748
rect 17129 16739 17187 16745
rect 17494 16736 17500 16748
rect 17552 16736 17558 16788
rect 18506 16736 18512 16788
rect 18564 16776 18570 16788
rect 18874 16776 18880 16788
rect 18564 16748 18880 16776
rect 18564 16736 18570 16748
rect 18874 16736 18880 16748
rect 18932 16736 18938 16788
rect 23474 16736 23480 16788
rect 23532 16776 23538 16788
rect 24762 16776 24768 16788
rect 23532 16748 24768 16776
rect 23532 16736 23538 16748
rect 24762 16736 24768 16748
rect 24820 16736 24826 16788
rect 24946 16736 24952 16788
rect 25004 16776 25010 16788
rect 26973 16779 27031 16785
rect 25004 16748 25912 16776
rect 25004 16736 25010 16748
rect 11606 16668 11612 16720
rect 11664 16708 11670 16720
rect 15580 16708 15608 16736
rect 11664 16680 15608 16708
rect 17313 16711 17371 16717
rect 11664 16668 11670 16680
rect 11072 16612 12388 16640
rect 11072 16584 11100 16612
rect 12360 16584 12388 16612
rect 10735 16544 10916 16572
rect 10735 16541 10747 16544
rect 10689 16535 10747 16541
rect 7791 16476 8892 16504
rect 9048 16476 9628 16504
rect 9769 16507 9827 16513
rect 7791 16473 7803 16476
rect 7745 16467 7803 16473
rect 3605 16439 3663 16445
rect 3605 16405 3617 16439
rect 3651 16405 3663 16439
rect 3605 16399 3663 16405
rect 6362 16396 6368 16448
rect 6420 16396 6426 16448
rect 6730 16396 6736 16448
rect 6788 16396 6794 16448
rect 7650 16396 7656 16448
rect 7708 16436 7714 16448
rect 9048 16436 9076 16476
rect 9769 16473 9781 16507
rect 9815 16504 9827 16507
rect 10781 16507 10839 16513
rect 10781 16504 10793 16507
rect 9815 16476 10793 16504
rect 9815 16473 9827 16476
rect 9769 16467 9827 16473
rect 10781 16473 10793 16476
rect 10827 16473 10839 16507
rect 10888 16504 10916 16544
rect 10964 16575 11022 16581
rect 10964 16541 10976 16575
rect 11010 16541 11022 16575
rect 10964 16535 11022 16541
rect 11054 16532 11060 16584
rect 11112 16532 11118 16584
rect 11698 16532 11704 16584
rect 11756 16532 11762 16584
rect 12250 16532 12256 16584
rect 12308 16532 12314 16584
rect 12342 16532 12348 16584
rect 12400 16532 12406 16584
rect 12452 16581 12480 16680
rect 17313 16677 17325 16711
rect 17359 16708 17371 16711
rect 17954 16708 17960 16720
rect 17359 16680 17960 16708
rect 17359 16677 17371 16680
rect 17313 16671 17371 16677
rect 17954 16668 17960 16680
rect 18012 16668 18018 16720
rect 18690 16668 18696 16720
rect 18748 16708 18754 16720
rect 18748 16680 20760 16708
rect 18748 16668 18754 16680
rect 14277 16643 14335 16649
rect 14277 16609 14289 16643
rect 14323 16640 14335 16643
rect 15378 16640 15384 16652
rect 14323 16612 15384 16640
rect 14323 16609 14335 16612
rect 14277 16603 14335 16609
rect 15378 16600 15384 16612
rect 15436 16640 15442 16652
rect 18141 16643 18199 16649
rect 15436 16612 15884 16640
rect 15436 16600 15442 16612
rect 15856 16584 15884 16612
rect 17420 16612 18092 16640
rect 17420 16584 17448 16612
rect 12437 16575 12495 16581
rect 12437 16541 12449 16575
rect 12483 16541 12495 16575
rect 12437 16535 12495 16541
rect 13446 16532 13452 16584
rect 13504 16532 13510 16584
rect 13538 16532 13544 16584
rect 13596 16532 13602 16584
rect 14366 16572 14372 16584
rect 13740 16544 14372 16572
rect 11716 16504 11744 16532
rect 12268 16504 12296 16532
rect 10888 16476 11008 16504
rect 11716 16476 12296 16504
rect 13464 16504 13492 16532
rect 13740 16513 13768 16544
rect 14366 16532 14372 16544
rect 14424 16532 14430 16584
rect 14458 16532 14464 16584
rect 14516 16572 14522 16584
rect 14740 16575 14798 16581
rect 14740 16572 14752 16575
rect 14516 16544 14752 16572
rect 14516 16532 14522 16544
rect 14740 16541 14752 16544
rect 14786 16541 14798 16575
rect 14740 16535 14798 16541
rect 15838 16532 15844 16584
rect 15896 16532 15902 16584
rect 17402 16572 17408 16584
rect 16960 16544 17408 16572
rect 16960 16516 16988 16544
rect 17402 16532 17408 16544
rect 17460 16532 17466 16584
rect 17681 16575 17739 16581
rect 17681 16541 17693 16575
rect 17727 16541 17739 16575
rect 18064 16572 18092 16612
rect 18141 16609 18153 16643
rect 18187 16640 18199 16643
rect 19978 16640 19984 16652
rect 18187 16612 19984 16640
rect 18187 16609 18199 16612
rect 18141 16603 18199 16609
rect 19978 16600 19984 16612
rect 20036 16600 20042 16652
rect 20732 16640 20760 16680
rect 20806 16668 20812 16720
rect 20864 16708 20870 16720
rect 22557 16711 22615 16717
rect 22557 16708 22569 16711
rect 20864 16680 22569 16708
rect 20864 16668 20870 16680
rect 22557 16677 22569 16680
rect 22603 16677 22615 16711
rect 22557 16671 22615 16677
rect 21821 16643 21879 16649
rect 21821 16640 21833 16643
rect 20732 16612 21833 16640
rect 21821 16609 21833 16612
rect 21867 16609 21879 16643
rect 21821 16603 21879 16609
rect 22204 16612 22600 16640
rect 18693 16575 18751 16581
rect 18064 16544 18552 16572
rect 17681 16535 17739 16541
rect 13725 16507 13783 16513
rect 13725 16504 13737 16507
rect 13464 16476 13737 16504
rect 10781 16467 10839 16473
rect 7708 16408 9076 16436
rect 9125 16439 9183 16445
rect 7708 16396 7714 16408
rect 9125 16405 9137 16439
rect 9171 16436 9183 16439
rect 9398 16436 9404 16448
rect 9171 16408 9404 16436
rect 9171 16405 9183 16408
rect 9125 16399 9183 16405
rect 9398 16396 9404 16408
rect 9456 16436 9462 16448
rect 9784 16436 9812 16467
rect 9456 16408 9812 16436
rect 9456 16396 9462 16408
rect 10134 16396 10140 16448
rect 10192 16396 10198 16448
rect 10226 16396 10232 16448
rect 10284 16436 10290 16448
rect 10413 16439 10471 16445
rect 10413 16436 10425 16439
rect 10284 16408 10425 16436
rect 10284 16396 10290 16408
rect 10413 16405 10425 16408
rect 10459 16405 10471 16439
rect 10980 16436 11008 16476
rect 13725 16473 13737 16476
rect 13771 16473 13783 16507
rect 13725 16467 13783 16473
rect 14642 16464 14648 16516
rect 14700 16504 14706 16516
rect 14700 16476 14780 16504
rect 14700 16464 14706 16476
rect 11974 16436 11980 16448
rect 10980 16408 11980 16436
rect 10413 16399 10471 16405
rect 11974 16396 11980 16408
rect 12032 16396 12038 16448
rect 13906 16396 13912 16448
rect 13964 16396 13970 16448
rect 14752 16445 14780 16476
rect 16942 16464 16948 16516
rect 17000 16464 17006 16516
rect 17218 16513 17224 16516
rect 17161 16507 17224 16513
rect 17161 16473 17173 16507
rect 17207 16473 17224 16507
rect 17161 16467 17224 16473
rect 17218 16464 17224 16467
rect 17276 16504 17282 16516
rect 17696 16504 17724 16535
rect 17276 16476 17724 16504
rect 17773 16507 17831 16513
rect 17276 16464 17282 16476
rect 17773 16473 17785 16507
rect 17819 16504 17831 16507
rect 18138 16504 18144 16516
rect 17819 16476 18144 16504
rect 17819 16473 17831 16476
rect 17773 16467 17831 16473
rect 18138 16464 18144 16476
rect 18196 16464 18202 16516
rect 18417 16507 18475 16513
rect 18417 16473 18429 16507
rect 18463 16473 18475 16507
rect 18417 16467 18475 16473
rect 14737 16439 14795 16445
rect 14737 16405 14749 16439
rect 14783 16405 14795 16439
rect 14737 16399 14795 16405
rect 14918 16396 14924 16448
rect 14976 16396 14982 16448
rect 17494 16396 17500 16448
rect 17552 16436 17558 16448
rect 17589 16439 17647 16445
rect 17589 16436 17601 16439
rect 17552 16408 17601 16436
rect 17552 16396 17558 16408
rect 17589 16405 17601 16408
rect 17635 16405 17647 16439
rect 17589 16399 17647 16405
rect 17678 16396 17684 16448
rect 17736 16436 17742 16448
rect 18432 16436 18460 16467
rect 17736 16408 18460 16436
rect 18524 16436 18552 16544
rect 18693 16541 18705 16575
rect 18739 16572 18751 16575
rect 19426 16572 19432 16584
rect 18739 16544 19432 16572
rect 18739 16541 18751 16544
rect 18693 16535 18751 16541
rect 19426 16532 19432 16544
rect 19484 16532 19490 16584
rect 22094 16572 22100 16584
rect 22055 16544 22100 16572
rect 22094 16532 22100 16544
rect 22152 16532 22158 16584
rect 22204 16581 22232 16612
rect 22572 16584 22600 16612
rect 22646 16600 22652 16652
rect 22704 16640 22710 16652
rect 24118 16640 24124 16652
rect 22704 16612 24124 16640
rect 22704 16600 22710 16612
rect 24118 16600 24124 16612
rect 24176 16600 24182 16652
rect 22189 16575 22247 16581
rect 22189 16541 22201 16575
rect 22235 16541 22247 16575
rect 22189 16535 22247 16541
rect 22278 16532 22284 16584
rect 22336 16532 22342 16584
rect 22465 16575 22523 16581
rect 22465 16541 22477 16575
rect 22511 16541 22523 16575
rect 22465 16535 22523 16541
rect 19610 16464 19616 16516
rect 19668 16504 19674 16516
rect 20898 16504 20904 16516
rect 19668 16476 20904 16504
rect 19668 16464 19674 16476
rect 20898 16464 20904 16476
rect 20956 16464 20962 16516
rect 22480 16436 22508 16535
rect 22554 16532 22560 16584
rect 22612 16532 22618 16584
rect 22830 16572 22836 16584
rect 22791 16544 22836 16572
rect 22830 16532 22836 16544
rect 22888 16532 22894 16584
rect 22925 16575 22983 16581
rect 22925 16541 22937 16575
rect 22971 16541 22983 16575
rect 22925 16535 22983 16541
rect 22572 16504 22600 16532
rect 22940 16504 22968 16535
rect 23014 16532 23020 16584
rect 23072 16532 23078 16584
rect 23198 16532 23204 16584
rect 23256 16532 23262 16584
rect 25884 16572 25912 16748
rect 26973 16745 26985 16779
rect 27019 16776 27031 16779
rect 27062 16776 27068 16788
rect 27019 16748 27068 16776
rect 27019 16745 27031 16748
rect 26973 16739 27031 16745
rect 27062 16736 27068 16748
rect 27120 16736 27126 16788
rect 29546 16736 29552 16788
rect 29604 16776 29610 16788
rect 30742 16776 30748 16788
rect 29604 16748 30748 16776
rect 29604 16736 29610 16748
rect 30742 16736 30748 16748
rect 30800 16736 30806 16788
rect 30926 16785 30932 16788
rect 30916 16779 30932 16785
rect 30916 16745 30928 16779
rect 30916 16739 30932 16745
rect 30926 16736 30932 16739
rect 30984 16736 30990 16788
rect 32214 16736 32220 16788
rect 32272 16776 32278 16788
rect 32401 16779 32459 16785
rect 32401 16776 32413 16779
rect 32272 16748 32413 16776
rect 32272 16736 32278 16748
rect 32401 16745 32413 16748
rect 32447 16745 32459 16779
rect 32401 16739 32459 16745
rect 32600 16748 34008 16776
rect 27614 16600 27620 16652
rect 27672 16640 27678 16652
rect 27672 16612 32076 16640
rect 27672 16600 27678 16612
rect 25961 16575 26019 16581
rect 25961 16572 25973 16575
rect 25884 16544 25973 16572
rect 25961 16541 25973 16544
rect 26007 16541 26019 16575
rect 25961 16535 26019 16541
rect 26326 16532 26332 16584
rect 26384 16572 26390 16584
rect 27154 16572 27160 16584
rect 26384 16544 27160 16572
rect 26384 16532 26390 16544
rect 27154 16532 27160 16544
rect 27212 16532 27218 16584
rect 30377 16575 30435 16581
rect 30377 16541 30389 16575
rect 30423 16541 30435 16575
rect 30377 16535 30435 16541
rect 30469 16575 30527 16581
rect 30469 16541 30481 16575
rect 30515 16572 30527 16575
rect 30653 16575 30711 16581
rect 30653 16572 30665 16575
rect 30515 16544 30665 16572
rect 30515 16541 30527 16544
rect 30469 16535 30527 16541
rect 30653 16541 30665 16544
rect 30699 16541 30711 16575
rect 32048 16572 32076 16612
rect 32600 16572 32628 16748
rect 32953 16643 33011 16649
rect 32953 16609 32965 16643
rect 32999 16640 33011 16643
rect 33042 16640 33048 16652
rect 32999 16612 33048 16640
rect 32999 16609 33011 16612
rect 32953 16603 33011 16609
rect 33042 16600 33048 16612
rect 33100 16600 33106 16652
rect 32048 16558 32628 16572
rect 32062 16544 32628 16558
rect 30653 16535 30711 16541
rect 22572 16476 22968 16504
rect 22646 16436 22652 16448
rect 18524 16408 22652 16436
rect 17736 16396 17742 16408
rect 22646 16396 22652 16408
rect 22704 16396 22710 16448
rect 22738 16396 22744 16448
rect 22796 16436 22802 16448
rect 23032 16436 23060 16532
rect 22796 16408 23060 16436
rect 23216 16436 23244 16532
rect 24118 16464 24124 16516
rect 24176 16504 24182 16516
rect 25682 16504 25688 16516
rect 24176 16476 25688 16504
rect 24176 16464 24182 16476
rect 25682 16464 25688 16476
rect 25740 16504 25746 16516
rect 26145 16507 26203 16513
rect 26145 16504 26157 16507
rect 25740 16476 26157 16504
rect 25740 16464 25746 16476
rect 26145 16473 26157 16476
rect 26191 16473 26203 16507
rect 26145 16467 26203 16473
rect 26237 16507 26295 16513
rect 26237 16473 26249 16507
rect 26283 16504 26295 16507
rect 26418 16504 26424 16516
rect 26283 16476 26424 16504
rect 26283 16473 26295 16476
rect 26237 16467 26295 16473
rect 26418 16464 26424 16476
rect 26476 16464 26482 16516
rect 26605 16507 26663 16513
rect 26605 16504 26617 16507
rect 26528 16476 26617 16504
rect 25498 16436 25504 16448
rect 23216 16408 25504 16436
rect 22796 16396 22802 16408
rect 25498 16396 25504 16408
rect 25556 16396 25562 16448
rect 25866 16396 25872 16448
rect 25924 16436 25930 16448
rect 26326 16436 26332 16448
rect 25924 16408 26332 16436
rect 25924 16396 25930 16408
rect 26326 16396 26332 16408
rect 26384 16396 26390 16448
rect 26528 16445 26556 16476
rect 26605 16473 26617 16476
rect 26651 16473 26663 16507
rect 26605 16467 26663 16473
rect 26786 16464 26792 16516
rect 26844 16464 26850 16516
rect 29178 16464 29184 16516
rect 29236 16504 29242 16516
rect 30098 16504 30104 16516
rect 29236 16476 30104 16504
rect 29236 16464 29242 16476
rect 30098 16464 30104 16476
rect 30156 16464 30162 16516
rect 30392 16504 30420 16535
rect 32674 16532 32680 16584
rect 32732 16532 32738 16584
rect 33980 16516 34008 16748
rect 30392 16476 31156 16504
rect 31128 16448 31156 16476
rect 33962 16464 33968 16516
rect 34020 16464 34026 16516
rect 26513 16439 26571 16445
rect 26513 16405 26525 16439
rect 26559 16405 26571 16439
rect 26513 16399 26571 16405
rect 27890 16396 27896 16448
rect 27948 16436 27954 16448
rect 30190 16436 30196 16448
rect 27948 16408 30196 16436
rect 27948 16396 27954 16408
rect 30190 16396 30196 16408
rect 30248 16396 30254 16448
rect 31110 16396 31116 16448
rect 31168 16396 31174 16448
rect 34422 16396 34428 16448
rect 34480 16396 34486 16448
rect 1104 16346 38272 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 38272 16346
rect 1104 16272 38272 16294
rect 1949 16235 2007 16241
rect 1949 16232 1961 16235
rect 1780 16204 1961 16232
rect 934 16124 940 16176
rect 992 16164 998 16176
rect 1780 16173 1808 16204
rect 1949 16201 1961 16204
rect 1995 16201 2007 16235
rect 1949 16195 2007 16201
rect 3970 16192 3976 16244
rect 4028 16192 4034 16244
rect 6362 16192 6368 16244
rect 6420 16192 6426 16244
rect 7282 16192 7288 16244
rect 7340 16192 7346 16244
rect 7837 16235 7895 16241
rect 7837 16201 7849 16235
rect 7883 16232 7895 16235
rect 7926 16232 7932 16244
rect 7883 16204 7932 16232
rect 7883 16201 7895 16204
rect 7837 16195 7895 16201
rect 7926 16192 7932 16204
rect 7984 16192 7990 16244
rect 8573 16235 8631 16241
rect 8573 16201 8585 16235
rect 8619 16232 8631 16235
rect 9214 16232 9220 16244
rect 8619 16204 9220 16232
rect 8619 16201 8631 16204
rect 8573 16195 8631 16201
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 9950 16232 9956 16244
rect 9554 16204 9956 16232
rect 1397 16167 1455 16173
rect 1397 16164 1409 16167
rect 992 16136 1409 16164
rect 992 16124 998 16136
rect 1397 16133 1409 16136
rect 1443 16133 1455 16167
rect 1397 16127 1455 16133
rect 1765 16167 1823 16173
rect 1765 16133 1777 16167
rect 1811 16133 1823 16167
rect 1765 16127 1823 16133
rect 2133 16099 2191 16105
rect 2133 16065 2145 16099
rect 2179 16065 2191 16099
rect 2133 16059 2191 16065
rect 3881 16099 3939 16105
rect 3881 16065 3893 16099
rect 3927 16096 3939 16099
rect 3988 16096 4016 16192
rect 3927 16068 4016 16096
rect 5445 16099 5503 16105
rect 3927 16065 3939 16068
rect 3881 16059 3939 16065
rect 5445 16065 5457 16099
rect 5491 16096 5503 16099
rect 6380 16096 6408 16192
rect 7300 16164 7328 16192
rect 9554 16164 9582 16204
rect 9692 16173 9720 16204
rect 9950 16192 9956 16204
rect 10008 16232 10014 16244
rect 10229 16235 10287 16241
rect 10229 16232 10241 16235
rect 10008 16204 10241 16232
rect 10008 16192 10014 16204
rect 10229 16201 10241 16204
rect 10275 16232 10287 16235
rect 11606 16232 11612 16244
rect 10275 16204 11612 16232
rect 10275 16201 10287 16204
rect 10229 16195 10287 16201
rect 11606 16192 11612 16204
rect 11664 16192 11670 16244
rect 11974 16192 11980 16244
rect 12032 16192 12038 16244
rect 12342 16192 12348 16244
rect 12400 16232 12406 16244
rect 13998 16232 14004 16244
rect 12400 16204 14004 16232
rect 12400 16192 12406 16204
rect 7208 16136 7328 16164
rect 7576 16136 9582 16164
rect 9677 16167 9735 16173
rect 7208 16105 7236 16136
rect 5491 16068 6408 16096
rect 7193 16099 7251 16105
rect 5491 16065 5503 16068
rect 5445 16059 5503 16065
rect 7193 16065 7205 16099
rect 7239 16065 7251 16099
rect 7193 16059 7251 16065
rect 7285 16099 7343 16105
rect 7285 16065 7297 16099
rect 7331 16096 7343 16099
rect 7576 16096 7604 16136
rect 9677 16133 9689 16167
rect 9723 16133 9735 16167
rect 9677 16127 9735 16133
rect 9766 16124 9772 16176
rect 9824 16124 9830 16176
rect 10686 16164 10692 16176
rect 10152 16136 10692 16164
rect 7331 16068 7604 16096
rect 7331 16065 7343 16068
rect 7285 16059 7343 16065
rect 2148 15960 2176 16059
rect 7650 16056 7656 16108
rect 7708 16056 7714 16108
rect 7742 16056 7748 16108
rect 7800 16056 7806 16108
rect 8110 16056 8116 16108
rect 8168 16096 8174 16108
rect 8168 16068 8340 16096
rect 8168 16056 8174 16068
rect 7760 16028 7788 16056
rect 8312 16037 8340 16068
rect 8386 16056 8392 16108
rect 8444 16056 8450 16108
rect 9398 16056 9404 16108
rect 9456 16086 9462 16108
rect 9560 16099 9618 16105
rect 9560 16096 9572 16099
rect 9556 16094 9572 16096
rect 9554 16086 9572 16094
rect 9456 16065 9572 16086
rect 9606 16065 9618 16099
rect 9456 16059 9618 16065
rect 9456 16058 9582 16059
rect 9456 16056 9462 16058
rect 9858 16056 9864 16108
rect 9916 16105 9922 16108
rect 10152 16105 10180 16136
rect 10686 16124 10692 16136
rect 10744 16124 10750 16176
rect 9916 16099 9955 16105
rect 9943 16065 9955 16099
rect 9916 16059 9955 16065
rect 10045 16099 10103 16105
rect 10045 16065 10057 16099
rect 10091 16065 10103 16099
rect 10045 16059 10103 16065
rect 10137 16099 10195 16105
rect 10137 16065 10149 16099
rect 10183 16065 10195 16099
rect 10137 16059 10195 16065
rect 9916 16056 9922 16059
rect 7929 16031 7987 16037
rect 7929 16028 7941 16031
rect 7760 16000 7941 16028
rect 7929 15997 7941 16000
rect 7975 15997 7987 16031
rect 7929 15991 7987 15997
rect 8297 16031 8355 16037
rect 8297 15997 8309 16031
rect 8343 15997 8355 16031
rect 8297 15991 8355 15997
rect 9674 15988 9680 16040
rect 9732 16028 9738 16040
rect 10060 16028 10088 16059
rect 10410 16056 10416 16108
rect 10468 16056 10474 16108
rect 10594 16056 10600 16108
rect 10652 16056 10658 16108
rect 11054 16056 11060 16108
rect 11112 16056 11118 16108
rect 11992 16096 12020 16192
rect 12544 16105 12572 16204
rect 13998 16192 14004 16204
rect 14056 16192 14062 16244
rect 14274 16192 14280 16244
rect 14332 16232 14338 16244
rect 14458 16232 14464 16244
rect 14332 16204 14464 16232
rect 14332 16192 14338 16204
rect 14458 16192 14464 16204
rect 14516 16232 14522 16244
rect 15378 16232 15384 16244
rect 14516 16204 15384 16232
rect 14516 16192 14522 16204
rect 15378 16192 15384 16204
rect 15436 16192 15442 16244
rect 17586 16192 17592 16244
rect 17644 16232 17650 16244
rect 19610 16232 19616 16244
rect 17644 16204 19616 16232
rect 17644 16192 17650 16204
rect 19610 16192 19616 16204
rect 19668 16192 19674 16244
rect 19702 16192 19708 16244
rect 19760 16192 19766 16244
rect 20640 16204 21588 16232
rect 12618 16124 12624 16176
rect 12676 16164 12682 16176
rect 15654 16164 15660 16176
rect 12676 16136 15660 16164
rect 12676 16124 12682 16136
rect 12728 16105 12756 16136
rect 15654 16124 15660 16136
rect 15712 16164 15718 16176
rect 19334 16164 19340 16176
rect 15712 16136 16068 16164
rect 15712 16124 15718 16136
rect 12345 16099 12403 16105
rect 12345 16096 12357 16099
rect 11992 16068 12357 16096
rect 12345 16065 12357 16068
rect 12391 16065 12403 16099
rect 12345 16059 12403 16065
rect 12529 16099 12587 16105
rect 12529 16065 12541 16099
rect 12575 16065 12587 16099
rect 12529 16059 12587 16065
rect 12713 16099 12771 16105
rect 12713 16065 12725 16099
rect 12759 16065 12771 16099
rect 12713 16059 12771 16065
rect 12805 16099 12863 16105
rect 12805 16065 12817 16099
rect 12851 16065 12863 16099
rect 12805 16059 12863 16065
rect 11072 16028 11100 16056
rect 12820 16028 12848 16059
rect 12986 16056 12992 16108
rect 13044 16096 13050 16108
rect 13173 16099 13231 16105
rect 13173 16096 13185 16099
rect 13044 16068 13185 16096
rect 13044 16056 13050 16068
rect 13173 16065 13185 16068
rect 13219 16096 13231 16099
rect 13262 16096 13268 16108
rect 13219 16068 13268 16096
rect 13219 16065 13231 16068
rect 13173 16059 13231 16065
rect 13262 16056 13268 16068
rect 13320 16056 13326 16108
rect 13354 16056 13360 16108
rect 13412 16056 13418 16108
rect 13906 16056 13912 16108
rect 13964 16096 13970 16108
rect 14274 16096 14280 16108
rect 13964 16068 14280 16096
rect 13964 16056 13970 16068
rect 14274 16056 14280 16068
rect 14332 16096 14338 16108
rect 14369 16099 14427 16105
rect 14369 16096 14381 16099
rect 14332 16068 14381 16096
rect 14332 16056 14338 16068
rect 14369 16065 14381 16068
rect 14415 16065 14427 16099
rect 14921 16099 14979 16105
rect 14921 16096 14933 16099
rect 14369 16059 14427 16065
rect 14476 16068 14933 16096
rect 9732 16000 11100 16028
rect 12452 16000 12848 16028
rect 13817 16031 13875 16037
rect 9732 15988 9738 16000
rect 12452 15972 12480 16000
rect 13817 15997 13829 16031
rect 13863 16028 13875 16031
rect 14090 16028 14096 16040
rect 13863 16000 14096 16028
rect 13863 15997 13875 16000
rect 13817 15991 13875 15997
rect 14090 15988 14096 16000
rect 14148 15988 14154 16040
rect 14182 15988 14188 16040
rect 14240 15988 14246 16040
rect 9858 15960 9864 15972
rect 2148 15932 9864 15960
rect 9858 15920 9864 15932
rect 9916 15920 9922 15972
rect 12434 15920 12440 15972
rect 12492 15920 12498 15972
rect 14476 15960 14504 16068
rect 14921 16065 14933 16068
rect 14967 16065 14979 16099
rect 14921 16059 14979 16065
rect 15749 16099 15807 16105
rect 15749 16065 15761 16099
rect 15795 16096 15807 16099
rect 15930 16096 15936 16108
rect 15795 16068 15936 16096
rect 15795 16065 15807 16068
rect 15749 16059 15807 16065
rect 15930 16056 15936 16068
rect 15988 16056 15994 16108
rect 16040 16105 16068 16136
rect 16132 16136 19340 16164
rect 16025 16099 16083 16105
rect 16025 16065 16037 16099
rect 16071 16065 16083 16099
rect 16025 16059 16083 16065
rect 14737 16031 14795 16037
rect 14737 16028 14749 16031
rect 12912 15932 14504 15960
rect 14568 16000 14749 16028
rect 12912 15904 12940 15932
rect 14568 15904 14596 16000
rect 14737 15997 14749 16000
rect 14783 15997 14795 16031
rect 14737 15991 14795 15997
rect 14826 15988 14832 16040
rect 14884 16028 14890 16040
rect 16132 16028 16160 16136
rect 19334 16124 19340 16136
rect 19392 16124 19398 16176
rect 19536 16136 20576 16164
rect 19536 16108 19564 16136
rect 20548 16108 20576 16136
rect 20640 16108 20668 16204
rect 20732 16136 21496 16164
rect 16206 16056 16212 16108
rect 16264 16056 16270 16108
rect 16485 16099 16543 16105
rect 16485 16065 16497 16099
rect 16531 16096 16543 16099
rect 17218 16096 17224 16108
rect 16531 16068 17224 16096
rect 16531 16065 16543 16068
rect 16485 16059 16543 16065
rect 17218 16056 17224 16068
rect 17276 16056 17282 16108
rect 17494 16056 17500 16108
rect 17552 16056 17558 16108
rect 18049 16099 18107 16105
rect 18049 16065 18061 16099
rect 18095 16096 18107 16099
rect 18598 16096 18604 16108
rect 18095 16068 18604 16096
rect 18095 16065 18107 16068
rect 18049 16059 18107 16065
rect 14884 16000 16160 16028
rect 16224 16028 16252 16056
rect 17310 16028 17316 16040
rect 16224 16000 17316 16028
rect 14884 15988 14890 16000
rect 17310 15988 17316 16000
rect 17368 16028 17374 16040
rect 18064 16028 18092 16059
rect 18598 16056 18604 16068
rect 18656 16056 18662 16108
rect 18785 16099 18843 16105
rect 18785 16065 18797 16099
rect 18831 16065 18843 16099
rect 18785 16059 18843 16065
rect 17368 16000 18092 16028
rect 17368 15988 17374 16000
rect 18322 15988 18328 16040
rect 18380 16028 18386 16040
rect 18509 16031 18567 16037
rect 18509 16028 18521 16031
rect 18380 16000 18521 16028
rect 18380 15988 18386 16000
rect 18509 15997 18521 16000
rect 18555 15997 18567 16031
rect 18509 15991 18567 15997
rect 14645 15963 14703 15969
rect 14645 15929 14657 15963
rect 14691 15960 14703 15963
rect 15562 15960 15568 15972
rect 14691 15932 15568 15960
rect 14691 15929 14703 15932
rect 14645 15923 14703 15929
rect 15562 15920 15568 15932
rect 15620 15920 15626 15972
rect 15838 15920 15844 15972
rect 15896 15920 15902 15972
rect 18141 15963 18199 15969
rect 18141 15929 18153 15963
rect 18187 15960 18199 15963
rect 18800 15960 18828 16059
rect 19518 16056 19524 16108
rect 19576 16056 19582 16108
rect 19610 16056 19616 16108
rect 19668 16105 19674 16108
rect 19668 16099 19701 16105
rect 19689 16065 19701 16099
rect 20436 16099 20494 16105
rect 20436 16096 20448 16099
rect 19668 16059 19701 16065
rect 19786 16068 20448 16096
rect 19668 16056 19674 16059
rect 19334 15988 19340 16040
rect 19392 16028 19398 16040
rect 19786 16028 19814 16068
rect 20436 16065 20448 16068
rect 20482 16065 20494 16099
rect 20436 16059 20494 16065
rect 19392 16000 19814 16028
rect 19392 15988 19398 16000
rect 19886 15988 19892 16040
rect 19944 15988 19950 16040
rect 20165 16031 20223 16037
rect 20165 15997 20177 16031
rect 20211 15997 20223 16031
rect 20451 16028 20479 16059
rect 20530 16056 20536 16108
rect 20588 16056 20594 16108
rect 20622 16056 20628 16108
rect 20680 16056 20686 16108
rect 20732 16028 20760 16136
rect 20808 16099 20866 16105
rect 20808 16065 20820 16099
rect 20854 16065 20866 16099
rect 20808 16059 20866 16065
rect 20451 16000 20760 16028
rect 20824 16028 20852 16059
rect 20898 16056 20904 16108
rect 20956 16096 20962 16108
rect 21358 16096 21364 16108
rect 20956 16068 21364 16096
rect 20956 16056 20962 16068
rect 21358 16056 21364 16068
rect 21416 16056 21422 16108
rect 20824 16000 20944 16028
rect 20165 15991 20223 15997
rect 18187 15932 18828 15960
rect 18187 15929 18199 15932
rect 18141 15923 18199 15929
rect 4062 15852 4068 15904
rect 4120 15852 4126 15904
rect 5074 15852 5080 15904
rect 5132 15892 5138 15904
rect 5261 15895 5319 15901
rect 5261 15892 5273 15895
rect 5132 15864 5273 15892
rect 5132 15852 5138 15864
rect 5261 15861 5273 15864
rect 5307 15861 5319 15895
rect 5261 15855 5319 15861
rect 7653 15895 7711 15901
rect 7653 15861 7665 15895
rect 7699 15892 7711 15895
rect 7742 15892 7748 15904
rect 7699 15864 7748 15892
rect 7699 15861 7711 15864
rect 7653 15855 7711 15861
rect 7742 15852 7748 15864
rect 7800 15852 7806 15904
rect 9401 15895 9459 15901
rect 9401 15861 9413 15895
rect 9447 15892 9459 15895
rect 9766 15892 9772 15904
rect 9447 15864 9772 15892
rect 9447 15861 9459 15864
rect 9401 15855 9459 15861
rect 9766 15852 9772 15864
rect 9824 15852 9830 15904
rect 9950 15852 9956 15904
rect 10008 15892 10014 15904
rect 10870 15892 10876 15904
rect 10008 15864 10876 15892
rect 10008 15852 10014 15864
rect 10870 15852 10876 15864
rect 10928 15852 10934 15904
rect 12894 15852 12900 15904
rect 12952 15852 12958 15904
rect 13630 15852 13636 15904
rect 13688 15892 13694 15904
rect 14550 15892 14556 15904
rect 13688 15864 14556 15892
rect 13688 15852 13694 15864
rect 14550 15852 14556 15864
rect 14608 15852 14614 15904
rect 15197 15895 15255 15901
rect 15197 15861 15209 15895
rect 15243 15892 15255 15895
rect 15654 15892 15660 15904
rect 15243 15864 15660 15892
rect 15243 15861 15255 15864
rect 15197 15855 15255 15861
rect 15654 15852 15660 15864
rect 15712 15852 15718 15904
rect 18800 15892 18828 15932
rect 19521 15963 19579 15969
rect 19521 15929 19533 15963
rect 19567 15960 19579 15963
rect 19904 15960 19932 15988
rect 19567 15932 19932 15960
rect 19567 15929 19579 15932
rect 19521 15923 19579 15929
rect 20070 15920 20076 15972
rect 20128 15920 20134 15972
rect 20180 15960 20208 15991
rect 20257 15963 20315 15969
rect 20257 15960 20269 15963
rect 20180 15932 20269 15960
rect 20257 15929 20269 15932
rect 20303 15929 20315 15963
rect 20257 15923 20315 15929
rect 20916 15904 20944 16000
rect 21468 15960 21496 16136
rect 21560 16028 21588 16204
rect 22370 16192 22376 16244
rect 22428 16232 22434 16244
rect 22557 16235 22615 16241
rect 22557 16232 22569 16235
rect 22428 16204 22569 16232
rect 22428 16192 22434 16204
rect 22557 16201 22569 16204
rect 22603 16201 22615 16235
rect 22557 16195 22615 16201
rect 24118 16192 24124 16244
rect 24176 16192 24182 16244
rect 24394 16232 24400 16244
rect 24228 16204 24400 16232
rect 21634 16124 21640 16176
rect 21692 16164 21698 16176
rect 24136 16164 24164 16192
rect 21692 16136 22416 16164
rect 21692 16124 21698 16136
rect 22094 16056 22100 16108
rect 22152 16056 22158 16108
rect 22186 16056 22192 16108
rect 22244 16056 22250 16108
rect 22388 16105 22416 16136
rect 24044 16136 24164 16164
rect 22373 16099 22431 16105
rect 22373 16065 22385 16099
rect 22419 16096 22431 16099
rect 23750 16096 23756 16108
rect 22419 16068 23756 16096
rect 22419 16065 22431 16068
rect 22373 16059 22431 16065
rect 23750 16056 23756 16068
rect 23808 16056 23814 16108
rect 24044 16105 24072 16136
rect 24228 16105 24256 16204
rect 24394 16192 24400 16204
rect 24452 16192 24458 16244
rect 25038 16192 25044 16244
rect 25096 16232 25102 16244
rect 25225 16235 25283 16241
rect 25225 16232 25237 16235
rect 25096 16204 25237 16232
rect 25096 16192 25102 16204
rect 25225 16201 25237 16204
rect 25271 16201 25283 16235
rect 25225 16195 25283 16201
rect 26421 16235 26479 16241
rect 26421 16201 26433 16235
rect 26467 16232 26479 16235
rect 26786 16232 26792 16244
rect 26467 16204 26792 16232
rect 26467 16201 26479 16204
rect 26421 16195 26479 16201
rect 26786 16192 26792 16204
rect 26844 16192 26850 16244
rect 27430 16192 27436 16244
rect 27488 16232 27494 16244
rect 29822 16232 29828 16244
rect 27488 16204 29828 16232
rect 27488 16192 27494 16204
rect 29822 16192 29828 16204
rect 29880 16192 29886 16244
rect 30024 16204 30328 16232
rect 24670 16164 24676 16176
rect 24320 16136 24676 16164
rect 24320 16105 24348 16136
rect 24670 16124 24676 16136
rect 24728 16164 24734 16176
rect 24728 16136 26285 16164
rect 24728 16124 24734 16136
rect 24029 16099 24087 16105
rect 24029 16065 24041 16099
rect 24075 16065 24087 16099
rect 24029 16059 24087 16065
rect 24177 16099 24256 16105
rect 24177 16065 24189 16099
rect 24223 16068 24256 16099
rect 24305 16099 24363 16105
rect 24223 16065 24235 16068
rect 24177 16059 24235 16065
rect 24305 16065 24317 16099
rect 24351 16065 24363 16099
rect 24305 16059 24363 16065
rect 24397 16099 24455 16105
rect 24397 16065 24409 16099
rect 24443 16065 24455 16099
rect 24397 16059 24455 16065
rect 24320 16028 24348 16059
rect 21560 16000 24348 16028
rect 24118 15960 24124 15972
rect 21468 15932 24124 15960
rect 24118 15920 24124 15932
rect 24176 15920 24182 15972
rect 24302 15920 24308 15972
rect 24360 15960 24366 15972
rect 24412 15960 24440 16059
rect 24486 16056 24492 16108
rect 24544 16105 24550 16108
rect 24544 16096 24552 16105
rect 24765 16099 24823 16105
rect 24544 16068 24589 16096
rect 24544 16059 24552 16068
rect 24765 16065 24777 16099
rect 24811 16065 24823 16099
rect 24765 16059 24823 16065
rect 24857 16099 24915 16105
rect 24857 16065 24869 16099
rect 24903 16096 24915 16099
rect 24903 16068 24992 16096
rect 24903 16065 24915 16068
rect 24857 16059 24915 16065
rect 24544 16056 24550 16059
rect 24780 15960 24808 16059
rect 24964 16040 24992 16068
rect 25038 16056 25044 16108
rect 25096 16056 25102 16108
rect 25130 16056 25136 16108
rect 25188 16096 25194 16108
rect 25774 16096 25780 16108
rect 25188 16068 25780 16096
rect 25188 16056 25194 16068
rect 25774 16056 25780 16068
rect 25832 16056 25838 16108
rect 25958 16105 25964 16108
rect 25925 16099 25964 16105
rect 25925 16065 25937 16099
rect 25925 16059 25964 16065
rect 25958 16056 25964 16059
rect 26016 16056 26022 16108
rect 26257 16105 26285 16136
rect 26326 16124 26332 16176
rect 26384 16164 26390 16176
rect 28534 16164 28540 16176
rect 26384 16136 28540 16164
rect 26384 16124 26390 16136
rect 28534 16124 28540 16136
rect 28592 16124 28598 16176
rect 30024 16164 30052 16204
rect 29564 16136 30052 16164
rect 26053 16099 26111 16105
rect 26053 16065 26065 16099
rect 26099 16065 26111 16099
rect 26053 16059 26111 16065
rect 26145 16099 26203 16105
rect 26145 16065 26157 16099
rect 26191 16065 26203 16099
rect 26145 16059 26203 16065
rect 26242 16099 26300 16105
rect 26242 16065 26254 16099
rect 26288 16065 26300 16099
rect 26242 16059 26300 16065
rect 24946 15988 24952 16040
rect 25004 15988 25010 16040
rect 25866 15960 25872 15972
rect 24360 15932 24440 15960
rect 24504 15932 25872 15960
rect 24360 15920 24366 15932
rect 19610 15892 19616 15904
rect 18800 15864 19616 15892
rect 19610 15852 19616 15864
rect 19668 15892 19674 15904
rect 19794 15892 19800 15904
rect 19668 15864 19800 15892
rect 19668 15852 19674 15864
rect 19794 15852 19800 15864
rect 19852 15852 19858 15904
rect 20898 15852 20904 15904
rect 20956 15852 20962 15904
rect 21450 15852 21456 15904
rect 21508 15892 21514 15904
rect 24504 15892 24532 15932
rect 25866 15920 25872 15932
rect 25924 15960 25930 15972
rect 26073 15960 26101 16059
rect 26160 16028 26188 16059
rect 26344 16028 26372 16124
rect 27893 16099 27951 16105
rect 27893 16096 27905 16099
rect 26160 16000 26372 16028
rect 26436 16068 27905 16096
rect 25924 15932 26101 15960
rect 25924 15920 25930 15932
rect 26326 15920 26332 15972
rect 26384 15960 26390 15972
rect 26436 15960 26464 16068
rect 27893 16065 27905 16068
rect 27939 16065 27951 16099
rect 27893 16059 27951 16065
rect 28626 16056 28632 16108
rect 28684 16056 28690 16108
rect 29086 16056 29092 16108
rect 29144 16056 29150 16108
rect 29564 16105 29592 16136
rect 30098 16124 30104 16176
rect 30156 16124 30162 16176
rect 30190 16124 30196 16176
rect 30248 16124 30254 16176
rect 30300 16164 30328 16204
rect 32674 16192 32680 16244
rect 32732 16232 32738 16244
rect 32861 16235 32919 16241
rect 32861 16232 32873 16235
rect 32732 16204 32873 16232
rect 32732 16192 32738 16204
rect 32861 16201 32873 16204
rect 32907 16201 32919 16235
rect 32861 16195 32919 16201
rect 33226 16192 33232 16244
rect 33284 16192 33290 16244
rect 33318 16192 33324 16244
rect 33376 16232 33382 16244
rect 33597 16235 33655 16241
rect 33597 16232 33609 16235
rect 33376 16204 33609 16232
rect 33376 16192 33382 16204
rect 33597 16201 33609 16204
rect 33643 16232 33655 16235
rect 33778 16232 33784 16244
rect 33643 16204 33784 16232
rect 33643 16201 33655 16204
rect 33597 16195 33655 16201
rect 33778 16192 33784 16204
rect 33836 16192 33842 16244
rect 34422 16192 34428 16244
rect 34480 16192 34486 16244
rect 31021 16167 31079 16173
rect 31021 16164 31033 16167
rect 30300 16136 31033 16164
rect 31021 16133 31033 16136
rect 31067 16133 31079 16167
rect 31021 16127 31079 16133
rect 33689 16167 33747 16173
rect 33689 16133 33701 16167
rect 33735 16164 33747 16167
rect 34440 16164 34468 16192
rect 33735 16136 34468 16164
rect 33735 16133 33747 16136
rect 33689 16127 33747 16133
rect 29549 16099 29607 16105
rect 29549 16065 29561 16099
rect 29595 16065 29607 16099
rect 29822 16096 29828 16108
rect 29549 16059 29607 16065
rect 29664 16068 29828 16096
rect 26602 15988 26608 16040
rect 26660 16028 26666 16040
rect 26660 16000 27798 16028
rect 26660 15988 26666 16000
rect 26384 15932 26464 15960
rect 27770 15960 27798 16000
rect 27982 15988 27988 16040
rect 28040 15988 28046 16040
rect 28074 15988 28080 16040
rect 28132 16028 28138 16040
rect 29664 16028 29692 16068
rect 29822 16056 29828 16068
rect 29880 16056 29886 16108
rect 30374 16105 30380 16108
rect 29973 16099 30031 16105
rect 29973 16065 29985 16099
rect 30019 16094 30031 16099
rect 30331 16099 30380 16105
rect 30019 16065 30052 16094
rect 29973 16059 30052 16065
rect 30331 16065 30343 16099
rect 30377 16065 30380 16099
rect 30331 16059 30380 16065
rect 28132 16000 29692 16028
rect 30024 16028 30052 16059
rect 30374 16056 30380 16059
rect 30432 16056 30438 16108
rect 30837 16099 30895 16105
rect 30837 16065 30849 16099
rect 30883 16065 30895 16099
rect 30837 16059 30895 16065
rect 30024 16000 30144 16028
rect 28132 15988 28138 16000
rect 28000 15960 28028 15988
rect 27770 15932 28028 15960
rect 26384 15920 26390 15932
rect 28350 15920 28356 15972
rect 28408 15960 28414 15972
rect 28408 15932 29408 15960
rect 28408 15920 28414 15932
rect 21508 15864 24532 15892
rect 24673 15895 24731 15901
rect 21508 15852 21514 15864
rect 24673 15861 24685 15895
rect 24719 15892 24731 15895
rect 25038 15892 25044 15904
rect 24719 15864 25044 15892
rect 24719 15861 24731 15864
rect 24673 15855 24731 15861
rect 25038 15852 25044 15864
rect 25096 15852 25102 15904
rect 25314 15852 25320 15904
rect 25372 15892 25378 15904
rect 27246 15892 27252 15904
rect 25372 15864 27252 15892
rect 25372 15852 25378 15864
rect 27246 15852 27252 15864
rect 27304 15892 27310 15904
rect 27893 15895 27951 15901
rect 27893 15892 27905 15895
rect 27304 15864 27905 15892
rect 27304 15852 27310 15864
rect 27893 15861 27905 15864
rect 27939 15861 27951 15895
rect 27893 15855 27951 15861
rect 28258 15852 28264 15904
rect 28316 15852 28322 15904
rect 28626 15852 28632 15904
rect 28684 15892 28690 15904
rect 29270 15892 29276 15904
rect 28684 15864 29276 15892
rect 28684 15852 28690 15864
rect 29270 15852 29276 15864
rect 29328 15852 29334 15904
rect 29380 15892 29408 15932
rect 29546 15920 29552 15972
rect 29604 15920 29610 15972
rect 30116 15960 30144 16000
rect 30558 15988 30564 16040
rect 30616 15988 30622 16040
rect 30650 15988 30656 16040
rect 30708 16028 30714 16040
rect 30852 16028 30880 16059
rect 32030 16056 32036 16108
rect 32088 16096 32094 16108
rect 32953 16099 33011 16105
rect 32953 16096 32965 16099
rect 32088 16068 32965 16096
rect 32088 16056 32094 16068
rect 32953 16065 32965 16068
rect 32999 16096 33011 16099
rect 33134 16096 33140 16108
rect 32999 16068 33140 16096
rect 32999 16065 33011 16068
rect 32953 16059 33011 16065
rect 33134 16056 33140 16068
rect 33192 16056 33198 16108
rect 30708 16000 30880 16028
rect 30708 15988 30714 16000
rect 33704 15960 33732 16127
rect 33870 15988 33876 16040
rect 33928 15988 33934 16040
rect 30116 15932 33732 15960
rect 30116 15892 30144 15932
rect 29380 15864 30144 15892
rect 30469 15895 30527 15901
rect 30469 15861 30481 15895
rect 30515 15892 30527 15895
rect 30653 15895 30711 15901
rect 30653 15892 30665 15895
rect 30515 15864 30665 15892
rect 30515 15861 30527 15864
rect 30469 15855 30527 15861
rect 30653 15861 30665 15864
rect 30699 15861 30711 15895
rect 30653 15855 30711 15861
rect 1104 15802 38272 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38272 15802
rect 1104 15728 38272 15750
rect 6730 15648 6736 15700
rect 6788 15648 6794 15700
rect 9766 15648 9772 15700
rect 9824 15648 9830 15700
rect 9858 15648 9864 15700
rect 9916 15688 9922 15700
rect 11241 15691 11299 15697
rect 11241 15688 11253 15691
rect 9916 15660 11253 15688
rect 9916 15648 9922 15660
rect 11241 15657 11253 15660
rect 11287 15657 11299 15691
rect 11241 15651 11299 15657
rect 12066 15648 12072 15700
rect 12124 15688 12130 15700
rect 12345 15691 12403 15697
rect 12345 15688 12357 15691
rect 12124 15660 12357 15688
rect 12124 15648 12130 15660
rect 12345 15657 12357 15660
rect 12391 15657 12403 15691
rect 12345 15651 12403 15657
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 12805 15691 12863 15697
rect 12805 15688 12817 15691
rect 12492 15660 12817 15688
rect 12492 15648 12498 15660
rect 12805 15657 12817 15660
rect 12851 15657 12863 15691
rect 12805 15651 12863 15657
rect 12894 15648 12900 15700
rect 12952 15648 12958 15700
rect 19334 15688 19340 15700
rect 14108 15660 16344 15688
rect 6748 15620 6776 15648
rect 14108 15632 14136 15660
rect 13081 15623 13139 15629
rect 6748 15592 12020 15620
rect 4985 15555 5043 15561
rect 4985 15521 4997 15555
rect 5031 15552 5043 15555
rect 5074 15552 5080 15564
rect 5031 15524 5080 15552
rect 5031 15521 5043 15524
rect 4985 15515 5043 15521
rect 5074 15512 5080 15524
rect 5132 15512 5138 15564
rect 6178 15552 6184 15564
rect 6104 15524 6184 15552
rect 3970 15444 3976 15496
rect 4028 15484 4034 15496
rect 4433 15487 4491 15493
rect 4433 15484 4445 15487
rect 4028 15456 4445 15484
rect 4028 15444 4034 15456
rect 4433 15453 4445 15456
rect 4479 15453 4491 15487
rect 4433 15447 4491 15453
rect 4525 15487 4583 15493
rect 4525 15453 4537 15487
rect 4571 15484 4583 15487
rect 4709 15487 4767 15493
rect 4709 15484 4721 15487
rect 4571 15456 4721 15484
rect 4571 15453 4583 15456
rect 4525 15447 4583 15453
rect 4709 15453 4721 15456
rect 4755 15453 4767 15487
rect 6104 15470 6132 15524
rect 6178 15512 6184 15524
rect 6236 15512 6242 15564
rect 6748 15561 6776 15592
rect 6733 15555 6791 15561
rect 6733 15521 6745 15555
rect 6779 15521 6791 15555
rect 6733 15515 6791 15521
rect 8938 15512 8944 15564
rect 8996 15552 9002 15564
rect 9306 15552 9312 15564
rect 8996 15524 9312 15552
rect 8996 15512 9002 15524
rect 9306 15512 9312 15524
rect 9364 15512 9370 15564
rect 9858 15512 9864 15564
rect 9916 15512 9922 15564
rect 10060 15524 10272 15552
rect 4709 15447 4767 15453
rect 6822 15444 6828 15496
rect 6880 15484 6886 15496
rect 7469 15487 7527 15493
rect 7469 15484 7481 15487
rect 6880 15456 7481 15484
rect 6880 15444 6886 15456
rect 7469 15453 7481 15456
rect 7515 15453 7527 15487
rect 7469 15447 7527 15453
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15484 7987 15487
rect 9122 15484 9128 15496
rect 7975 15456 9128 15484
rect 7975 15453 7987 15456
rect 7929 15447 7987 15453
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 9950 15444 9956 15496
rect 10008 15484 10014 15496
rect 10060 15493 10088 15524
rect 10244 15496 10272 15524
rect 11238 15512 11244 15564
rect 11296 15552 11302 15564
rect 11992 15552 12020 15592
rect 13081 15589 13093 15623
rect 13127 15620 13139 15623
rect 13354 15620 13360 15632
rect 13127 15592 13360 15620
rect 13127 15589 13139 15592
rect 13081 15583 13139 15589
rect 13354 15580 13360 15592
rect 13412 15580 13418 15632
rect 13630 15580 13636 15632
rect 13688 15620 13694 15632
rect 14090 15620 14096 15632
rect 13688 15592 14096 15620
rect 13688 15580 13694 15592
rect 14090 15580 14096 15592
rect 14148 15580 14154 15632
rect 14550 15580 14556 15632
rect 14608 15580 14614 15632
rect 14918 15580 14924 15632
rect 14976 15620 14982 15632
rect 16209 15623 16267 15629
rect 16209 15620 16221 15623
rect 14976 15592 16221 15620
rect 14976 15580 14982 15592
rect 16209 15589 16221 15592
rect 16255 15589 16267 15623
rect 16209 15583 16267 15589
rect 12897 15555 12955 15561
rect 11296 15524 11560 15552
rect 11992 15524 12112 15552
rect 11296 15512 11302 15524
rect 10045 15487 10103 15493
rect 10045 15484 10057 15487
rect 10008 15456 10057 15484
rect 10008 15444 10014 15456
rect 10045 15453 10057 15456
rect 10091 15453 10103 15487
rect 10045 15447 10103 15453
rect 10134 15444 10140 15496
rect 10192 15444 10198 15496
rect 10226 15444 10232 15496
rect 10284 15444 10290 15496
rect 11532 15493 11560 15524
rect 12084 15496 12112 15524
rect 12897 15521 12909 15555
rect 12943 15552 12955 15555
rect 12986 15552 12992 15564
rect 12943 15524 12992 15552
rect 12943 15521 12955 15524
rect 12897 15515 12955 15521
rect 12986 15512 12992 15524
rect 13044 15512 13050 15564
rect 14182 15512 14188 15564
rect 14240 15512 14246 15564
rect 11425 15487 11483 15493
rect 11425 15453 11437 15487
rect 11471 15453 11483 15487
rect 11425 15447 11483 15453
rect 11517 15487 11575 15493
rect 11517 15453 11529 15487
rect 11563 15453 11575 15487
rect 11517 15447 11575 15453
rect 9769 15419 9827 15425
rect 9769 15385 9781 15419
rect 9815 15416 9827 15419
rect 10152 15416 10180 15444
rect 9815 15388 10180 15416
rect 9815 15385 9827 15388
rect 9769 15379 9827 15385
rect 7190 15308 7196 15360
rect 7248 15348 7254 15360
rect 7377 15351 7435 15357
rect 7377 15348 7389 15351
rect 7248 15320 7389 15348
rect 7248 15308 7254 15320
rect 7377 15317 7389 15320
rect 7423 15317 7435 15351
rect 7377 15311 7435 15317
rect 7742 15308 7748 15360
rect 7800 15308 7806 15360
rect 10226 15308 10232 15360
rect 10284 15308 10290 15360
rect 11440 15348 11468 15447
rect 11532 15416 11560 15447
rect 11606 15444 11612 15496
rect 11664 15484 11670 15496
rect 11701 15487 11759 15493
rect 11701 15484 11713 15487
rect 11664 15456 11713 15484
rect 11664 15444 11670 15456
rect 11701 15453 11713 15456
rect 11747 15453 11759 15487
rect 11701 15447 11759 15453
rect 11882 15444 11888 15496
rect 11940 15444 11946 15496
rect 11974 15444 11980 15496
rect 12032 15444 12038 15496
rect 12066 15444 12072 15496
rect 12124 15444 12130 15496
rect 12618 15444 12624 15496
rect 12676 15484 12682 15496
rect 12713 15487 12771 15493
rect 12713 15484 12725 15487
rect 12676 15456 12725 15484
rect 12676 15444 12682 15456
rect 12713 15453 12725 15456
rect 12759 15453 12771 15487
rect 12713 15447 12771 15453
rect 14274 15444 14280 15496
rect 14332 15444 14338 15496
rect 14568 15484 14596 15580
rect 14645 15487 14703 15493
rect 14645 15484 14657 15487
rect 14568 15456 14657 15484
rect 14645 15453 14657 15456
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 15378 15444 15384 15496
rect 15436 15444 15442 15496
rect 15749 15487 15807 15493
rect 15749 15453 15761 15487
rect 15795 15484 15807 15487
rect 15838 15484 15844 15496
rect 15795 15456 15844 15484
rect 15795 15453 15807 15456
rect 15749 15447 15807 15453
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 16022 15444 16028 15496
rect 16080 15444 16086 15496
rect 16316 15484 16344 15660
rect 18524 15660 19340 15688
rect 18049 15623 18107 15629
rect 18049 15589 18061 15623
rect 18095 15620 18107 15623
rect 18414 15620 18420 15632
rect 18095 15592 18420 15620
rect 18095 15589 18107 15592
rect 18049 15583 18107 15589
rect 18414 15580 18420 15592
rect 18472 15580 18478 15632
rect 17218 15512 17224 15564
rect 17276 15512 17282 15564
rect 18524 15561 18552 15660
rect 19334 15648 19340 15660
rect 19392 15648 19398 15700
rect 21450 15688 21456 15700
rect 19536 15660 21456 15688
rect 19058 15580 19064 15632
rect 19116 15620 19122 15632
rect 19426 15620 19432 15632
rect 19116 15592 19432 15620
rect 19116 15580 19122 15592
rect 19426 15580 19432 15592
rect 19484 15620 19490 15632
rect 19536 15620 19564 15660
rect 21450 15648 21456 15660
rect 21508 15648 21514 15700
rect 21545 15691 21603 15697
rect 21545 15657 21557 15691
rect 21591 15688 21603 15691
rect 21818 15688 21824 15700
rect 21591 15660 21824 15688
rect 21591 15657 21603 15660
rect 21545 15651 21603 15657
rect 21818 15648 21824 15660
rect 21876 15648 21882 15700
rect 22186 15648 22192 15700
rect 22244 15688 22250 15700
rect 22281 15691 22339 15697
rect 22281 15688 22293 15691
rect 22244 15660 22293 15688
rect 22244 15648 22250 15660
rect 22281 15657 22293 15660
rect 22327 15657 22339 15691
rect 22281 15651 22339 15657
rect 22370 15648 22376 15700
rect 22428 15688 22434 15700
rect 22465 15691 22523 15697
rect 22465 15688 22477 15691
rect 22428 15660 22477 15688
rect 22428 15648 22434 15660
rect 22465 15657 22477 15660
rect 22511 15688 22523 15691
rect 25314 15688 25320 15700
rect 22511 15660 25320 15688
rect 22511 15657 22523 15660
rect 22465 15651 22523 15657
rect 25314 15648 25320 15660
rect 25372 15648 25378 15700
rect 26050 15648 26056 15700
rect 26108 15688 26114 15700
rect 26145 15691 26203 15697
rect 26145 15688 26157 15691
rect 26108 15660 26157 15688
rect 26108 15648 26114 15660
rect 26145 15657 26157 15660
rect 26191 15657 26203 15691
rect 26145 15651 26203 15657
rect 26418 15648 26424 15700
rect 26476 15648 26482 15700
rect 26878 15648 26884 15700
rect 26936 15648 26942 15700
rect 28350 15688 28356 15700
rect 27632 15660 28356 15688
rect 19484 15592 19564 15620
rect 19797 15623 19855 15629
rect 19484 15580 19490 15592
rect 19797 15589 19809 15623
rect 19843 15589 19855 15623
rect 19797 15583 19855 15589
rect 18509 15555 18567 15561
rect 18509 15552 18521 15555
rect 17420 15524 18092 15552
rect 17420 15496 17448 15524
rect 16485 15487 16543 15493
rect 16485 15484 16497 15487
rect 16316 15456 16497 15484
rect 16485 15453 16497 15456
rect 16531 15453 16543 15487
rect 16485 15447 16543 15453
rect 17402 15444 17408 15496
rect 17460 15444 17466 15496
rect 17494 15444 17500 15496
rect 17552 15444 17558 15496
rect 17954 15444 17960 15496
rect 18012 15444 18018 15496
rect 18064 15493 18092 15524
rect 18345 15524 18521 15552
rect 18049 15487 18107 15493
rect 18049 15453 18061 15487
rect 18095 15453 18107 15487
rect 18049 15447 18107 15453
rect 18233 15487 18291 15493
rect 18233 15453 18245 15487
rect 18279 15453 18291 15487
rect 18233 15447 18291 15453
rect 11532 15388 11744 15416
rect 11716 15360 11744 15388
rect 15102 15376 15108 15428
rect 15160 15376 15166 15428
rect 15562 15376 15568 15428
rect 15620 15416 15626 15428
rect 16393 15419 16451 15425
rect 16393 15416 16405 15419
rect 15620 15388 16405 15416
rect 15620 15376 15626 15388
rect 16393 15385 16405 15388
rect 16439 15385 16451 15419
rect 16393 15379 16451 15385
rect 16942 15376 16948 15428
rect 17000 15376 17006 15428
rect 17126 15376 17132 15428
rect 17184 15376 17190 15428
rect 17972 15416 18000 15444
rect 18248 15416 18276 15447
rect 17972 15388 18276 15416
rect 11514 15348 11520 15360
rect 11440 15320 11520 15348
rect 11514 15308 11520 15320
rect 11572 15308 11578 15360
rect 11698 15308 11704 15360
rect 11756 15308 11762 15360
rect 17144 15348 17172 15376
rect 18345 15348 18373 15524
rect 18509 15521 18521 15524
rect 18555 15521 18567 15555
rect 18509 15515 18567 15521
rect 18616 15524 19288 15552
rect 18616 15496 18644 15524
rect 18414 15444 18420 15496
rect 18472 15444 18478 15496
rect 18598 15444 18604 15496
rect 18656 15444 18662 15496
rect 19260 15493 19288 15524
rect 19444 15493 19472 15580
rect 19812 15552 19840 15583
rect 20070 15580 20076 15632
rect 20128 15580 20134 15632
rect 20441 15623 20499 15629
rect 20441 15589 20453 15623
rect 20487 15589 20499 15623
rect 20441 15583 20499 15589
rect 20088 15552 20116 15580
rect 19536 15524 19748 15552
rect 19812 15524 20116 15552
rect 19536 15493 19564 15524
rect 18877 15487 18935 15493
rect 18877 15453 18889 15487
rect 18923 15453 18935 15487
rect 18877 15447 18935 15453
rect 19245 15487 19303 15493
rect 19245 15453 19257 15487
rect 19291 15453 19303 15487
rect 19245 15447 19303 15453
rect 19429 15487 19487 15493
rect 19429 15453 19441 15487
rect 19475 15453 19487 15487
rect 19429 15447 19487 15453
rect 19521 15487 19579 15493
rect 19521 15453 19533 15487
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 18432 15416 18460 15444
rect 18892 15416 18920 15447
rect 18432 15388 18920 15416
rect 19260 15416 19288 15447
rect 19610 15444 19616 15496
rect 19668 15444 19674 15496
rect 19720 15484 19748 15524
rect 19886 15484 19892 15496
rect 19720 15456 19892 15484
rect 19886 15444 19892 15456
rect 19944 15444 19950 15496
rect 20165 15487 20223 15493
rect 20165 15484 20177 15487
rect 19996 15456 20177 15484
rect 19996 15416 20024 15456
rect 20165 15453 20177 15456
rect 20211 15453 20223 15487
rect 20165 15447 20223 15453
rect 20254 15444 20260 15496
rect 20312 15444 20318 15496
rect 20456 15484 20484 15583
rect 21358 15580 21364 15632
rect 21416 15620 21422 15632
rect 25958 15620 25964 15632
rect 21416 15592 25176 15620
rect 21416 15580 21422 15592
rect 25148 15564 25176 15592
rect 25424 15592 25964 15620
rect 20530 15512 20536 15564
rect 20588 15552 20594 15564
rect 20588 15524 21312 15552
rect 20588 15512 20594 15524
rect 21284 15496 21312 15524
rect 22554 15512 22560 15564
rect 22612 15552 22618 15564
rect 23382 15552 23388 15564
rect 22612 15524 23388 15552
rect 22612 15512 22618 15524
rect 23382 15512 23388 15524
rect 23440 15512 23446 15564
rect 25130 15512 25136 15564
rect 25188 15552 25194 15564
rect 25314 15552 25320 15564
rect 25188 15524 25320 15552
rect 25188 15512 25194 15524
rect 25314 15512 25320 15524
rect 25372 15512 25378 15564
rect 25424 15561 25452 15592
rect 25958 15580 25964 15592
rect 26016 15580 26022 15632
rect 26436 15620 26464 15648
rect 27632 15620 27660 15660
rect 28350 15648 28356 15660
rect 28408 15648 28414 15700
rect 28534 15648 28540 15700
rect 28592 15688 28598 15700
rect 28592 15660 28994 15688
rect 28592 15648 28598 15660
rect 26160 15592 27660 15620
rect 25409 15555 25467 15561
rect 25409 15521 25421 15555
rect 25455 15521 25467 15555
rect 26160 15552 26188 15592
rect 28258 15580 28264 15632
rect 28316 15580 28322 15632
rect 28445 15623 28503 15629
rect 28445 15589 28457 15623
rect 28491 15620 28503 15623
rect 28813 15623 28871 15629
rect 28813 15620 28825 15623
rect 28491 15592 28825 15620
rect 28491 15589 28503 15592
rect 28445 15583 28503 15589
rect 28813 15589 28825 15592
rect 28859 15589 28871 15623
rect 28813 15583 28871 15589
rect 25409 15515 25467 15521
rect 25885 15524 26188 15552
rect 26252 15524 26740 15552
rect 20901 15487 20959 15493
rect 20901 15484 20913 15487
rect 20456 15456 20913 15484
rect 20901 15453 20913 15456
rect 20947 15453 20959 15487
rect 20901 15447 20959 15453
rect 20994 15487 21052 15493
rect 20994 15453 21006 15487
rect 21040 15453 21052 15487
rect 20994 15447 21052 15453
rect 19260 15388 20024 15416
rect 20070 15376 20076 15428
rect 20128 15376 20134 15428
rect 20530 15376 20536 15428
rect 20588 15416 20594 15428
rect 20714 15416 20720 15428
rect 20588 15388 20720 15416
rect 20588 15376 20594 15388
rect 20714 15376 20720 15388
rect 20772 15376 20778 15428
rect 21008 15416 21036 15447
rect 21266 15444 21272 15496
rect 21324 15444 21330 15496
rect 21407 15487 21465 15493
rect 21407 15453 21419 15487
rect 21453 15484 21465 15487
rect 22278 15484 22284 15496
rect 21453 15456 22284 15484
rect 21453 15453 21465 15456
rect 21407 15447 21465 15453
rect 22278 15444 22284 15456
rect 22336 15444 22342 15496
rect 22649 15487 22707 15493
rect 22649 15453 22661 15487
rect 22695 15453 22707 15487
rect 22649 15447 22707 15453
rect 24857 15487 24915 15493
rect 24857 15453 24869 15487
rect 24903 15484 24915 15487
rect 25501 15487 25559 15493
rect 25501 15484 25513 15487
rect 24903 15456 25513 15484
rect 24903 15453 24915 15456
rect 24857 15447 24915 15453
rect 25501 15453 25513 15456
rect 25547 15453 25559 15487
rect 25501 15447 25559 15453
rect 20916 15388 21036 15416
rect 21177 15419 21235 15425
rect 20916 15360 20944 15388
rect 21177 15385 21189 15419
rect 21223 15385 21235 15419
rect 22664 15416 22692 15447
rect 25590 15444 25596 15496
rect 25648 15484 25654 15496
rect 25885 15493 25913 15524
rect 26050 15493 26056 15496
rect 25869 15487 25927 15493
rect 25648 15456 25693 15484
rect 25648 15444 25654 15456
rect 25869 15453 25881 15487
rect 25915 15453 25927 15487
rect 25869 15447 25927 15453
rect 26007 15487 26056 15493
rect 26007 15453 26019 15487
rect 26053 15453 26056 15487
rect 26007 15447 26056 15453
rect 26050 15444 26056 15447
rect 26108 15444 26114 15496
rect 26252 15493 26280 15524
rect 26712 15496 26740 15524
rect 26786 15512 26792 15564
rect 26844 15552 26850 15564
rect 27157 15555 27215 15561
rect 27157 15552 27169 15555
rect 26844 15524 27169 15552
rect 26844 15512 26850 15524
rect 27157 15521 27169 15524
rect 27203 15552 27215 15555
rect 28276 15552 28304 15580
rect 28966 15552 28994 15660
rect 29086 15648 29092 15700
rect 29144 15648 29150 15700
rect 29270 15648 29276 15700
rect 29328 15648 29334 15700
rect 30101 15691 30159 15697
rect 30101 15657 30113 15691
rect 30147 15688 30159 15691
rect 30558 15688 30564 15700
rect 30147 15660 30564 15688
rect 30147 15657 30159 15660
rect 30101 15651 30159 15657
rect 30558 15648 30564 15660
rect 30616 15648 30622 15700
rect 29288 15620 29316 15648
rect 30374 15620 30380 15632
rect 29288 15592 30380 15620
rect 30374 15580 30380 15592
rect 30432 15580 30438 15632
rect 33502 15552 33508 15564
rect 27203 15524 27660 15552
rect 28276 15524 28672 15552
rect 27203 15521 27215 15524
rect 27157 15515 27215 15521
rect 26237 15487 26295 15493
rect 26237 15453 26249 15487
rect 26283 15453 26295 15487
rect 26237 15447 26295 15453
rect 26326 15444 26332 15496
rect 26384 15444 26390 15496
rect 26418 15444 26424 15496
rect 26476 15444 26482 15496
rect 26513 15487 26571 15493
rect 26513 15453 26525 15487
rect 26559 15453 26571 15487
rect 26513 15447 26571 15453
rect 22830 15416 22836 15428
rect 21177 15379 21235 15385
rect 21468 15388 22094 15416
rect 22664 15388 22836 15416
rect 17144 15320 18373 15348
rect 18969 15351 19027 15357
rect 18969 15317 18981 15351
rect 19015 15348 19027 15351
rect 19610 15348 19616 15360
rect 19015 15320 19616 15348
rect 19015 15317 19027 15320
rect 18969 15311 19027 15317
rect 19610 15308 19616 15320
rect 19668 15308 19674 15360
rect 19794 15308 19800 15360
rect 19852 15348 19858 15360
rect 20625 15351 20683 15357
rect 20625 15348 20637 15351
rect 19852 15320 20637 15348
rect 19852 15308 19858 15320
rect 20625 15317 20637 15320
rect 20671 15317 20683 15351
rect 20625 15311 20683 15317
rect 20898 15308 20904 15360
rect 20956 15308 20962 15360
rect 21192 15348 21220 15379
rect 21468 15348 21496 15388
rect 21192 15320 21496 15348
rect 22066 15348 22094 15388
rect 22830 15376 22836 15388
rect 22888 15376 22894 15428
rect 23290 15376 23296 15428
rect 23348 15416 23354 15428
rect 24026 15416 24032 15428
rect 23348 15388 24032 15416
rect 23348 15376 23354 15388
rect 24026 15376 24032 15388
rect 24084 15376 24090 15428
rect 25038 15376 25044 15428
rect 25096 15376 25102 15428
rect 25774 15376 25780 15428
rect 25832 15416 25838 15428
rect 26344 15416 26372 15444
rect 26528 15416 26556 15447
rect 26602 15444 26608 15496
rect 26660 15444 26666 15496
rect 26694 15444 26700 15496
rect 26752 15444 26758 15496
rect 27062 15444 27068 15496
rect 27120 15484 27126 15496
rect 27525 15487 27583 15493
rect 27525 15484 27537 15487
rect 27120 15456 27537 15484
rect 27120 15444 27126 15456
rect 27525 15453 27537 15456
rect 27571 15453 27583 15487
rect 27525 15447 27583 15453
rect 25832 15388 26004 15416
rect 26344 15388 26556 15416
rect 27433 15419 27491 15425
rect 25832 15376 25838 15388
rect 25976 15360 26004 15388
rect 27433 15385 27445 15419
rect 27479 15416 27491 15419
rect 27479 15388 27568 15416
rect 27479 15385 27491 15388
rect 27433 15379 27491 15385
rect 27540 15360 27568 15388
rect 23842 15348 23848 15360
rect 22066 15320 23848 15348
rect 23842 15308 23848 15320
rect 23900 15348 23906 15360
rect 24762 15348 24768 15360
rect 23900 15320 24768 15348
rect 23900 15308 23906 15320
rect 24762 15308 24768 15320
rect 24820 15308 24826 15360
rect 25130 15308 25136 15360
rect 25188 15308 25194 15360
rect 25225 15351 25283 15357
rect 25225 15317 25237 15351
rect 25271 15348 25283 15351
rect 25498 15348 25504 15360
rect 25271 15320 25504 15348
rect 25271 15317 25283 15320
rect 25225 15311 25283 15317
rect 25498 15308 25504 15320
rect 25556 15308 25562 15360
rect 25958 15308 25964 15360
rect 26016 15308 26022 15360
rect 27246 15308 27252 15360
rect 27304 15348 27310 15360
rect 27341 15351 27399 15357
rect 27341 15348 27353 15351
rect 27304 15320 27353 15348
rect 27304 15308 27310 15320
rect 27341 15317 27353 15320
rect 27387 15317 27399 15351
rect 27341 15311 27399 15317
rect 27522 15308 27528 15360
rect 27580 15308 27586 15360
rect 27632 15348 27660 15524
rect 27709 15487 27767 15493
rect 27709 15453 27721 15487
rect 27755 15484 27767 15487
rect 27801 15487 27859 15493
rect 27801 15484 27813 15487
rect 27755 15456 27813 15484
rect 27755 15453 27767 15456
rect 27709 15447 27767 15453
rect 27801 15453 27813 15456
rect 27847 15453 27859 15487
rect 27801 15447 27859 15453
rect 27890 15444 27896 15496
rect 27948 15484 27954 15496
rect 27948 15456 27993 15484
rect 27948 15444 27954 15456
rect 28166 15444 28172 15496
rect 28224 15444 28230 15496
rect 28258 15444 28264 15496
rect 28316 15493 28322 15496
rect 28644 15493 28672 15524
rect 28828 15524 29592 15552
rect 28828 15496 28856 15524
rect 28316 15447 28324 15493
rect 28629 15487 28687 15493
rect 28629 15453 28641 15487
rect 28675 15453 28687 15487
rect 28629 15447 28687 15453
rect 28316 15444 28322 15447
rect 28718 15444 28724 15496
rect 28776 15444 28782 15496
rect 28810 15444 28816 15496
rect 28868 15444 28874 15496
rect 28902 15444 28908 15496
rect 28960 15444 28966 15496
rect 29564 15493 29592 15524
rect 29840 15524 33508 15552
rect 29840 15493 29868 15524
rect 33502 15512 33508 15524
rect 33560 15512 33566 15564
rect 29549 15487 29607 15493
rect 29549 15453 29561 15487
rect 29595 15453 29607 15487
rect 29549 15447 29607 15453
rect 29825 15487 29883 15493
rect 29825 15453 29837 15487
rect 29871 15453 29883 15487
rect 29825 15447 29883 15453
rect 29917 15487 29975 15493
rect 29917 15453 29929 15487
rect 29963 15484 29975 15487
rect 30190 15484 30196 15496
rect 29963 15456 30196 15484
rect 29963 15453 29975 15456
rect 29917 15447 29975 15453
rect 28074 15376 28080 15428
rect 28132 15416 28138 15428
rect 28442 15416 28448 15428
rect 28132 15388 28448 15416
rect 28132 15376 28138 15388
rect 28442 15376 28448 15388
rect 28500 15376 28506 15428
rect 29086 15376 29092 15428
rect 29144 15416 29150 15428
rect 29733 15419 29791 15425
rect 29733 15416 29745 15419
rect 29144 15388 29745 15416
rect 29144 15376 29150 15388
rect 29733 15385 29745 15388
rect 29779 15385 29791 15419
rect 29733 15379 29791 15385
rect 29840 15348 29868 15447
rect 30190 15444 30196 15456
rect 30248 15444 30254 15496
rect 30558 15444 30564 15496
rect 30616 15444 30622 15496
rect 30834 15444 30840 15496
rect 30892 15444 30898 15496
rect 32398 15444 32404 15496
rect 32456 15484 32462 15496
rect 33597 15487 33655 15493
rect 33597 15484 33609 15487
rect 32456 15456 33609 15484
rect 32456 15444 32462 15456
rect 33597 15453 33609 15456
rect 33643 15453 33655 15487
rect 33597 15447 33655 15453
rect 31113 15419 31171 15425
rect 31113 15416 31125 15419
rect 30760 15388 31125 15416
rect 30760 15357 30788 15388
rect 31113 15385 31125 15388
rect 31159 15385 31171 15419
rect 33962 15416 33968 15428
rect 32338 15388 33968 15416
rect 31113 15379 31171 15385
rect 33962 15376 33968 15388
rect 34020 15376 34026 15428
rect 27632 15320 29868 15348
rect 30745 15351 30803 15357
rect 30745 15317 30757 15351
rect 30791 15317 30803 15351
rect 30745 15311 30803 15317
rect 32582 15308 32588 15360
rect 32640 15308 32646 15360
rect 33318 15308 33324 15360
rect 33376 15348 33382 15360
rect 33505 15351 33563 15357
rect 33505 15348 33517 15351
rect 33376 15320 33517 15348
rect 33376 15308 33382 15320
rect 33505 15317 33517 15320
rect 33551 15317 33563 15351
rect 33505 15311 33563 15317
rect 1104 15258 38272 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 38272 15258
rect 1104 15184 38272 15206
rect 1762 15104 1768 15156
rect 1820 15104 1826 15156
rect 9122 15104 9128 15156
rect 9180 15104 9186 15156
rect 9493 15147 9551 15153
rect 9493 15113 9505 15147
rect 9539 15144 9551 15147
rect 11146 15144 11152 15156
rect 9539 15116 11152 15144
rect 9539 15113 9551 15116
rect 9493 15107 9551 15113
rect 7469 15079 7527 15085
rect 7469 15045 7481 15079
rect 7515 15076 7527 15079
rect 7742 15076 7748 15088
rect 7515 15048 7748 15076
rect 7515 15045 7527 15048
rect 7469 15039 7527 15045
rect 7742 15036 7748 15048
rect 7800 15036 7806 15088
rect 9030 15076 9036 15088
rect 8694 15048 9036 15076
rect 9030 15036 9036 15048
rect 9088 15036 9094 15088
rect 1946 14968 1952 15020
rect 2004 14968 2010 15020
rect 9508 15008 9536 15107
rect 11146 15104 11152 15116
rect 11204 15104 11210 15156
rect 11882 15104 11888 15156
rect 11940 15144 11946 15156
rect 11977 15147 12035 15153
rect 11977 15144 11989 15147
rect 11940 15116 11989 15144
rect 11940 15104 11946 15116
rect 11977 15113 11989 15116
rect 12023 15113 12035 15147
rect 11977 15107 12035 15113
rect 15013 15147 15071 15153
rect 15013 15113 15025 15147
rect 15059 15144 15071 15147
rect 16850 15144 16856 15156
rect 15059 15116 16856 15144
rect 15059 15113 15071 15116
rect 15013 15107 15071 15113
rect 16850 15104 16856 15116
rect 16908 15104 16914 15156
rect 17678 15104 17684 15156
rect 17736 15104 17742 15156
rect 17954 15104 17960 15156
rect 18012 15144 18018 15156
rect 18012 15116 18644 15144
rect 18012 15104 18018 15116
rect 11698 15076 11704 15088
rect 8680 14980 9536 15008
rect 9600 15048 11704 15076
rect 7190 14900 7196 14952
rect 7248 14900 7254 14952
rect 8018 14900 8024 14952
rect 8076 14940 8082 14952
rect 8680 14940 8708 14980
rect 9600 14949 9628 15048
rect 11698 15036 11704 15048
rect 11756 15036 11762 15088
rect 15381 15079 15439 15085
rect 12176 15048 12940 15076
rect 10226 14968 10232 15020
rect 10284 14968 10290 15020
rect 12176 15017 12204 15048
rect 12161 15011 12219 15017
rect 12161 14977 12173 15011
rect 12207 14977 12219 15011
rect 12161 14971 12219 14977
rect 12250 14968 12256 15020
rect 12308 14968 12314 15020
rect 12434 14968 12440 15020
rect 12492 14968 12498 15020
rect 12529 15011 12587 15017
rect 12529 14977 12541 15011
rect 12575 15008 12587 15011
rect 12802 15008 12808 15020
rect 12575 14980 12808 15008
rect 12575 14977 12587 14980
rect 12529 14971 12587 14977
rect 12802 14968 12808 14980
rect 12860 14968 12866 15020
rect 8076 14912 8708 14940
rect 8941 14943 8999 14949
rect 8076 14900 8082 14912
rect 8941 14909 8953 14943
rect 8987 14940 8999 14943
rect 9585 14943 9643 14949
rect 9585 14940 9597 14943
rect 8987 14912 9597 14940
rect 8987 14909 8999 14912
rect 8941 14903 8999 14909
rect 9585 14909 9597 14912
rect 9631 14909 9643 14943
rect 9585 14903 9643 14909
rect 9677 14943 9735 14949
rect 9677 14909 9689 14943
rect 9723 14909 9735 14943
rect 9677 14903 9735 14909
rect 10413 14943 10471 14949
rect 10413 14909 10425 14943
rect 10459 14909 10471 14943
rect 10413 14903 10471 14909
rect 9692 14872 9720 14903
rect 9646 14844 9720 14872
rect 10428 14872 10456 14903
rect 11054 14872 11060 14884
rect 10428 14844 11060 14872
rect 9646 14816 9674 14844
rect 11054 14832 11060 14844
rect 11112 14832 11118 14884
rect 12268 14872 12296 14968
rect 12912 14952 12940 15048
rect 15381 15045 15393 15079
rect 15427 15045 15439 15079
rect 15381 15039 15439 15045
rect 17405 15079 17463 15085
rect 17405 15045 17417 15079
rect 17451 15076 17463 15079
rect 17696 15076 17724 15104
rect 17451 15048 17724 15076
rect 17880 15048 18368 15076
rect 17451 15045 17463 15048
rect 17405 15039 17463 15045
rect 14550 14968 14556 15020
rect 14608 15008 14614 15020
rect 14737 15011 14795 15017
rect 14737 15008 14749 15011
rect 14608 14980 14749 15008
rect 14608 14968 14614 14980
rect 14737 14977 14749 14980
rect 14783 14977 14795 15011
rect 14737 14971 14795 14977
rect 14918 14968 14924 15020
rect 14976 15008 14982 15020
rect 15197 15011 15255 15017
rect 15197 15008 15209 15011
rect 14976 14980 15209 15008
rect 14976 14968 14982 14980
rect 15197 14977 15209 14980
rect 15243 14977 15255 15011
rect 15197 14971 15255 14977
rect 12894 14900 12900 14952
rect 12952 14900 12958 14952
rect 15396 14940 15424 15039
rect 15473 15011 15531 15017
rect 15473 14977 15485 15011
rect 15519 15008 15531 15011
rect 15654 15008 15660 15020
rect 15519 14980 15660 15008
rect 15519 14977 15531 14980
rect 15473 14971 15531 14977
rect 15654 14968 15660 14980
rect 15712 14968 15718 15020
rect 17126 14968 17132 15020
rect 17184 14968 17190 15020
rect 17222 15011 17280 15017
rect 17222 14977 17234 15011
rect 17268 14977 17280 15011
rect 17222 14971 17280 14977
rect 17497 15011 17555 15017
rect 17497 14977 17509 15011
rect 17543 14977 17555 15011
rect 17497 14971 17555 14977
rect 17635 15011 17693 15017
rect 17635 14977 17647 15011
rect 17681 15008 17693 15011
rect 17770 15008 17776 15020
rect 17681 14980 17776 15008
rect 17681 14977 17693 14980
rect 17635 14971 17693 14977
rect 15562 14940 15568 14952
rect 15396 14912 15568 14940
rect 15562 14900 15568 14912
rect 15620 14900 15626 14952
rect 15933 14943 15991 14949
rect 15933 14909 15945 14943
rect 15979 14940 15991 14943
rect 16390 14940 16396 14952
rect 15979 14912 16396 14940
rect 15979 14909 15991 14912
rect 15933 14903 15991 14909
rect 16390 14900 16396 14912
rect 16448 14900 16454 14952
rect 17236 14884 17264 14971
rect 17218 14872 17224 14884
rect 12268 14844 17224 14872
rect 17218 14832 17224 14844
rect 17276 14832 17282 14884
rect 9582 14764 9588 14816
rect 9640 14776 9674 14816
rect 9640 14764 9646 14776
rect 12158 14764 12164 14816
rect 12216 14804 12222 14816
rect 17512 14804 17540 14971
rect 17770 14968 17776 14980
rect 17828 14968 17834 15020
rect 17880 15017 17908 15048
rect 18340 15020 18368 15048
rect 17865 15011 17923 15017
rect 17865 14977 17877 15011
rect 17911 14977 17923 15011
rect 17865 14971 17923 14977
rect 17954 14968 17960 15020
rect 18012 14968 18018 15020
rect 18141 15011 18199 15017
rect 18141 14977 18153 15011
rect 18187 14977 18199 15011
rect 18141 14971 18199 14977
rect 18156 14940 18184 14971
rect 18230 14968 18236 15020
rect 18288 14968 18294 15020
rect 18322 14968 18328 15020
rect 18380 14968 18386 15020
rect 18414 14968 18420 15020
rect 18472 14968 18478 15020
rect 18509 15011 18567 15017
rect 18509 14977 18521 15011
rect 18555 14977 18567 15011
rect 18509 14971 18567 14977
rect 17788 14912 18184 14940
rect 17788 14881 17816 14912
rect 17773 14875 17831 14881
rect 17773 14841 17785 14875
rect 17819 14841 17831 14875
rect 18248 14872 18276 14968
rect 18524 14940 18552 14971
rect 18432 14912 18552 14940
rect 18325 14875 18383 14881
rect 18325 14872 18337 14875
rect 18248 14844 18337 14872
rect 17773 14835 17831 14841
rect 18325 14841 18337 14844
rect 18371 14841 18383 14875
rect 18325 14835 18383 14841
rect 18432 14804 18460 14912
rect 18616 14872 18644 15116
rect 19702 15104 19708 15156
rect 19760 15144 19766 15156
rect 20257 15147 20315 15153
rect 20257 15144 20269 15147
rect 19760 15116 20269 15144
rect 19760 15104 19766 15116
rect 20257 15113 20269 15116
rect 20303 15113 20315 15147
rect 20257 15107 20315 15113
rect 20346 15104 20352 15156
rect 20404 15144 20410 15156
rect 20622 15144 20628 15156
rect 20404 15116 20628 15144
rect 20404 15104 20410 15116
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 20990 15144 20996 15156
rect 20916 15116 20996 15144
rect 18690 15036 18696 15088
rect 18748 15036 18754 15088
rect 18785 15079 18843 15085
rect 18785 15045 18797 15079
rect 18831 15076 18843 15079
rect 19518 15076 19524 15088
rect 18831 15048 19524 15076
rect 18831 15045 18843 15048
rect 18785 15039 18843 15045
rect 19518 15036 19524 15048
rect 19576 15036 19582 15088
rect 19889 15079 19947 15085
rect 19889 15045 19901 15079
rect 19935 15076 19947 15079
rect 19935 15048 20208 15076
rect 19935 15045 19947 15048
rect 19889 15039 19947 15045
rect 20180 15020 20208 15048
rect 20806 15036 20812 15088
rect 20864 15036 20870 15088
rect 20916 15085 20944 15116
rect 20990 15104 20996 15116
rect 21048 15104 21054 15156
rect 24394 15104 24400 15156
rect 24452 15104 24458 15156
rect 24762 15104 24768 15156
rect 24820 15144 24826 15156
rect 24820 15116 25084 15144
rect 24820 15104 24826 15116
rect 20901 15079 20959 15085
rect 20901 15045 20913 15079
rect 20947 15045 20959 15079
rect 24412 15076 24440 15104
rect 25056 15085 25084 15116
rect 25222 15104 25228 15156
rect 25280 15104 25286 15156
rect 25409 15147 25467 15153
rect 25409 15113 25421 15147
rect 25455 15113 25467 15147
rect 25409 15107 25467 15113
rect 24489 15079 24547 15085
rect 24489 15076 24501 15079
rect 20901 15039 20959 15045
rect 22296 15048 24348 15076
rect 24412 15048 24501 15076
rect 22296 15020 22324 15048
rect 18877 15011 18935 15017
rect 18877 14977 18889 15011
rect 18923 15008 18935 15011
rect 19426 15008 19432 15020
rect 18923 14980 19432 15008
rect 18923 14977 18935 14980
rect 18877 14971 18935 14977
rect 19426 14968 19432 14980
rect 19484 14968 19490 15020
rect 19610 14968 19616 15020
rect 19668 14968 19674 15020
rect 19794 15017 19800 15020
rect 19771 15011 19800 15017
rect 19771 14977 19783 15011
rect 19771 14971 19800 14977
rect 19794 14968 19800 14971
rect 19852 14968 19858 15020
rect 19981 15011 20039 15017
rect 19981 14977 19993 15011
rect 20027 14977 20039 15011
rect 19981 14971 20039 14977
rect 20073 15011 20131 15017
rect 20073 14977 20085 15011
rect 20119 14977 20131 15011
rect 20073 14971 20131 14977
rect 18969 14943 19027 14949
rect 18969 14909 18981 14943
rect 19015 14940 19027 14943
rect 19996 14940 20024 14971
rect 19015 14912 20024 14940
rect 20088 14940 20116 14971
rect 20162 14968 20168 15020
rect 20220 14968 20226 15020
rect 20530 14968 20536 15020
rect 20588 14968 20594 15020
rect 20622 14968 20628 15020
rect 20680 14968 20686 15020
rect 20993 15011 21051 15017
rect 20993 14977 21005 15011
rect 21039 15008 21051 15011
rect 21726 15008 21732 15020
rect 21039 14980 21732 15008
rect 21039 14977 21051 14980
rect 20993 14971 21051 14977
rect 21726 14968 21732 14980
rect 21784 14968 21790 15020
rect 21910 14968 21916 15020
rect 21968 15008 21974 15020
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21968 14980 22017 15008
rect 21968 14968 21974 14980
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 22278 14968 22284 15020
rect 22336 14968 22342 15020
rect 23382 14968 23388 15020
rect 23440 14968 23446 15020
rect 24213 15011 24271 15017
rect 24213 14977 24225 15011
rect 24259 14977 24271 15011
rect 24213 14971 24271 14977
rect 20640 14940 20668 14968
rect 21174 14940 21180 14952
rect 20088 14912 20576 14940
rect 20640 14912 21180 14940
rect 19015 14909 19027 14912
rect 18969 14903 19027 14909
rect 19702 14872 19708 14884
rect 18616 14844 19708 14872
rect 19702 14832 19708 14844
rect 19760 14832 19766 14884
rect 20548 14881 20576 14912
rect 21174 14900 21180 14912
rect 21232 14900 21238 14952
rect 21266 14900 21272 14952
rect 21324 14940 21330 14952
rect 21821 14943 21879 14949
rect 21821 14940 21833 14943
rect 21324 14912 21833 14940
rect 21324 14900 21330 14912
rect 21821 14909 21833 14912
rect 21867 14909 21879 14943
rect 23566 14940 23572 14952
rect 21821 14903 21879 14909
rect 21928 14912 23572 14940
rect 20533 14875 20591 14881
rect 20533 14841 20545 14875
rect 20579 14841 20591 14875
rect 20533 14835 20591 14841
rect 20714 14832 20720 14884
rect 20772 14872 20778 14884
rect 21928 14872 21956 14912
rect 23566 14900 23572 14912
rect 23624 14900 23630 14952
rect 24228 14872 24256 14971
rect 24320 14940 24348 15048
rect 24489 15045 24501 15048
rect 24535 15076 24547 15079
rect 25041 15079 25099 15085
rect 24535 15048 24900 15076
rect 24535 15045 24547 15048
rect 24489 15039 24547 15045
rect 24394 14968 24400 15020
rect 24452 14968 24458 15020
rect 24578 14968 24584 15020
rect 24636 14968 24642 15020
rect 24872 15017 24900 15048
rect 25041 15045 25053 15079
rect 25087 15045 25099 15079
rect 25041 15039 25099 15045
rect 25133 15079 25191 15085
rect 25133 15045 25145 15079
rect 25179 15076 25191 15079
rect 25240 15076 25268 15104
rect 25179 15048 25268 15076
rect 25424 15076 25452 15107
rect 25682 15104 25688 15156
rect 25740 15144 25746 15156
rect 26142 15144 26148 15156
rect 25740 15116 26148 15144
rect 25740 15104 25746 15116
rect 26142 15104 26148 15116
rect 26200 15104 26206 15156
rect 26418 15104 26424 15156
rect 26476 15144 26482 15156
rect 26513 15147 26571 15153
rect 26513 15144 26525 15147
rect 26476 15116 26525 15144
rect 26476 15104 26482 15116
rect 26513 15113 26525 15116
rect 26559 15113 26571 15147
rect 28534 15144 28540 15156
rect 26513 15107 26571 15113
rect 28092 15116 28540 15144
rect 28092 15076 28120 15116
rect 28534 15104 28540 15116
rect 28592 15104 28598 15156
rect 28629 15147 28687 15153
rect 28629 15113 28641 15147
rect 28675 15144 28687 15147
rect 28718 15144 28724 15156
rect 28675 15116 28724 15144
rect 28675 15113 28687 15116
rect 28629 15107 28687 15113
rect 28718 15104 28724 15116
rect 28776 15104 28782 15156
rect 30558 15104 30564 15156
rect 30616 15144 30622 15156
rect 30745 15147 30803 15153
rect 30745 15144 30757 15147
rect 30616 15116 30757 15144
rect 30616 15104 30622 15116
rect 30745 15113 30757 15116
rect 30791 15113 30803 15147
rect 30745 15107 30803 15113
rect 30834 15104 30840 15156
rect 30892 15144 30898 15156
rect 31021 15147 31079 15153
rect 31021 15144 31033 15147
rect 30892 15116 31033 15144
rect 30892 15104 30898 15116
rect 31021 15113 31033 15116
rect 31067 15113 31079 15147
rect 31021 15107 31079 15113
rect 33229 15147 33287 15153
rect 33229 15113 33241 15147
rect 33275 15144 33287 15147
rect 33275 15116 33640 15144
rect 33275 15113 33287 15116
rect 33229 15107 33287 15113
rect 33612 15085 33640 15116
rect 33962 15104 33968 15156
rect 34020 15104 34026 15156
rect 25424 15048 26096 15076
rect 25179 15045 25191 15048
rect 25133 15039 25191 15045
rect 24857 15011 24915 15017
rect 24857 14977 24869 15011
rect 24903 14977 24915 15011
rect 24857 14971 24915 14977
rect 25225 15011 25283 15017
rect 25225 14977 25237 15011
rect 25271 15008 25283 15011
rect 25498 15008 25504 15020
rect 25271 14980 25504 15008
rect 25271 14977 25283 14980
rect 25225 14971 25283 14977
rect 25498 14968 25504 14980
rect 25556 14968 25562 15020
rect 26068 15017 26096 15048
rect 26157 15048 28120 15076
rect 25951 15011 26009 15017
rect 25951 14977 25963 15011
rect 25997 14977 26009 15011
rect 25951 14971 26009 14977
rect 26053 15011 26111 15017
rect 26053 14977 26065 15011
rect 26099 14977 26111 15011
rect 26053 14971 26111 14977
rect 25966 14940 25994 14971
rect 26157 14940 26185 15048
rect 28092 15017 28120 15048
rect 28261 15079 28319 15085
rect 28261 15045 28273 15079
rect 28307 15076 28319 15079
rect 29089 15079 29147 15085
rect 29089 15076 29101 15079
rect 28307 15048 29101 15076
rect 28307 15045 28319 15048
rect 28261 15039 28319 15045
rect 29089 15045 29101 15048
rect 29135 15045 29147 15079
rect 29089 15039 29147 15045
rect 33597 15079 33655 15085
rect 33597 15045 33609 15079
rect 33643 15045 33655 15079
rect 33980 15076 34008 15104
rect 33980 15048 34086 15076
rect 33597 15039 33655 15045
rect 26237 15011 26295 15017
rect 26237 14977 26249 15011
rect 26283 14977 26295 15011
rect 26237 14971 26295 14977
rect 26329 15011 26387 15017
rect 26329 14977 26341 15011
rect 26375 14977 26387 15011
rect 26329 14971 26387 14977
rect 28077 15011 28135 15017
rect 28077 14977 28089 15011
rect 28123 14977 28135 15011
rect 28077 14971 28135 14977
rect 24320 14912 26185 14940
rect 24946 14872 24952 14884
rect 20772 14844 21956 14872
rect 22066 14844 22508 14872
rect 24228 14844 24952 14872
rect 20772 14832 20778 14844
rect 18506 14804 18512 14816
rect 12216 14776 18512 14804
rect 12216 14764 12222 14776
rect 18506 14764 18512 14776
rect 18564 14764 18570 14816
rect 19426 14764 19432 14816
rect 19484 14804 19490 14816
rect 22066 14804 22094 14844
rect 22480 14816 22508 14844
rect 24946 14832 24952 14844
rect 25004 14872 25010 14884
rect 25590 14872 25596 14884
rect 25004 14844 25596 14872
rect 25004 14832 25010 14844
rect 25590 14832 25596 14844
rect 25648 14872 25654 14884
rect 26252 14872 26280 14971
rect 26344 14940 26372 14971
rect 28350 14968 28356 15020
rect 28408 14968 28414 15020
rect 28445 15011 28503 15017
rect 28445 14977 28457 15011
rect 28491 14977 28503 15011
rect 28445 14971 28503 14977
rect 26418 14940 26424 14952
rect 26344 14912 26424 14940
rect 26418 14900 26424 14912
rect 26476 14900 26482 14952
rect 28166 14900 28172 14952
rect 28224 14940 28230 14952
rect 28460 14940 28488 14971
rect 28534 14968 28540 15020
rect 28592 15008 28598 15020
rect 28721 15011 28779 15017
rect 28721 15008 28733 15011
rect 28592 14980 28733 15008
rect 28592 14968 28598 14980
rect 28721 14977 28733 14980
rect 28767 14977 28779 15011
rect 28721 14971 28779 14977
rect 28810 14968 28816 15020
rect 28868 15008 28874 15020
rect 28905 15011 28963 15017
rect 28905 15008 28917 15011
rect 28868 14980 28917 15008
rect 28868 14968 28874 14980
rect 28905 14977 28917 14980
rect 28951 14977 28963 15011
rect 30377 15011 30435 15017
rect 28905 14971 28963 14977
rect 29012 14980 30328 15008
rect 29012 14940 29040 14980
rect 28224 14912 28488 14940
rect 28552 14912 29040 14940
rect 28224 14900 28230 14912
rect 28552 14872 28580 14912
rect 30098 14900 30104 14952
rect 30156 14900 30162 14952
rect 30300 14949 30328 14980
rect 30377 14977 30389 15011
rect 30423 15008 30435 15011
rect 30466 15008 30472 15020
rect 30423 14980 30472 15008
rect 30423 14977 30435 14980
rect 30377 14971 30435 14977
rect 30466 14968 30472 14980
rect 30524 14968 30530 15020
rect 31110 14968 31116 15020
rect 31168 15008 31174 15020
rect 31662 15008 31668 15020
rect 31168 14980 31668 15008
rect 31168 14968 31174 14980
rect 31662 14968 31668 14980
rect 31720 15008 31726 15020
rect 32398 15008 32404 15020
rect 31720 14980 32404 15008
rect 31720 14968 31726 14980
rect 32398 14968 32404 14980
rect 32456 14968 32462 15020
rect 33042 14968 33048 15020
rect 33100 14968 33106 15020
rect 30285 14943 30343 14949
rect 30285 14909 30297 14943
rect 30331 14940 30343 14943
rect 32582 14940 32588 14952
rect 30331 14912 32588 14940
rect 30331 14909 30343 14912
rect 30285 14903 30343 14909
rect 32582 14900 32588 14912
rect 32640 14900 32646 14952
rect 33318 14900 33324 14952
rect 33376 14900 33382 14952
rect 25648 14844 28580 14872
rect 25648 14832 25654 14844
rect 28902 14832 28908 14884
rect 28960 14832 28966 14884
rect 19484 14776 22094 14804
rect 19484 14764 19490 14776
rect 22186 14764 22192 14816
rect 22244 14764 22250 14816
rect 22462 14764 22468 14816
rect 22520 14764 22526 14816
rect 23198 14764 23204 14816
rect 23256 14764 23262 14816
rect 24765 14807 24823 14813
rect 24765 14773 24777 14807
rect 24811 14804 24823 14807
rect 28920 14804 28948 14832
rect 24811 14776 28948 14804
rect 24811 14773 24823 14776
rect 24765 14767 24823 14773
rect 29822 14764 29828 14816
rect 29880 14804 29886 14816
rect 31110 14804 31116 14816
rect 29880 14776 31116 14804
rect 29880 14764 29886 14776
rect 31110 14764 31116 14776
rect 31168 14764 31174 14816
rect 33594 14764 33600 14816
rect 33652 14804 33658 14816
rect 35069 14807 35127 14813
rect 35069 14804 35081 14807
rect 33652 14776 35081 14804
rect 33652 14764 33658 14776
rect 35069 14773 35081 14776
rect 35115 14773 35127 14807
rect 35069 14767 35127 14773
rect 1104 14714 38272 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38272 14714
rect 1104 14640 38272 14662
rect 1946 14560 1952 14612
rect 2004 14600 2010 14612
rect 4157 14603 4215 14609
rect 4157 14600 4169 14603
rect 2004 14572 4169 14600
rect 2004 14560 2010 14572
rect 4157 14569 4169 14572
rect 4203 14569 4215 14603
rect 12250 14600 12256 14612
rect 4157 14563 4215 14569
rect 7024 14572 12256 14600
rect 5350 14464 5356 14476
rect 4356 14436 5356 14464
rect 4356 14405 4384 14436
rect 5350 14424 5356 14436
rect 5408 14424 5414 14476
rect 7024 14473 7052 14572
rect 12250 14560 12256 14572
rect 12308 14560 12314 14612
rect 12434 14560 12440 14612
rect 12492 14600 12498 14612
rect 12529 14603 12587 14609
rect 12529 14600 12541 14603
rect 12492 14572 12541 14600
rect 12492 14560 12498 14572
rect 12529 14569 12541 14572
rect 12575 14569 12587 14603
rect 12529 14563 12587 14569
rect 13906 14560 13912 14612
rect 13964 14600 13970 14612
rect 17034 14600 17040 14612
rect 13964 14572 17040 14600
rect 13964 14560 13970 14572
rect 17034 14560 17040 14572
rect 17092 14560 17098 14612
rect 17954 14600 17960 14612
rect 17149 14572 17960 14600
rect 7208 14504 8524 14532
rect 7208 14476 7236 14504
rect 6365 14467 6423 14473
rect 6365 14433 6377 14467
rect 6411 14464 6423 14467
rect 7009 14467 7067 14473
rect 7009 14464 7021 14467
rect 6411 14436 7021 14464
rect 6411 14433 6423 14436
rect 6365 14427 6423 14433
rect 7009 14433 7021 14436
rect 7055 14433 7067 14467
rect 7009 14427 7067 14433
rect 7190 14424 7196 14476
rect 7248 14424 7254 14476
rect 8018 14424 8024 14476
rect 8076 14424 8082 14476
rect 8202 14424 8208 14476
rect 8260 14424 8266 14476
rect 8496 14464 8524 14504
rect 9858 14492 9864 14544
rect 9916 14532 9922 14544
rect 10045 14535 10103 14541
rect 10045 14532 10057 14535
rect 9916 14504 10057 14532
rect 9916 14492 9922 14504
rect 10045 14501 10057 14504
rect 10091 14501 10103 14535
rect 10045 14495 10103 14501
rect 11698 14492 11704 14544
rect 11756 14532 11762 14544
rect 17149 14532 17177 14572
rect 17954 14560 17960 14572
rect 18012 14560 18018 14612
rect 18141 14603 18199 14609
rect 18141 14569 18153 14603
rect 18187 14600 18199 14603
rect 18414 14600 18420 14612
rect 18187 14572 18420 14600
rect 18187 14569 18199 14572
rect 18141 14563 18199 14569
rect 18414 14560 18420 14572
rect 18472 14560 18478 14612
rect 19886 14560 19892 14612
rect 19944 14600 19950 14612
rect 20990 14600 20996 14612
rect 19944 14572 20996 14600
rect 19944 14560 19950 14572
rect 20990 14560 20996 14572
rect 21048 14560 21054 14612
rect 21726 14560 21732 14612
rect 21784 14560 21790 14612
rect 24213 14603 24271 14609
rect 24213 14569 24225 14603
rect 24259 14600 24271 14603
rect 24302 14600 24308 14612
rect 24259 14572 24308 14600
rect 24259 14569 24271 14572
rect 24213 14563 24271 14569
rect 24302 14560 24308 14572
rect 24360 14560 24366 14612
rect 25958 14560 25964 14612
rect 26016 14600 26022 14612
rect 26510 14600 26516 14612
rect 26016 14572 26516 14600
rect 26016 14560 26022 14572
rect 26510 14560 26516 14572
rect 26568 14560 26574 14612
rect 28810 14560 28816 14612
rect 28868 14600 28874 14612
rect 32490 14600 32496 14612
rect 28868 14572 32496 14600
rect 28868 14560 28874 14572
rect 32490 14560 32496 14572
rect 32548 14600 32554 14612
rect 32861 14603 32919 14609
rect 32861 14600 32873 14603
rect 32548 14572 32873 14600
rect 32548 14560 32554 14572
rect 32861 14569 32873 14572
rect 32907 14569 32919 14603
rect 32861 14563 32919 14569
rect 33042 14560 33048 14612
rect 33100 14600 33106 14612
rect 33229 14603 33287 14609
rect 33229 14600 33241 14603
rect 33100 14572 33241 14600
rect 33100 14560 33106 14572
rect 33229 14569 33241 14572
rect 33275 14569 33287 14603
rect 33229 14563 33287 14569
rect 37829 14603 37887 14609
rect 37829 14569 37841 14603
rect 37875 14600 37887 14603
rect 37875 14572 38332 14600
rect 37875 14569 37887 14572
rect 37829 14563 37887 14569
rect 11756 14504 17177 14532
rect 11756 14492 11762 14504
rect 11054 14464 11060 14476
rect 8496 14436 11060 14464
rect 11054 14424 11060 14436
rect 11112 14424 11118 14476
rect 12158 14464 12164 14476
rect 11992 14436 12164 14464
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14365 4399 14399
rect 4341 14359 4399 14365
rect 4522 14356 4528 14408
rect 4580 14356 4586 14408
rect 4614 14356 4620 14408
rect 4672 14356 4678 14408
rect 6917 14399 6975 14405
rect 6917 14365 6929 14399
rect 6963 14396 6975 14399
rect 7098 14396 7104 14408
rect 6963 14368 7104 14396
rect 6963 14365 6975 14368
rect 6917 14359 6975 14365
rect 7098 14356 7104 14368
rect 7156 14396 7162 14408
rect 8036 14396 8064 14424
rect 7156 14368 8064 14396
rect 9861 14399 9919 14405
rect 7156 14356 7162 14368
rect 9861 14365 9873 14399
rect 9907 14396 9919 14399
rect 10042 14396 10048 14408
rect 9907 14368 10048 14396
rect 9907 14365 9919 14368
rect 9861 14359 9919 14365
rect 10042 14356 10048 14368
rect 10100 14356 10106 14408
rect 10134 14356 10140 14408
rect 10192 14396 10198 14408
rect 10505 14399 10563 14405
rect 10505 14396 10517 14399
rect 10192 14368 10517 14396
rect 10192 14356 10198 14368
rect 10505 14365 10517 14368
rect 10551 14365 10563 14399
rect 10505 14359 10563 14365
rect 11149 14399 11207 14405
rect 11149 14365 11161 14399
rect 11195 14396 11207 14399
rect 11606 14396 11612 14408
rect 11195 14368 11612 14396
rect 11195 14365 11207 14368
rect 11149 14359 11207 14365
rect 11606 14356 11612 14368
rect 11664 14356 11670 14408
rect 11992 14405 12020 14436
rect 12158 14424 12164 14436
rect 12216 14424 12222 14476
rect 12268 14405 12296 14504
rect 17218 14492 17224 14544
rect 17276 14532 17282 14544
rect 20530 14532 20536 14544
rect 17276 14504 20536 14532
rect 17276 14492 17282 14504
rect 20530 14492 20536 14504
rect 20588 14492 20594 14544
rect 14642 14424 14648 14476
rect 14700 14464 14706 14476
rect 19886 14464 19892 14476
rect 14700 14436 19892 14464
rect 14700 14424 14706 14436
rect 19886 14424 19892 14436
rect 19944 14424 19950 14476
rect 20162 14424 20168 14476
rect 20220 14424 20226 14476
rect 11977 14399 12035 14405
rect 11977 14365 11989 14399
rect 12023 14365 12035 14399
rect 11977 14359 12035 14365
rect 12253 14399 12311 14405
rect 12253 14365 12265 14399
rect 12299 14365 12311 14399
rect 12253 14359 12311 14365
rect 12345 14399 12403 14405
rect 12345 14365 12357 14399
rect 12391 14396 12403 14399
rect 12618 14396 12624 14408
rect 12391 14368 12624 14396
rect 12391 14365 12403 14368
rect 12345 14359 12403 14365
rect 4893 14331 4951 14337
rect 4893 14297 4905 14331
rect 4939 14297 4951 14331
rect 6178 14328 6184 14340
rect 6118 14300 6184 14328
rect 4893 14291 4951 14297
rect 4908 14260 4936 14291
rect 6178 14288 6184 14300
rect 6236 14328 6242 14340
rect 7929 14331 7987 14337
rect 6236 14300 7696 14328
rect 6236 14288 6242 14300
rect 5258 14260 5264 14272
rect 4908 14232 5264 14260
rect 5258 14220 5264 14232
rect 5316 14220 5322 14272
rect 6546 14220 6552 14272
rect 6604 14220 6610 14272
rect 7558 14220 7564 14272
rect 7616 14220 7622 14272
rect 7668 14260 7696 14300
rect 7929 14297 7941 14331
rect 7975 14328 7987 14331
rect 8478 14328 8484 14340
rect 7975 14300 8484 14328
rect 7975 14297 7987 14300
rect 7929 14291 7987 14297
rect 8478 14288 8484 14300
rect 8536 14328 8542 14340
rect 11992 14328 12020 14359
rect 12618 14356 12624 14368
rect 12676 14356 12682 14408
rect 15010 14356 15016 14408
rect 15068 14356 15074 14408
rect 17310 14356 17316 14408
rect 17368 14396 17374 14408
rect 17773 14399 17831 14405
rect 17773 14396 17785 14399
rect 17368 14368 17785 14396
rect 17368 14356 17374 14368
rect 17773 14365 17785 14368
rect 17819 14365 17831 14399
rect 17773 14359 17831 14365
rect 17862 14356 17868 14408
rect 17920 14356 17926 14408
rect 17954 14356 17960 14408
rect 18012 14396 18018 14408
rect 18138 14396 18144 14408
rect 18012 14368 18144 14396
rect 18012 14356 18018 14368
rect 18138 14356 18144 14368
rect 18196 14396 18202 14408
rect 19242 14396 19248 14408
rect 18196 14368 19248 14396
rect 18196 14356 18202 14368
rect 19242 14356 19248 14368
rect 19300 14356 19306 14408
rect 19334 14356 19340 14408
rect 19392 14396 19398 14408
rect 19978 14396 19984 14408
rect 19392 14368 19984 14396
rect 19392 14356 19398 14368
rect 19978 14356 19984 14368
rect 20036 14399 20042 14408
rect 20257 14399 20315 14405
rect 20036 14393 20095 14399
rect 20036 14359 20049 14393
rect 20083 14359 20095 14393
rect 20257 14365 20269 14399
rect 20303 14396 20315 14399
rect 20714 14396 20720 14408
rect 20303 14368 20720 14396
rect 20303 14365 20315 14368
rect 20257 14359 20315 14365
rect 20036 14356 20095 14359
rect 20714 14356 20720 14368
rect 20772 14356 20778 14408
rect 21008 14405 21036 14560
rect 38304 14544 38332 14572
rect 21376 14504 22416 14532
rect 21376 14405 21404 14504
rect 20993 14399 21051 14405
rect 20993 14365 21005 14399
rect 21039 14365 21051 14399
rect 21361 14399 21419 14405
rect 21361 14396 21373 14399
rect 20993 14359 21051 14365
rect 21100 14368 21373 14396
rect 20037 14353 20095 14356
rect 8536 14300 12020 14328
rect 12161 14331 12219 14337
rect 8536 14288 8542 14300
rect 12161 14297 12173 14331
rect 12207 14328 12219 14331
rect 12526 14328 12532 14340
rect 12207 14300 12532 14328
rect 12207 14297 12219 14300
rect 12161 14291 12219 14297
rect 12526 14288 12532 14300
rect 12584 14288 12590 14340
rect 16482 14288 16488 14340
rect 16540 14328 16546 14340
rect 17589 14331 17647 14337
rect 17589 14328 17601 14331
rect 16540 14300 17601 14328
rect 16540 14288 16546 14300
rect 17589 14297 17601 14300
rect 17635 14328 17647 14331
rect 18598 14328 18604 14340
rect 17635 14300 18604 14328
rect 17635 14297 17647 14300
rect 17589 14291 17647 14297
rect 18598 14288 18604 14300
rect 18656 14288 18662 14340
rect 20165 14331 20223 14337
rect 20165 14297 20177 14331
rect 20211 14297 20223 14331
rect 20165 14291 20223 14297
rect 9030 14260 9036 14272
rect 7668 14232 9036 14260
rect 9030 14220 9036 14232
rect 9088 14260 9094 14272
rect 14274 14260 14280 14272
rect 9088 14232 14280 14260
rect 9088 14220 9094 14232
rect 14274 14220 14280 14232
rect 14332 14220 14338 14272
rect 14918 14220 14924 14272
rect 14976 14220 14982 14272
rect 17678 14220 17684 14272
rect 17736 14260 17742 14272
rect 17862 14260 17868 14272
rect 17736 14232 17868 14260
rect 17736 14220 17742 14232
rect 17862 14220 17868 14232
rect 17920 14220 17926 14272
rect 20180 14260 20208 14291
rect 20438 14288 20444 14340
rect 20496 14288 20502 14340
rect 20530 14288 20536 14340
rect 20588 14328 20594 14340
rect 21100 14328 21128 14368
rect 21361 14365 21373 14368
rect 21407 14365 21419 14399
rect 21361 14359 21419 14365
rect 21910 14356 21916 14408
rect 21968 14356 21974 14408
rect 22005 14399 22063 14405
rect 22005 14365 22017 14399
rect 22051 14396 22063 14399
rect 22186 14396 22192 14408
rect 22051 14368 22192 14396
rect 22051 14365 22063 14368
rect 22005 14359 22063 14365
rect 22186 14356 22192 14368
rect 22244 14356 22250 14408
rect 20588 14300 21128 14328
rect 20588 14288 20594 14300
rect 21174 14288 21180 14340
rect 21232 14288 21238 14340
rect 21266 14288 21272 14340
rect 21324 14288 21330 14340
rect 21729 14331 21787 14337
rect 21729 14328 21741 14331
rect 21560 14300 21741 14328
rect 20898 14260 20904 14272
rect 20180 14232 20904 14260
rect 20898 14220 20904 14232
rect 20956 14260 20962 14272
rect 21358 14260 21364 14272
rect 20956 14232 21364 14260
rect 20956 14220 20962 14232
rect 21358 14220 21364 14232
rect 21416 14220 21422 14272
rect 21560 14269 21588 14300
rect 21729 14297 21741 14300
rect 21775 14297 21787 14331
rect 21729 14291 21787 14297
rect 22094 14288 22100 14340
rect 22152 14288 22158 14340
rect 21545 14263 21603 14269
rect 21545 14229 21557 14263
rect 21591 14229 21603 14263
rect 22112 14260 22140 14288
rect 22189 14263 22247 14269
rect 22189 14260 22201 14263
rect 22112 14232 22201 14260
rect 21545 14223 21603 14229
rect 22189 14229 22201 14232
rect 22235 14229 22247 14263
rect 22388 14260 22416 14504
rect 23934 14492 23940 14544
rect 23992 14532 23998 14544
rect 26418 14532 26424 14544
rect 23992 14504 26424 14532
rect 23992 14492 23998 14504
rect 26418 14492 26424 14504
rect 26476 14532 26482 14544
rect 29270 14532 29276 14544
rect 26476 14504 29276 14532
rect 26476 14492 26482 14504
rect 29270 14492 29276 14504
rect 29328 14532 29334 14544
rect 30190 14532 30196 14544
rect 29328 14504 30196 14532
rect 29328 14492 29334 14504
rect 30190 14492 30196 14504
rect 30248 14492 30254 14544
rect 32508 14504 34008 14532
rect 22741 14467 22799 14473
rect 22741 14433 22753 14467
rect 22787 14464 22799 14467
rect 23198 14464 23204 14476
rect 22787 14436 23204 14464
rect 22787 14433 22799 14436
rect 22741 14427 22799 14433
rect 23198 14424 23204 14436
rect 23256 14424 23262 14476
rect 24670 14424 24676 14476
rect 24728 14464 24734 14476
rect 25682 14464 25688 14476
rect 24728 14436 25688 14464
rect 24728 14424 24734 14436
rect 25682 14424 25688 14436
rect 25740 14424 25746 14476
rect 27522 14424 27528 14476
rect 27580 14464 27586 14476
rect 29638 14464 29644 14476
rect 27580 14436 29644 14464
rect 27580 14424 27586 14436
rect 29638 14424 29644 14436
rect 29696 14424 29702 14476
rect 22462 14356 22468 14408
rect 22520 14356 22526 14408
rect 27706 14356 27712 14408
rect 27764 14356 27770 14408
rect 28258 14356 28264 14408
rect 28316 14356 28322 14408
rect 29362 14356 29368 14408
rect 29420 14396 29426 14408
rect 30282 14396 30288 14408
rect 29420 14368 30288 14396
rect 29420 14356 29426 14368
rect 30282 14356 30288 14368
rect 30340 14356 30346 14408
rect 30837 14399 30895 14405
rect 30837 14396 30849 14399
rect 30668 14368 30849 14396
rect 23198 14288 23204 14340
rect 23256 14288 23262 14340
rect 24762 14288 24768 14340
rect 24820 14328 24826 14340
rect 27982 14328 27988 14340
rect 24820 14300 27988 14328
rect 24820 14288 24826 14300
rect 27982 14288 27988 14300
rect 28040 14288 28046 14340
rect 24780 14260 24808 14288
rect 30668 14272 30696 14368
rect 30837 14365 30849 14368
rect 30883 14365 30895 14399
rect 30837 14359 30895 14365
rect 30929 14399 30987 14405
rect 30929 14365 30941 14399
rect 30975 14396 30987 14399
rect 31113 14399 31171 14405
rect 31113 14396 31125 14399
rect 30975 14368 31125 14396
rect 30975 14365 30987 14368
rect 30929 14359 30987 14365
rect 31113 14365 31125 14368
rect 31159 14365 31171 14399
rect 32508 14382 32536 14504
rect 33980 14476 34008 14504
rect 38286 14492 38292 14544
rect 38344 14492 38350 14544
rect 33134 14424 33140 14476
rect 33192 14424 33198 14476
rect 33318 14424 33324 14476
rect 33376 14464 33382 14476
rect 33781 14467 33839 14473
rect 33781 14464 33793 14467
rect 33376 14436 33793 14464
rect 33376 14424 33382 14436
rect 33781 14433 33793 14436
rect 33827 14433 33839 14467
rect 33781 14427 33839 14433
rect 33962 14424 33968 14476
rect 34020 14424 34026 14476
rect 33152 14396 33180 14424
rect 35345 14399 35403 14405
rect 35345 14396 35357 14399
rect 33152 14368 35357 14396
rect 31113 14359 31171 14365
rect 35345 14365 35357 14368
rect 35391 14365 35403 14399
rect 35345 14359 35403 14365
rect 37642 14356 37648 14408
rect 37700 14356 37706 14408
rect 31386 14288 31392 14340
rect 31444 14288 31450 14340
rect 33502 14288 33508 14340
rect 33560 14288 33566 14340
rect 22388 14232 24808 14260
rect 22189 14223 22247 14229
rect 24854 14220 24860 14272
rect 24912 14260 24918 14272
rect 27801 14263 27859 14269
rect 27801 14260 27813 14263
rect 24912 14232 27813 14260
rect 24912 14220 24918 14232
rect 27801 14229 27813 14232
rect 27847 14260 27859 14263
rect 29086 14260 29092 14272
rect 27847 14232 29092 14260
rect 27847 14229 27859 14232
rect 27801 14223 27859 14229
rect 29086 14220 29092 14232
rect 29144 14220 29150 14272
rect 30650 14220 30656 14272
rect 30708 14220 30714 14272
rect 33520 14260 33548 14288
rect 33597 14263 33655 14269
rect 33597 14260 33609 14263
rect 33520 14232 33609 14260
rect 33597 14229 33609 14232
rect 33643 14229 33655 14263
rect 33597 14223 33655 14229
rect 33689 14263 33747 14269
rect 33689 14229 33701 14263
rect 33735 14260 33747 14263
rect 33778 14260 33784 14272
rect 33735 14232 33784 14260
rect 33735 14229 33747 14232
rect 33689 14223 33747 14229
rect 33778 14220 33784 14232
rect 33836 14220 33842 14272
rect 35434 14220 35440 14272
rect 35492 14220 35498 14272
rect 1104 14170 38272 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 38272 14170
rect 1104 14096 38272 14118
rect 4614 14016 4620 14068
rect 4672 14056 4678 14068
rect 4801 14059 4859 14065
rect 4801 14056 4813 14059
rect 4672 14028 4813 14056
rect 4672 14016 4678 14028
rect 4801 14025 4813 14028
rect 4847 14025 4859 14059
rect 4801 14019 4859 14025
rect 5169 14059 5227 14065
rect 5169 14025 5181 14059
rect 5215 14056 5227 14059
rect 5258 14056 5264 14068
rect 5215 14028 5264 14056
rect 5215 14025 5227 14028
rect 5169 14019 5227 14025
rect 5258 14016 5264 14028
rect 5316 14016 5322 14068
rect 6546 14016 6552 14068
rect 6604 14016 6610 14068
rect 7558 14016 7564 14068
rect 7616 14016 7622 14068
rect 7668 14028 11560 14056
rect 1765 13991 1823 13997
rect 1765 13957 1777 13991
rect 1811 13988 1823 13991
rect 6454 13988 6460 14000
rect 1811 13960 6460 13988
rect 1811 13957 1823 13960
rect 1765 13951 1823 13957
rect 6454 13948 6460 13960
rect 6512 13948 6518 14000
rect 4893 13923 4951 13929
rect 4893 13920 4905 13923
rect 4816 13892 4905 13920
rect 1486 13812 1492 13864
rect 1544 13812 1550 13864
rect 4816 13796 4844 13892
rect 4893 13889 4905 13892
rect 4939 13889 4951 13923
rect 4893 13883 4951 13889
rect 5353 13923 5411 13929
rect 5353 13889 5365 13923
rect 5399 13920 5411 13923
rect 6564 13920 6592 14016
rect 5399 13892 6592 13920
rect 7469 13923 7527 13929
rect 5399 13889 5411 13892
rect 5353 13883 5411 13889
rect 7469 13889 7481 13923
rect 7515 13920 7527 13923
rect 7576 13920 7604 14016
rect 7515 13892 7604 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 7668 13852 7696 14028
rect 9582 13948 9588 14000
rect 9640 13988 9646 14000
rect 11149 13991 11207 13997
rect 11149 13988 11161 13991
rect 9640 13960 11161 13988
rect 9640 13948 9646 13960
rect 11149 13957 11161 13960
rect 11195 13957 11207 13991
rect 11149 13951 11207 13957
rect 9766 13880 9772 13932
rect 9824 13880 9830 13932
rect 9861 13923 9919 13929
rect 9861 13889 9873 13923
rect 9907 13920 9919 13923
rect 9950 13920 9956 13932
rect 9907 13892 9956 13920
rect 9907 13889 9919 13892
rect 9861 13883 9919 13889
rect 9950 13880 9956 13892
rect 10008 13880 10014 13932
rect 10045 13923 10103 13929
rect 10045 13889 10057 13923
rect 10091 13889 10103 13923
rect 10045 13883 10103 13889
rect 9784 13852 9812 13880
rect 10060 13852 10088 13883
rect 10134 13880 10140 13932
rect 10192 13880 10198 13932
rect 10318 13880 10324 13932
rect 10376 13880 10382 13932
rect 10502 13880 10508 13932
rect 10560 13920 10566 13932
rect 10873 13923 10931 13929
rect 10873 13920 10885 13923
rect 10560 13892 10885 13920
rect 10560 13880 10566 13892
rect 10873 13889 10885 13892
rect 10919 13889 10931 13923
rect 10873 13883 10931 13889
rect 5736 13824 7696 13852
rect 9692 13824 10088 13852
rect 4798 13744 4804 13796
rect 4856 13744 4862 13796
rect 4522 13676 4528 13728
rect 4580 13716 4586 13728
rect 5258 13716 5264 13728
rect 4580 13688 5264 13716
rect 4580 13676 4586 13688
rect 5258 13676 5264 13688
rect 5316 13716 5322 13728
rect 5736 13716 5764 13824
rect 9122 13744 9128 13796
rect 9180 13784 9186 13796
rect 9692 13784 9720 13824
rect 10226 13812 10232 13864
rect 10284 13852 10290 13864
rect 10689 13855 10747 13861
rect 10689 13852 10701 13855
rect 10284 13824 10701 13852
rect 10284 13812 10290 13824
rect 10689 13821 10701 13824
rect 10735 13821 10747 13855
rect 10689 13815 10747 13821
rect 9180 13756 9720 13784
rect 9180 13744 9186 13756
rect 10594 13744 10600 13796
rect 10652 13744 10658 13796
rect 10888 13784 10916 13883
rect 11532 13852 11560 14028
rect 11790 14016 11796 14068
rect 11848 14056 11854 14068
rect 11885 14059 11943 14065
rect 11885 14056 11897 14059
rect 11848 14028 11897 14056
rect 11848 14016 11854 14028
rect 11885 14025 11897 14028
rect 11931 14025 11943 14059
rect 13909 14059 13967 14065
rect 11885 14019 11943 14025
rect 11992 14028 12572 14056
rect 11992 13988 12020 14028
rect 11624 13960 12020 13988
rect 12084 13960 12296 13988
rect 11624 13932 11652 13960
rect 11606 13880 11612 13932
rect 11664 13880 11670 13932
rect 11974 13880 11980 13932
rect 12032 13920 12038 13932
rect 12084 13920 12112 13960
rect 12268 13929 12296 13960
rect 12032 13892 12112 13920
rect 12161 13923 12219 13929
rect 12032 13880 12038 13892
rect 12161 13889 12173 13923
rect 12207 13889 12219 13923
rect 12161 13883 12219 13889
rect 12253 13923 12311 13929
rect 12253 13889 12265 13923
rect 12299 13889 12311 13923
rect 12253 13883 12311 13889
rect 12176 13852 12204 13883
rect 12342 13880 12348 13932
rect 12400 13880 12406 13932
rect 12544 13929 12572 14028
rect 13909 14025 13921 14059
rect 13955 14025 13967 14059
rect 13909 14019 13967 14025
rect 14277 14059 14335 14065
rect 14277 14025 14289 14059
rect 14323 14056 14335 14059
rect 14734 14056 14740 14068
rect 14323 14028 14740 14056
rect 14323 14025 14335 14028
rect 14277 14019 14335 14025
rect 12529 13923 12587 13929
rect 12529 13889 12541 13923
rect 12575 13889 12587 13923
rect 12529 13883 12587 13889
rect 13725 13923 13783 13929
rect 13725 13889 13737 13923
rect 13771 13920 13783 13923
rect 13924 13920 13952 14019
rect 14734 14016 14740 14028
rect 14792 14016 14798 14068
rect 14918 14016 14924 14068
rect 14976 14016 14982 14068
rect 15286 14016 15292 14068
rect 15344 14056 15350 14068
rect 16390 14056 16396 14068
rect 15344 14028 16396 14056
rect 15344 14016 15350 14028
rect 16390 14016 16396 14028
rect 16448 14056 16454 14068
rect 16448 14028 18367 14056
rect 16448 14016 16454 14028
rect 14369 13991 14427 13997
rect 14369 13957 14381 13991
rect 14415 13988 14427 13991
rect 14936 13988 14964 14016
rect 14415 13960 14688 13988
rect 14415 13957 14427 13960
rect 14369 13951 14427 13957
rect 14660 13932 14688 13960
rect 14752 13960 14964 13988
rect 14550 13920 14556 13932
rect 13771 13892 13952 13920
rect 14476 13892 14556 13920
rect 13771 13889 13783 13892
rect 13725 13883 13783 13889
rect 14476 13861 14504 13892
rect 14550 13880 14556 13892
rect 14608 13880 14614 13932
rect 14642 13880 14648 13932
rect 14700 13880 14706 13932
rect 14752 13929 14780 13960
rect 17494 13948 17500 14000
rect 17552 13948 17558 14000
rect 17972 13960 18276 13988
rect 14737 13923 14795 13929
rect 14737 13889 14749 13923
rect 14783 13889 14795 13923
rect 14737 13883 14795 13889
rect 16114 13880 16120 13932
rect 16172 13880 16178 13932
rect 17972 13929 18000 13960
rect 18248 13932 18276 13960
rect 17772 13923 17830 13929
rect 17772 13920 17784 13923
rect 16224 13892 17784 13920
rect 14461 13855 14519 13861
rect 11532 13824 14376 13852
rect 14348 13784 14376 13824
rect 14461 13821 14473 13855
rect 14507 13821 14519 13855
rect 16224 13852 16252 13892
rect 17772 13889 17784 13892
rect 17818 13889 17830 13923
rect 17772 13883 17830 13889
rect 17865 13923 17923 13929
rect 17865 13889 17877 13923
rect 17911 13889 17923 13923
rect 17865 13883 17923 13889
rect 17957 13923 18015 13929
rect 17957 13889 17969 13923
rect 18003 13889 18015 13923
rect 17957 13883 18015 13889
rect 14461 13815 14519 13821
rect 14568 13824 16252 13852
rect 14568 13784 14596 13824
rect 17793 13796 17821 13883
rect 10888 13756 13676 13784
rect 14348 13756 14596 13784
rect 5316 13688 5764 13716
rect 5316 13676 5322 13688
rect 7098 13676 7104 13728
rect 7156 13716 7162 13728
rect 7285 13719 7343 13725
rect 7285 13716 7297 13719
rect 7156 13688 7297 13716
rect 7156 13676 7162 13688
rect 7285 13685 7297 13688
rect 7331 13685 7343 13719
rect 7285 13679 7343 13685
rect 9674 13676 9680 13728
rect 9732 13716 9738 13728
rect 9950 13716 9956 13728
rect 9732 13688 9956 13716
rect 9732 13676 9738 13688
rect 9950 13676 9956 13688
rect 10008 13676 10014 13728
rect 10042 13676 10048 13728
rect 10100 13676 10106 13728
rect 13354 13676 13360 13728
rect 13412 13716 13418 13728
rect 13541 13719 13599 13725
rect 13541 13716 13553 13719
rect 13412 13688 13553 13716
rect 13412 13676 13418 13688
rect 13541 13685 13553 13688
rect 13587 13685 13599 13719
rect 13648 13716 13676 13756
rect 17770 13744 17776 13796
rect 17828 13744 17834 13796
rect 17880 13784 17908 13883
rect 18138 13880 18144 13932
rect 18196 13880 18202 13932
rect 18230 13880 18236 13932
rect 18288 13880 18294 13932
rect 18339 13852 18367 14028
rect 18690 14016 18696 14068
rect 18748 14056 18754 14068
rect 19429 14059 19487 14065
rect 18748 14028 19380 14056
rect 18748 14016 18754 14028
rect 18598 13948 18604 14000
rect 18656 13988 18662 14000
rect 19153 13991 19211 13997
rect 19153 13988 19165 13991
rect 18656 13960 19165 13988
rect 18656 13948 18662 13960
rect 19153 13957 19165 13960
rect 19199 13957 19211 13991
rect 19352 13988 19380 14028
rect 19429 14025 19441 14059
rect 19475 14056 19487 14059
rect 21726 14056 21732 14068
rect 19475 14028 21732 14056
rect 19475 14025 19487 14028
rect 19429 14019 19487 14025
rect 21726 14016 21732 14028
rect 21784 14016 21790 14068
rect 21821 14059 21879 14065
rect 21821 14025 21833 14059
rect 21867 14056 21879 14059
rect 21910 14056 21916 14068
rect 21867 14028 21916 14056
rect 21867 14025 21879 14028
rect 21821 14019 21879 14025
rect 21910 14016 21916 14028
rect 21968 14016 21974 14068
rect 22462 14016 22468 14068
rect 22520 14056 22526 14068
rect 22649 14059 22707 14065
rect 22649 14056 22661 14059
rect 22520 14028 22661 14056
rect 22520 14016 22526 14028
rect 22649 14025 22661 14028
rect 22695 14025 22707 14059
rect 22649 14019 22707 14025
rect 23382 14016 23388 14068
rect 23440 14016 23446 14068
rect 23474 14016 23480 14068
rect 23532 14016 23538 14068
rect 23753 14059 23811 14065
rect 23753 14025 23765 14059
rect 23799 14056 23811 14059
rect 24302 14056 24308 14068
rect 23799 14028 24308 14056
rect 23799 14025 23811 14028
rect 23753 14019 23811 14025
rect 24302 14016 24308 14028
rect 24360 14016 24366 14068
rect 25498 14016 25504 14068
rect 25556 14056 25562 14068
rect 29178 14056 29184 14068
rect 25556 14028 29184 14056
rect 25556 14016 25562 14028
rect 29178 14016 29184 14028
rect 29236 14016 29242 14068
rect 31386 14016 31392 14068
rect 31444 14016 31450 14068
rect 32125 14059 32183 14065
rect 32125 14056 32137 14059
rect 31726 14028 32137 14056
rect 20162 13988 20168 14000
rect 19352 13960 20168 13988
rect 19153 13951 19211 13957
rect 20162 13948 20168 13960
rect 20220 13948 20226 14000
rect 20438 13948 20444 14000
rect 20496 13988 20502 14000
rect 21453 13991 21511 13997
rect 20496 13960 21036 13988
rect 20496 13948 20502 13960
rect 18506 13880 18512 13932
rect 18564 13920 18570 13932
rect 18877 13923 18935 13929
rect 18877 13920 18889 13923
rect 18564 13892 18889 13920
rect 18564 13880 18570 13892
rect 18877 13889 18889 13892
rect 18923 13889 18935 13923
rect 18877 13883 18935 13889
rect 19058 13880 19064 13932
rect 19116 13880 19122 13932
rect 19245 13923 19303 13929
rect 19245 13889 19257 13923
rect 19291 13920 19303 13923
rect 20898 13920 20904 13932
rect 19291 13892 20904 13920
rect 19291 13889 19303 13892
rect 19245 13883 19303 13889
rect 20898 13880 20904 13892
rect 20956 13880 20962 13932
rect 20530 13852 20536 13864
rect 18339 13824 20536 13852
rect 20530 13812 20536 13824
rect 20588 13812 20594 13864
rect 18598 13784 18604 13796
rect 17880 13756 18604 13784
rect 18598 13744 18604 13756
rect 18656 13784 18662 13796
rect 18874 13784 18880 13796
rect 18656 13756 18880 13784
rect 18656 13744 18662 13756
rect 18874 13744 18880 13756
rect 18932 13744 18938 13796
rect 21008 13784 21036 13960
rect 21453 13957 21465 13991
rect 21499 13988 21511 13991
rect 22189 13991 22247 13997
rect 22189 13988 22201 13991
rect 21499 13960 22201 13988
rect 21499 13957 21511 13960
rect 21453 13951 21511 13957
rect 22189 13957 22201 13960
rect 22235 13957 22247 13991
rect 23492 13988 23520 14016
rect 23845 13991 23903 13997
rect 23845 13988 23857 13991
rect 23492 13960 23857 13988
rect 22189 13951 22247 13957
rect 23845 13957 23857 13960
rect 23891 13957 23903 13991
rect 23845 13951 23903 13957
rect 24118 13948 24124 14000
rect 24176 13988 24182 14000
rect 25516 13988 25544 14016
rect 24176 13960 25544 13988
rect 24176 13948 24182 13960
rect 26326 13948 26332 14000
rect 26384 13948 26390 14000
rect 26694 13948 26700 14000
rect 26752 13988 26758 14000
rect 26752 13960 27936 13988
rect 26752 13948 26758 13960
rect 21082 13880 21088 13932
rect 21140 13880 21146 13932
rect 21269 13923 21327 13929
rect 21269 13889 21281 13923
rect 21315 13920 21327 13923
rect 21358 13920 21364 13932
rect 21315 13892 21364 13920
rect 21315 13889 21327 13892
rect 21269 13883 21327 13889
rect 21358 13880 21364 13892
rect 21416 13880 21422 13932
rect 21910 13880 21916 13932
rect 21968 13920 21974 13932
rect 22005 13923 22063 13929
rect 22005 13920 22017 13923
rect 21968 13892 22017 13920
rect 21968 13880 21974 13892
rect 22005 13889 22017 13892
rect 22051 13889 22063 13923
rect 22005 13883 22063 13889
rect 22097 13923 22155 13929
rect 22097 13889 22109 13923
rect 22143 13889 22155 13923
rect 22097 13883 22155 13889
rect 22112 13784 22140 13883
rect 22278 13880 22284 13932
rect 22336 13920 22342 13932
rect 22373 13923 22431 13929
rect 22373 13920 22385 13923
rect 22336 13892 22385 13920
rect 22336 13880 22342 13892
rect 22373 13889 22385 13892
rect 22419 13920 22431 13923
rect 22462 13920 22468 13932
rect 22419 13892 22468 13920
rect 22419 13889 22431 13892
rect 22373 13883 22431 13889
rect 22462 13880 22468 13892
rect 22520 13880 22526 13932
rect 22646 13880 22652 13932
rect 22704 13920 22710 13932
rect 22741 13923 22799 13929
rect 22741 13920 22753 13923
rect 22704 13892 22753 13920
rect 22704 13880 22710 13892
rect 22741 13889 22753 13892
rect 22787 13889 22799 13923
rect 26344 13920 26372 13948
rect 27525 13923 27583 13929
rect 27525 13920 27537 13923
rect 26344 13892 27537 13920
rect 22741 13883 22799 13889
rect 27525 13889 27537 13892
rect 27571 13920 27583 13923
rect 27908 13920 27936 13960
rect 27982 13948 27988 14000
rect 28040 13988 28046 14000
rect 29917 13991 29975 13997
rect 28040 13960 28994 13988
rect 28040 13948 28046 13960
rect 28810 13920 28816 13932
rect 27571 13892 27844 13920
rect 27908 13892 28816 13920
rect 27571 13889 27583 13892
rect 27525 13883 27583 13889
rect 23937 13855 23995 13861
rect 23937 13821 23949 13855
rect 23983 13821 23995 13855
rect 27617 13855 27675 13861
rect 27617 13852 27629 13855
rect 23937 13815 23995 13821
rect 24872 13824 27629 13852
rect 21008 13756 22140 13784
rect 23474 13744 23480 13796
rect 23532 13784 23538 13796
rect 23952 13784 23980 13815
rect 23532 13756 23980 13784
rect 23532 13744 23538 13756
rect 24302 13744 24308 13796
rect 24360 13784 24366 13796
rect 24872 13784 24900 13824
rect 27617 13821 27629 13824
rect 27663 13821 27675 13855
rect 27816 13852 27844 13892
rect 28810 13880 28816 13892
rect 28868 13880 28874 13932
rect 28258 13852 28264 13864
rect 27816 13824 28264 13852
rect 27617 13815 27675 13821
rect 28258 13812 28264 13824
rect 28316 13812 28322 13864
rect 24360 13756 24900 13784
rect 24360 13744 24366 13756
rect 24946 13744 24952 13796
rect 25004 13744 25010 13796
rect 28350 13784 28356 13796
rect 27540 13756 28356 13784
rect 14826 13716 14832 13728
rect 13648 13688 14832 13716
rect 13541 13679 13599 13685
rect 14826 13676 14832 13688
rect 14884 13676 14890 13728
rect 15000 13719 15058 13725
rect 15000 13685 15012 13719
rect 15046 13716 15058 13719
rect 15194 13716 15200 13728
rect 15046 13688 15200 13716
rect 15046 13685 15058 13688
rect 15000 13679 15058 13685
rect 15194 13676 15200 13688
rect 15252 13676 15258 13728
rect 16482 13676 16488 13728
rect 16540 13676 16546 13728
rect 17034 13676 17040 13728
rect 17092 13716 17098 13728
rect 24670 13716 24676 13728
rect 17092 13688 24676 13716
rect 17092 13676 17098 13688
rect 24670 13676 24676 13688
rect 24728 13676 24734 13728
rect 24964 13716 24992 13744
rect 26786 13716 26792 13728
rect 24964 13688 26792 13716
rect 26786 13676 26792 13688
rect 26844 13676 26850 13728
rect 27246 13676 27252 13728
rect 27304 13716 27310 13728
rect 27540 13725 27568 13756
rect 28350 13744 28356 13756
rect 28408 13744 28414 13796
rect 28966 13784 28994 13960
rect 29917 13957 29929 13991
rect 29963 13957 29975 13991
rect 29917 13951 29975 13957
rect 29178 13880 29184 13932
rect 29236 13880 29242 13932
rect 29270 13880 29276 13932
rect 29328 13920 29334 13932
rect 29687 13923 29745 13929
rect 29687 13920 29699 13923
rect 29328 13892 29699 13920
rect 29328 13880 29334 13892
rect 29687 13889 29699 13892
rect 29733 13889 29745 13923
rect 29687 13883 29745 13889
rect 29822 13880 29828 13932
rect 29880 13880 29886 13932
rect 29932 13920 29960 13951
rect 30101 13923 30159 13929
rect 29932 13892 30016 13920
rect 29196 13852 29224 13880
rect 29988 13852 30016 13892
rect 30101 13889 30113 13923
rect 30147 13889 30159 13923
rect 30101 13883 30159 13889
rect 31573 13923 31631 13929
rect 31573 13889 31585 13923
rect 31619 13920 31631 13923
rect 31726 13920 31754 14028
rect 32125 14025 32137 14028
rect 32171 14025 32183 14059
rect 32125 14019 32183 14025
rect 32490 14016 32496 14068
rect 32548 14016 32554 14068
rect 32585 14059 32643 14065
rect 32585 14025 32597 14059
rect 32631 14056 32643 14059
rect 33778 14056 33784 14068
rect 32631 14028 33784 14056
rect 32631 14025 32643 14028
rect 32585 14019 32643 14025
rect 33778 14016 33784 14028
rect 33836 14016 33842 14068
rect 35434 14016 35440 14068
rect 35492 14016 35498 14068
rect 31619 13892 31754 13920
rect 31864 13892 33640 13920
rect 31619 13889 31631 13892
rect 31573 13883 31631 13889
rect 29196 13824 30016 13852
rect 30116 13852 30144 13883
rect 31864 13852 31892 13892
rect 33612 13864 33640 13892
rect 33962 13880 33968 13932
rect 34020 13880 34026 13932
rect 35345 13923 35403 13929
rect 35345 13889 35357 13923
rect 35391 13920 35403 13923
rect 35452 13920 35480 14016
rect 35391 13892 35480 13920
rect 35391 13889 35403 13892
rect 35345 13883 35403 13889
rect 30116 13824 31892 13852
rect 32677 13855 32735 13861
rect 28966 13756 29692 13784
rect 27525 13719 27583 13725
rect 27525 13716 27537 13719
rect 27304 13688 27537 13716
rect 27304 13676 27310 13688
rect 27525 13685 27537 13688
rect 27571 13685 27583 13719
rect 27525 13679 27583 13685
rect 27798 13676 27804 13728
rect 27856 13716 27862 13728
rect 27893 13719 27951 13725
rect 27893 13716 27905 13719
rect 27856 13688 27905 13716
rect 27856 13676 27862 13688
rect 27893 13685 27905 13688
rect 27939 13685 27951 13719
rect 27893 13679 27951 13685
rect 29546 13676 29552 13728
rect 29604 13676 29610 13728
rect 29664 13716 29692 13756
rect 30116 13716 30144 13824
rect 32677 13821 32689 13855
rect 32723 13821 32735 13855
rect 32677 13815 32735 13821
rect 30374 13744 30380 13796
rect 30432 13784 30438 13796
rect 31294 13784 31300 13796
rect 30432 13756 31300 13784
rect 30432 13744 30438 13756
rect 31294 13744 31300 13756
rect 31352 13784 31358 13796
rect 32692 13784 32720 13815
rect 33594 13812 33600 13864
rect 33652 13812 33658 13864
rect 31352 13756 32720 13784
rect 31352 13744 31358 13756
rect 32692 13728 32720 13756
rect 29664 13688 30144 13716
rect 32674 13676 32680 13728
rect 32732 13676 32738 13728
rect 34054 13676 34060 13728
rect 34112 13716 34118 13728
rect 35081 13719 35139 13725
rect 35081 13716 35093 13719
rect 34112 13688 35093 13716
rect 34112 13676 34118 13688
rect 35081 13685 35093 13688
rect 35127 13685 35139 13719
rect 35081 13679 35139 13685
rect 1104 13626 38272 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38272 13626
rect 1104 13552 38272 13574
rect 8478 13472 8484 13524
rect 8536 13472 8542 13524
rect 9861 13515 9919 13521
rect 9861 13481 9873 13515
rect 9907 13512 9919 13515
rect 9907 13484 11376 13512
rect 9907 13481 9919 13484
rect 9861 13475 9919 13481
rect 10042 13404 10048 13456
rect 10100 13404 10106 13456
rect 10502 13404 10508 13456
rect 10560 13404 10566 13456
rect 10594 13404 10600 13456
rect 10652 13444 10658 13456
rect 10652 13416 11284 13444
rect 10652 13404 10658 13416
rect 5445 13379 5503 13385
rect 5445 13345 5457 13379
rect 5491 13376 5503 13379
rect 5534 13376 5540 13388
rect 5491 13348 5540 13376
rect 5491 13345 5503 13348
rect 5445 13339 5503 13345
rect 5534 13336 5540 13348
rect 5592 13336 5598 13388
rect 7009 13379 7067 13385
rect 7009 13345 7021 13379
rect 7055 13376 7067 13379
rect 7098 13376 7104 13388
rect 7055 13348 7104 13376
rect 7055 13345 7067 13348
rect 7009 13339 7067 13345
rect 7098 13336 7104 13348
rect 7156 13336 7162 13388
rect 9490 13336 9496 13388
rect 9548 13376 9554 13388
rect 10060 13376 10088 13404
rect 9548 13348 9812 13376
rect 10060 13348 10916 13376
rect 9548 13336 9554 13348
rect 3970 13268 3976 13320
rect 4028 13268 4034 13320
rect 5258 13268 5264 13320
rect 5316 13268 5322 13320
rect 6454 13268 6460 13320
rect 6512 13268 6518 13320
rect 6549 13311 6607 13317
rect 6549 13277 6561 13311
rect 6595 13308 6607 13311
rect 6733 13311 6791 13317
rect 6733 13308 6745 13311
rect 6595 13280 6745 13308
rect 6595 13277 6607 13280
rect 6549 13271 6607 13277
rect 6733 13277 6745 13280
rect 6779 13277 6791 13311
rect 9030 13308 9036 13320
rect 8142 13280 9036 13308
rect 6733 13271 6791 13277
rect 9030 13268 9036 13280
rect 9088 13268 9094 13320
rect 9784 13317 9812 13348
rect 10244 13317 10272 13348
rect 9585 13311 9643 13317
rect 9585 13277 9597 13311
rect 9631 13277 9643 13311
rect 9585 13271 9643 13277
rect 9769 13311 9827 13317
rect 9769 13277 9781 13311
rect 9815 13308 9827 13311
rect 10045 13311 10103 13317
rect 10045 13308 10057 13311
rect 9815 13280 10057 13308
rect 9815 13277 9827 13280
rect 9769 13271 9827 13277
rect 10045 13277 10057 13280
rect 10091 13277 10103 13311
rect 10045 13271 10103 13277
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 5353 13243 5411 13249
rect 5353 13209 5365 13243
rect 5399 13240 5411 13243
rect 6914 13240 6920 13252
rect 5399 13212 6920 13240
rect 5399 13209 5411 13212
rect 5353 13203 5411 13209
rect 6914 13200 6920 13212
rect 6972 13200 6978 13252
rect 9600 13184 9628 13271
rect 10318 13268 10324 13320
rect 10376 13308 10382 13320
rect 10888 13317 10916 13348
rect 11256 13317 11284 13416
rect 11348 13385 11376 13484
rect 12342 13472 12348 13524
rect 12400 13512 12406 13524
rect 12805 13515 12863 13521
rect 12805 13512 12817 13515
rect 12400 13484 12817 13512
rect 12400 13472 12406 13484
rect 12805 13481 12817 13484
rect 12851 13481 12863 13515
rect 12805 13475 12863 13481
rect 13078 13472 13084 13524
rect 13136 13512 13142 13524
rect 13262 13512 13268 13524
rect 13136 13484 13268 13512
rect 13136 13472 13142 13484
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 15194 13472 15200 13524
rect 15252 13472 15258 13524
rect 17957 13515 18015 13521
rect 15304 13484 15884 13512
rect 12621 13447 12679 13453
rect 12621 13413 12633 13447
rect 12667 13444 12679 13447
rect 14550 13444 14556 13456
rect 12667 13416 14556 13444
rect 12667 13413 12679 13416
rect 12621 13407 12679 13413
rect 14550 13404 14556 13416
rect 14608 13404 14614 13456
rect 14734 13404 14740 13456
rect 14792 13444 14798 13456
rect 15304 13444 15332 13484
rect 14792 13416 15332 13444
rect 15565 13447 15623 13453
rect 14792 13404 14798 13416
rect 15565 13413 15577 13447
rect 15611 13413 15623 13447
rect 15565 13407 15623 13413
rect 11333 13379 11391 13385
rect 11333 13345 11345 13379
rect 11379 13376 11391 13379
rect 11379 13348 12020 13376
rect 11379 13345 11391 13348
rect 11333 13339 11391 13345
rect 10689 13311 10747 13317
rect 10689 13308 10701 13311
rect 10376 13280 10701 13308
rect 10376 13268 10382 13280
rect 10689 13277 10701 13280
rect 10735 13277 10747 13311
rect 10689 13271 10747 13277
rect 10873 13311 10931 13317
rect 10873 13277 10885 13311
rect 10919 13277 10931 13311
rect 10873 13271 10931 13277
rect 11241 13311 11299 13317
rect 11241 13277 11253 13311
rect 11287 13277 11299 13311
rect 11241 13271 11299 13277
rect 11882 13268 11888 13320
rect 11940 13268 11946 13320
rect 11992 13317 12020 13348
rect 12084 13348 12664 13376
rect 11977 13311 12035 13317
rect 11977 13277 11989 13311
rect 12023 13277 12035 13311
rect 11977 13271 12035 13277
rect 10597 13243 10655 13249
rect 10597 13209 10609 13243
rect 10643 13209 10655 13243
rect 10597 13203 10655 13209
rect 3878 13132 3884 13184
rect 3936 13132 3942 13184
rect 4706 13132 4712 13184
rect 4764 13172 4770 13184
rect 4893 13175 4951 13181
rect 4893 13172 4905 13175
rect 4764 13144 4905 13172
rect 4764 13132 4770 13144
rect 4893 13141 4905 13144
rect 4939 13141 4951 13175
rect 4893 13135 4951 13141
rect 9582 13132 9588 13184
rect 9640 13132 9646 13184
rect 9766 13132 9772 13184
rect 9824 13172 9830 13184
rect 10612 13172 10640 13203
rect 12084 13172 12112 13348
rect 12636 13317 12664 13348
rect 12802 13336 12808 13388
rect 12860 13376 12866 13388
rect 12860 13348 13400 13376
rect 12860 13336 12866 13348
rect 12621 13311 12679 13317
rect 12621 13277 12633 13311
rect 12667 13277 12679 13311
rect 12989 13311 13047 13317
rect 12989 13308 13001 13311
rect 12621 13271 12679 13277
rect 12912 13280 13001 13308
rect 12912 13184 12940 13280
rect 12989 13277 13001 13280
rect 13035 13277 13047 13311
rect 12989 13271 13047 13277
rect 13081 13311 13139 13317
rect 13081 13277 13093 13311
rect 13127 13277 13139 13311
rect 13081 13271 13139 13277
rect 13096 13240 13124 13271
rect 13262 13268 13268 13320
rect 13320 13268 13326 13320
rect 13372 13317 13400 13348
rect 13357 13311 13415 13317
rect 13357 13277 13369 13311
rect 13403 13308 13415 13311
rect 13446 13308 13452 13320
rect 13403 13280 13452 13308
rect 13403 13277 13415 13280
rect 13357 13271 13415 13277
rect 13446 13268 13452 13280
rect 13504 13268 13510 13320
rect 13633 13311 13691 13317
rect 13633 13277 13645 13311
rect 13679 13277 13691 13311
rect 13633 13271 13691 13277
rect 15381 13311 15439 13317
rect 15381 13277 15393 13311
rect 15427 13308 15439 13311
rect 15580 13308 15608 13407
rect 15746 13336 15752 13388
rect 15804 13336 15810 13388
rect 15427 13280 15608 13308
rect 15427 13277 15439 13280
rect 15381 13271 15439 13277
rect 13004 13212 13124 13240
rect 13004 13184 13032 13212
rect 13538 13200 13544 13252
rect 13596 13200 13602 13252
rect 13648 13240 13676 13271
rect 15764 13240 15792 13336
rect 13648 13212 15792 13240
rect 15856 13240 15884 13484
rect 17957 13481 17969 13515
rect 18003 13512 18015 13515
rect 18138 13512 18144 13524
rect 18003 13484 18144 13512
rect 18003 13481 18015 13484
rect 17957 13475 18015 13481
rect 18138 13472 18144 13484
rect 18196 13472 18202 13524
rect 18322 13472 18328 13524
rect 18380 13512 18386 13524
rect 20714 13512 20720 13524
rect 18380 13484 20720 13512
rect 18380 13472 18386 13484
rect 20714 13472 20720 13484
rect 20772 13512 20778 13524
rect 22922 13512 22928 13524
rect 20772 13484 22928 13512
rect 20772 13472 20778 13484
rect 22922 13472 22928 13484
rect 22980 13472 22986 13524
rect 26237 13515 26295 13521
rect 25608 13484 26188 13512
rect 25608 13456 25636 13484
rect 16022 13404 16028 13456
rect 16080 13444 16086 13456
rect 16942 13444 16948 13456
rect 16080 13416 16948 13444
rect 16080 13404 16086 13416
rect 16942 13404 16948 13416
rect 17000 13404 17006 13456
rect 17865 13447 17923 13453
rect 17421 13416 17724 13444
rect 16114 13336 16120 13388
rect 16172 13336 16178 13388
rect 16758 13336 16764 13388
rect 16816 13376 16822 13388
rect 17421 13376 17449 13416
rect 16816 13348 17449 13376
rect 16816 13336 16822 13348
rect 17586 13336 17592 13388
rect 17644 13336 17650 13388
rect 17696 13376 17724 13416
rect 17865 13413 17877 13447
rect 17911 13444 17923 13447
rect 17911 13416 18184 13444
rect 17911 13413 17923 13416
rect 17865 13407 17923 13413
rect 17696 13348 18092 13376
rect 15933 13311 15991 13317
rect 15933 13277 15945 13311
rect 15979 13308 15991 13311
rect 16482 13308 16488 13320
rect 15979 13280 16488 13308
rect 15979 13277 15991 13280
rect 15933 13271 15991 13277
rect 16482 13268 16488 13280
rect 16540 13268 16546 13320
rect 16025 13243 16083 13249
rect 16025 13240 16037 13243
rect 15856 13212 16037 13240
rect 16025 13209 16037 13212
rect 16071 13240 16083 13243
rect 16776 13240 16804 13336
rect 17126 13268 17132 13320
rect 17184 13308 17190 13320
rect 17221 13311 17279 13317
rect 17221 13308 17233 13311
rect 17184 13280 17233 13308
rect 17184 13268 17190 13280
rect 17221 13277 17233 13280
rect 17267 13277 17279 13311
rect 17221 13271 17279 13277
rect 17310 13268 17316 13320
rect 17368 13308 17374 13320
rect 17497 13311 17555 13317
rect 17368 13280 17413 13308
rect 17368 13268 17374 13280
rect 17497 13277 17509 13311
rect 17543 13308 17555 13311
rect 17604 13308 17632 13336
rect 17543 13280 17632 13308
rect 17686 13311 17744 13317
rect 17543 13277 17555 13280
rect 17497 13271 17555 13277
rect 17686 13277 17698 13311
rect 17732 13308 17744 13311
rect 17732 13280 17816 13308
rect 17732 13277 17744 13280
rect 17686 13271 17744 13277
rect 16071 13212 16804 13240
rect 16071 13209 16083 13212
rect 16025 13203 16083 13209
rect 16942 13200 16948 13252
rect 17000 13240 17006 13252
rect 17589 13243 17647 13249
rect 17589 13240 17601 13243
rect 17000 13212 17601 13240
rect 17000 13200 17006 13212
rect 17589 13209 17601 13212
rect 17635 13209 17647 13243
rect 17788 13240 17816 13280
rect 17862 13240 17868 13252
rect 17788 13212 17868 13240
rect 17589 13203 17647 13209
rect 17862 13200 17868 13212
rect 17920 13200 17926 13252
rect 18064 13240 18092 13348
rect 18156 13317 18184 13416
rect 18230 13404 18236 13456
rect 18288 13444 18294 13456
rect 25406 13444 25412 13456
rect 18288 13416 25412 13444
rect 18288 13404 18294 13416
rect 25406 13404 25412 13416
rect 25464 13404 25470 13456
rect 25590 13404 25596 13456
rect 25648 13404 25654 13456
rect 25682 13404 25688 13456
rect 25740 13444 25746 13456
rect 25958 13444 25964 13456
rect 25740 13416 25964 13444
rect 25740 13404 25746 13416
rect 25958 13404 25964 13416
rect 26016 13444 26022 13456
rect 26016 13416 26101 13444
rect 26016 13404 26022 13416
rect 20073 13379 20131 13385
rect 20073 13376 20085 13379
rect 18339 13348 20085 13376
rect 18141 13311 18199 13317
rect 18141 13277 18153 13311
rect 18187 13277 18199 13311
rect 18141 13271 18199 13277
rect 18339 13240 18367 13348
rect 20073 13345 20085 13348
rect 20119 13345 20131 13379
rect 20073 13339 20131 13345
rect 20162 13336 20168 13388
rect 20220 13336 20226 13388
rect 24486 13376 24492 13388
rect 20272 13348 24492 13376
rect 18414 13268 18420 13320
rect 18472 13268 18478 13320
rect 20272 13308 20300 13348
rect 24486 13336 24492 13348
rect 24544 13376 24550 13388
rect 24544 13348 24716 13376
rect 24544 13336 24550 13348
rect 19076 13280 20300 13308
rect 20625 13311 20683 13317
rect 18064 13212 18367 13240
rect 18432 13240 18460 13268
rect 18966 13240 18972 13252
rect 18432 13212 18972 13240
rect 18966 13200 18972 13212
rect 19024 13200 19030 13252
rect 9824 13144 12112 13172
rect 9824 13132 9830 13144
rect 12894 13132 12900 13184
rect 12952 13132 12958 13184
rect 12986 13132 12992 13184
rect 13044 13172 13050 13184
rect 17310 13172 17316 13184
rect 13044 13144 17316 13172
rect 13044 13132 13050 13144
rect 17310 13132 17316 13144
rect 17368 13172 17374 13184
rect 18230 13172 18236 13184
rect 17368 13144 18236 13172
rect 17368 13132 17374 13144
rect 18230 13132 18236 13144
rect 18288 13132 18294 13184
rect 18322 13132 18328 13184
rect 18380 13172 18386 13184
rect 19076 13172 19104 13280
rect 20625 13277 20637 13311
rect 20671 13308 20683 13311
rect 22646 13308 22652 13320
rect 20671 13280 22652 13308
rect 20671 13277 20683 13280
rect 20625 13271 20683 13277
rect 22646 13268 22652 13280
rect 22704 13268 22710 13320
rect 24688 13317 24716 13348
rect 24964 13348 25913 13376
rect 24964 13317 24992 13348
rect 24673 13311 24731 13317
rect 24673 13277 24685 13311
rect 24719 13277 24731 13311
rect 24673 13271 24731 13277
rect 24949 13311 25007 13317
rect 24949 13277 24961 13311
rect 24995 13277 25007 13311
rect 24949 13271 25007 13277
rect 25041 13311 25099 13317
rect 25041 13277 25053 13311
rect 25087 13277 25099 13311
rect 25041 13271 25099 13277
rect 19981 13243 20039 13249
rect 19981 13209 19993 13243
rect 20027 13240 20039 13243
rect 21358 13240 21364 13252
rect 20027 13212 21364 13240
rect 20027 13209 20039 13212
rect 19981 13203 20039 13209
rect 21358 13200 21364 13212
rect 21416 13200 21422 13252
rect 24854 13240 24860 13252
rect 22066 13212 24860 13240
rect 18380 13144 19104 13172
rect 18380 13132 18386 13144
rect 19426 13132 19432 13184
rect 19484 13172 19490 13184
rect 19613 13175 19671 13181
rect 19613 13172 19625 13175
rect 19484 13144 19625 13172
rect 19484 13132 19490 13144
rect 19613 13141 19625 13144
rect 19659 13141 19671 13175
rect 19613 13135 19671 13141
rect 19702 13132 19708 13184
rect 19760 13172 19766 13184
rect 20533 13175 20591 13181
rect 20533 13172 20545 13175
rect 19760 13144 20545 13172
rect 19760 13132 19766 13144
rect 20533 13141 20545 13144
rect 20579 13141 20591 13175
rect 20533 13135 20591 13141
rect 20806 13132 20812 13184
rect 20864 13172 20870 13184
rect 22066 13172 22094 13212
rect 24854 13200 24860 13212
rect 24912 13200 24918 13252
rect 25056 13240 25084 13271
rect 25222 13268 25228 13320
rect 25280 13308 25286 13320
rect 25593 13311 25651 13317
rect 25593 13308 25605 13311
rect 25280 13280 25605 13308
rect 25280 13268 25286 13280
rect 25593 13277 25605 13280
rect 25639 13277 25651 13311
rect 25593 13271 25651 13277
rect 25682 13268 25688 13320
rect 25740 13308 25746 13320
rect 25885 13308 25913 13348
rect 26073 13317 26101 13416
rect 26160 13376 26188 13484
rect 26237 13481 26249 13515
rect 26283 13512 26295 13515
rect 27249 13515 27307 13521
rect 26283 13484 27200 13512
rect 26283 13481 26295 13484
rect 26237 13475 26295 13481
rect 26881 13447 26939 13453
rect 26881 13413 26893 13447
rect 26927 13444 26939 13447
rect 26927 13416 27108 13444
rect 26927 13413 26939 13416
rect 26881 13407 26939 13413
rect 26160 13348 26832 13376
rect 25961 13311 26019 13317
rect 25961 13308 25973 13311
rect 25740 13280 25785 13308
rect 25885 13280 25973 13308
rect 25740 13268 25746 13280
rect 25961 13277 25973 13280
rect 26007 13277 26019 13311
rect 25961 13271 26019 13277
rect 26058 13311 26116 13317
rect 26058 13277 26070 13311
rect 26104 13277 26116 13311
rect 26160 13308 26188 13348
rect 26329 13311 26387 13317
rect 26329 13308 26341 13311
rect 26160 13280 26341 13308
rect 26058 13271 26116 13277
rect 26329 13277 26341 13280
rect 26375 13277 26387 13311
rect 26329 13271 26387 13277
rect 26697 13311 26755 13317
rect 26697 13277 26709 13311
rect 26743 13277 26755 13311
rect 26804 13308 26832 13348
rect 26973 13311 27031 13317
rect 26804 13280 26924 13308
rect 26697 13271 26755 13277
rect 25498 13240 25504 13252
rect 25056 13212 25504 13240
rect 25498 13200 25504 13212
rect 25556 13200 25562 13252
rect 25866 13200 25872 13252
rect 25924 13200 25930 13252
rect 20864 13144 22094 13172
rect 25225 13175 25283 13181
rect 20864 13132 20870 13144
rect 25225 13141 25237 13175
rect 25271 13172 25283 13175
rect 25774 13172 25780 13184
rect 25271 13144 25780 13172
rect 25271 13141 25283 13144
rect 25225 13135 25283 13141
rect 25774 13132 25780 13144
rect 25832 13132 25838 13184
rect 25976 13172 26004 13271
rect 26142 13200 26148 13252
rect 26200 13240 26206 13252
rect 26513 13243 26571 13249
rect 26513 13240 26525 13243
rect 26200 13212 26525 13240
rect 26200 13200 26206 13212
rect 26513 13209 26525 13212
rect 26559 13209 26571 13243
rect 26513 13203 26571 13209
rect 26602 13200 26608 13252
rect 26660 13200 26666 13252
rect 26418 13172 26424 13184
rect 25976 13144 26424 13172
rect 26418 13132 26424 13144
rect 26476 13132 26482 13184
rect 26712 13172 26740 13271
rect 26896 13240 26924 13280
rect 26973 13277 26985 13311
rect 27019 13308 27031 13311
rect 27080 13308 27108 13416
rect 27172 13317 27200 13484
rect 27249 13481 27261 13515
rect 27295 13512 27307 13515
rect 27338 13512 27344 13524
rect 27295 13484 27344 13512
rect 27295 13481 27307 13484
rect 27249 13475 27307 13481
rect 27338 13472 27344 13484
rect 27396 13472 27402 13524
rect 28810 13472 28816 13524
rect 28868 13512 28874 13524
rect 31113 13515 31171 13521
rect 31113 13512 31125 13515
rect 28868 13484 30144 13512
rect 28868 13472 28874 13484
rect 27985 13447 28043 13453
rect 27985 13413 27997 13447
rect 28031 13444 28043 13447
rect 28353 13447 28411 13453
rect 28353 13444 28365 13447
rect 28031 13416 28365 13444
rect 28031 13413 28043 13416
rect 27985 13407 28043 13413
rect 28353 13413 28365 13416
rect 28399 13413 28411 13447
rect 28353 13407 28411 13413
rect 28844 13416 28994 13444
rect 27338 13336 27344 13388
rect 27396 13376 27402 13388
rect 28261 13379 28319 13385
rect 27396 13348 28120 13376
rect 27396 13336 27402 13348
rect 27019 13280 27108 13308
rect 27157 13311 27215 13317
rect 27019 13277 27031 13280
rect 26973 13271 27031 13277
rect 27157 13277 27169 13311
rect 27203 13277 27215 13311
rect 27157 13271 27215 13277
rect 27798 13268 27804 13320
rect 27856 13268 27862 13320
rect 27890 13268 27896 13320
rect 27948 13268 27954 13320
rect 28092 13317 28120 13348
rect 28261 13345 28273 13379
rect 28307 13376 28319 13379
rect 28844 13376 28872 13416
rect 28307 13348 28872 13376
rect 28966 13376 28994 13416
rect 29546 13404 29552 13456
rect 29604 13444 29610 13456
rect 29604 13416 30052 13444
rect 29604 13404 29610 13416
rect 28966 13348 29960 13376
rect 28307 13345 28319 13348
rect 28261 13339 28319 13345
rect 28077 13311 28135 13317
rect 28077 13277 28089 13311
rect 28123 13277 28135 13311
rect 28077 13271 28135 13277
rect 28442 13268 28448 13320
rect 28500 13308 28506 13320
rect 28537 13311 28595 13317
rect 28537 13308 28549 13311
rect 28500 13280 28549 13308
rect 28500 13268 28506 13280
rect 28537 13277 28549 13280
rect 28583 13277 28595 13311
rect 28537 13271 28595 13277
rect 28629 13311 28687 13317
rect 28629 13277 28641 13311
rect 28675 13308 28687 13311
rect 28675 13280 28856 13308
rect 28675 13277 28687 13280
rect 28629 13271 28687 13277
rect 28644 13240 28672 13271
rect 26896 13212 28672 13240
rect 28718 13200 28724 13252
rect 28776 13200 28782 13252
rect 28828 13240 28856 13280
rect 28902 13268 28908 13320
rect 28960 13268 28966 13320
rect 29362 13268 29368 13320
rect 29420 13308 29426 13320
rect 29932 13317 29960 13348
rect 29917 13311 29975 13317
rect 29420 13280 29776 13308
rect 29420 13268 29426 13280
rect 28994 13240 29000 13252
rect 28828 13212 29000 13240
rect 28994 13200 29000 13212
rect 29052 13240 29058 13252
rect 29638 13240 29644 13252
rect 29052 13212 29644 13240
rect 29052 13200 29058 13212
rect 29638 13200 29644 13212
rect 29696 13200 29702 13252
rect 29748 13240 29776 13280
rect 29917 13277 29929 13311
rect 29963 13277 29975 13311
rect 30024 13308 30052 13416
rect 30116 13376 30144 13484
rect 30392 13484 31125 13512
rect 30282 13404 30288 13456
rect 30340 13404 30346 13456
rect 30193 13379 30251 13385
rect 30193 13376 30205 13379
rect 30116 13348 30205 13376
rect 30193 13345 30205 13348
rect 30239 13345 30251 13379
rect 30193 13339 30251 13345
rect 30098 13308 30104 13320
rect 30024 13280 30104 13308
rect 29917 13271 29975 13277
rect 30098 13268 30104 13280
rect 30156 13268 30162 13320
rect 30282 13268 30288 13320
rect 30340 13268 30346 13320
rect 30392 13240 30420 13484
rect 31113 13481 31125 13484
rect 31159 13481 31171 13515
rect 31113 13475 31171 13481
rect 33229 13515 33287 13521
rect 33229 13481 33241 13515
rect 33275 13512 33287 13515
rect 34054 13512 34060 13524
rect 33275 13484 34060 13512
rect 33275 13481 33287 13484
rect 33229 13475 33287 13481
rect 34054 13472 34060 13484
rect 34112 13472 34118 13524
rect 30650 13404 30656 13456
rect 30708 13444 30714 13456
rect 33321 13447 33379 13453
rect 30708 13416 32260 13444
rect 30708 13404 30714 13416
rect 30466 13336 30472 13388
rect 30524 13376 30530 13388
rect 30524 13348 30788 13376
rect 30524 13336 30530 13348
rect 30558 13268 30564 13320
rect 30616 13308 30622 13320
rect 30653 13311 30711 13317
rect 30653 13308 30665 13311
rect 30616 13280 30665 13308
rect 30616 13268 30622 13280
rect 30653 13277 30665 13280
rect 30699 13277 30711 13311
rect 30760 13308 30788 13348
rect 31297 13311 31355 13317
rect 31297 13308 31309 13311
rect 30760 13280 31309 13308
rect 30653 13271 30711 13277
rect 31297 13277 31309 13280
rect 31343 13277 31355 13311
rect 31297 13271 31355 13277
rect 31389 13311 31447 13317
rect 31389 13277 31401 13311
rect 31435 13277 31447 13311
rect 31389 13271 31447 13277
rect 29748 13212 30420 13240
rect 30742 13200 30748 13252
rect 30800 13240 30806 13252
rect 31404 13240 31432 13271
rect 31478 13268 31484 13320
rect 31536 13268 31542 13320
rect 31573 13311 31631 13317
rect 31573 13277 31585 13311
rect 31619 13277 31631 13311
rect 31573 13271 31631 13277
rect 31757 13311 31815 13317
rect 31757 13277 31769 13311
rect 31803 13308 31815 13311
rect 31938 13308 31944 13320
rect 31803 13280 31944 13308
rect 31803 13277 31815 13280
rect 31757 13271 31815 13277
rect 30800 13212 31432 13240
rect 30800 13200 30806 13212
rect 27154 13172 27160 13184
rect 26712 13144 27160 13172
rect 27154 13132 27160 13144
rect 27212 13132 27218 13184
rect 31110 13132 31116 13184
rect 31168 13172 31174 13184
rect 31588 13172 31616 13271
rect 31938 13268 31944 13280
rect 31996 13268 32002 13320
rect 32232 13317 32260 13416
rect 33321 13413 33333 13447
rect 33367 13413 33379 13447
rect 33321 13407 33379 13413
rect 32217 13311 32275 13317
rect 32217 13277 32229 13311
rect 32263 13277 32275 13311
rect 32217 13271 32275 13277
rect 33045 13311 33103 13317
rect 33045 13277 33057 13311
rect 33091 13308 33103 13311
rect 33336 13308 33364 13407
rect 33594 13336 33600 13388
rect 33652 13376 33658 13388
rect 33781 13379 33839 13385
rect 33781 13376 33793 13379
rect 33652 13348 33793 13376
rect 33652 13336 33658 13348
rect 33781 13345 33793 13348
rect 33827 13345 33839 13379
rect 33781 13339 33839 13345
rect 33870 13336 33876 13388
rect 33928 13336 33934 13388
rect 33091 13280 33364 13308
rect 33091 13277 33103 13280
rect 33045 13271 33103 13277
rect 33226 13200 33232 13252
rect 33284 13240 33290 13252
rect 33888 13240 33916 13336
rect 33284 13212 33916 13240
rect 33284 13200 33290 13212
rect 31168 13144 31616 13172
rect 31941 13175 31999 13181
rect 31168 13132 31174 13144
rect 31941 13141 31953 13175
rect 31987 13172 31999 13175
rect 32030 13172 32036 13184
rect 31987 13144 32036 13172
rect 31987 13141 31999 13144
rect 31941 13135 31999 13141
rect 32030 13132 32036 13144
rect 32088 13132 32094 13184
rect 32306 13132 32312 13184
rect 32364 13132 32370 13184
rect 33686 13132 33692 13184
rect 33744 13132 33750 13184
rect 1104 13082 38272 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 38272 13082
rect 1104 13008 38272 13030
rect 3878 12928 3884 12980
rect 3936 12928 3942 12980
rect 9674 12968 9680 12980
rect 8956 12940 9680 12968
rect 3896 12900 3924 12928
rect 3528 12872 3924 12900
rect 3528 12841 3556 12872
rect 5258 12860 5264 12912
rect 5316 12900 5322 12912
rect 5537 12903 5595 12909
rect 5537 12900 5549 12903
rect 5316 12872 5549 12900
rect 5316 12860 5322 12872
rect 5537 12869 5549 12872
rect 5583 12869 5595 12903
rect 5537 12863 5595 12869
rect 6178 12860 6184 12912
rect 6236 12860 6242 12912
rect 3513 12835 3571 12841
rect 3513 12801 3525 12835
rect 3559 12801 3571 12835
rect 6196 12832 6224 12860
rect 8956 12841 8984 12940
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 9766 12928 9772 12980
rect 9824 12928 9830 12980
rect 12526 12968 12532 12980
rect 12360 12940 12532 12968
rect 9125 12903 9183 12909
rect 9125 12869 9137 12903
rect 9171 12900 9183 12903
rect 9582 12900 9588 12912
rect 9171 12872 9588 12900
rect 9171 12869 9183 12872
rect 9125 12863 9183 12869
rect 9582 12860 9588 12872
rect 9640 12900 9646 12912
rect 12360 12909 12388 12940
rect 12526 12928 12532 12940
rect 12584 12928 12590 12980
rect 12713 12971 12771 12977
rect 12713 12937 12725 12971
rect 12759 12968 12771 12971
rect 13078 12968 13084 12980
rect 12759 12940 13084 12968
rect 12759 12937 12771 12940
rect 12713 12931 12771 12937
rect 13078 12928 13084 12940
rect 13136 12928 13142 12980
rect 13538 12968 13544 12980
rect 13183 12940 13544 12968
rect 12345 12903 12403 12909
rect 9640 12872 10364 12900
rect 9640 12860 9646 12872
rect 4922 12804 6224 12832
rect 8481 12835 8539 12841
rect 3513 12795 3571 12801
rect 8481 12801 8493 12835
rect 8527 12801 8539 12835
rect 8481 12795 8539 12801
rect 8665 12835 8723 12841
rect 8665 12801 8677 12835
rect 8711 12832 8723 12835
rect 8849 12835 8907 12841
rect 8849 12832 8861 12835
rect 8711 12804 8861 12832
rect 8711 12801 8723 12804
rect 8665 12795 8723 12801
rect 8849 12801 8861 12804
rect 8895 12801 8907 12835
rect 8849 12795 8907 12801
rect 8941 12835 8999 12841
rect 8941 12801 8953 12835
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12801 9091 12835
rect 9033 12795 9091 12801
rect 9217 12835 9275 12841
rect 9217 12801 9229 12835
rect 9263 12801 9275 12835
rect 9217 12795 9275 12801
rect 3789 12767 3847 12773
rect 3789 12733 3801 12767
rect 3835 12764 3847 12767
rect 4430 12764 4436 12776
rect 3835 12736 4436 12764
rect 3835 12733 3847 12736
rect 3789 12727 3847 12733
rect 4430 12724 4436 12736
rect 4488 12724 4494 12776
rect 8496 12628 8524 12795
rect 8864 12764 8892 12795
rect 9048 12764 9076 12795
rect 8864 12736 9076 12764
rect 9122 12724 9128 12776
rect 9180 12764 9186 12776
rect 9232 12764 9260 12795
rect 9490 12792 9496 12844
rect 9548 12792 9554 12844
rect 9858 12792 9864 12844
rect 9916 12792 9922 12844
rect 10042 12792 10048 12844
rect 10100 12792 10106 12844
rect 10137 12835 10195 12841
rect 10137 12801 10149 12835
rect 10183 12832 10195 12835
rect 10226 12832 10232 12844
rect 10183 12804 10232 12832
rect 10183 12801 10195 12804
rect 10137 12795 10195 12801
rect 10226 12792 10232 12804
rect 10284 12792 10290 12844
rect 10336 12841 10364 12872
rect 12345 12869 12357 12903
rect 12391 12869 12403 12903
rect 13183 12900 13211 12940
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 14642 12928 14648 12980
rect 14700 12968 14706 12980
rect 14737 12971 14795 12977
rect 14737 12968 14749 12971
rect 14700 12940 14749 12968
rect 14700 12928 14706 12940
rect 14737 12937 14749 12940
rect 14783 12937 14795 12971
rect 18322 12968 18328 12980
rect 14737 12931 14795 12937
rect 16592 12940 18328 12968
rect 12345 12863 12403 12869
rect 13004 12872 13211 12900
rect 13265 12903 13323 12909
rect 10321 12835 10379 12841
rect 10321 12801 10333 12835
rect 10367 12801 10379 12835
rect 10321 12795 10379 12801
rect 10594 12792 10600 12844
rect 10652 12832 10658 12844
rect 10781 12835 10839 12841
rect 10781 12832 10793 12835
rect 10652 12804 10793 12832
rect 10652 12792 10658 12804
rect 10781 12801 10793 12804
rect 10827 12801 10839 12835
rect 11974 12832 11980 12844
rect 10781 12795 10839 12801
rect 10888 12804 11980 12832
rect 9180 12736 9260 12764
rect 9309 12767 9367 12773
rect 9180 12724 9186 12736
rect 9309 12733 9321 12767
rect 9355 12733 9367 12767
rect 10060 12764 10088 12792
rect 10888 12764 10916 12804
rect 11974 12792 11980 12804
rect 12032 12832 12038 12844
rect 12161 12835 12219 12841
rect 12161 12832 12173 12835
rect 12032 12804 12173 12832
rect 12032 12792 12038 12804
rect 12161 12801 12173 12804
rect 12207 12801 12219 12835
rect 12161 12795 12219 12801
rect 12437 12835 12495 12841
rect 12437 12801 12449 12835
rect 12483 12801 12495 12835
rect 12437 12795 12495 12801
rect 12529 12835 12587 12841
rect 12529 12801 12541 12835
rect 12575 12832 12587 12835
rect 12618 12832 12624 12844
rect 12575 12804 12624 12832
rect 12575 12801 12587 12804
rect 12529 12795 12587 12801
rect 10060 12736 10916 12764
rect 9309 12727 9367 12733
rect 8573 12699 8631 12705
rect 8573 12665 8585 12699
rect 8619 12696 8631 12699
rect 9030 12696 9036 12708
rect 8619 12668 9036 12696
rect 8619 12665 8631 12668
rect 8573 12659 8631 12665
rect 9030 12656 9036 12668
rect 9088 12696 9094 12708
rect 9324 12696 9352 12727
rect 10962 12724 10968 12776
rect 11020 12724 11026 12776
rect 12452 12764 12480 12795
rect 12618 12792 12624 12804
rect 12676 12832 12682 12844
rect 12802 12832 12808 12844
rect 12676 12804 12808 12832
rect 12676 12792 12682 12804
rect 12802 12792 12808 12804
rect 12860 12792 12866 12844
rect 13004 12841 13032 12872
rect 13265 12869 13277 12903
rect 13311 12900 13323 12903
rect 13354 12900 13360 12912
rect 13311 12872 13360 12900
rect 13311 12869 13323 12872
rect 13265 12863 13323 12869
rect 13354 12860 13360 12872
rect 13412 12860 13418 12912
rect 16206 12860 16212 12912
rect 16264 12860 16270 12912
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 14274 12792 14280 12844
rect 14332 12832 14338 12844
rect 16224 12832 16252 12860
rect 14332 12804 16252 12832
rect 14332 12792 14338 12804
rect 16592 12764 16620 12940
rect 18322 12928 18328 12940
rect 18380 12928 18386 12980
rect 19426 12968 19432 12980
rect 19352 12940 19432 12968
rect 19352 12841 19380 12940
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 19521 12971 19579 12977
rect 19521 12937 19533 12971
rect 19567 12968 19579 12971
rect 19567 12940 19748 12968
rect 19567 12937 19579 12940
rect 19521 12931 19579 12937
rect 19720 12900 19748 12940
rect 21358 12928 21364 12980
rect 21416 12928 21422 12980
rect 24302 12928 24308 12980
rect 24360 12968 24366 12980
rect 24360 12940 25268 12968
rect 24360 12928 24366 12940
rect 19889 12903 19947 12909
rect 19889 12900 19901 12903
rect 19720 12872 19901 12900
rect 19889 12869 19901 12872
rect 19935 12869 19947 12903
rect 23198 12900 23204 12912
rect 21114 12872 23204 12900
rect 19889 12863 19947 12869
rect 23198 12860 23204 12872
rect 23256 12860 23262 12912
rect 24857 12903 24915 12909
rect 24857 12900 24869 12903
rect 24320 12872 24869 12900
rect 19337 12835 19395 12841
rect 19337 12801 19349 12835
rect 19383 12801 19395 12835
rect 19337 12795 19395 12801
rect 22278 12792 22284 12844
rect 22336 12792 22342 12844
rect 24320 12776 24348 12872
rect 24857 12869 24869 12872
rect 24903 12869 24915 12903
rect 24857 12863 24915 12869
rect 24581 12835 24639 12841
rect 24581 12801 24593 12835
rect 24627 12801 24639 12835
rect 24581 12795 24639 12801
rect 12406 12736 16620 12764
rect 9088 12668 9352 12696
rect 9088 12656 9094 12668
rect 9766 12656 9772 12708
rect 9824 12696 9830 12708
rect 12406 12696 12434 12736
rect 18230 12724 18236 12776
rect 18288 12764 18294 12776
rect 18782 12764 18788 12776
rect 18288 12736 18788 12764
rect 18288 12724 18294 12736
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 19610 12724 19616 12776
rect 19668 12724 19674 12776
rect 24302 12724 24308 12776
rect 24360 12724 24366 12776
rect 19518 12696 19524 12708
rect 9824 12668 12434 12696
rect 16224 12668 19524 12696
rect 9824 12656 9830 12668
rect 9122 12628 9128 12640
rect 8496 12600 9128 12628
rect 9122 12588 9128 12600
rect 9180 12588 9186 12640
rect 14366 12588 14372 12640
rect 14424 12628 14430 12640
rect 15102 12628 15108 12640
rect 14424 12600 15108 12628
rect 14424 12588 14430 12600
rect 15102 12588 15108 12600
rect 15160 12628 15166 12640
rect 16224 12628 16252 12668
rect 19518 12656 19524 12668
rect 19576 12656 19582 12708
rect 24596 12696 24624 12795
rect 24670 12792 24676 12844
rect 24728 12832 24734 12844
rect 24949 12835 25007 12841
rect 24728 12804 24773 12832
rect 24728 12792 24734 12804
rect 24949 12801 24961 12835
rect 24995 12801 25007 12835
rect 24949 12795 25007 12801
rect 24964 12764 24992 12795
rect 25038 12792 25044 12844
rect 25096 12841 25102 12844
rect 25096 12832 25104 12841
rect 25096 12804 25141 12832
rect 25096 12795 25104 12804
rect 25096 12792 25102 12795
rect 25240 12764 25268 12940
rect 25314 12928 25320 12980
rect 25372 12928 25378 12980
rect 25406 12928 25412 12980
rect 25464 12968 25470 12980
rect 25464 12940 26648 12968
rect 25464 12928 25470 12940
rect 25332 12841 25360 12928
rect 26510 12860 26516 12912
rect 26568 12860 26574 12912
rect 26620 12900 26648 12940
rect 26970 12928 26976 12980
rect 27028 12968 27034 12980
rect 27028 12940 27752 12968
rect 27028 12928 27034 12940
rect 27724 12900 27752 12940
rect 27890 12928 27896 12980
rect 27948 12928 27954 12980
rect 28353 12971 28411 12977
rect 28353 12937 28365 12971
rect 28399 12968 28411 12971
rect 28718 12968 28724 12980
rect 28399 12940 28724 12968
rect 28399 12937 28411 12940
rect 28353 12931 28411 12937
rect 28718 12928 28724 12940
rect 28776 12928 28782 12980
rect 28902 12928 28908 12980
rect 28960 12968 28966 12980
rect 29917 12971 29975 12977
rect 28960 12940 29776 12968
rect 28960 12928 28966 12940
rect 27985 12903 28043 12909
rect 26620 12872 27384 12900
rect 27724 12872 27936 12900
rect 25317 12835 25375 12841
rect 25317 12801 25329 12835
rect 25363 12801 25375 12835
rect 25317 12795 25375 12801
rect 25593 12835 25651 12841
rect 25593 12801 25605 12835
rect 25639 12832 25651 12835
rect 25639 12804 25912 12832
rect 25639 12801 25651 12804
rect 25593 12795 25651 12801
rect 25501 12767 25559 12773
rect 25501 12764 25513 12767
rect 24964 12736 25176 12764
rect 25240 12736 25513 12764
rect 25038 12696 25044 12708
rect 24596 12668 25044 12696
rect 25038 12656 25044 12668
rect 25096 12656 25102 12708
rect 15160 12600 16252 12628
rect 15160 12588 15166 12600
rect 16850 12588 16856 12640
rect 16908 12628 16914 12640
rect 22186 12628 22192 12640
rect 16908 12600 22192 12628
rect 16908 12588 16914 12600
rect 22186 12588 22192 12600
rect 22244 12588 22250 12640
rect 23382 12588 23388 12640
rect 23440 12628 23446 12640
rect 23569 12631 23627 12637
rect 23569 12628 23581 12631
rect 23440 12600 23581 12628
rect 23440 12588 23446 12600
rect 23569 12597 23581 12600
rect 23615 12597 23627 12631
rect 25148 12628 25176 12736
rect 25501 12733 25513 12736
rect 25547 12733 25559 12767
rect 25501 12727 25559 12733
rect 25685 12767 25743 12773
rect 25685 12733 25697 12767
rect 25731 12733 25743 12767
rect 25685 12727 25743 12733
rect 25225 12699 25283 12705
rect 25225 12665 25237 12699
rect 25271 12696 25283 12699
rect 25700 12696 25728 12727
rect 25774 12724 25780 12776
rect 25832 12724 25838 12776
rect 25271 12668 25728 12696
rect 25884 12696 25912 12804
rect 26050 12792 26056 12844
rect 26108 12832 26114 12844
rect 26620 12841 26648 12872
rect 26283 12835 26341 12841
rect 26283 12832 26295 12835
rect 26108 12804 26295 12832
rect 26108 12792 26114 12804
rect 26283 12801 26295 12804
rect 26329 12801 26341 12835
rect 26283 12795 26341 12801
rect 26421 12835 26479 12841
rect 26421 12801 26433 12835
rect 26467 12832 26479 12835
rect 26620 12835 26699 12841
rect 26467 12804 26556 12832
rect 26620 12804 26653 12835
rect 26467 12801 26479 12804
rect 26421 12795 26479 12801
rect 25961 12767 26019 12773
rect 25961 12733 25973 12767
rect 26007 12764 26019 12767
rect 26528 12764 26556 12804
rect 26641 12801 26653 12804
rect 26687 12801 26699 12835
rect 26641 12795 26699 12801
rect 26786 12792 26792 12844
rect 26844 12832 26850 12844
rect 26970 12832 26976 12844
rect 26844 12804 26976 12832
rect 26844 12792 26850 12804
rect 26970 12792 26976 12804
rect 27028 12792 27034 12844
rect 27246 12792 27252 12844
rect 27304 12792 27310 12844
rect 27356 12841 27384 12872
rect 27798 12841 27804 12844
rect 27342 12835 27400 12841
rect 27342 12801 27354 12835
rect 27388 12801 27400 12835
rect 27342 12795 27400 12801
rect 27525 12835 27583 12841
rect 27525 12801 27537 12835
rect 27571 12801 27583 12835
rect 27525 12795 27583 12801
rect 27617 12835 27675 12841
rect 27617 12801 27629 12835
rect 27663 12801 27675 12835
rect 27617 12795 27675 12801
rect 27755 12835 27804 12841
rect 27755 12801 27767 12835
rect 27801 12801 27804 12835
rect 27755 12795 27804 12801
rect 27540 12764 27568 12795
rect 26007 12736 26280 12764
rect 26528 12736 26648 12764
rect 26007 12733 26019 12736
rect 25961 12727 26019 12733
rect 26252 12708 26280 12736
rect 26620 12708 26648 12736
rect 26804 12736 27568 12764
rect 26804 12708 26832 12736
rect 26145 12699 26203 12705
rect 26145 12696 26157 12699
rect 25884 12668 26157 12696
rect 25271 12665 25283 12668
rect 25225 12659 25283 12665
rect 26145 12665 26157 12668
rect 26191 12665 26203 12699
rect 26145 12659 26203 12665
rect 26234 12656 26240 12708
rect 26292 12656 26298 12708
rect 26602 12656 26608 12708
rect 26660 12656 26666 12708
rect 26786 12656 26792 12708
rect 26844 12656 26850 12708
rect 26878 12656 26884 12708
rect 26936 12696 26942 12708
rect 27338 12696 27344 12708
rect 26936 12668 27344 12696
rect 26936 12656 26942 12668
rect 27338 12656 27344 12668
rect 27396 12656 27402 12708
rect 27632 12696 27660 12795
rect 27798 12792 27804 12795
rect 27856 12792 27862 12844
rect 27908 12832 27936 12872
rect 27985 12869 27997 12903
rect 28031 12900 28043 12903
rect 28534 12900 28540 12912
rect 28031 12872 28540 12900
rect 28031 12869 28043 12872
rect 27985 12863 28043 12869
rect 28534 12860 28540 12872
rect 28592 12860 28598 12912
rect 28994 12860 29000 12912
rect 29052 12900 29058 12912
rect 29052 12872 29592 12900
rect 29052 12860 29058 12872
rect 28169 12835 28227 12841
rect 28169 12832 28181 12835
rect 27908 12804 28181 12832
rect 28169 12801 28181 12804
rect 28215 12832 28227 12835
rect 28215 12804 28994 12832
rect 28215 12801 28227 12804
rect 28169 12795 28227 12801
rect 28966 12764 28994 12804
rect 29362 12792 29368 12844
rect 29420 12792 29426 12844
rect 29564 12841 29592 12872
rect 29748 12841 29776 12940
rect 29917 12937 29929 12971
rect 29963 12968 29975 12971
rect 30282 12968 30288 12980
rect 29963 12940 30288 12968
rect 29963 12937 29975 12940
rect 29917 12931 29975 12937
rect 30282 12928 30288 12940
rect 30340 12928 30346 12980
rect 31938 12928 31944 12980
rect 31996 12928 32002 12980
rect 32030 12928 32036 12980
rect 32088 12928 32094 12980
rect 32306 12928 32312 12980
rect 32364 12928 32370 12980
rect 31478 12860 31484 12912
rect 31536 12860 31542 12912
rect 29457 12835 29515 12841
rect 29457 12801 29469 12835
rect 29503 12801 29515 12835
rect 29564 12835 29626 12841
rect 29564 12804 29580 12835
rect 29457 12795 29515 12801
rect 29568 12801 29580 12804
rect 29614 12801 29626 12835
rect 29568 12795 29626 12801
rect 29733 12835 29791 12841
rect 29733 12801 29745 12835
rect 29779 12801 29791 12835
rect 29733 12795 29791 12801
rect 29472 12764 29500 12795
rect 30098 12792 30104 12844
rect 30156 12792 30162 12844
rect 31496 12832 31524 12860
rect 31573 12835 31631 12841
rect 31573 12832 31585 12835
rect 31404 12804 31585 12832
rect 30116 12764 30144 12792
rect 28966 12736 29408 12764
rect 29472 12736 30144 12764
rect 28994 12696 29000 12708
rect 27632 12668 29000 12696
rect 25590 12628 25596 12640
rect 25148 12600 25596 12628
rect 23569 12591 23627 12597
rect 25590 12588 25596 12600
rect 25648 12588 25654 12640
rect 25682 12588 25688 12640
rect 25740 12628 25746 12640
rect 27632 12628 27660 12668
rect 28994 12656 29000 12668
rect 29052 12656 29058 12708
rect 29380 12696 29408 12736
rect 31294 12724 31300 12776
rect 31352 12724 31358 12776
rect 31404 12696 31432 12804
rect 31573 12801 31585 12804
rect 31619 12801 31631 12835
rect 31573 12795 31631 12801
rect 31481 12767 31539 12773
rect 31481 12733 31493 12767
rect 31527 12733 31539 12767
rect 31481 12727 31539 12733
rect 29380 12668 31432 12696
rect 25740 12600 27660 12628
rect 25740 12588 25746 12600
rect 27890 12588 27896 12640
rect 27948 12628 27954 12640
rect 28534 12628 28540 12640
rect 27948 12600 28540 12628
rect 27948 12588 27954 12600
rect 28534 12588 28540 12600
rect 28592 12588 28598 12640
rect 30282 12588 30288 12640
rect 30340 12628 30346 12640
rect 31386 12628 31392 12640
rect 30340 12600 31392 12628
rect 30340 12588 30346 12600
rect 31386 12588 31392 12600
rect 31444 12628 31450 12640
rect 31496 12628 31524 12727
rect 31444 12600 31524 12628
rect 31588 12628 31616 12795
rect 32048 12764 32076 12928
rect 32324 12900 32352 12928
rect 32140 12872 32352 12900
rect 32140 12841 32168 12872
rect 32125 12835 32183 12841
rect 32125 12801 32137 12835
rect 32171 12801 32183 12835
rect 33962 12832 33968 12844
rect 33534 12804 33968 12832
rect 32125 12795 32183 12801
rect 33962 12792 33968 12804
rect 34020 12792 34026 12844
rect 32401 12767 32459 12773
rect 32401 12764 32413 12767
rect 32048 12736 32413 12764
rect 32401 12733 32413 12736
rect 32447 12733 32459 12767
rect 32401 12727 32459 12733
rect 33873 12631 33931 12637
rect 33873 12628 33885 12631
rect 31588 12600 33885 12628
rect 31444 12588 31450 12600
rect 33873 12597 33885 12600
rect 33919 12597 33931 12631
rect 33873 12591 33931 12597
rect 1104 12538 38272 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38272 12538
rect 1104 12464 38272 12486
rect 4157 12427 4215 12433
rect 4157 12393 4169 12427
rect 4203 12424 4215 12427
rect 4614 12424 4620 12436
rect 4203 12396 4620 12424
rect 4203 12393 4215 12396
rect 4157 12387 4215 12393
rect 4614 12384 4620 12396
rect 4672 12384 4678 12436
rect 9122 12384 9128 12436
rect 9180 12424 9186 12436
rect 9180 12396 11376 12424
rect 9180 12384 9186 12396
rect 10042 12356 10048 12368
rect 9646 12328 10048 12356
rect 4798 12248 4804 12300
rect 4856 12288 4862 12300
rect 4856 12260 6500 12288
rect 4856 12248 4862 12260
rect 4341 12223 4399 12229
rect 4341 12189 4353 12223
rect 4387 12220 4399 12223
rect 4706 12220 4712 12232
rect 4387 12192 4712 12220
rect 4387 12189 4399 12192
rect 4341 12183 4399 12189
rect 4706 12180 4712 12192
rect 4764 12180 4770 12232
rect 4908 12229 4936 12260
rect 6472 12232 6500 12260
rect 9122 12248 9128 12300
rect 9180 12288 9186 12300
rect 9646 12288 9674 12328
rect 10042 12316 10048 12328
rect 10100 12316 10106 12368
rect 10686 12316 10692 12368
rect 10744 12356 10750 12368
rect 10962 12356 10968 12368
rect 10744 12328 10968 12356
rect 10744 12316 10750 12328
rect 10962 12316 10968 12328
rect 11020 12316 11026 12368
rect 9180 12260 9674 12288
rect 9876 12260 11008 12288
rect 9180 12248 9186 12260
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12189 4951 12223
rect 4893 12183 4951 12189
rect 4985 12223 5043 12229
rect 4985 12189 4997 12223
rect 5031 12220 5043 12223
rect 5169 12223 5227 12229
rect 5169 12220 5181 12223
rect 5031 12192 5181 12220
rect 5031 12189 5043 12192
rect 4985 12183 5043 12189
rect 5169 12189 5181 12192
rect 5215 12189 5227 12223
rect 5169 12183 5227 12189
rect 6454 12180 6460 12232
rect 6512 12180 6518 12232
rect 9876 12229 9904 12260
rect 10980 12232 11008 12260
rect 9861 12223 9919 12229
rect 9861 12189 9873 12223
rect 9907 12189 9919 12223
rect 9861 12183 9919 12189
rect 9950 12180 9956 12232
rect 10008 12220 10014 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 10008 12192 10149 12220
rect 10008 12180 10014 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10778 12180 10784 12232
rect 10836 12180 10842 12232
rect 10873 12223 10931 12229
rect 10873 12189 10885 12223
rect 10919 12189 10931 12223
rect 10873 12183 10931 12189
rect 5442 12112 5448 12164
rect 5500 12112 5506 12164
rect 6178 12112 6184 12164
rect 6236 12112 6242 12164
rect 6822 12112 6828 12164
rect 6880 12152 6886 12164
rect 7193 12155 7251 12161
rect 7193 12152 7205 12155
rect 6880 12124 7205 12152
rect 6880 12112 6886 12124
rect 7193 12121 7205 12124
rect 7239 12152 7251 12155
rect 7239 12124 9628 12152
rect 7239 12121 7251 12124
rect 7193 12115 7251 12121
rect 9600 12084 9628 12124
rect 9674 12112 9680 12164
rect 9732 12152 9738 12164
rect 10888 12152 10916 12183
rect 10962 12180 10968 12232
rect 11020 12220 11026 12232
rect 11348 12229 11376 12396
rect 15378 12384 15384 12436
rect 15436 12384 15442 12436
rect 15654 12384 15660 12436
rect 15712 12424 15718 12436
rect 15838 12424 15844 12436
rect 15712 12396 15844 12424
rect 15712 12384 15718 12396
rect 15838 12384 15844 12396
rect 15896 12384 15902 12436
rect 15930 12384 15936 12436
rect 15988 12424 15994 12436
rect 16298 12424 16304 12436
rect 15988 12396 16304 12424
rect 15988 12384 15994 12396
rect 16298 12384 16304 12396
rect 16356 12384 16362 12436
rect 16390 12384 16396 12436
rect 16448 12424 16454 12436
rect 16577 12427 16635 12433
rect 16577 12424 16589 12427
rect 16448 12396 16589 12424
rect 16448 12384 16454 12396
rect 16577 12393 16589 12396
rect 16623 12393 16635 12427
rect 16577 12387 16635 12393
rect 16850 12384 16856 12436
rect 16908 12384 16914 12436
rect 21174 12424 21180 12436
rect 17328 12396 21180 12424
rect 15396 12288 15424 12384
rect 15212 12260 15424 12288
rect 15488 12328 16712 12356
rect 11241 12223 11299 12229
rect 11241 12220 11253 12223
rect 11020 12192 11253 12220
rect 11020 12180 11026 12192
rect 11241 12189 11253 12192
rect 11287 12189 11299 12223
rect 11241 12183 11299 12189
rect 11333 12223 11391 12229
rect 11333 12189 11345 12223
rect 11379 12189 11391 12223
rect 11333 12183 11391 12189
rect 11974 12180 11980 12232
rect 12032 12220 12038 12232
rect 15212 12229 15240 12260
rect 15488 12229 15516 12328
rect 15841 12291 15899 12297
rect 15841 12257 15853 12291
rect 15887 12288 15899 12291
rect 15887 12260 16068 12288
rect 15887 12257 15899 12260
rect 15841 12251 15899 12257
rect 12529 12223 12587 12229
rect 12529 12220 12541 12223
rect 12032 12192 12541 12220
rect 12032 12180 12038 12192
rect 12529 12189 12541 12192
rect 12575 12189 12587 12223
rect 12529 12183 12587 12189
rect 15197 12223 15255 12229
rect 15197 12189 15209 12223
rect 15243 12189 15255 12223
rect 15197 12183 15255 12189
rect 15381 12223 15439 12229
rect 15381 12189 15393 12223
rect 15427 12189 15439 12223
rect 15381 12183 15439 12189
rect 15473 12223 15531 12229
rect 15473 12189 15485 12223
rect 15519 12189 15531 12223
rect 15473 12183 15531 12189
rect 15565 12223 15623 12229
rect 15565 12189 15577 12223
rect 15611 12220 15623 12223
rect 15654 12220 15660 12232
rect 15611 12192 15660 12220
rect 15611 12189 15623 12192
rect 15565 12183 15623 12189
rect 12986 12152 12992 12164
rect 9732 12124 10916 12152
rect 12360 12124 12992 12152
rect 9732 12112 9738 12124
rect 12360 12084 12388 12124
rect 12986 12112 12992 12124
rect 13044 12112 13050 12164
rect 15102 12112 15108 12164
rect 15160 12152 15166 12164
rect 15396 12152 15424 12183
rect 15160 12124 15424 12152
rect 15488 12152 15516 12183
rect 15654 12180 15660 12192
rect 15712 12180 15718 12232
rect 16040 12229 16068 12260
rect 16114 12248 16120 12300
rect 16172 12288 16178 12300
rect 16684 12288 16712 12328
rect 17328 12300 17356 12396
rect 21174 12384 21180 12396
rect 21232 12384 21238 12436
rect 22097 12427 22155 12433
rect 22097 12393 22109 12427
rect 22143 12393 22155 12427
rect 22097 12387 22155 12393
rect 24320 12396 25820 12424
rect 17586 12316 17592 12368
rect 17644 12316 17650 12368
rect 18046 12316 18052 12368
rect 18104 12316 18110 12368
rect 19518 12316 19524 12368
rect 19576 12356 19582 12368
rect 22112 12356 22140 12387
rect 19576 12328 22140 12356
rect 19576 12316 19582 12328
rect 16172 12260 16344 12288
rect 16684 12260 17080 12288
rect 16172 12248 16178 12260
rect 16316 12229 16344 12260
rect 15933 12223 15991 12229
rect 15933 12220 15945 12223
rect 15856 12192 15945 12220
rect 15856 12164 15884 12192
rect 15933 12189 15945 12192
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 16025 12223 16083 12229
rect 16025 12189 16037 12223
rect 16071 12189 16083 12223
rect 16025 12183 16083 12189
rect 16301 12223 16359 12229
rect 16301 12189 16313 12223
rect 16347 12189 16359 12223
rect 16301 12183 16359 12189
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12220 16451 12223
rect 16482 12220 16488 12232
rect 16439 12192 16488 12220
rect 16439 12189 16451 12192
rect 16393 12183 16451 12189
rect 16482 12180 16488 12192
rect 16540 12180 16546 12232
rect 16942 12180 16948 12232
rect 17000 12180 17006 12232
rect 17052 12229 17080 12260
rect 17310 12248 17316 12300
rect 17368 12248 17374 12300
rect 17037 12223 17095 12229
rect 17037 12189 17049 12223
rect 17083 12189 17095 12223
rect 17037 12183 17095 12189
rect 17218 12180 17224 12232
rect 17276 12220 17282 12232
rect 17604 12220 17632 12316
rect 18598 12288 18604 12300
rect 18432 12260 18604 12288
rect 18432 12229 18460 12260
rect 18598 12248 18604 12260
rect 18656 12288 18662 12300
rect 18656 12260 18828 12288
rect 18656 12248 18662 12260
rect 18800 12232 18828 12260
rect 19702 12248 19708 12300
rect 19760 12288 19766 12300
rect 20806 12288 20812 12300
rect 19760 12260 20812 12288
rect 19760 12248 19766 12260
rect 20806 12248 20812 12260
rect 20864 12248 20870 12300
rect 22112 12288 22140 12328
rect 22922 12316 22928 12368
rect 22980 12356 22986 12368
rect 23569 12359 23627 12365
rect 23569 12356 23581 12359
rect 22980 12328 23581 12356
rect 22980 12316 22986 12328
rect 23569 12325 23581 12328
rect 23615 12356 23627 12359
rect 23934 12356 23940 12368
rect 23615 12328 23940 12356
rect 23615 12325 23627 12328
rect 23569 12319 23627 12325
rect 23934 12316 23940 12328
rect 23992 12316 23998 12368
rect 24320 12300 24348 12396
rect 24670 12316 24676 12368
rect 24728 12316 24734 12368
rect 24949 12359 25007 12365
rect 24949 12325 24961 12359
rect 24995 12325 25007 12359
rect 24949 12319 25007 12325
rect 24302 12288 24308 12300
rect 22112 12260 24308 12288
rect 22572 12232 22600 12260
rect 24302 12248 24308 12260
rect 24360 12248 24366 12300
rect 24688 12288 24716 12316
rect 24412 12260 24716 12288
rect 24964 12288 24992 12319
rect 25038 12316 25044 12368
rect 25096 12316 25102 12368
rect 25593 12359 25651 12365
rect 25593 12325 25605 12359
rect 25639 12356 25651 12359
rect 25682 12356 25688 12368
rect 25639 12328 25688 12356
rect 25639 12325 25651 12328
rect 25593 12319 25651 12325
rect 25682 12316 25688 12328
rect 25740 12316 25746 12368
rect 24964 12260 25729 12288
rect 17276 12192 17632 12220
rect 18324 12223 18382 12229
rect 17276 12180 17282 12192
rect 18324 12189 18336 12223
rect 18370 12189 18382 12223
rect 18324 12183 18382 12189
rect 18417 12223 18475 12229
rect 18417 12189 18429 12223
rect 18463 12189 18475 12223
rect 18417 12183 18475 12189
rect 18509 12223 18567 12229
rect 18509 12189 18521 12223
rect 18555 12189 18567 12223
rect 18509 12183 18567 12189
rect 15488 12124 15608 12152
rect 15160 12112 15166 12124
rect 15580 12096 15608 12124
rect 15838 12112 15844 12164
rect 15896 12112 15902 12164
rect 16209 12155 16267 12161
rect 16209 12121 16221 12155
rect 16255 12152 16267 12155
rect 16960 12152 16988 12180
rect 18339 12152 18367 12183
rect 16255 12124 16896 12152
rect 16960 12124 18367 12152
rect 18524 12152 18552 12183
rect 18690 12180 18696 12232
rect 18748 12180 18754 12232
rect 18782 12180 18788 12232
rect 18840 12220 18846 12232
rect 18840 12192 20944 12220
rect 18840 12180 18846 12192
rect 20916 12164 20944 12192
rect 21266 12180 21272 12232
rect 21324 12220 21330 12232
rect 22370 12220 22376 12232
rect 21324 12192 22376 12220
rect 21324 12180 21330 12192
rect 22370 12180 22376 12192
rect 22428 12180 22434 12232
rect 22554 12180 22560 12232
rect 22612 12180 22618 12232
rect 23661 12223 23719 12229
rect 23661 12189 23673 12223
rect 23707 12220 23719 12223
rect 24118 12220 24124 12232
rect 23707 12192 24124 12220
rect 23707 12189 23719 12192
rect 23661 12183 23719 12189
rect 20714 12152 20720 12164
rect 18524 12124 20720 12152
rect 16255 12121 16267 12124
rect 16209 12115 16267 12121
rect 9600 12056 12388 12084
rect 12434 12044 12440 12096
rect 12492 12044 12498 12096
rect 13354 12044 13360 12096
rect 13412 12084 13418 12096
rect 15010 12084 15016 12096
rect 13412 12056 15016 12084
rect 13412 12044 13418 12056
rect 15010 12044 15016 12056
rect 15068 12044 15074 12096
rect 15562 12044 15568 12096
rect 15620 12044 15626 12096
rect 16482 12044 16488 12096
rect 16540 12084 16546 12096
rect 16669 12087 16727 12093
rect 16669 12084 16681 12087
rect 16540 12056 16681 12084
rect 16540 12044 16546 12056
rect 16669 12053 16681 12056
rect 16715 12053 16727 12087
rect 16868 12084 16896 12124
rect 20714 12112 20720 12124
rect 20772 12112 20778 12164
rect 20898 12112 20904 12164
rect 20956 12112 20962 12164
rect 21174 12112 21180 12164
rect 21232 12152 21238 12164
rect 21913 12155 21971 12161
rect 21913 12152 21925 12155
rect 21232 12124 21925 12152
rect 21232 12112 21238 12124
rect 21913 12121 21925 12124
rect 21959 12121 21971 12155
rect 21913 12115 21971 12121
rect 22186 12112 22192 12164
rect 22244 12152 22250 12164
rect 23676 12152 23704 12183
rect 24118 12180 24124 12192
rect 24176 12180 24182 12232
rect 24412 12229 24440 12260
rect 24397 12223 24455 12229
rect 24397 12189 24409 12223
rect 24443 12189 24455 12223
rect 24397 12183 24455 12189
rect 24486 12180 24492 12232
rect 24544 12220 24550 12232
rect 24673 12223 24731 12229
rect 24673 12220 24685 12223
rect 24544 12192 24685 12220
rect 24544 12180 24550 12192
rect 24673 12189 24685 12192
rect 24719 12189 24731 12223
rect 24673 12183 24731 12189
rect 24765 12223 24823 12229
rect 24765 12189 24777 12223
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 22244 12124 23704 12152
rect 22244 12112 22250 12124
rect 23934 12112 23940 12164
rect 23992 12152 23998 12164
rect 24578 12152 24584 12164
rect 23992 12124 24584 12152
rect 23992 12112 23998 12124
rect 24578 12112 24584 12124
rect 24636 12112 24642 12164
rect 24780 12152 24808 12183
rect 24854 12180 24860 12232
rect 24912 12220 24918 12232
rect 24912 12192 25544 12220
rect 24912 12180 24918 12192
rect 25406 12152 25412 12164
rect 24688 12124 24808 12152
rect 24872 12124 25412 12152
rect 24688 12096 24716 12124
rect 24872 12096 24900 12124
rect 25406 12112 25412 12124
rect 25464 12112 25470 12164
rect 25516 12096 25544 12192
rect 25701 12152 25729 12260
rect 25792 12220 25820 12396
rect 25866 12384 25872 12436
rect 25924 12424 25930 12436
rect 26694 12424 26700 12436
rect 25924 12396 26700 12424
rect 25924 12384 25930 12396
rect 26694 12384 26700 12396
rect 26752 12384 26758 12436
rect 27065 12427 27123 12433
rect 27065 12393 27077 12427
rect 27111 12424 27123 12427
rect 27246 12424 27252 12436
rect 27111 12396 27252 12424
rect 27111 12393 27123 12396
rect 27065 12387 27123 12393
rect 27246 12384 27252 12396
rect 27304 12384 27310 12436
rect 29638 12384 29644 12436
rect 29696 12424 29702 12436
rect 31294 12424 31300 12436
rect 29696 12396 31300 12424
rect 29696 12384 29702 12396
rect 31294 12384 31300 12396
rect 31352 12424 31358 12436
rect 31757 12427 31815 12433
rect 31757 12424 31769 12427
rect 31352 12396 31769 12424
rect 31352 12384 31358 12396
rect 31757 12393 31769 12396
rect 31803 12393 31815 12427
rect 31757 12387 31815 12393
rect 26602 12316 26608 12368
rect 26660 12356 26666 12368
rect 27617 12359 27675 12365
rect 27617 12356 27629 12359
rect 26660 12328 27629 12356
rect 26660 12316 26666 12328
rect 27617 12325 27629 12328
rect 27663 12356 27675 12359
rect 27982 12356 27988 12368
rect 27663 12328 27988 12356
rect 27663 12325 27675 12328
rect 27617 12319 27675 12325
rect 27982 12316 27988 12328
rect 28040 12316 28046 12368
rect 31386 12316 31392 12368
rect 31444 12356 31450 12368
rect 33686 12356 33692 12368
rect 31444 12328 33692 12356
rect 31444 12316 31450 12328
rect 29270 12248 29276 12300
rect 29328 12288 29334 12300
rect 29638 12288 29644 12300
rect 29328 12260 29644 12288
rect 29328 12248 29334 12260
rect 29638 12248 29644 12260
rect 29696 12248 29702 12300
rect 30834 12288 30840 12300
rect 29748 12260 30840 12288
rect 27338 12220 27344 12232
rect 25792 12192 27344 12220
rect 27338 12180 27344 12192
rect 27396 12180 27402 12232
rect 29748 12229 29776 12260
rect 30834 12248 30840 12260
rect 30892 12248 30898 12300
rect 33410 12248 33416 12300
rect 33468 12248 33474 12300
rect 33520 12297 33548 12328
rect 33686 12316 33692 12328
rect 33744 12316 33750 12368
rect 33505 12291 33563 12297
rect 33505 12257 33517 12291
rect 33551 12257 33563 12291
rect 33505 12251 33563 12257
rect 27433 12223 27491 12229
rect 27433 12189 27445 12223
rect 27479 12220 27491 12223
rect 29733 12223 29791 12229
rect 27479 12192 27936 12220
rect 27479 12189 27491 12192
rect 27433 12183 27491 12189
rect 27908 12164 27936 12192
rect 29733 12189 29745 12223
rect 29779 12189 29791 12223
rect 29733 12183 29791 12189
rect 29825 12223 29883 12229
rect 29825 12189 29837 12223
rect 29871 12220 29883 12223
rect 30009 12223 30067 12229
rect 30009 12220 30021 12223
rect 29871 12192 30021 12220
rect 29871 12189 29883 12192
rect 29825 12183 29883 12189
rect 30009 12189 30021 12192
rect 30055 12189 30067 12223
rect 34057 12223 34115 12229
rect 34057 12220 34069 12223
rect 30009 12183 30067 12189
rect 31680 12192 34069 12220
rect 31680 12164 31708 12192
rect 34057 12189 34069 12192
rect 34103 12189 34115 12223
rect 34057 12183 34115 12189
rect 34333 12223 34391 12229
rect 34333 12189 34345 12223
rect 34379 12189 34391 12223
rect 34333 12183 34391 12189
rect 26878 12152 26884 12164
rect 25701 12124 26884 12152
rect 26878 12112 26884 12124
rect 26936 12112 26942 12164
rect 27062 12112 27068 12164
rect 27120 12152 27126 12164
rect 27249 12155 27307 12161
rect 27249 12152 27261 12155
rect 27120 12124 27261 12152
rect 27120 12112 27126 12124
rect 27249 12121 27261 12124
rect 27295 12121 27307 12155
rect 27249 12115 27307 12121
rect 27890 12112 27896 12164
rect 27948 12112 27954 12164
rect 30282 12112 30288 12164
rect 30340 12112 30346 12164
rect 31018 12112 31024 12164
rect 31076 12112 31082 12164
rect 31662 12112 31668 12164
rect 31720 12112 31726 12164
rect 33594 12112 33600 12164
rect 33652 12112 33658 12164
rect 34348 12152 34376 12183
rect 33980 12124 34376 12152
rect 17402 12084 17408 12096
rect 16868 12056 17408 12084
rect 16669 12047 16727 12053
rect 17402 12044 17408 12056
rect 17460 12044 17466 12096
rect 18506 12044 18512 12096
rect 18564 12084 18570 12096
rect 22097 12087 22155 12093
rect 22097 12084 22109 12087
rect 18564 12056 22109 12084
rect 18564 12044 18570 12056
rect 22097 12053 22109 12056
rect 22143 12084 22155 12087
rect 23290 12084 23296 12096
rect 22143 12056 23296 12084
rect 22143 12053 22155 12056
rect 22097 12047 22155 12053
rect 23290 12044 23296 12056
rect 23348 12044 23354 12096
rect 24670 12044 24676 12096
rect 24728 12044 24734 12096
rect 24854 12044 24860 12096
rect 24912 12044 24918 12096
rect 25038 12044 25044 12096
rect 25096 12084 25102 12096
rect 25225 12087 25283 12093
rect 25225 12084 25237 12087
rect 25096 12056 25237 12084
rect 25096 12044 25102 12056
rect 25225 12053 25237 12056
rect 25271 12053 25283 12087
rect 25225 12047 25283 12053
rect 25317 12087 25375 12093
rect 25317 12053 25329 12087
rect 25363 12084 25375 12087
rect 25498 12084 25504 12096
rect 25363 12056 25504 12084
rect 25363 12053 25375 12056
rect 25317 12047 25375 12053
rect 25498 12044 25504 12056
rect 25556 12044 25562 12096
rect 33980 12093 34008 12124
rect 33965 12087 34023 12093
rect 33965 12053 33977 12087
rect 34011 12053 34023 12087
rect 33965 12047 34023 12053
rect 34146 12044 34152 12096
rect 34204 12044 34210 12096
rect 34514 12044 34520 12096
rect 34572 12044 34578 12096
rect 1104 11994 38272 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 38272 11994
rect 1104 11920 38272 11942
rect 1949 11883 2007 11889
rect 1949 11880 1961 11883
rect 1780 11852 1961 11880
rect 1780 11821 1808 11852
rect 1949 11849 1961 11852
rect 1995 11849 2007 11883
rect 1949 11843 2007 11849
rect 5442 11840 5448 11892
rect 5500 11880 5506 11892
rect 5629 11883 5687 11889
rect 5629 11880 5641 11883
rect 5500 11852 5641 11880
rect 5500 11840 5506 11852
rect 5629 11849 5641 11852
rect 5675 11849 5687 11883
rect 5629 11843 5687 11849
rect 6822 11840 6828 11892
rect 6880 11840 6886 11892
rect 8938 11840 8944 11892
rect 8996 11880 9002 11892
rect 9861 11883 9919 11889
rect 9861 11880 9873 11883
rect 8996 11852 9873 11880
rect 8996 11840 9002 11852
rect 9861 11849 9873 11852
rect 9907 11880 9919 11883
rect 11241 11883 11299 11889
rect 9907 11852 11192 11880
rect 9907 11849 9919 11852
rect 9861 11843 9919 11849
rect 1765 11815 1823 11821
rect 1765 11781 1777 11815
rect 1811 11781 1823 11815
rect 1765 11775 1823 11781
rect 6733 11815 6791 11821
rect 6733 11781 6745 11815
rect 6779 11812 6791 11815
rect 6914 11812 6920 11824
rect 6779 11784 6920 11812
rect 6779 11781 6791 11784
rect 6733 11775 6791 11781
rect 6914 11772 6920 11784
rect 6972 11812 6978 11824
rect 9217 11815 9275 11821
rect 6972 11784 8064 11812
rect 6972 11772 6978 11784
rect 8036 11756 8064 11784
rect 9217 11781 9229 11815
rect 9263 11812 9275 11815
rect 9263 11784 10180 11812
rect 9263 11781 9275 11784
rect 9217 11775 9275 11781
rect 10152 11756 10180 11784
rect 10962 11772 10968 11824
rect 11020 11772 11026 11824
rect 11164 11812 11192 11852
rect 11241 11849 11253 11883
rect 11287 11880 11299 11883
rect 11287 11852 13952 11880
rect 11287 11849 11299 11852
rect 11241 11843 11299 11849
rect 12434 11812 12440 11824
rect 11164 11784 11560 11812
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 992 11716 1409 11744
rect 992 11704 998 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 2130 11704 2136 11756
rect 2188 11704 2194 11756
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11744 5871 11747
rect 5859 11716 6408 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 6380 11617 6408 11716
rect 7374 11704 7380 11756
rect 7432 11704 7438 11756
rect 8018 11704 8024 11756
rect 8076 11704 8082 11756
rect 9030 11704 9036 11756
rect 9088 11704 9094 11756
rect 9401 11747 9459 11753
rect 9401 11713 9413 11747
rect 9447 11744 9459 11747
rect 9490 11744 9496 11756
rect 9447 11716 9496 11744
rect 9447 11713 9459 11716
rect 9401 11707 9459 11713
rect 9490 11704 9496 11716
rect 9548 11704 9554 11756
rect 9677 11747 9735 11753
rect 9677 11713 9689 11747
rect 9723 11744 9735 11747
rect 9723 11716 10088 11744
rect 9723 11713 9735 11716
rect 9677 11707 9735 11713
rect 6638 11636 6644 11688
rect 6696 11636 6702 11688
rect 6914 11636 6920 11688
rect 6972 11636 6978 11688
rect 8849 11679 8907 11685
rect 8849 11645 8861 11679
rect 8895 11645 8907 11679
rect 8849 11639 8907 11645
rect 6365 11611 6423 11617
rect 6365 11577 6377 11611
rect 6411 11577 6423 11611
rect 6656 11608 6684 11636
rect 6932 11608 6960 11636
rect 6656 11580 6960 11608
rect 6365 11571 6423 11577
rect 7098 11500 7104 11552
rect 7156 11540 7162 11552
rect 7193 11543 7251 11549
rect 7193 11540 7205 11543
rect 7156 11512 7205 11540
rect 7156 11500 7162 11512
rect 7193 11509 7205 11512
rect 7239 11509 7251 11543
rect 8864 11540 8892 11639
rect 8938 11636 8944 11688
rect 8996 11676 9002 11688
rect 9214 11676 9220 11688
rect 8996 11648 9220 11676
rect 8996 11636 9002 11648
rect 9214 11636 9220 11648
rect 9272 11636 9278 11688
rect 9508 11608 9536 11704
rect 9950 11636 9956 11688
rect 10008 11636 10014 11688
rect 10060 11676 10088 11716
rect 10134 11704 10140 11756
rect 10192 11704 10198 11756
rect 10781 11747 10839 11753
rect 10781 11744 10793 11747
rect 10244 11716 10793 11744
rect 10244 11676 10272 11716
rect 10781 11713 10793 11716
rect 10827 11744 10839 11747
rect 10980 11744 11008 11772
rect 11532 11753 11560 11784
rect 12268 11784 12440 11812
rect 12268 11753 12296 11784
rect 12434 11772 12440 11784
rect 12492 11772 12498 11824
rect 12986 11772 12992 11824
rect 13044 11772 13050 11824
rect 13924 11812 13952 11852
rect 13998 11840 14004 11892
rect 14056 11880 14062 11892
rect 18506 11880 18512 11892
rect 14056 11852 15976 11880
rect 14056 11840 14062 11852
rect 14182 11812 14188 11824
rect 13924 11784 14188 11812
rect 14182 11772 14188 11784
rect 14240 11772 14246 11824
rect 14458 11772 14464 11824
rect 14516 11812 14522 11824
rect 15010 11812 15016 11824
rect 14516 11784 15016 11812
rect 14516 11772 14522 11784
rect 15010 11772 15016 11784
rect 15068 11812 15074 11824
rect 15068 11784 15332 11812
rect 15068 11772 15074 11784
rect 10827 11716 11008 11744
rect 11149 11747 11207 11753
rect 10827 11713 10839 11716
rect 10781 11707 10839 11713
rect 11149 11713 11161 11747
rect 11195 11713 11207 11747
rect 11149 11707 11207 11713
rect 11517 11747 11575 11753
rect 11517 11713 11529 11747
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 12253 11747 12311 11753
rect 12253 11713 12265 11747
rect 12299 11713 12311 11747
rect 12253 11707 12311 11713
rect 10060 11648 10272 11676
rect 10502 11636 10508 11688
rect 10560 11636 10566 11688
rect 10686 11636 10692 11688
rect 10744 11676 10750 11688
rect 11164 11676 11192 11707
rect 14274 11704 14280 11756
rect 14332 11744 14338 11756
rect 14642 11744 14648 11756
rect 14332 11716 14648 11744
rect 14332 11704 14338 11716
rect 14642 11704 14648 11716
rect 14700 11704 14706 11756
rect 10744 11648 11192 11676
rect 12529 11679 12587 11685
rect 10744 11636 10750 11648
rect 12529 11645 12541 11679
rect 12575 11676 12587 11679
rect 12618 11676 12624 11688
rect 12575 11648 12624 11676
rect 12575 11645 12587 11648
rect 12529 11639 12587 11645
rect 12618 11636 12624 11648
rect 12676 11636 12682 11688
rect 12986 11636 12992 11688
rect 13044 11676 13050 11688
rect 14461 11679 14519 11685
rect 14461 11676 14473 11679
rect 13044 11648 14473 11676
rect 13044 11636 13050 11648
rect 14461 11645 14473 11648
rect 14507 11645 14519 11679
rect 15304 11676 15332 11784
rect 15396 11784 15884 11812
rect 15396 11753 15424 11784
rect 15381 11747 15439 11753
rect 15381 11713 15393 11747
rect 15427 11713 15439 11747
rect 15381 11707 15439 11713
rect 15470 11704 15476 11756
rect 15528 11704 15534 11756
rect 15856 11753 15884 11784
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11713 15623 11747
rect 15565 11707 15623 11713
rect 15841 11747 15899 11753
rect 15841 11713 15853 11747
rect 15887 11713 15899 11747
rect 15948 11744 15976 11852
rect 16132 11852 18512 11880
rect 16132 11821 16160 11852
rect 18506 11840 18512 11852
rect 18564 11840 18570 11892
rect 18601 11883 18659 11889
rect 18601 11849 18613 11883
rect 18647 11880 18659 11883
rect 18690 11880 18696 11892
rect 18647 11852 18696 11880
rect 18647 11849 18659 11852
rect 18601 11843 18659 11849
rect 18690 11840 18696 11852
rect 18748 11840 18754 11892
rect 22462 11840 22468 11892
rect 22520 11840 22526 11892
rect 24397 11883 24455 11889
rect 23400 11852 24256 11880
rect 16117 11815 16175 11821
rect 16117 11781 16129 11815
rect 16163 11781 16175 11815
rect 16853 11815 16911 11821
rect 16853 11812 16865 11815
rect 16117 11775 16175 11781
rect 16224 11784 16865 11812
rect 16224 11744 16252 11784
rect 16853 11781 16865 11784
rect 16899 11812 16911 11815
rect 16899 11784 17448 11812
rect 16899 11781 16911 11784
rect 16853 11775 16911 11781
rect 15948 11716 16252 11744
rect 17037 11747 17095 11753
rect 15841 11707 15899 11713
rect 17037 11713 17049 11747
rect 17083 11744 17095 11747
rect 17310 11744 17316 11756
rect 17083 11716 17316 11744
rect 17083 11713 17095 11716
rect 17037 11707 17095 11713
rect 15580 11676 15608 11707
rect 15304 11648 15608 11676
rect 15856 11676 15884 11707
rect 15930 11676 15936 11688
rect 15856 11648 15936 11676
rect 14461 11639 14519 11645
rect 15930 11636 15936 11648
rect 15988 11676 15994 11688
rect 15988 11648 16528 11676
rect 15988 11636 15994 11648
rect 16500 11620 16528 11648
rect 16574 11636 16580 11688
rect 16632 11676 16638 11688
rect 17052 11676 17080 11707
rect 17310 11704 17316 11716
rect 17368 11704 17374 11756
rect 16632 11648 17080 11676
rect 17420 11676 17448 11784
rect 17770 11772 17776 11824
rect 17828 11812 17834 11824
rect 18141 11815 18199 11821
rect 18141 11812 18153 11815
rect 17828 11784 18153 11812
rect 17828 11772 17834 11784
rect 18141 11781 18153 11784
rect 18187 11781 18199 11815
rect 18141 11775 18199 11781
rect 18230 11772 18236 11824
rect 18288 11772 18294 11824
rect 18414 11772 18420 11824
rect 18472 11812 18478 11824
rect 20809 11815 20867 11821
rect 18472 11784 19334 11812
rect 18472 11772 18478 11784
rect 17494 11704 17500 11756
rect 17552 11744 17558 11756
rect 17678 11744 17684 11756
rect 17552 11716 17684 11744
rect 17552 11704 17558 11716
rect 17678 11704 17684 11716
rect 17736 11744 17742 11756
rect 18046 11753 18052 11756
rect 17865 11747 17923 11753
rect 17865 11744 17877 11747
rect 17736 11716 17877 11744
rect 17736 11704 17742 11716
rect 17865 11713 17877 11716
rect 17911 11713 17923 11747
rect 17865 11707 17923 11713
rect 18013 11747 18052 11753
rect 18013 11713 18025 11747
rect 18013 11707 18052 11713
rect 18028 11704 18052 11707
rect 18104 11704 18110 11756
rect 18330 11747 18388 11753
rect 18330 11713 18342 11747
rect 18376 11713 18388 11747
rect 18330 11707 18388 11713
rect 18785 11747 18843 11753
rect 18785 11713 18797 11747
rect 18831 11713 18843 11747
rect 18785 11707 18843 11713
rect 18028 11676 18056 11704
rect 17420 11648 18056 11676
rect 16632 11636 16638 11648
rect 11514 11608 11520 11620
rect 9508 11580 11520 11608
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 15749 11611 15807 11617
rect 15749 11608 15761 11611
rect 14476 11580 15761 11608
rect 10502 11540 10508 11552
rect 8864 11512 10508 11540
rect 7193 11503 7251 11509
rect 10502 11500 10508 11512
rect 10560 11500 10566 11552
rect 11701 11543 11759 11549
rect 11701 11509 11713 11543
rect 11747 11540 11759 11543
rect 12250 11540 12256 11552
rect 11747 11512 12256 11540
rect 11747 11509 11759 11512
rect 11701 11503 11759 11509
rect 12250 11500 12256 11512
rect 12308 11500 12314 11552
rect 13078 11500 13084 11552
rect 13136 11540 13142 11552
rect 14476 11540 14504 11580
rect 15749 11577 15761 11580
rect 15795 11577 15807 11611
rect 15749 11571 15807 11577
rect 13136 11512 14504 11540
rect 13136 11500 13142 11512
rect 15194 11500 15200 11552
rect 15252 11500 15258 11552
rect 15764 11540 15792 11571
rect 16482 11568 16488 11620
rect 16540 11568 16546 11620
rect 17402 11608 17408 11620
rect 16592 11580 17408 11608
rect 16592 11540 16620 11580
rect 17402 11568 17408 11580
rect 17460 11568 17466 11620
rect 18345 11608 18373 11707
rect 18414 11636 18420 11688
rect 18472 11676 18478 11688
rect 18800 11676 18828 11707
rect 18966 11704 18972 11756
rect 19024 11704 19030 11756
rect 19061 11747 19119 11753
rect 19061 11713 19073 11747
rect 19107 11713 19119 11747
rect 19306 11744 19334 11784
rect 20809 11781 20821 11815
rect 20855 11812 20867 11815
rect 20898 11812 20904 11824
rect 20855 11784 20904 11812
rect 20855 11781 20867 11784
rect 20809 11775 20867 11781
rect 20898 11772 20904 11784
rect 20956 11772 20962 11824
rect 20993 11815 21051 11821
rect 20993 11781 21005 11815
rect 21039 11812 21051 11815
rect 21542 11812 21548 11824
rect 21039 11784 21548 11812
rect 21039 11781 21051 11784
rect 20993 11775 21051 11781
rect 21542 11772 21548 11784
rect 21600 11812 21606 11824
rect 22094 11812 22100 11824
rect 21600 11784 22100 11812
rect 21600 11772 21606 11784
rect 22094 11772 22100 11784
rect 22152 11772 22158 11824
rect 22186 11772 22192 11824
rect 22244 11772 22250 11824
rect 22278 11772 22284 11824
rect 22336 11812 22342 11824
rect 23400 11812 23428 11852
rect 22336 11784 23428 11812
rect 22336 11772 22342 11784
rect 23474 11772 23480 11824
rect 23532 11812 23538 11824
rect 23661 11815 23719 11821
rect 23661 11812 23673 11815
rect 23532 11784 23673 11812
rect 23532 11772 23538 11784
rect 23661 11781 23673 11784
rect 23707 11781 23719 11815
rect 23661 11775 23719 11781
rect 23845 11815 23903 11821
rect 23845 11781 23857 11815
rect 23891 11812 23903 11815
rect 24118 11812 24124 11824
rect 23891 11784 24124 11812
rect 23891 11781 23903 11784
rect 23845 11775 23903 11781
rect 24118 11772 24124 11784
rect 24176 11772 24182 11824
rect 24228 11821 24256 11852
rect 24397 11849 24409 11883
rect 24443 11880 24455 11883
rect 24949 11883 25007 11889
rect 24949 11880 24961 11883
rect 24443 11852 24961 11880
rect 24443 11849 24455 11852
rect 24397 11843 24455 11849
rect 24949 11849 24961 11852
rect 24995 11880 25007 11883
rect 27062 11880 27068 11892
rect 24995 11852 27068 11880
rect 24995 11849 25007 11852
rect 24949 11843 25007 11849
rect 24213 11815 24271 11821
rect 24213 11781 24225 11815
rect 24259 11781 24271 11815
rect 24213 11775 24271 11781
rect 22204 11744 22232 11772
rect 19306 11716 22232 11744
rect 22833 11747 22891 11753
rect 19061 11707 19119 11713
rect 22833 11713 22845 11747
rect 22879 11713 22891 11747
rect 22833 11707 22891 11713
rect 18472 11648 18828 11676
rect 18472 11636 18478 11648
rect 18874 11636 18880 11688
rect 18932 11676 18938 11688
rect 19076 11676 19104 11707
rect 18932 11648 19104 11676
rect 22848 11676 22876 11707
rect 23290 11704 23296 11756
rect 23348 11744 23354 11756
rect 23385 11747 23443 11753
rect 23385 11744 23397 11747
rect 23348 11716 23397 11744
rect 23348 11704 23354 11716
rect 23385 11713 23397 11716
rect 23431 11744 23443 11747
rect 24412 11744 24440 11843
rect 27062 11840 27068 11852
rect 27120 11840 27126 11892
rect 28442 11840 28448 11892
rect 28500 11880 28506 11892
rect 30006 11880 30012 11892
rect 28500 11852 30012 11880
rect 28500 11840 28506 11852
rect 30006 11840 30012 11852
rect 30064 11840 30070 11892
rect 30101 11883 30159 11889
rect 30101 11849 30113 11883
rect 30147 11880 30159 11883
rect 30282 11880 30288 11892
rect 30147 11852 30288 11880
rect 30147 11849 30159 11852
rect 30101 11843 30159 11849
rect 30282 11840 30288 11852
rect 30340 11840 30346 11892
rect 34146 11840 34152 11892
rect 34204 11880 34210 11892
rect 34204 11852 35112 11880
rect 34204 11840 34210 11852
rect 24765 11815 24823 11821
rect 24765 11781 24777 11815
rect 24811 11781 24823 11815
rect 24765 11775 24823 11781
rect 23431 11716 24440 11744
rect 23431 11713 23443 11716
rect 23385 11707 23443 11713
rect 24780 11688 24808 11775
rect 25130 11772 25136 11824
rect 25188 11812 25194 11824
rect 25314 11812 25320 11824
rect 25188 11784 25320 11812
rect 25188 11772 25194 11784
rect 25314 11772 25320 11784
rect 25372 11772 25378 11824
rect 29362 11772 29368 11824
rect 29420 11772 29426 11824
rect 30745 11815 30803 11821
rect 30745 11812 30757 11815
rect 29564 11784 30757 11812
rect 25225 11747 25283 11753
rect 25225 11713 25237 11747
rect 25271 11744 25283 11747
rect 26786 11744 26792 11756
rect 25271 11716 26792 11744
rect 25271 11713 25283 11716
rect 25225 11707 25283 11713
rect 25516 11688 25544 11716
rect 26786 11704 26792 11716
rect 26844 11744 26850 11756
rect 27982 11744 27988 11756
rect 26844 11716 27988 11744
rect 26844 11704 26850 11716
rect 27982 11704 27988 11716
rect 28040 11704 28046 11756
rect 22848 11648 23152 11676
rect 18932 11636 18938 11648
rect 17926 11580 18373 11608
rect 15764 11512 16620 11540
rect 16669 11543 16727 11549
rect 16669 11509 16681 11543
rect 16715 11540 16727 11543
rect 16850 11540 16856 11552
rect 16715 11512 16856 11540
rect 16715 11509 16727 11512
rect 16669 11503 16727 11509
rect 16850 11500 16856 11512
rect 16908 11500 16914 11552
rect 17126 11500 17132 11552
rect 17184 11540 17190 11552
rect 17310 11540 17316 11552
rect 17184 11512 17316 11540
rect 17184 11500 17190 11512
rect 17310 11500 17316 11512
rect 17368 11540 17374 11552
rect 17926 11540 17954 11580
rect 18598 11568 18604 11620
rect 18656 11608 18662 11620
rect 22848 11608 22876 11648
rect 18656 11580 22876 11608
rect 18656 11568 18662 11580
rect 23124 11552 23152 11648
rect 23474 11636 23480 11688
rect 23532 11676 23538 11688
rect 24762 11676 24768 11688
rect 23532 11648 24768 11676
rect 23532 11636 23538 11648
rect 24762 11636 24768 11648
rect 24820 11636 24826 11688
rect 25498 11636 25504 11688
rect 25556 11636 25562 11688
rect 27338 11636 27344 11688
rect 27396 11676 27402 11688
rect 27614 11676 27620 11688
rect 27396 11648 27620 11676
rect 27396 11636 27402 11648
rect 27614 11636 27620 11648
rect 27672 11676 27678 11688
rect 28534 11676 28540 11688
rect 27672 11648 28540 11676
rect 27672 11636 27678 11648
rect 28534 11636 28540 11648
rect 28592 11636 28598 11688
rect 29380 11676 29408 11772
rect 29564 11753 29592 11784
rect 30745 11781 30757 11784
rect 30791 11781 30803 11815
rect 30745 11775 30803 11781
rect 34054 11772 34060 11824
rect 34112 11772 34118 11824
rect 34514 11772 34520 11824
rect 34572 11812 34578 11824
rect 34793 11815 34851 11821
rect 34793 11812 34805 11815
rect 34572 11784 34805 11812
rect 34572 11772 34578 11784
rect 34793 11781 34805 11784
rect 34839 11781 34851 11815
rect 34793 11775 34851 11781
rect 29549 11747 29607 11753
rect 29549 11713 29561 11747
rect 29595 11713 29607 11747
rect 29549 11707 29607 11713
rect 29733 11747 29791 11753
rect 29733 11713 29745 11747
rect 29779 11713 29791 11747
rect 29733 11707 29791 11713
rect 29748 11676 29776 11707
rect 29822 11704 29828 11756
rect 29880 11704 29886 11756
rect 29914 11704 29920 11756
rect 29972 11744 29978 11756
rect 30282 11744 30288 11756
rect 29972 11716 30288 11744
rect 29972 11704 29978 11716
rect 30282 11704 30288 11716
rect 30340 11704 30346 11756
rect 31294 11704 31300 11756
rect 31352 11704 31358 11756
rect 35084 11753 35112 11852
rect 35069 11747 35127 11753
rect 35069 11713 35081 11747
rect 35115 11713 35127 11747
rect 35069 11707 35127 11713
rect 37642 11704 37648 11756
rect 37700 11704 37706 11756
rect 29380 11648 29776 11676
rect 29840 11676 29868 11704
rect 30190 11676 30196 11688
rect 29840 11648 30196 11676
rect 30190 11636 30196 11648
rect 30248 11636 30254 11688
rect 33321 11679 33379 11685
rect 33321 11645 33333 11679
rect 33367 11676 33379 11679
rect 33594 11676 33600 11688
rect 33367 11648 33600 11676
rect 33367 11645 33379 11648
rect 33321 11639 33379 11645
rect 33594 11636 33600 11648
rect 33652 11636 33658 11688
rect 23860 11580 24992 11608
rect 17368 11512 17954 11540
rect 17368 11500 17374 11512
rect 18506 11500 18512 11552
rect 18564 11500 18570 11552
rect 20806 11500 20812 11552
rect 20864 11540 20870 11552
rect 21085 11543 21143 11549
rect 21085 11540 21097 11543
rect 20864 11512 21097 11540
rect 20864 11500 20870 11512
rect 21085 11509 21097 11512
rect 21131 11540 21143 11543
rect 22094 11540 22100 11552
rect 21131 11512 22100 11540
rect 21131 11509 21143 11512
rect 21085 11503 21143 11509
rect 22094 11500 22100 11512
rect 22152 11500 22158 11552
rect 23106 11500 23112 11552
rect 23164 11540 23170 11552
rect 23860 11549 23888 11580
rect 23845 11543 23903 11549
rect 23845 11540 23857 11543
rect 23164 11512 23857 11540
rect 23164 11500 23170 11512
rect 23845 11509 23857 11512
rect 23891 11509 23903 11543
rect 23845 11503 23903 11509
rect 23934 11500 23940 11552
rect 23992 11540 23998 11552
rect 24029 11543 24087 11549
rect 24029 11540 24041 11543
rect 23992 11512 24041 11540
rect 23992 11500 23998 11512
rect 24029 11509 24041 11512
rect 24075 11509 24087 11543
rect 24029 11503 24087 11509
rect 24302 11500 24308 11552
rect 24360 11540 24366 11552
rect 24397 11543 24455 11549
rect 24397 11540 24409 11543
rect 24360 11512 24409 11540
rect 24360 11500 24366 11512
rect 24397 11509 24409 11512
rect 24443 11509 24455 11543
rect 24397 11503 24455 11509
rect 24486 11500 24492 11552
rect 24544 11540 24550 11552
rect 24964 11549 24992 11580
rect 27062 11568 27068 11620
rect 27120 11608 27126 11620
rect 30374 11608 30380 11620
rect 27120 11580 30380 11608
rect 27120 11568 27126 11580
rect 30374 11568 30380 11580
rect 30432 11568 30438 11620
rect 37826 11568 37832 11620
rect 37884 11568 37890 11620
rect 24581 11543 24639 11549
rect 24581 11540 24593 11543
rect 24544 11512 24593 11540
rect 24544 11500 24550 11512
rect 24581 11509 24593 11512
rect 24627 11509 24639 11543
rect 24581 11503 24639 11509
rect 24949 11543 25007 11549
rect 24949 11509 24961 11543
rect 24995 11540 25007 11543
rect 27706 11540 27712 11552
rect 24995 11512 27712 11540
rect 24995 11509 25007 11512
rect 24949 11503 25007 11509
rect 27706 11500 27712 11512
rect 27764 11500 27770 11552
rect 1104 11450 38272 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38272 11450
rect 1104 11376 38272 11398
rect 2130 11296 2136 11348
rect 2188 11336 2194 11348
rect 4709 11339 4767 11345
rect 4709 11336 4721 11339
rect 2188 11308 4721 11336
rect 2188 11296 2194 11308
rect 4709 11305 4721 11308
rect 4755 11305 4767 11339
rect 4709 11299 4767 11305
rect 10134 11296 10140 11348
rect 10192 11296 10198 11348
rect 12618 11296 12624 11348
rect 12676 11336 12682 11348
rect 12805 11339 12863 11345
rect 12805 11336 12817 11339
rect 12676 11308 12817 11336
rect 12676 11296 12682 11308
rect 12805 11305 12817 11308
rect 12851 11305 12863 11339
rect 12805 11299 12863 11305
rect 12894 11296 12900 11348
rect 12952 11336 12958 11348
rect 14829 11339 14887 11345
rect 12952 11308 14228 11336
rect 12952 11296 12958 11308
rect 7009 11203 7067 11209
rect 7009 11169 7021 11203
rect 7055 11200 7067 11203
rect 7098 11200 7104 11212
rect 7055 11172 7104 11200
rect 7055 11169 7067 11172
rect 7009 11163 7067 11169
rect 7098 11160 7104 11172
rect 7156 11160 7162 11212
rect 4893 11135 4951 11141
rect 4893 11101 4905 11135
rect 4939 11101 4951 11135
rect 4893 11095 4951 11101
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11132 5135 11135
rect 5626 11132 5632 11144
rect 5123 11104 5632 11132
rect 5123 11101 5135 11104
rect 5077 11095 5135 11101
rect 4908 11064 4936 11095
rect 5626 11092 5632 11104
rect 5684 11092 5690 11144
rect 6454 11092 6460 11144
rect 6512 11092 6518 11144
rect 10152 11141 10180 11296
rect 12912 11268 12940 11296
rect 11900 11240 12940 11268
rect 13173 11271 13231 11277
rect 10870 11160 10876 11212
rect 10928 11160 10934 11212
rect 6549 11135 6607 11141
rect 6549 11101 6561 11135
rect 6595 11132 6607 11135
rect 6733 11135 6791 11141
rect 6733 11132 6745 11135
rect 6595 11104 6745 11132
rect 6595 11101 6607 11104
rect 6549 11095 6607 11101
rect 6733 11101 6745 11104
rect 6779 11101 6791 11135
rect 6733 11095 6791 11101
rect 10137 11135 10195 11141
rect 10137 11101 10149 11135
rect 10183 11101 10195 11135
rect 10137 11095 10195 11101
rect 10686 11092 10692 11144
rect 10744 11092 10750 11144
rect 11698 11092 11704 11144
rect 11756 11132 11762 11144
rect 11900 11141 11928 11240
rect 13173 11237 13185 11271
rect 13219 11237 13231 11271
rect 13173 11231 13231 11237
rect 13078 11200 13084 11212
rect 11992 11172 13084 11200
rect 11992 11141 12020 11172
rect 13078 11160 13084 11172
rect 13136 11160 13142 11212
rect 11885 11135 11943 11141
rect 11885 11132 11897 11135
rect 11756 11104 11897 11132
rect 11756 11092 11762 11104
rect 11885 11101 11897 11104
rect 11931 11101 11943 11135
rect 11885 11095 11943 11101
rect 11977 11135 12035 11141
rect 11977 11101 11989 11135
rect 12023 11101 12035 11135
rect 11977 11095 12035 11101
rect 5442 11064 5448 11076
rect 4908 11036 5448 11064
rect 5442 11024 5448 11036
rect 5500 11024 5506 11076
rect 6472 11064 6500 11092
rect 6914 11064 6920 11076
rect 6472 11036 6920 11064
rect 6914 11024 6920 11036
rect 6972 11024 6978 11076
rect 7742 11024 7748 11076
rect 7800 11024 7806 11076
rect 11992 11064 12020 11095
rect 12158 11092 12164 11144
rect 12216 11092 12222 11144
rect 12253 11135 12311 11141
rect 12253 11101 12265 11135
rect 12299 11132 12311 11135
rect 12989 11135 13047 11141
rect 12299 11104 12434 11132
rect 12299 11101 12311 11104
rect 12253 11095 12311 11101
rect 8496 11036 12020 11064
rect 12406 11064 12434 11104
rect 12989 11101 13001 11135
rect 13035 11132 13047 11135
rect 13188 11132 13216 11231
rect 13725 11203 13783 11209
rect 13725 11169 13737 11203
rect 13771 11200 13783 11203
rect 13814 11200 13820 11212
rect 13771 11172 13820 11200
rect 13771 11169 13783 11172
rect 13725 11163 13783 11169
rect 13814 11160 13820 11172
rect 13872 11200 13878 11212
rect 14090 11200 14096 11212
rect 13872 11172 14096 11200
rect 13872 11160 13878 11172
rect 14090 11160 14096 11172
rect 14148 11160 14154 11212
rect 14200 11200 14228 11308
rect 14829 11305 14841 11339
rect 14875 11336 14887 11339
rect 15102 11336 15108 11348
rect 14875 11308 15108 11336
rect 14875 11305 14887 11308
rect 14829 11299 14887 11305
rect 15102 11296 15108 11308
rect 15160 11296 15166 11348
rect 15654 11296 15660 11348
rect 15712 11296 15718 11348
rect 16022 11336 16028 11348
rect 15856 11308 16028 11336
rect 14200 11172 14734 11200
rect 13035 11104 13216 11132
rect 13035 11101 13047 11104
rect 12989 11095 13047 11101
rect 13446 11092 13452 11144
rect 13504 11092 13510 11144
rect 13541 11135 13599 11141
rect 13541 11101 13553 11135
rect 13587 11132 13599 11135
rect 13998 11132 14004 11144
rect 13587 11104 14004 11132
rect 13587 11101 13599 11104
rect 13541 11095 13599 11101
rect 13998 11092 14004 11104
rect 14056 11092 14062 11144
rect 14182 11092 14188 11144
rect 14240 11092 14246 11144
rect 14274 11092 14280 11144
rect 14332 11132 14338 11144
rect 14706 11141 14734 11172
rect 15194 11160 15200 11212
rect 15252 11160 15258 11212
rect 14691 11135 14749 11141
rect 14332 11104 14377 11132
rect 14332 11092 14338 11104
rect 14691 11101 14703 11135
rect 14737 11132 14749 11135
rect 14918 11132 14924 11144
rect 14737 11104 14924 11132
rect 14737 11101 14749 11104
rect 14691 11095 14749 11101
rect 14918 11092 14924 11104
rect 14976 11092 14982 11144
rect 15212 11132 15240 11160
rect 15289 11135 15347 11141
rect 15289 11132 15301 11135
rect 15212 11104 15301 11132
rect 15289 11101 15301 11104
rect 15335 11101 15347 11135
rect 15289 11095 15347 11101
rect 15382 11135 15440 11141
rect 15382 11101 15394 11135
rect 15428 11101 15440 11135
rect 15382 11095 15440 11101
rect 13464 11064 13492 11092
rect 12406 11036 13492 11064
rect 13633 11067 13691 11073
rect 8496 11008 8524 11036
rect 13633 11033 13645 11067
rect 13679 11064 13691 11067
rect 13814 11064 13820 11076
rect 13679 11036 13820 11064
rect 13679 11033 13691 11036
rect 13633 11027 13691 11033
rect 13814 11024 13820 11036
rect 13872 11024 13878 11076
rect 14090 11024 14096 11076
rect 14148 11064 14154 11076
rect 14458 11064 14464 11076
rect 14148 11036 14464 11064
rect 14148 11024 14154 11036
rect 14458 11024 14464 11036
rect 14516 11024 14522 11076
rect 14550 11024 14556 11076
rect 14608 11024 14614 11076
rect 15396 11064 15424 11095
rect 15562 11092 15568 11144
rect 15620 11092 15626 11144
rect 15672 11141 15700 11296
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11101 15715 11135
rect 15657 11095 15715 11101
rect 15754 11135 15812 11141
rect 15754 11101 15766 11135
rect 15800 11132 15812 11135
rect 15856 11132 15884 11308
rect 16022 11296 16028 11308
rect 16080 11296 16086 11348
rect 16206 11296 16212 11348
rect 16264 11336 16270 11348
rect 16264 11308 16712 11336
rect 16264 11296 16270 11308
rect 15933 11271 15991 11277
rect 15933 11237 15945 11271
rect 15979 11268 15991 11271
rect 16684 11268 16712 11308
rect 16758 11296 16764 11348
rect 16816 11296 16822 11348
rect 17957 11339 18015 11345
rect 17957 11305 17969 11339
rect 18003 11336 18015 11339
rect 18414 11336 18420 11348
rect 18003 11308 18420 11336
rect 18003 11305 18015 11308
rect 17957 11299 18015 11305
rect 18414 11296 18420 11308
rect 18472 11296 18478 11348
rect 18877 11339 18935 11345
rect 18877 11305 18889 11339
rect 18923 11336 18935 11339
rect 19150 11336 19156 11348
rect 18923 11308 19156 11336
rect 18923 11305 18935 11308
rect 18877 11299 18935 11305
rect 19150 11296 19156 11308
rect 19208 11296 19214 11348
rect 20162 11296 20168 11348
rect 20220 11336 20226 11348
rect 20220 11308 23060 11336
rect 20220 11296 20226 11308
rect 16945 11271 17003 11277
rect 16945 11268 16957 11271
rect 15979 11240 16344 11268
rect 16684 11240 16957 11268
rect 15979 11237 15991 11240
rect 15933 11231 15991 11237
rect 16206 11160 16212 11212
rect 16264 11160 16270 11212
rect 16316 11200 16344 11240
rect 16945 11237 16957 11240
rect 16991 11237 17003 11271
rect 16945 11231 17003 11237
rect 18340 11240 20024 11268
rect 18340 11212 18368 11240
rect 16669 11203 16727 11209
rect 16669 11200 16681 11203
rect 16316 11172 16681 11200
rect 16669 11169 16681 11172
rect 16715 11169 16727 11203
rect 16669 11163 16727 11169
rect 17144 11172 17724 11200
rect 15800 11104 15884 11132
rect 16025 11135 16083 11141
rect 15800 11101 15812 11104
rect 15754 11095 15812 11101
rect 16025 11101 16037 11135
rect 16071 11101 16083 11135
rect 16025 11095 16083 11101
rect 16577 11135 16635 11141
rect 16577 11101 16589 11135
rect 16623 11101 16635 11135
rect 16577 11095 16635 11101
rect 15028 11036 15424 11064
rect 8478 10956 8484 11008
rect 8536 10956 8542 11008
rect 11606 10956 11612 11008
rect 11664 10996 11670 11008
rect 11701 10999 11759 11005
rect 11701 10996 11713 10999
rect 11664 10968 11713 10996
rect 11664 10956 11670 10968
rect 11701 10965 11713 10968
rect 11747 10965 11759 10999
rect 11701 10959 11759 10965
rect 11974 10956 11980 11008
rect 12032 10996 12038 11008
rect 12526 10996 12532 11008
rect 12032 10968 12532 10996
rect 12032 10956 12038 10968
rect 12526 10956 12532 10968
rect 12584 10956 12590 11008
rect 14274 10956 14280 11008
rect 14332 10996 14338 11008
rect 15028 10996 15056 11036
rect 14332 10968 15056 10996
rect 14332 10956 14338 10968
rect 15102 10956 15108 11008
rect 15160 10996 15166 11008
rect 15470 10996 15476 11008
rect 15160 10968 15476 10996
rect 15160 10956 15166 10968
rect 15470 10956 15476 10968
rect 15528 10996 15534 11008
rect 16040 10996 16068 11095
rect 16592 11064 16620 11095
rect 17034 11064 17040 11076
rect 16592 11036 17040 11064
rect 17034 11024 17040 11036
rect 17092 11024 17098 11076
rect 15528 10968 16068 10996
rect 15528 10956 15534 10968
rect 16574 10956 16580 11008
rect 16632 10996 16638 11008
rect 17144 10996 17172 11172
rect 17310 11092 17316 11144
rect 17368 11092 17374 11144
rect 17402 11092 17408 11144
rect 17460 11132 17466 11144
rect 17460 11104 17505 11132
rect 17460 11092 17466 11104
rect 17218 11024 17224 11076
rect 17276 11064 17282 11076
rect 17696 11073 17724 11172
rect 18322 11160 18328 11212
rect 18380 11160 18386 11212
rect 18414 11160 18420 11212
rect 18472 11160 18478 11212
rect 18524 11172 18736 11200
rect 18524 11144 18552 11172
rect 17770 11092 17776 11144
rect 17828 11141 17834 11144
rect 17828 11132 17836 11141
rect 17828 11104 17873 11132
rect 17828 11095 17836 11104
rect 17828 11092 17834 11095
rect 18506 11092 18512 11144
rect 18564 11092 18570 11144
rect 18598 11092 18604 11144
rect 18656 11092 18662 11144
rect 18708 11141 18736 11172
rect 18966 11160 18972 11212
rect 19024 11200 19030 11212
rect 19996 11200 20024 11240
rect 20070 11228 20076 11280
rect 20128 11228 20134 11280
rect 21634 11268 21640 11280
rect 20823 11240 21640 11268
rect 19024 11172 19840 11200
rect 19996 11172 20576 11200
rect 19024 11160 19030 11172
rect 18693 11135 18751 11141
rect 18693 11101 18705 11135
rect 18739 11101 18751 11135
rect 18693 11095 18751 11101
rect 19426 11092 19432 11144
rect 19484 11092 19490 11144
rect 19812 11141 19840 11172
rect 19797 11135 19855 11141
rect 19797 11101 19809 11135
rect 19843 11101 19855 11135
rect 19797 11095 19855 11101
rect 20441 11135 20499 11141
rect 20441 11101 20453 11135
rect 20487 11101 20499 11135
rect 20548 11132 20576 11172
rect 20714 11160 20720 11212
rect 20772 11160 20778 11212
rect 20823 11132 20851 11240
rect 21634 11228 21640 11240
rect 21692 11228 21698 11280
rect 21729 11271 21787 11277
rect 21729 11237 21741 11271
rect 21775 11237 21787 11271
rect 21729 11231 21787 11237
rect 20898 11160 20904 11212
rect 20956 11200 20962 11212
rect 21744 11200 21772 11231
rect 21818 11228 21824 11280
rect 21876 11268 21882 11280
rect 22922 11268 22928 11280
rect 21876 11240 22928 11268
rect 21876 11228 21882 11240
rect 22922 11228 22928 11240
rect 22980 11228 22986 11280
rect 23032 11268 23060 11308
rect 24486 11296 24492 11348
rect 24544 11336 24550 11348
rect 26789 11339 26847 11345
rect 24544 11308 26740 11336
rect 24544 11296 24550 11308
rect 23658 11268 23664 11280
rect 23032 11240 23664 11268
rect 20956 11172 21036 11200
rect 21744 11172 21864 11200
rect 20956 11160 20962 11172
rect 21008 11141 21036 11172
rect 21836 11144 21864 11172
rect 20548 11104 20851 11132
rect 20993 11135 21051 11141
rect 20441 11095 20499 11101
rect 20993 11101 21005 11135
rect 21039 11101 21051 11135
rect 20993 11095 21051 11101
rect 17589 11067 17647 11073
rect 17589 11064 17601 11067
rect 17276 11036 17601 11064
rect 17276 11024 17282 11036
rect 17589 11033 17601 11036
rect 17635 11033 17647 11067
rect 17589 11027 17647 11033
rect 17681 11067 17739 11073
rect 17681 11033 17693 11067
rect 17727 11033 17739 11067
rect 17681 11027 17739 11033
rect 18230 11024 18236 11076
rect 18288 11064 18294 11076
rect 19521 11067 19579 11073
rect 19521 11064 19533 11067
rect 18288 11036 19533 11064
rect 18288 11024 18294 11036
rect 19521 11033 19533 11036
rect 19567 11033 19579 11067
rect 19521 11027 19579 11033
rect 19613 11067 19671 11073
rect 19613 11033 19625 11067
rect 19659 11064 19671 11067
rect 19702 11064 19708 11076
rect 19659 11036 19708 11064
rect 19659 11033 19671 11036
rect 19613 11027 19671 11033
rect 19702 11024 19708 11036
rect 19760 11024 19766 11076
rect 20456 11064 20484 11095
rect 20898 11064 20904 11076
rect 20456 11036 20904 11064
rect 20898 11024 20904 11036
rect 20956 11024 20962 11076
rect 21008 11064 21036 11095
rect 21266 11092 21272 11144
rect 21324 11132 21330 11144
rect 21361 11135 21419 11141
rect 21361 11132 21373 11135
rect 21324 11104 21373 11132
rect 21324 11092 21330 11104
rect 21361 11101 21373 11104
rect 21407 11101 21419 11135
rect 21361 11095 21419 11101
rect 21818 11092 21824 11144
rect 21876 11132 21882 11144
rect 21876 11104 22140 11132
rect 21876 11092 21882 11104
rect 22112 11064 22140 11104
rect 22186 11092 22192 11144
rect 22244 11092 22250 11144
rect 22554 11092 22560 11144
rect 22612 11092 22618 11144
rect 23032 11142 23060 11240
rect 23658 11228 23664 11240
rect 23716 11228 23722 11280
rect 23753 11271 23811 11277
rect 23753 11237 23765 11271
rect 23799 11268 23811 11271
rect 24210 11268 24216 11280
rect 23799 11240 24216 11268
rect 23799 11237 23811 11240
rect 23753 11231 23811 11237
rect 24210 11228 24216 11240
rect 24268 11228 24274 11280
rect 25317 11271 25375 11277
rect 25317 11237 25329 11271
rect 25363 11237 25375 11271
rect 26712 11268 26740 11308
rect 26789 11305 26801 11339
rect 26835 11336 26847 11339
rect 27522 11336 27528 11348
rect 26835 11308 27528 11336
rect 26835 11305 26847 11308
rect 26789 11299 26847 11305
rect 27522 11296 27528 11308
rect 27580 11296 27586 11348
rect 28350 11296 28356 11348
rect 28408 11296 28414 11348
rect 28442 11296 28448 11348
rect 28500 11296 28506 11348
rect 28534 11296 28540 11348
rect 28592 11336 28598 11348
rect 28592 11308 28994 11336
rect 28592 11296 28598 11308
rect 27614 11268 27620 11280
rect 26712 11240 27620 11268
rect 25317 11231 25375 11237
rect 25332 11200 25360 11231
rect 27614 11228 27620 11240
rect 27672 11228 27678 11280
rect 28261 11271 28319 11277
rect 28261 11237 28273 11271
rect 28307 11268 28319 11271
rect 28460 11268 28488 11296
rect 28307 11240 28488 11268
rect 28721 11271 28779 11277
rect 28307 11237 28319 11240
rect 28261 11231 28319 11237
rect 28721 11237 28733 11271
rect 28767 11237 28779 11271
rect 28721 11231 28779 11237
rect 26145 11203 26203 11209
rect 23493 11172 25268 11200
rect 25332 11172 26004 11200
rect 23097 11145 23155 11151
rect 23097 11142 23109 11145
rect 23032 11114 23109 11142
rect 23097 11111 23109 11114
rect 23143 11111 23155 11145
rect 23097 11105 23155 11111
rect 23290 11092 23296 11144
rect 23348 11092 23354 11144
rect 23385 11135 23443 11141
rect 23385 11101 23397 11135
rect 23431 11101 23443 11135
rect 23493 11119 23521 11172
rect 23385 11095 23443 11101
rect 23478 11113 23536 11119
rect 22830 11064 22836 11076
rect 21008 11036 21496 11064
rect 22112 11036 22836 11064
rect 16632 10968 17172 10996
rect 16632 10956 16638 10968
rect 17494 10956 17500 11008
rect 17552 10996 17558 11008
rect 18874 10996 18880 11008
rect 17552 10968 18880 10996
rect 17552 10956 17558 10968
rect 18874 10956 18880 10968
rect 18932 10956 18938 11008
rect 19242 10956 19248 11008
rect 19300 10956 19306 11008
rect 21468 10996 21496 11036
rect 22830 11024 22836 11036
rect 22888 11064 22894 11076
rect 23400 11064 23428 11095
rect 23478 11079 23490 11113
rect 23524 11079 23536 11113
rect 23750 11092 23756 11144
rect 23808 11132 23814 11144
rect 23934 11132 23940 11144
rect 23808 11104 23940 11132
rect 23808 11092 23814 11104
rect 23934 11092 23940 11104
rect 23992 11092 23998 11144
rect 24765 11135 24823 11141
rect 24765 11101 24777 11135
rect 24811 11101 24823 11135
rect 24765 11095 24823 11101
rect 23478 11076 23536 11079
rect 22888 11036 23428 11064
rect 22888 11024 22894 11036
rect 23474 11024 23480 11076
rect 23532 11024 23538 11076
rect 24026 11024 24032 11076
rect 24084 11064 24090 11076
rect 24780 11064 24808 11095
rect 24946 11092 24952 11144
rect 25004 11092 25010 11144
rect 25130 11092 25136 11144
rect 25188 11092 25194 11144
rect 24084 11036 24808 11064
rect 25041 11067 25099 11073
rect 24084 11024 24090 11036
rect 25041 11033 25053 11067
rect 25087 11033 25099 11067
rect 25240 11064 25268 11172
rect 25498 11092 25504 11144
rect 25556 11092 25562 11144
rect 25685 11135 25743 11141
rect 25685 11101 25697 11135
rect 25731 11101 25743 11135
rect 25685 11095 25743 11101
rect 25700 11064 25728 11095
rect 25774 11092 25780 11144
rect 25832 11092 25838 11144
rect 25866 11092 25872 11144
rect 25924 11092 25930 11144
rect 25976 11141 26004 11172
rect 26145 11169 26157 11203
rect 26191 11200 26203 11203
rect 26329 11203 26387 11209
rect 26329 11200 26341 11203
rect 26191 11172 26341 11200
rect 26191 11169 26203 11172
rect 26145 11163 26203 11169
rect 26329 11169 26341 11172
rect 26375 11169 26387 11203
rect 28445 11203 28503 11209
rect 28445 11200 28457 11203
rect 26329 11163 26387 11169
rect 27586 11172 28457 11200
rect 25961 11135 26019 11141
rect 25961 11101 25973 11135
rect 26007 11101 26019 11135
rect 25961 11095 26019 11101
rect 26237 11135 26295 11141
rect 26237 11101 26249 11135
rect 26283 11132 26295 11135
rect 26418 11132 26424 11144
rect 26283 11104 26424 11132
rect 26283 11101 26295 11104
rect 26237 11095 26295 11101
rect 26418 11092 26424 11104
rect 26476 11092 26482 11144
rect 26510 11092 26516 11144
rect 26568 11092 26574 11144
rect 26602 11092 26608 11144
rect 26660 11092 26666 11144
rect 27586 11064 27614 11172
rect 28445 11169 28457 11172
rect 28491 11169 28503 11203
rect 28445 11163 28503 11169
rect 27798 11092 27804 11144
rect 27856 11092 27862 11144
rect 28077 11135 28135 11141
rect 28077 11132 28089 11135
rect 27908 11104 28089 11132
rect 27908 11064 27936 11104
rect 28077 11101 28089 11104
rect 28123 11101 28135 11135
rect 28077 11095 28135 11101
rect 28258 11092 28264 11144
rect 28316 11132 28322 11144
rect 28353 11135 28411 11141
rect 28353 11132 28365 11135
rect 28316 11104 28365 11132
rect 28316 11092 28322 11104
rect 28353 11101 28365 11104
rect 28399 11101 28411 11135
rect 28736 11132 28764 11231
rect 28966 11200 28994 11308
rect 29454 11296 29460 11348
rect 29512 11336 29518 11348
rect 29549 11339 29607 11345
rect 29549 11336 29561 11339
rect 29512 11308 29561 11336
rect 29512 11296 29518 11308
rect 29549 11305 29561 11308
rect 29595 11305 29607 11339
rect 29549 11299 29607 11305
rect 30558 11268 30564 11280
rect 30300 11240 30564 11268
rect 29917 11203 29975 11209
rect 28966 11172 29316 11200
rect 28353 11095 28411 11101
rect 28460 11104 28764 11132
rect 28460 11064 28488 11104
rect 25240 11036 27614 11064
rect 27816 11036 27936 11064
rect 28000 11036 28488 11064
rect 29288 11064 29316 11172
rect 29917 11169 29929 11203
rect 29963 11200 29975 11203
rect 30193 11203 30251 11209
rect 30193 11200 30205 11203
rect 29963 11172 30205 11200
rect 29963 11169 29975 11172
rect 29917 11163 29975 11169
rect 30193 11169 30205 11172
rect 30239 11169 30251 11203
rect 30193 11163 30251 11169
rect 29730 11092 29736 11144
rect 29788 11092 29794 11144
rect 29822 11092 29828 11144
rect 29880 11092 29886 11144
rect 30009 11135 30067 11141
rect 30009 11101 30021 11135
rect 30055 11132 30067 11135
rect 30300 11132 30328 11240
rect 30558 11228 30564 11240
rect 30616 11228 30622 11280
rect 30374 11160 30380 11212
rect 30432 11160 30438 11212
rect 30742 11200 30748 11212
rect 30484 11172 30748 11200
rect 30484 11141 30512 11172
rect 30742 11160 30748 11172
rect 30800 11160 30806 11212
rect 30055 11104 30328 11132
rect 30469 11135 30527 11141
rect 30055 11101 30067 11104
rect 30009 11095 30067 11101
rect 30469 11101 30481 11135
rect 30515 11101 30527 11135
rect 30469 11095 30527 11101
rect 30561 11135 30619 11141
rect 30561 11101 30573 11135
rect 30607 11101 30619 11135
rect 30561 11095 30619 11101
rect 30653 11135 30711 11141
rect 30653 11101 30665 11135
rect 30699 11132 30711 11135
rect 30834 11132 30840 11144
rect 30699 11104 30840 11132
rect 30699 11101 30711 11104
rect 30653 11095 30711 11101
rect 30484 11064 30512 11095
rect 29288 11036 30512 11064
rect 25041 11027 25099 11033
rect 24946 10996 24952 11008
rect 21468 10968 24952 10996
rect 24946 10956 24952 10968
rect 25004 10956 25010 11008
rect 25056 10996 25084 11027
rect 25682 10996 25688 11008
rect 25056 10968 25688 10996
rect 25682 10956 25688 10968
rect 25740 10956 25746 11008
rect 26418 10956 26424 11008
rect 26476 10996 26482 11008
rect 27816 10996 27844 11036
rect 26476 10968 27844 10996
rect 27893 10999 27951 11005
rect 26476 10956 26482 10968
rect 27893 10965 27905 10999
rect 27939 10996 27951 10999
rect 28000 10996 28028 11036
rect 27939 10968 28028 10996
rect 27939 10965 27951 10968
rect 27893 10959 27951 10965
rect 28166 10956 28172 11008
rect 28224 10996 28230 11008
rect 30576 10996 30604 11095
rect 30834 11092 30840 11104
rect 30892 11132 30898 11144
rect 31110 11132 31116 11144
rect 30892 11104 31116 11132
rect 30892 11092 30898 11104
rect 31110 11092 31116 11104
rect 31168 11092 31174 11144
rect 32490 10996 32496 11008
rect 28224 10968 32496 10996
rect 28224 10956 28230 10968
rect 32490 10956 32496 10968
rect 32548 10956 32554 11008
rect 1104 10906 38272 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 38272 10906
rect 1104 10832 38272 10854
rect 5261 10795 5319 10801
rect 5261 10761 5273 10795
rect 5307 10761 5319 10795
rect 5261 10755 5319 10761
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10656 5135 10659
rect 5276 10656 5304 10755
rect 7374 10752 7380 10804
rect 7432 10792 7438 10804
rect 7561 10795 7619 10801
rect 7561 10792 7573 10795
rect 7432 10764 7573 10792
rect 7432 10752 7438 10764
rect 7561 10761 7573 10764
rect 7607 10761 7619 10795
rect 7561 10755 7619 10761
rect 8021 10795 8079 10801
rect 8021 10761 8033 10795
rect 8067 10792 8079 10795
rect 8478 10792 8484 10804
rect 8067 10764 8484 10792
rect 8067 10761 8079 10764
rect 8021 10755 8079 10761
rect 8478 10752 8484 10764
rect 8536 10752 8542 10804
rect 8570 10752 8576 10804
rect 8628 10792 8634 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 8628 10764 8953 10792
rect 8628 10752 8634 10764
rect 8941 10761 8953 10764
rect 8987 10761 8999 10795
rect 8941 10755 8999 10761
rect 11790 10752 11796 10804
rect 11848 10752 11854 10804
rect 12158 10752 12164 10804
rect 12216 10792 12222 10804
rect 12253 10795 12311 10801
rect 12253 10792 12265 10795
rect 12216 10764 12265 10792
rect 12216 10752 12222 10764
rect 12253 10761 12265 10764
rect 12299 10761 12311 10795
rect 12802 10792 12808 10804
rect 12253 10755 12311 10761
rect 12452 10764 12808 10792
rect 6914 10684 6920 10736
rect 6972 10724 6978 10736
rect 11146 10724 11152 10736
rect 6972 10696 11152 10724
rect 6972 10684 6978 10696
rect 5123 10628 5304 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 5626 10616 5632 10668
rect 5684 10616 5690 10668
rect 5721 10659 5779 10665
rect 5721 10625 5733 10659
rect 5767 10656 5779 10659
rect 7929 10659 7987 10665
rect 7929 10656 7941 10659
rect 5767 10628 7941 10656
rect 5767 10625 5779 10628
rect 5721 10619 5779 10625
rect 7929 10625 7941 10628
rect 7975 10656 7987 10659
rect 8662 10656 8668 10668
rect 7975 10628 8668 10656
rect 7975 10625 7987 10628
rect 7929 10619 7987 10625
rect 8662 10616 8668 10628
rect 8720 10616 8726 10668
rect 9968 10665 9996 10696
rect 11146 10684 11152 10696
rect 11204 10684 11210 10736
rect 11606 10684 11612 10736
rect 11664 10724 11670 10736
rect 11808 10724 11836 10752
rect 12342 10724 12348 10736
rect 11664 10696 11744 10724
rect 11664 10684 11670 10696
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10625 9367 10659
rect 9309 10619 9367 10625
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10656 10011 10659
rect 9999 10628 10033 10656
rect 9999 10625 10011 10628
rect 9953 10619 10011 10625
rect 5644 10588 5672 10616
rect 5905 10591 5963 10597
rect 5644 10560 5764 10588
rect 4706 10412 4712 10464
rect 4764 10452 4770 10464
rect 4893 10455 4951 10461
rect 4893 10452 4905 10455
rect 4764 10424 4905 10452
rect 4764 10412 4770 10424
rect 4893 10421 4905 10424
rect 4939 10421 4951 10455
rect 5736 10452 5764 10560
rect 5905 10557 5917 10591
rect 5951 10557 5963 10591
rect 5905 10551 5963 10557
rect 5810 10480 5816 10532
rect 5868 10520 5874 10532
rect 5920 10520 5948 10551
rect 6638 10548 6644 10600
rect 6696 10588 6702 10600
rect 8113 10591 8171 10597
rect 8113 10588 8125 10591
rect 6696 10560 8125 10588
rect 6696 10548 6702 10560
rect 8113 10557 8125 10560
rect 8159 10557 8171 10591
rect 8680 10588 8708 10616
rect 9324 10588 9352 10619
rect 11514 10616 11520 10668
rect 11572 10616 11578 10668
rect 11716 10665 11744 10696
rect 11808 10696 12348 10724
rect 11808 10665 11836 10696
rect 12342 10684 12348 10696
rect 12400 10684 12406 10736
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 11793 10659 11851 10665
rect 11793 10625 11805 10659
rect 11839 10625 11851 10659
rect 11793 10619 11851 10625
rect 8680 10560 9352 10588
rect 8113 10551 8171 10557
rect 9398 10548 9404 10600
rect 9456 10548 9462 10600
rect 9490 10548 9496 10600
rect 9548 10548 9554 10600
rect 9858 10548 9864 10600
rect 9916 10548 9922 10600
rect 11238 10548 11244 10600
rect 11296 10588 11302 10600
rect 11808 10588 11836 10619
rect 11882 10616 11888 10668
rect 11940 10616 11946 10668
rect 12452 10665 12480 10764
rect 12802 10752 12808 10764
rect 12860 10792 12866 10804
rect 14090 10792 14096 10804
rect 12860 10764 14096 10792
rect 12860 10752 12866 10764
rect 14090 10752 14096 10764
rect 14148 10752 14154 10804
rect 14182 10752 14188 10804
rect 14240 10792 14246 10804
rect 14369 10795 14427 10801
rect 14369 10792 14381 10795
rect 14240 10764 14381 10792
rect 14240 10752 14246 10764
rect 14369 10761 14381 10764
rect 14415 10761 14427 10795
rect 15470 10792 15476 10804
rect 14369 10755 14427 10761
rect 14476 10764 15476 10792
rect 12529 10727 12587 10733
rect 12529 10693 12541 10727
rect 12575 10724 12587 10727
rect 12894 10724 12900 10736
rect 12575 10696 12900 10724
rect 12575 10693 12587 10696
rect 12529 10687 12587 10693
rect 12894 10684 12900 10696
rect 12952 10724 12958 10736
rect 14476 10724 14504 10764
rect 15470 10752 15476 10764
rect 15528 10792 15534 10804
rect 15657 10795 15715 10801
rect 15528 10764 15608 10792
rect 15528 10752 15534 10764
rect 12952 10696 14504 10724
rect 15381 10727 15439 10733
rect 12952 10684 12958 10696
rect 15381 10693 15393 10727
rect 15427 10724 15439 10727
rect 15580 10724 15608 10764
rect 15657 10761 15669 10795
rect 15703 10792 15715 10795
rect 16301 10795 16359 10801
rect 15703 10764 16160 10792
rect 15703 10761 15715 10764
rect 15657 10755 15715 10761
rect 15427 10696 15608 10724
rect 16132 10724 16160 10764
rect 16301 10761 16313 10795
rect 16347 10792 16359 10795
rect 17034 10792 17040 10804
rect 16347 10764 17040 10792
rect 16347 10761 16359 10764
rect 16301 10755 16359 10761
rect 17034 10752 17040 10764
rect 17092 10752 17098 10804
rect 17126 10752 17132 10804
rect 17184 10792 17190 10804
rect 17310 10792 17316 10804
rect 17184 10764 17316 10792
rect 17184 10752 17190 10764
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 17402 10752 17408 10804
rect 17460 10752 17466 10804
rect 17589 10795 17647 10801
rect 17589 10761 17601 10795
rect 17635 10761 17647 10795
rect 17589 10755 17647 10761
rect 18325 10795 18383 10801
rect 18325 10761 18337 10795
rect 18371 10792 18383 10795
rect 18414 10792 18420 10804
rect 18371 10764 18420 10792
rect 18371 10761 18383 10764
rect 18325 10755 18383 10761
rect 16758 10724 16764 10736
rect 16132 10696 16764 10724
rect 15427 10693 15439 10696
rect 15381 10687 15439 10693
rect 16758 10684 16764 10696
rect 16816 10684 16822 10736
rect 17218 10684 17224 10736
rect 17276 10684 17282 10736
rect 17420 10724 17448 10752
rect 17604 10724 17632 10755
rect 18414 10752 18420 10764
rect 18472 10752 18478 10804
rect 18598 10752 18604 10804
rect 18656 10752 18662 10804
rect 18874 10752 18880 10804
rect 18932 10792 18938 10804
rect 20530 10792 20536 10804
rect 18932 10764 20536 10792
rect 18932 10752 18938 10764
rect 20530 10752 20536 10764
rect 20588 10752 20594 10804
rect 20898 10752 20904 10804
rect 20956 10752 20962 10804
rect 22005 10795 22063 10801
rect 22005 10792 22017 10795
rect 21008 10764 22017 10792
rect 18616 10724 18644 10752
rect 20806 10724 20812 10736
rect 17420 10696 17540 10724
rect 17604 10696 18644 10724
rect 18984 10696 20812 10724
rect 12437 10659 12495 10665
rect 12437 10625 12449 10659
rect 12483 10625 12495 10659
rect 12437 10619 12495 10625
rect 12618 10616 12624 10668
rect 12676 10616 12682 10668
rect 12805 10659 12863 10665
rect 12805 10625 12817 10659
rect 12851 10656 12863 10659
rect 13909 10659 13967 10665
rect 12851 10628 13860 10656
rect 12851 10625 12863 10628
rect 12805 10619 12863 10625
rect 12820 10588 12848 10619
rect 11296 10560 11836 10588
rect 12268 10560 12848 10588
rect 11296 10548 11302 10560
rect 6822 10520 6828 10532
rect 5868 10492 6828 10520
rect 5868 10480 5874 10492
rect 6822 10480 6828 10492
rect 6880 10480 6886 10532
rect 8202 10480 8208 10532
rect 8260 10520 8266 10532
rect 12268 10520 12296 10560
rect 13630 10548 13636 10600
rect 13688 10548 13694 10600
rect 8260 10492 12296 10520
rect 8260 10480 8266 10492
rect 12342 10480 12348 10532
rect 12400 10520 12406 10532
rect 13078 10520 13084 10532
rect 12400 10492 13084 10520
rect 12400 10480 12406 10492
rect 13078 10480 13084 10492
rect 13136 10480 13142 10532
rect 6362 10452 6368 10464
rect 5736 10424 6368 10452
rect 4893 10415 4951 10421
rect 6362 10412 6368 10424
rect 6420 10452 6426 10464
rect 11606 10452 11612 10464
rect 6420 10424 11612 10452
rect 6420 10412 6426 10424
rect 11606 10412 11612 10424
rect 11664 10412 11670 10464
rect 11790 10412 11796 10464
rect 11848 10452 11854 10464
rect 12161 10455 12219 10461
rect 12161 10452 12173 10455
rect 11848 10424 12173 10452
rect 11848 10412 11854 10424
rect 12161 10421 12173 10424
rect 12207 10421 12219 10455
rect 13648 10452 13676 10548
rect 13832 10520 13860 10628
rect 13909 10625 13921 10659
rect 13955 10656 13967 10659
rect 13998 10656 14004 10668
rect 13955 10628 14004 10656
rect 13955 10625 13967 10628
rect 13909 10619 13967 10625
rect 13998 10616 14004 10628
rect 14056 10616 14062 10668
rect 14185 10659 14243 10665
rect 14185 10625 14197 10659
rect 14231 10656 14243 10659
rect 14366 10656 14372 10668
rect 14231 10628 14372 10656
rect 14231 10625 14243 10628
rect 14185 10619 14243 10625
rect 14366 10616 14372 10628
rect 14424 10616 14430 10668
rect 14550 10616 14556 10668
rect 14608 10656 14614 10668
rect 15105 10659 15163 10665
rect 15105 10656 15117 10659
rect 14608 10628 15117 10656
rect 14608 10616 14614 10628
rect 15105 10625 15117 10628
rect 15151 10625 15163 10659
rect 15105 10619 15163 10625
rect 15194 10616 15200 10668
rect 15252 10659 15258 10668
rect 15562 10665 15568 10668
rect 15289 10659 15347 10665
rect 15252 10631 15301 10659
rect 15252 10616 15258 10631
rect 15289 10625 15301 10631
rect 15335 10625 15347 10659
rect 15289 10619 15347 10625
rect 15519 10659 15568 10665
rect 15519 10625 15531 10659
rect 15565 10625 15568 10659
rect 15519 10619 15568 10625
rect 15562 10616 15568 10619
rect 15620 10616 15626 10668
rect 15749 10659 15807 10665
rect 15749 10656 15761 10659
rect 15672 10628 15761 10656
rect 14090 10548 14096 10600
rect 14148 10588 14154 10600
rect 14458 10588 14464 10600
rect 14148 10560 14464 10588
rect 14148 10548 14154 10560
rect 14458 10548 14464 10560
rect 14516 10548 14522 10600
rect 15672 10520 15700 10628
rect 15749 10625 15761 10628
rect 15795 10625 15807 10659
rect 15749 10619 15807 10625
rect 15930 10616 15936 10668
rect 15988 10616 15994 10668
rect 16025 10659 16083 10665
rect 16025 10625 16037 10659
rect 16071 10625 16083 10659
rect 16025 10619 16083 10625
rect 16040 10588 16068 10619
rect 16114 10616 16120 10668
rect 16172 10616 16178 10668
rect 16206 10616 16212 10668
rect 16264 10656 16270 10668
rect 17034 10656 17040 10668
rect 16264 10628 17040 10656
rect 16264 10616 16270 10628
rect 17034 10616 17040 10628
rect 17092 10616 17098 10668
rect 16224 10588 16252 10616
rect 16040 10560 16252 10588
rect 16850 10548 16856 10600
rect 16908 10588 16914 10600
rect 17236 10588 17264 10684
rect 17310 10616 17316 10668
rect 17368 10616 17374 10668
rect 17402 10616 17408 10668
rect 17460 10616 17466 10668
rect 17512 10656 17540 10696
rect 17681 10659 17739 10665
rect 17681 10656 17693 10659
rect 17512 10628 17693 10656
rect 17681 10625 17693 10628
rect 17727 10625 17739 10659
rect 17681 10619 17739 10625
rect 17865 10659 17923 10665
rect 17865 10625 17877 10659
rect 17911 10625 17923 10659
rect 17865 10619 17923 10625
rect 17880 10588 17908 10619
rect 17954 10616 17960 10668
rect 18012 10616 18018 10668
rect 18049 10659 18107 10665
rect 18049 10625 18061 10659
rect 18095 10656 18107 10659
rect 18138 10656 18144 10668
rect 18095 10628 18144 10656
rect 18095 10625 18107 10628
rect 18049 10619 18107 10625
rect 18138 10616 18144 10628
rect 18196 10616 18202 10668
rect 18506 10616 18512 10668
rect 18564 10616 18570 10668
rect 18598 10616 18604 10668
rect 18656 10656 18662 10668
rect 18984 10665 19012 10696
rect 20806 10684 20812 10696
rect 20864 10684 20870 10736
rect 21008 10724 21036 10764
rect 22005 10761 22017 10764
rect 22051 10792 22063 10795
rect 22738 10792 22744 10804
rect 22051 10764 22744 10792
rect 22051 10761 22063 10764
rect 22005 10755 22063 10761
rect 22738 10752 22744 10764
rect 22796 10752 22802 10804
rect 22922 10752 22928 10804
rect 22980 10752 22986 10804
rect 23290 10752 23296 10804
rect 23348 10752 23354 10804
rect 24486 10752 24492 10804
rect 24544 10792 24550 10804
rect 25406 10792 25412 10804
rect 24544 10764 25412 10792
rect 24544 10752 24550 10764
rect 25406 10752 25412 10764
rect 25464 10752 25470 10804
rect 26237 10795 26295 10801
rect 25701 10764 26197 10792
rect 20916 10696 21036 10724
rect 21192 10696 21496 10724
rect 18969 10659 19027 10665
rect 18969 10656 18981 10659
rect 18656 10628 18981 10656
rect 18656 10616 18662 10628
rect 18969 10625 18981 10628
rect 19015 10625 19027 10659
rect 18969 10619 19027 10625
rect 19058 10616 19064 10668
rect 19116 10616 19122 10668
rect 19242 10616 19248 10668
rect 19300 10616 19306 10668
rect 20714 10616 20720 10668
rect 20772 10656 20778 10668
rect 20916 10656 20944 10696
rect 20772 10628 20944 10656
rect 20772 10616 20778 10628
rect 21082 10616 21088 10668
rect 21140 10616 21146 10668
rect 18693 10591 18751 10597
rect 18693 10588 18705 10591
rect 16908 10560 17264 10588
rect 17328 10560 17908 10588
rect 18248 10560 18705 10588
rect 16908 10548 16914 10560
rect 13832 10492 15700 10520
rect 14001 10455 14059 10461
rect 14001 10452 14013 10455
rect 13648 10424 14013 10452
rect 12161 10415 12219 10421
rect 14001 10421 14013 10424
rect 14047 10452 14059 10455
rect 14182 10452 14188 10464
rect 14047 10424 14188 10452
rect 14047 10421 14059 10424
rect 14001 10415 14059 10421
rect 14182 10412 14188 10424
rect 14240 10412 14246 10464
rect 15672 10452 15700 10492
rect 17218 10480 17224 10532
rect 17276 10520 17282 10532
rect 17328 10520 17356 10560
rect 17276 10492 17356 10520
rect 17276 10480 17282 10492
rect 17586 10480 17592 10532
rect 17644 10520 17650 10532
rect 17954 10520 17960 10532
rect 17644 10492 17960 10520
rect 17644 10480 17650 10492
rect 17954 10480 17960 10492
rect 18012 10480 18018 10532
rect 18248 10529 18276 10560
rect 18693 10557 18705 10560
rect 18739 10557 18751 10591
rect 18693 10551 18751 10557
rect 18785 10591 18843 10597
rect 18785 10557 18797 10591
rect 18831 10588 18843 10591
rect 18874 10588 18880 10600
rect 18831 10560 18880 10588
rect 18831 10557 18843 10560
rect 18785 10551 18843 10557
rect 18874 10548 18880 10560
rect 18932 10548 18938 10600
rect 19260 10588 19288 10616
rect 19168 10560 19288 10588
rect 18233 10523 18291 10529
rect 18233 10489 18245 10523
rect 18279 10489 18291 10523
rect 18233 10483 18291 10489
rect 18601 10523 18659 10529
rect 18601 10489 18613 10523
rect 18647 10520 18659 10523
rect 19168 10520 19196 10560
rect 19518 10548 19524 10600
rect 19576 10588 19582 10600
rect 20809 10591 20867 10597
rect 20809 10588 20821 10591
rect 19576 10560 20821 10588
rect 19576 10548 19582 10560
rect 20809 10557 20821 10560
rect 20855 10588 20867 10591
rect 21192 10588 21220 10696
rect 21269 10659 21327 10665
rect 21269 10625 21281 10659
rect 21315 10625 21327 10659
rect 21269 10619 21327 10625
rect 20855 10560 21220 10588
rect 20855 10557 20867 10560
rect 20809 10551 20867 10557
rect 18647 10492 19196 10520
rect 19306 10492 20479 10520
rect 18647 10489 18659 10492
rect 18601 10483 18659 10489
rect 16574 10452 16580 10464
rect 15672 10424 16580 10452
rect 16574 10412 16580 10424
rect 16632 10452 16638 10464
rect 17770 10452 17776 10464
rect 16632 10424 17776 10452
rect 16632 10412 16638 10424
rect 17770 10412 17776 10424
rect 17828 10412 17834 10464
rect 17972 10452 18000 10480
rect 19306 10452 19334 10492
rect 17972 10424 19334 10452
rect 20451 10452 20479 10492
rect 20530 10480 20536 10532
rect 20588 10520 20594 10532
rect 21284 10520 21312 10619
rect 21358 10616 21364 10668
rect 21416 10616 21422 10668
rect 21468 10588 21496 10696
rect 21542 10684 21548 10736
rect 21600 10724 21606 10736
rect 21821 10727 21879 10733
rect 21821 10724 21833 10727
rect 21600 10696 21833 10724
rect 21600 10684 21606 10696
rect 21821 10693 21833 10696
rect 21867 10693 21879 10727
rect 21821 10687 21879 10693
rect 22462 10684 22468 10736
rect 22520 10724 22526 10736
rect 22940 10724 22968 10752
rect 22520 10696 22784 10724
rect 22940 10696 23152 10724
rect 22520 10684 22526 10696
rect 21726 10616 21732 10668
rect 21784 10656 21790 10668
rect 22756 10665 22784 10696
rect 22281 10659 22339 10665
rect 22281 10656 22293 10659
rect 21784 10628 22293 10656
rect 21784 10616 21790 10628
rect 22281 10625 22293 10628
rect 22327 10625 22339 10659
rect 22281 10619 22339 10625
rect 22741 10659 22799 10665
rect 22741 10625 22753 10659
rect 22787 10625 22799 10659
rect 22741 10619 22799 10625
rect 22830 10616 22836 10668
rect 22888 10616 22894 10668
rect 22922 10616 22928 10668
rect 22980 10656 22986 10668
rect 23124 10665 23152 10696
rect 25701 10668 25729 10764
rect 25869 10727 25927 10733
rect 25869 10693 25881 10727
rect 25915 10693 25927 10727
rect 26169 10724 26197 10764
rect 26237 10761 26249 10795
rect 26283 10792 26295 10795
rect 26602 10792 26608 10804
rect 26283 10764 26608 10792
rect 26283 10761 26295 10764
rect 26237 10755 26295 10761
rect 26602 10752 26608 10764
rect 26660 10752 26666 10804
rect 27709 10795 27767 10801
rect 27709 10761 27721 10795
rect 27755 10792 27767 10795
rect 27798 10792 27804 10804
rect 27755 10764 27804 10792
rect 27755 10761 27767 10764
rect 27709 10755 27767 10761
rect 27798 10752 27804 10764
rect 27856 10752 27862 10804
rect 29178 10752 29184 10804
rect 29236 10792 29242 10804
rect 29236 10764 29500 10792
rect 29236 10752 29242 10764
rect 27433 10727 27491 10733
rect 27433 10724 27445 10727
rect 26169 10696 27445 10724
rect 25869 10687 25927 10693
rect 27433 10693 27445 10696
rect 27479 10724 27491 10727
rect 28166 10724 28172 10736
rect 27479 10696 28172 10724
rect 27479 10693 27491 10696
rect 27433 10687 27491 10693
rect 23017 10659 23075 10665
rect 23017 10656 23029 10659
rect 22980 10628 23029 10656
rect 22980 10616 22986 10628
rect 23017 10625 23029 10628
rect 23063 10625 23075 10659
rect 23017 10619 23075 10625
rect 23109 10659 23167 10665
rect 23109 10625 23121 10659
rect 23155 10625 23167 10659
rect 23109 10619 23167 10625
rect 23385 10659 23443 10665
rect 23385 10625 23397 10659
rect 23431 10625 23443 10659
rect 23385 10619 23443 10625
rect 23400 10588 23428 10619
rect 25222 10616 25228 10668
rect 25280 10656 25286 10668
rect 25593 10659 25651 10665
rect 25593 10656 25605 10659
rect 25280 10628 25605 10656
rect 25280 10616 25286 10628
rect 25593 10625 25605 10628
rect 25639 10625 25651 10659
rect 25593 10619 25651 10625
rect 25682 10616 25688 10668
rect 25740 10656 25746 10668
rect 25740 10628 25785 10656
rect 25740 10616 25746 10628
rect 21468 10560 23428 10588
rect 23474 10548 23480 10600
rect 23532 10588 23538 10600
rect 24118 10588 24124 10600
rect 23532 10560 24124 10588
rect 23532 10548 23538 10560
rect 24118 10548 24124 10560
rect 24176 10548 24182 10600
rect 24762 10548 24768 10600
rect 24820 10588 24826 10600
rect 25133 10591 25191 10597
rect 25133 10588 25145 10591
rect 24820 10560 25145 10588
rect 24820 10548 24826 10560
rect 25133 10557 25145 10560
rect 25179 10588 25191 10591
rect 25179 10560 25452 10588
rect 25179 10557 25191 10560
rect 25133 10551 25191 10557
rect 25424 10532 25452 10560
rect 25498 10548 25504 10600
rect 25556 10588 25562 10600
rect 25884 10588 25912 10687
rect 28166 10684 28172 10696
rect 28224 10684 28230 10736
rect 28810 10684 28816 10736
rect 28868 10684 28874 10736
rect 29472 10733 29500 10764
rect 29822 10752 29828 10804
rect 29880 10752 29886 10804
rect 31018 10752 31024 10804
rect 31076 10792 31082 10804
rect 31570 10792 31576 10804
rect 31076 10764 31576 10792
rect 31076 10752 31082 10764
rect 31570 10752 31576 10764
rect 31628 10752 31634 10804
rect 32125 10795 32183 10801
rect 32125 10761 32137 10795
rect 32171 10761 32183 10795
rect 32125 10755 32183 10761
rect 33873 10795 33931 10801
rect 33873 10761 33885 10795
rect 33919 10761 33931 10795
rect 33873 10755 33931 10761
rect 29457 10727 29515 10733
rect 29457 10693 29469 10727
rect 29503 10724 29515 10727
rect 29503 10696 30052 10724
rect 29503 10693 29515 10696
rect 29457 10687 29515 10693
rect 30024 10668 30052 10696
rect 25958 10616 25964 10668
rect 26016 10616 26022 10668
rect 26142 10665 26148 10668
rect 26099 10659 26148 10665
rect 26099 10625 26111 10659
rect 26145 10625 26148 10659
rect 26099 10619 26148 10625
rect 26142 10616 26148 10619
rect 26200 10616 26206 10668
rect 27249 10659 27307 10665
rect 27249 10625 27261 10659
rect 27295 10656 27307 10659
rect 27706 10656 27712 10668
rect 27295 10628 27712 10656
rect 27295 10625 27307 10628
rect 27249 10619 27307 10625
rect 27706 10616 27712 10628
rect 27764 10616 27770 10668
rect 28350 10665 28356 10668
rect 28307 10659 28356 10665
rect 28307 10625 28319 10659
rect 28353 10625 28356 10659
rect 28307 10619 28356 10625
rect 28350 10616 28356 10619
rect 28408 10616 28414 10668
rect 28718 10665 28724 10668
rect 28445 10662 28503 10665
rect 28445 10659 28580 10662
rect 28445 10625 28457 10659
rect 28491 10634 28580 10659
rect 28491 10625 28503 10634
rect 28445 10619 28503 10625
rect 28552 10600 28580 10634
rect 28675 10659 28724 10665
rect 28675 10625 28687 10659
rect 28721 10625 28724 10659
rect 28675 10619 28724 10625
rect 28718 10616 28724 10619
rect 28776 10616 28782 10668
rect 28905 10659 28963 10665
rect 28905 10625 28917 10659
rect 28951 10625 28963 10659
rect 28905 10619 28963 10625
rect 25556 10560 25912 10588
rect 25556 10548 25562 10560
rect 28074 10548 28080 10600
rect 28132 10548 28138 10600
rect 28534 10548 28540 10600
rect 28592 10548 28598 10600
rect 28920 10588 28948 10619
rect 28994 10616 29000 10668
rect 29052 10656 29058 10668
rect 29089 10659 29147 10665
rect 29089 10656 29101 10659
rect 29052 10628 29101 10656
rect 29052 10616 29058 10628
rect 29089 10625 29101 10628
rect 29135 10625 29147 10659
rect 29089 10619 29147 10625
rect 29273 10659 29331 10665
rect 29273 10625 29285 10659
rect 29319 10656 29331 10659
rect 29319 10628 29500 10656
rect 29319 10625 29331 10628
rect 29273 10619 29331 10625
rect 28920 10560 29316 10588
rect 24026 10520 24032 10532
rect 20588 10492 24032 10520
rect 20588 10480 20594 10492
rect 24026 10480 24032 10492
rect 24084 10480 24090 10532
rect 25406 10480 25412 10532
rect 25464 10480 25470 10532
rect 27985 10523 28043 10529
rect 27985 10489 27997 10523
rect 28031 10520 28043 10523
rect 28031 10492 28304 10520
rect 28031 10489 28043 10492
rect 27985 10483 28043 10489
rect 22005 10455 22063 10461
rect 22005 10452 22017 10455
rect 20451 10424 22017 10452
rect 22005 10421 22017 10424
rect 22051 10421 22063 10455
rect 22005 10415 22063 10421
rect 22462 10412 22468 10464
rect 22520 10452 22526 10464
rect 23198 10452 23204 10464
rect 22520 10424 23204 10452
rect 22520 10412 22526 10424
rect 23198 10412 23204 10424
rect 23256 10412 23262 10464
rect 25130 10412 25136 10464
rect 25188 10452 25194 10464
rect 26878 10452 26884 10464
rect 25188 10424 26884 10452
rect 25188 10412 25194 10424
rect 26878 10412 26884 10424
rect 26936 10412 26942 10464
rect 27617 10455 27675 10461
rect 27617 10421 27629 10455
rect 27663 10452 27675 10455
rect 27890 10452 27896 10464
rect 27663 10424 27896 10452
rect 27663 10421 27675 10424
rect 27617 10415 27675 10421
rect 27890 10412 27896 10424
rect 27948 10412 27954 10464
rect 28166 10412 28172 10464
rect 28224 10412 28230 10464
rect 28276 10452 28304 10492
rect 28537 10455 28595 10461
rect 28537 10452 28549 10455
rect 28276 10424 28549 10452
rect 28537 10421 28549 10424
rect 28583 10421 28595 10455
rect 28537 10415 28595 10421
rect 28626 10412 28632 10464
rect 28684 10452 28690 10464
rect 29288 10452 29316 10560
rect 29472 10532 29500 10628
rect 29546 10616 29552 10668
rect 29604 10616 29610 10668
rect 29638 10616 29644 10668
rect 29696 10616 29702 10668
rect 30006 10616 30012 10668
rect 30064 10616 30070 10668
rect 31389 10659 31447 10665
rect 31389 10625 31401 10659
rect 31435 10656 31447 10659
rect 32140 10656 32168 10755
rect 32582 10684 32588 10736
rect 32640 10724 32646 10736
rect 33505 10727 33563 10733
rect 33505 10724 33517 10727
rect 32640 10696 33517 10724
rect 32640 10684 32646 10696
rect 33505 10693 33517 10696
rect 33551 10693 33563 10727
rect 33505 10687 33563 10693
rect 31435 10628 32168 10656
rect 31435 10625 31447 10628
rect 31389 10619 31447 10625
rect 32490 10616 32496 10668
rect 32548 10616 32554 10668
rect 33888 10656 33916 10755
rect 33965 10659 34023 10665
rect 33965 10656 33977 10659
rect 33888 10628 33977 10656
rect 33965 10625 33977 10628
rect 34011 10625 34023 10659
rect 33965 10619 34023 10625
rect 32582 10548 32588 10600
rect 32640 10548 32646 10600
rect 32674 10548 32680 10600
rect 32732 10548 32738 10600
rect 33226 10548 33232 10600
rect 33284 10548 33290 10600
rect 33318 10548 33324 10600
rect 33376 10588 33382 10600
rect 33413 10591 33471 10597
rect 33413 10588 33425 10591
rect 33376 10560 33425 10588
rect 33376 10548 33382 10560
rect 33413 10557 33425 10560
rect 33459 10557 33471 10591
rect 33413 10551 33471 10557
rect 29454 10480 29460 10532
rect 29512 10520 29518 10532
rect 33336 10520 33364 10548
rect 29512 10492 33364 10520
rect 29512 10480 29518 10492
rect 28684 10424 29316 10452
rect 31205 10455 31263 10461
rect 28684 10412 28690 10424
rect 31205 10421 31217 10455
rect 31251 10452 31263 10455
rect 31294 10452 31300 10464
rect 31251 10424 31300 10452
rect 31251 10421 31263 10424
rect 31205 10415 31263 10421
rect 31294 10412 31300 10424
rect 31352 10412 31358 10464
rect 34149 10455 34207 10461
rect 34149 10421 34161 10455
rect 34195 10452 34207 10455
rect 34514 10452 34520 10464
rect 34195 10424 34520 10452
rect 34195 10421 34207 10424
rect 34149 10415 34207 10421
rect 34514 10412 34520 10424
rect 34572 10412 34578 10464
rect 1104 10362 38272 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38272 10362
rect 1104 10288 38272 10310
rect 4604 10251 4662 10257
rect 4604 10217 4616 10251
rect 4650 10248 4662 10251
rect 4706 10248 4712 10260
rect 4650 10220 4712 10248
rect 4650 10217 4662 10220
rect 4604 10211 4662 10217
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 8662 10248 8668 10260
rect 7760 10220 8668 10248
rect 3970 10072 3976 10124
rect 4028 10112 4034 10124
rect 4614 10112 4620 10124
rect 4028 10084 4620 10112
rect 4028 10072 4034 10084
rect 4080 10053 4108 10084
rect 4614 10072 4620 10084
rect 4672 10072 4678 10124
rect 6362 10072 6368 10124
rect 6420 10072 6426 10124
rect 6730 10072 6736 10124
rect 6788 10072 6794 10124
rect 7760 10121 7788 10220
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 9398 10208 9404 10260
rect 9456 10248 9462 10260
rect 10689 10251 10747 10257
rect 10689 10248 10701 10251
rect 9456 10220 10701 10248
rect 9456 10208 9462 10220
rect 10689 10217 10701 10220
rect 10735 10248 10747 10251
rect 12894 10248 12900 10260
rect 10735 10220 12900 10248
rect 10735 10217 10747 10220
rect 10689 10211 10747 10217
rect 12894 10208 12900 10220
rect 12952 10208 12958 10260
rect 13078 10208 13084 10260
rect 13136 10248 13142 10260
rect 15194 10248 15200 10260
rect 13136 10220 15200 10248
rect 13136 10208 13142 10220
rect 15194 10208 15200 10220
rect 15252 10208 15258 10260
rect 15378 10208 15384 10260
rect 15436 10208 15442 10260
rect 15746 10208 15752 10260
rect 15804 10248 15810 10260
rect 15933 10251 15991 10257
rect 15933 10248 15945 10251
rect 15804 10220 15945 10248
rect 15804 10208 15810 10220
rect 15933 10217 15945 10220
rect 15979 10217 15991 10251
rect 15933 10211 15991 10217
rect 18138 10208 18144 10260
rect 18196 10248 18202 10260
rect 19334 10248 19340 10260
rect 18196 10220 19340 10248
rect 18196 10208 18202 10220
rect 19334 10208 19340 10220
rect 19392 10208 19398 10260
rect 20625 10251 20683 10257
rect 20625 10217 20637 10251
rect 20671 10248 20683 10251
rect 21082 10248 21088 10260
rect 20671 10220 21088 10248
rect 20671 10217 20683 10220
rect 20625 10211 20683 10217
rect 21082 10208 21088 10220
rect 21140 10208 21146 10260
rect 22094 10208 22100 10260
rect 22152 10208 22158 10260
rect 22830 10208 22836 10260
rect 22888 10248 22894 10260
rect 23569 10251 23627 10257
rect 23569 10248 23581 10251
rect 22888 10220 23581 10248
rect 22888 10208 22894 10220
rect 23569 10217 23581 10220
rect 23615 10217 23627 10251
rect 23569 10211 23627 10217
rect 23842 10208 23848 10260
rect 23900 10248 23906 10260
rect 24118 10248 24124 10260
rect 23900 10220 24124 10248
rect 23900 10208 23906 10220
rect 24118 10208 24124 10220
rect 24176 10208 24182 10260
rect 25593 10251 25651 10257
rect 25593 10217 25605 10251
rect 25639 10248 25651 10251
rect 25866 10248 25872 10260
rect 25639 10220 25872 10248
rect 25639 10217 25651 10220
rect 25593 10211 25651 10217
rect 25866 10208 25872 10220
rect 25924 10208 25930 10260
rect 28074 10208 28080 10260
rect 28132 10248 28138 10260
rect 28445 10251 28503 10257
rect 28445 10248 28457 10251
rect 28132 10220 28457 10248
rect 28132 10208 28138 10220
rect 28445 10217 28457 10220
rect 28491 10217 28503 10251
rect 28445 10211 28503 10217
rect 28534 10208 28540 10260
rect 28592 10248 28598 10260
rect 28813 10251 28871 10257
rect 28813 10248 28825 10251
rect 28592 10220 28825 10248
rect 28592 10208 28598 10220
rect 28813 10217 28825 10220
rect 28859 10217 28871 10251
rect 28813 10211 28871 10217
rect 28997 10251 29055 10257
rect 28997 10217 29009 10251
rect 29043 10248 29055 10251
rect 29730 10248 29736 10260
rect 29043 10220 29736 10248
rect 29043 10217 29055 10220
rect 28997 10211 29055 10217
rect 29730 10208 29736 10220
rect 29788 10208 29794 10260
rect 32490 10208 32496 10260
rect 32548 10248 32554 10260
rect 32769 10251 32827 10257
rect 32769 10248 32781 10251
rect 32548 10220 32781 10248
rect 32548 10208 32554 10220
rect 32769 10217 32781 10220
rect 32815 10217 32827 10251
rect 32769 10211 32827 10217
rect 11606 10140 11612 10192
rect 11664 10180 11670 10192
rect 11882 10180 11888 10192
rect 11664 10152 11888 10180
rect 11664 10140 11670 10152
rect 11882 10140 11888 10152
rect 11940 10180 11946 10192
rect 16942 10180 16948 10192
rect 11940 10152 16948 10180
rect 11940 10140 11946 10152
rect 16942 10140 16948 10152
rect 17000 10140 17006 10192
rect 17034 10140 17040 10192
rect 17092 10180 17098 10192
rect 17497 10183 17555 10189
rect 17497 10180 17509 10183
rect 17092 10152 17509 10180
rect 17092 10140 17098 10152
rect 17497 10149 17509 10152
rect 17543 10149 17555 10183
rect 17497 10143 17555 10149
rect 17954 10140 17960 10192
rect 18012 10140 18018 10192
rect 21542 10180 21548 10192
rect 18432 10152 21548 10180
rect 7745 10115 7803 10121
rect 7745 10081 7757 10115
rect 7791 10081 7803 10115
rect 7745 10075 7803 10081
rect 7929 10115 7987 10121
rect 7929 10081 7941 10115
rect 7975 10112 7987 10115
rect 8110 10112 8116 10124
rect 7975 10084 8116 10112
rect 7975 10081 7987 10084
rect 7929 10075 7987 10081
rect 8110 10072 8116 10084
rect 8168 10072 8174 10124
rect 15746 10112 15752 10124
rect 8772 10084 12664 10112
rect 4065 10047 4123 10053
rect 4065 10013 4077 10047
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4341 10047 4399 10053
rect 4341 10044 4353 10047
rect 4203 10016 4353 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 4341 10013 4353 10016
rect 4387 10013 4399 10047
rect 4341 10007 4399 10013
rect 6641 10047 6699 10053
rect 6641 10013 6653 10047
rect 6687 10044 6699 10047
rect 6748 10044 6776 10072
rect 6687 10016 6776 10044
rect 7009 10047 7067 10053
rect 6687 10013 6699 10016
rect 6641 10007 6699 10013
rect 7009 10013 7021 10047
rect 7055 10044 7067 10047
rect 8297 10047 8355 10053
rect 7055 10016 7328 10044
rect 7055 10013 7067 10016
rect 7009 10007 7067 10013
rect 6178 9976 6184 9988
rect 5842 9948 6184 9976
rect 6178 9936 6184 9948
rect 6236 9936 6242 9988
rect 6546 9868 6552 9920
rect 6604 9868 6610 9920
rect 6822 9868 6828 9920
rect 6880 9868 6886 9920
rect 7300 9917 7328 10016
rect 8297 10013 8309 10047
rect 8343 10044 8355 10047
rect 8570 10044 8576 10056
rect 8343 10016 8576 10044
rect 8343 10013 8355 10016
rect 8297 10007 8355 10013
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 8772 10053 8800 10084
rect 12636 10056 12664 10084
rect 12912 10084 15752 10112
rect 8757 10047 8815 10053
rect 8757 10013 8769 10047
rect 8803 10013 8815 10047
rect 8757 10007 8815 10013
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 8665 9979 8723 9985
rect 8665 9945 8677 9979
rect 8711 9976 8723 9979
rect 8956 9976 8984 10007
rect 12618 10004 12624 10056
rect 12676 10044 12682 10056
rect 12912 10053 12940 10084
rect 15746 10072 15752 10084
rect 15804 10072 15810 10124
rect 17310 10112 17316 10124
rect 16960 10084 17316 10112
rect 16960 10056 16988 10084
rect 17310 10072 17316 10084
rect 17368 10072 17374 10124
rect 17972 10112 18000 10140
rect 17788 10084 18000 10112
rect 12897 10047 12955 10053
rect 12897 10044 12909 10047
rect 12676 10016 12909 10044
rect 12676 10004 12682 10016
rect 12897 10013 12909 10016
rect 12943 10013 12955 10047
rect 12897 10007 12955 10013
rect 13538 10004 13544 10056
rect 13596 10044 13602 10056
rect 14550 10044 14556 10056
rect 13596 10016 14556 10044
rect 13596 10004 13602 10016
rect 14550 10004 14556 10016
rect 14608 10044 14614 10056
rect 14734 10044 14740 10056
rect 14608 10016 14740 10044
rect 14608 10004 14614 10016
rect 14734 10004 14740 10016
rect 14792 10004 14798 10056
rect 15194 10004 15200 10056
rect 15252 10004 15258 10056
rect 15289 10047 15347 10053
rect 15289 10013 15301 10047
rect 15335 10013 15347 10047
rect 15289 10007 15347 10013
rect 8711 9948 8984 9976
rect 9217 9979 9275 9985
rect 8711 9945 8723 9948
rect 8665 9939 8723 9945
rect 9217 9945 9229 9979
rect 9263 9945 9275 9979
rect 10962 9976 10968 9988
rect 10442 9948 10968 9976
rect 9217 9939 9275 9945
rect 7285 9911 7343 9917
rect 7285 9877 7297 9911
rect 7331 9877 7343 9911
rect 7285 9871 7343 9877
rect 7653 9911 7711 9917
rect 7653 9877 7665 9911
rect 7699 9908 7711 9911
rect 8202 9908 8208 9920
rect 7699 9880 8208 9908
rect 7699 9877 7711 9880
rect 7653 9871 7711 9877
rect 8202 9868 8208 9880
rect 8260 9868 8266 9920
rect 8481 9911 8539 9917
rect 8481 9877 8493 9911
rect 8527 9908 8539 9911
rect 9232 9908 9260 9939
rect 10962 9936 10968 9948
rect 11020 9936 11026 9988
rect 11330 9936 11336 9988
rect 11388 9976 11394 9988
rect 11606 9976 11612 9988
rect 11388 9948 11612 9976
rect 11388 9936 11394 9948
rect 11606 9936 11612 9948
rect 11664 9936 11670 9988
rect 15304 9976 15332 10007
rect 16942 10004 16948 10056
rect 17000 10004 17006 10056
rect 17402 10004 17408 10056
rect 17460 10004 17466 10056
rect 17788 10053 17816 10084
rect 17773 10047 17831 10053
rect 17773 10044 17785 10047
rect 17604 10016 17785 10044
rect 15304 9948 15424 9976
rect 15396 9920 15424 9948
rect 17310 9936 17316 9988
rect 17368 9976 17374 9988
rect 17604 9976 17632 10016
rect 17773 10013 17785 10016
rect 17819 10013 17831 10047
rect 17773 10007 17831 10013
rect 17862 10004 17868 10056
rect 17920 10004 17926 10056
rect 18046 10004 18052 10056
rect 18104 10004 18110 10056
rect 17368 9948 17632 9976
rect 17681 9979 17739 9985
rect 17368 9936 17374 9948
rect 17681 9945 17693 9979
rect 17727 9976 17739 9979
rect 17954 9976 17960 9988
rect 17727 9948 17960 9976
rect 17727 9945 17739 9948
rect 17681 9939 17739 9945
rect 17954 9936 17960 9948
rect 18012 9976 18018 9988
rect 18432 9976 18460 10152
rect 21542 10140 21548 10152
rect 21600 10140 21606 10192
rect 22922 10140 22928 10192
rect 22980 10180 22986 10192
rect 26234 10180 26240 10192
rect 22980 10152 26240 10180
rect 22980 10140 22986 10152
rect 26234 10140 26240 10152
rect 26292 10140 26298 10192
rect 27246 10140 27252 10192
rect 27304 10180 27310 10192
rect 28166 10180 28172 10192
rect 27304 10152 28172 10180
rect 27304 10140 27310 10152
rect 28166 10140 28172 10152
rect 28224 10140 28230 10192
rect 29546 10180 29552 10192
rect 28368 10152 29552 10180
rect 18874 10072 18880 10124
rect 18932 10112 18938 10124
rect 23382 10112 23388 10124
rect 18932 10084 23388 10112
rect 18932 10072 18938 10084
rect 23382 10072 23388 10084
rect 23440 10112 23446 10124
rect 23440 10084 26096 10112
rect 23440 10072 23446 10084
rect 19518 10044 19524 10056
rect 18012 9948 18460 9976
rect 19306 10016 19524 10044
rect 18012 9936 18018 9948
rect 8527 9880 9260 9908
rect 8527 9877 8539 9880
rect 8481 9871 8539 9877
rect 9490 9868 9496 9920
rect 9548 9908 9554 9920
rect 10226 9908 10232 9920
rect 9548 9880 10232 9908
rect 9548 9868 9554 9880
rect 10226 9868 10232 9880
rect 10284 9868 10290 9920
rect 11514 9868 11520 9920
rect 11572 9908 11578 9920
rect 11882 9908 11888 9920
rect 11572 9880 11888 9908
rect 11572 9868 11578 9880
rect 11882 9868 11888 9880
rect 11940 9868 11946 9920
rect 12158 9868 12164 9920
rect 12216 9908 12222 9920
rect 12805 9911 12863 9917
rect 12805 9908 12817 9911
rect 12216 9880 12817 9908
rect 12216 9868 12222 9880
rect 12805 9877 12817 9880
rect 12851 9877 12863 9911
rect 12805 9871 12863 9877
rect 15378 9868 15384 9920
rect 15436 9868 15442 9920
rect 15562 9868 15568 9920
rect 15620 9868 15626 9920
rect 15746 9868 15752 9920
rect 15804 9908 15810 9920
rect 15930 9908 15936 9920
rect 15804 9880 15936 9908
rect 15804 9868 15810 9880
rect 15930 9868 15936 9880
rect 15988 9908 15994 9920
rect 19058 9908 19064 9920
rect 15988 9880 19064 9908
rect 15988 9868 15994 9880
rect 19058 9868 19064 9880
rect 19116 9868 19122 9920
rect 19150 9868 19156 9920
rect 19208 9908 19214 9920
rect 19306 9908 19334 10016
rect 19518 10004 19524 10016
rect 19576 10004 19582 10056
rect 19610 10004 19616 10056
rect 19668 10004 19674 10056
rect 19886 10004 19892 10056
rect 19944 10044 19950 10056
rect 19981 10047 20039 10053
rect 19981 10044 19993 10047
rect 19944 10016 19993 10044
rect 19944 10004 19950 10016
rect 19981 10013 19993 10016
rect 20027 10013 20039 10047
rect 19981 10007 20039 10013
rect 20074 10047 20132 10053
rect 20074 10013 20086 10047
rect 20120 10013 20132 10047
rect 20349 10047 20407 10053
rect 20349 10044 20361 10047
rect 20074 10007 20132 10013
rect 20180 10016 20361 10044
rect 19628 9976 19656 10004
rect 20088 9976 20116 10007
rect 19628 9948 20116 9976
rect 19208 9880 19334 9908
rect 19208 9868 19214 9880
rect 19518 9868 19524 9920
rect 19576 9908 19582 9920
rect 20180 9908 20208 10016
rect 20349 10013 20361 10016
rect 20395 10013 20407 10047
rect 20349 10007 20407 10013
rect 20257 9979 20315 9985
rect 20257 9945 20269 9979
rect 20303 9945 20315 9979
rect 20364 9976 20392 10007
rect 20438 10004 20444 10056
rect 20496 10053 20502 10056
rect 20496 10044 20504 10053
rect 20496 10016 20541 10044
rect 20496 10007 20504 10016
rect 20496 10004 20502 10007
rect 21634 10004 21640 10056
rect 21692 10044 21698 10056
rect 22094 10044 22100 10056
rect 21692 10016 22100 10044
rect 21692 10004 21698 10016
rect 22094 10004 22100 10016
rect 22152 10044 22158 10056
rect 22281 10047 22339 10053
rect 22281 10044 22293 10047
rect 22152 10016 22293 10044
rect 22152 10004 22158 10016
rect 22281 10013 22293 10016
rect 22327 10013 22339 10047
rect 22281 10007 22339 10013
rect 22554 10004 22560 10056
rect 22612 10004 22618 10056
rect 23474 10004 23480 10056
rect 23532 10044 23538 10056
rect 23753 10047 23811 10053
rect 23753 10044 23765 10047
rect 23532 10016 23765 10044
rect 23532 10004 23538 10016
rect 23753 10013 23765 10016
rect 23799 10013 23811 10047
rect 23753 10007 23811 10013
rect 23842 10004 23848 10056
rect 23900 10004 23906 10056
rect 24026 10044 24032 10056
rect 23952 10016 24032 10044
rect 23658 9976 23664 9988
rect 20364 9948 23664 9976
rect 20257 9939 20315 9945
rect 19576 9880 20208 9908
rect 20272 9908 20300 9939
rect 23658 9936 23664 9948
rect 23716 9936 23722 9988
rect 23952 9985 23980 10016
rect 24026 10004 24032 10016
rect 24084 10004 24090 10056
rect 24121 10047 24179 10053
rect 24121 10013 24133 10047
rect 24167 10013 24179 10047
rect 24121 10007 24179 10013
rect 23937 9979 23995 9985
rect 23937 9945 23949 9979
rect 23983 9945 23995 9979
rect 23937 9939 23995 9945
rect 24136 9976 24164 10007
rect 24946 10004 24952 10056
rect 25004 10004 25010 10056
rect 25042 10047 25100 10053
rect 25042 10013 25054 10047
rect 25088 10013 25100 10047
rect 25042 10007 25100 10013
rect 25455 10047 25513 10053
rect 25455 10013 25467 10047
rect 25501 10044 25513 10047
rect 25682 10044 25688 10056
rect 25501 10016 25688 10044
rect 25501 10013 25513 10016
rect 25455 10007 25513 10013
rect 25056 9976 25084 10007
rect 25682 10004 25688 10016
rect 25740 10004 25746 10056
rect 26068 10053 26096 10084
rect 26053 10047 26111 10053
rect 26053 10013 26065 10047
rect 26099 10013 26111 10047
rect 26252 10044 26280 10140
rect 27614 10072 27620 10124
rect 27672 10112 27678 10124
rect 27798 10112 27804 10124
rect 27672 10084 27804 10112
rect 27672 10072 27678 10084
rect 27798 10072 27804 10084
rect 27856 10112 27862 10124
rect 27856 10084 28304 10112
rect 27856 10072 27862 10084
rect 27893 10047 27951 10053
rect 27893 10044 27905 10047
rect 26252 10016 27905 10044
rect 26053 10007 26111 10013
rect 27893 10013 27905 10016
rect 27939 10013 27951 10047
rect 27893 10007 27951 10013
rect 27982 10004 27988 10056
rect 28040 10044 28046 10056
rect 28276 10053 28304 10084
rect 28077 10047 28135 10053
rect 28077 10044 28089 10047
rect 28040 10016 28089 10044
rect 28040 10004 28046 10016
rect 28077 10013 28089 10016
rect 28123 10013 28135 10047
rect 28077 10007 28135 10013
rect 28261 10047 28319 10053
rect 28261 10013 28273 10047
rect 28307 10013 28319 10047
rect 28261 10007 28319 10013
rect 24136 9948 25084 9976
rect 25225 9979 25283 9985
rect 20438 9908 20444 9920
rect 20272 9880 20444 9908
rect 19576 9868 19582 9880
rect 20438 9868 20444 9880
rect 20496 9868 20502 9920
rect 22462 9868 22468 9920
rect 22520 9868 22526 9920
rect 23676 9908 23704 9936
rect 24136 9908 24164 9948
rect 25225 9945 25237 9979
rect 25271 9945 25283 9979
rect 25225 9939 25283 9945
rect 25317 9979 25375 9985
rect 25317 9945 25329 9979
rect 25363 9976 25375 9979
rect 25958 9976 25964 9988
rect 25363 9948 25964 9976
rect 25363 9945 25375 9948
rect 25317 9939 25375 9945
rect 23676 9880 24164 9908
rect 25240 9908 25268 9939
rect 25958 9936 25964 9948
rect 26016 9976 26022 9988
rect 26016 9948 28120 9976
rect 26016 9936 26022 9948
rect 25590 9908 25596 9920
rect 25240 9880 25596 9908
rect 25590 9868 25596 9880
rect 25648 9868 25654 9920
rect 27525 9911 27583 9917
rect 27525 9877 27537 9911
rect 27571 9908 27583 9911
rect 27614 9908 27620 9920
rect 27571 9880 27620 9908
rect 27571 9877 27583 9880
rect 27525 9871 27583 9877
rect 27614 9868 27620 9880
rect 27672 9868 27678 9920
rect 28092 9908 28120 9948
rect 28166 9936 28172 9988
rect 28224 9976 28230 9988
rect 28368 9976 28396 10152
rect 29546 10140 29552 10152
rect 29604 10140 29610 10192
rect 28442 10072 28448 10124
rect 28500 10112 28506 10124
rect 28500 10084 28948 10112
rect 28500 10072 28506 10084
rect 28810 10004 28816 10056
rect 28868 10004 28874 10056
rect 28920 10044 28948 10084
rect 28994 10072 29000 10124
rect 29052 10112 29058 10124
rect 29730 10112 29736 10124
rect 29052 10084 29736 10112
rect 29052 10072 29058 10084
rect 29730 10072 29736 10084
rect 29788 10072 29794 10124
rect 30374 10072 30380 10124
rect 30432 10112 30438 10124
rect 30650 10112 30656 10124
rect 30432 10084 30656 10112
rect 30432 10072 30438 10084
rect 30650 10072 30656 10084
rect 30708 10072 30714 10124
rect 31294 10072 31300 10124
rect 31352 10072 31358 10124
rect 31846 10072 31852 10124
rect 31904 10112 31910 10124
rect 31904 10084 33180 10112
rect 31904 10072 31910 10084
rect 29178 10044 29184 10056
rect 28920 10016 29184 10044
rect 29178 10004 29184 10016
rect 29236 10004 29242 10056
rect 30668 10044 30696 10072
rect 33152 10056 33180 10084
rect 30745 10047 30803 10053
rect 30745 10044 30757 10047
rect 30668 10016 30757 10044
rect 30745 10013 30757 10016
rect 30791 10013 30803 10047
rect 30745 10007 30803 10013
rect 30837 10047 30895 10053
rect 30837 10013 30849 10047
rect 30883 10044 30895 10047
rect 31021 10047 31079 10053
rect 31021 10044 31033 10047
rect 30883 10016 31033 10044
rect 30883 10013 30895 10016
rect 30837 10007 30895 10013
rect 31021 10013 31033 10016
rect 31067 10013 31079 10047
rect 31021 10007 31079 10013
rect 33134 10004 33140 10056
rect 33192 10044 33198 10056
rect 33413 10047 33471 10053
rect 33413 10044 33425 10047
rect 33192 10016 33425 10044
rect 33192 10004 33198 10016
rect 33413 10013 33425 10016
rect 33459 10013 33471 10047
rect 33413 10007 33471 10013
rect 28224 9948 28396 9976
rect 28629 9979 28687 9985
rect 28224 9936 28230 9948
rect 28629 9945 28641 9979
rect 28675 9976 28687 9979
rect 28828 9976 28856 10004
rect 31294 9976 31300 9988
rect 28675 9948 31300 9976
rect 28675 9945 28687 9948
rect 28629 9939 28687 9945
rect 28644 9908 28672 9939
rect 31294 9936 31300 9948
rect 31352 9936 31358 9988
rect 31570 9936 31576 9988
rect 31628 9976 31634 9988
rect 31628 9948 31786 9976
rect 31628 9936 31634 9948
rect 28092 9880 28672 9908
rect 28810 9868 28816 9920
rect 28868 9917 28874 9920
rect 28868 9911 28887 9917
rect 28875 9877 28887 9911
rect 28868 9871 28887 9877
rect 28868 9868 28874 9871
rect 29546 9868 29552 9920
rect 29604 9908 29610 9920
rect 32766 9908 32772 9920
rect 29604 9880 32772 9908
rect 29604 9868 29610 9880
rect 32766 9868 32772 9880
rect 32824 9868 32830 9920
rect 33505 9911 33563 9917
rect 33505 9877 33517 9911
rect 33551 9908 33563 9911
rect 35066 9908 35072 9920
rect 33551 9880 35072 9908
rect 33551 9877 33563 9880
rect 33505 9871 33563 9877
rect 35066 9868 35072 9880
rect 35124 9868 35130 9920
rect 1104 9818 38272 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 38272 9818
rect 1104 9744 38272 9766
rect 6546 9664 6552 9716
rect 6604 9664 6610 9716
rect 6822 9704 6828 9716
rect 6656 9676 6828 9704
rect 6564 9636 6592 9664
rect 6656 9645 6684 9676
rect 6822 9664 6828 9676
rect 6880 9664 6886 9716
rect 6914 9664 6920 9716
rect 6972 9704 6978 9716
rect 8113 9707 8171 9713
rect 6972 9676 8064 9704
rect 6972 9664 6978 9676
rect 6380 9608 6592 9636
rect 6641 9639 6699 9645
rect 6380 9577 6408 9608
rect 6641 9605 6653 9639
rect 6687 9605 6699 9639
rect 8036 9636 8064 9676
rect 8113 9673 8125 9707
rect 8159 9704 8171 9707
rect 8202 9704 8208 9716
rect 8159 9676 8208 9704
rect 8159 9673 8171 9676
rect 8113 9667 8171 9673
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 10778 9704 10784 9716
rect 8312 9676 10784 9704
rect 8312 9636 8340 9676
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 11606 9704 11612 9716
rect 11348 9676 11612 9704
rect 9858 9636 9864 9648
rect 8036 9608 8340 9636
rect 9600 9608 9864 9636
rect 6641 9599 6699 9605
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9537 6423 9571
rect 6365 9531 6423 9537
rect 7742 9528 7748 9580
rect 7800 9568 7806 9580
rect 7926 9568 7932 9580
rect 7800 9540 7932 9568
rect 7800 9528 7806 9540
rect 7926 9528 7932 9540
rect 7984 9528 7990 9580
rect 9600 9577 9628 9608
rect 9858 9596 9864 9608
rect 9916 9596 9922 9648
rect 11348 9636 11376 9676
rect 11606 9664 11612 9676
rect 11664 9664 11670 9716
rect 11882 9664 11888 9716
rect 11940 9704 11946 9716
rect 16485 9707 16543 9713
rect 11940 9676 16436 9704
rect 11940 9664 11946 9676
rect 12158 9636 12164 9648
rect 11164 9608 11376 9636
rect 11992 9608 12164 9636
rect 9585 9571 9643 9577
rect 9585 9537 9597 9571
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 10962 9528 10968 9580
rect 11020 9528 11026 9580
rect 6178 9460 6184 9512
rect 6236 9500 6242 9512
rect 7760 9500 7788 9528
rect 6236 9472 7788 9500
rect 6236 9460 6242 9472
rect 9858 9460 9864 9512
rect 9916 9460 9922 9512
rect 10594 9460 10600 9512
rect 10652 9500 10658 9512
rect 11164 9500 11192 9608
rect 11992 9577 12020 9608
rect 12158 9596 12164 9608
rect 12216 9596 12222 9648
rect 13906 9596 13912 9648
rect 13964 9596 13970 9648
rect 15562 9596 15568 9648
rect 15620 9636 15626 9648
rect 16408 9636 16436 9676
rect 16485 9673 16497 9707
rect 16531 9704 16543 9707
rect 16666 9704 16672 9716
rect 16531 9676 16672 9704
rect 16531 9673 16543 9676
rect 16485 9667 16543 9673
rect 16666 9664 16672 9676
rect 16724 9664 16730 9716
rect 16776 9676 17724 9704
rect 16776 9636 16804 9676
rect 15620 9608 16344 9636
rect 16408 9608 16804 9636
rect 15620 9596 15626 9608
rect 11977 9571 12035 9577
rect 11977 9537 11989 9571
rect 12023 9537 12035 9571
rect 11977 9531 12035 9537
rect 13354 9528 13360 9580
rect 13412 9528 13418 9580
rect 15286 9528 15292 9580
rect 15344 9568 15350 9580
rect 15654 9568 15660 9580
rect 15344 9540 15660 9568
rect 15344 9528 15350 9540
rect 15654 9528 15660 9540
rect 15712 9528 15718 9580
rect 15838 9528 15844 9580
rect 15896 9528 15902 9580
rect 15930 9528 15936 9580
rect 15988 9528 15994 9580
rect 16114 9528 16120 9580
rect 16172 9528 16178 9580
rect 16316 9577 16344 9608
rect 16942 9596 16948 9648
rect 17000 9636 17006 9648
rect 17037 9639 17095 9645
rect 17037 9636 17049 9639
rect 17000 9608 17049 9636
rect 17000 9596 17006 9608
rect 17037 9605 17049 9608
rect 17083 9605 17095 9639
rect 17494 9636 17500 9648
rect 17037 9599 17095 9605
rect 17144 9608 17500 9636
rect 16209 9571 16267 9577
rect 16209 9537 16221 9571
rect 16255 9537 16267 9571
rect 16209 9531 16267 9537
rect 16301 9571 16359 9577
rect 16301 9537 16313 9571
rect 16347 9537 16359 9571
rect 16301 9531 16359 9537
rect 11514 9500 11520 9512
rect 10652 9472 11192 9500
rect 11256 9472 11520 9500
rect 10652 9460 10658 9472
rect 10870 9392 10876 9444
rect 10928 9432 10934 9444
rect 11256 9432 11284 9472
rect 11514 9460 11520 9472
rect 11572 9460 11578 9512
rect 12986 9460 12992 9512
rect 13044 9500 13050 9512
rect 13372 9500 13400 9528
rect 13044 9472 13400 9500
rect 13648 9472 15792 9500
rect 13044 9460 13050 9472
rect 10928 9404 11284 9432
rect 10928 9392 10934 9404
rect 13262 9392 13268 9444
rect 13320 9432 13326 9444
rect 13648 9432 13676 9472
rect 13320 9404 13676 9432
rect 13725 9435 13783 9441
rect 13320 9392 13326 9404
rect 13725 9401 13737 9435
rect 13771 9432 13783 9435
rect 14274 9432 14280 9444
rect 13771 9404 14280 9432
rect 13771 9401 13783 9404
rect 13725 9395 13783 9401
rect 14274 9392 14280 9404
rect 14332 9392 14338 9444
rect 10410 9324 10416 9376
rect 10468 9364 10474 9376
rect 11333 9367 11391 9373
rect 11333 9364 11345 9367
rect 10468 9336 11345 9364
rect 10468 9324 10474 9336
rect 11333 9333 11345 9336
rect 11379 9333 11391 9367
rect 11333 9327 11391 9333
rect 11514 9324 11520 9376
rect 11572 9364 11578 9376
rect 11790 9364 11796 9376
rect 11572 9336 11796 9364
rect 11572 9324 11578 9336
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 12240 9367 12298 9373
rect 12240 9333 12252 9367
rect 12286 9364 12298 9367
rect 12342 9364 12348 9376
rect 12286 9336 12348 9364
rect 12286 9333 12298 9336
rect 12240 9327 12298 9333
rect 12342 9324 12348 9336
rect 12400 9324 12406 9376
rect 14458 9324 14464 9376
rect 14516 9364 14522 9376
rect 15197 9367 15255 9373
rect 15197 9364 15209 9367
rect 14516 9336 15209 9364
rect 14516 9324 14522 9336
rect 15197 9333 15209 9336
rect 15243 9333 15255 9367
rect 15764 9364 15792 9472
rect 15856 9432 15884 9528
rect 16224 9500 16252 9531
rect 16666 9528 16672 9580
rect 16724 9568 16730 9580
rect 17144 9568 17172 9608
rect 17328 9577 17356 9608
rect 17494 9596 17500 9608
rect 17552 9596 17558 9648
rect 17696 9636 17724 9676
rect 17770 9664 17776 9716
rect 17828 9664 17834 9716
rect 18417 9707 18475 9713
rect 18417 9673 18429 9707
rect 18463 9704 18475 9707
rect 18506 9704 18512 9716
rect 18463 9676 18512 9704
rect 18463 9673 18475 9676
rect 18417 9667 18475 9673
rect 18506 9664 18512 9676
rect 18564 9664 18570 9716
rect 20162 9704 20168 9716
rect 18984 9676 20168 9704
rect 18984 9636 19012 9676
rect 20162 9664 20168 9676
rect 20220 9664 20226 9716
rect 20898 9664 20904 9716
rect 20956 9704 20962 9716
rect 21358 9704 21364 9716
rect 20956 9676 21364 9704
rect 20956 9664 20962 9676
rect 21358 9664 21364 9676
rect 21416 9664 21422 9716
rect 21542 9664 21548 9716
rect 21600 9704 21606 9716
rect 21600 9676 22600 9704
rect 21600 9664 21606 9676
rect 17696 9608 19012 9636
rect 19058 9596 19064 9648
rect 19116 9636 19122 9648
rect 21266 9636 21272 9648
rect 19116 9608 21272 9636
rect 19116 9596 19122 9608
rect 21266 9596 21272 9608
rect 21324 9596 21330 9648
rect 22572 9636 22600 9676
rect 22646 9664 22652 9716
rect 22704 9704 22710 9716
rect 24210 9704 24216 9716
rect 22704 9676 24216 9704
rect 22704 9664 22710 9676
rect 24210 9664 24216 9676
rect 24268 9664 24274 9716
rect 24946 9704 24952 9716
rect 24596 9676 24952 9704
rect 24596 9674 24624 9676
rect 23198 9636 23204 9648
rect 22572 9608 23204 9636
rect 23198 9596 23204 9608
rect 23256 9596 23262 9648
rect 23934 9596 23940 9648
rect 23992 9596 23998 9648
rect 24504 9646 24624 9674
rect 24946 9664 24952 9676
rect 25004 9664 25010 9716
rect 28166 9704 28172 9716
rect 26620 9676 28172 9704
rect 16724 9540 17172 9568
rect 17221 9571 17279 9577
rect 16724 9528 16730 9540
rect 17221 9537 17233 9571
rect 17267 9537 17279 9571
rect 17221 9531 17279 9537
rect 17313 9571 17371 9577
rect 17313 9537 17325 9571
rect 17359 9537 17371 9571
rect 17313 9531 17371 9537
rect 16758 9500 16764 9512
rect 16224 9472 16764 9500
rect 16758 9460 16764 9472
rect 16816 9460 16822 9512
rect 16482 9432 16488 9444
rect 15856 9404 16488 9432
rect 16482 9392 16488 9404
rect 16540 9392 16546 9444
rect 17034 9432 17040 9444
rect 16868 9404 17040 9432
rect 16868 9364 16896 9404
rect 17034 9392 17040 9404
rect 17092 9392 17098 9444
rect 15764 9336 16896 9364
rect 15197 9327 15255 9333
rect 16942 9324 16948 9376
rect 17000 9364 17006 9376
rect 17236 9364 17264 9531
rect 17402 9528 17408 9580
rect 17460 9528 17466 9580
rect 17681 9571 17739 9577
rect 17681 9537 17693 9571
rect 17727 9537 17739 9571
rect 17681 9531 17739 9537
rect 17957 9571 18015 9577
rect 17957 9537 17969 9571
rect 18003 9568 18015 9571
rect 18046 9568 18052 9580
rect 18003 9540 18052 9568
rect 18003 9537 18015 9540
rect 17957 9531 18015 9537
rect 17696 9500 17724 9531
rect 18046 9528 18052 9540
rect 18104 9528 18110 9580
rect 19334 9528 19340 9580
rect 19392 9528 19398 9580
rect 20070 9528 20076 9580
rect 20128 9568 20134 9580
rect 20128 9540 20484 9568
rect 20128 9528 20134 9540
rect 20456 9512 20484 9540
rect 21818 9528 21824 9580
rect 21876 9568 21882 9580
rect 22097 9571 22155 9577
rect 22097 9568 22109 9571
rect 21876 9540 22109 9568
rect 21876 9528 21882 9540
rect 22097 9537 22109 9540
rect 22143 9537 22155 9571
rect 22097 9531 22155 9537
rect 22741 9571 22799 9577
rect 22741 9537 22753 9571
rect 22787 9568 22799 9571
rect 22830 9568 22836 9580
rect 22787 9540 22836 9568
rect 22787 9537 22799 9540
rect 22741 9531 22799 9537
rect 22830 9528 22836 9540
rect 22888 9528 22894 9580
rect 23566 9528 23572 9580
rect 23624 9528 23630 9580
rect 23658 9528 23664 9580
rect 23716 9528 23722 9580
rect 23750 9528 23756 9580
rect 23808 9568 23814 9580
rect 24504 9577 24532 9646
rect 24670 9596 24676 9648
rect 24728 9596 24734 9648
rect 24854 9596 24860 9648
rect 24912 9596 24918 9648
rect 25041 9639 25099 9645
rect 25041 9605 25053 9639
rect 25087 9636 25099 9639
rect 26620 9636 26648 9676
rect 25087 9608 26648 9636
rect 25087 9605 25099 9608
rect 25041 9599 25099 9605
rect 26694 9596 26700 9648
rect 26752 9636 26758 9648
rect 27341 9639 27399 9645
rect 27341 9636 27353 9639
rect 26752 9608 27353 9636
rect 26752 9596 26758 9608
rect 27341 9605 27353 9608
rect 27387 9605 27399 9639
rect 27341 9599 27399 9605
rect 25866 9577 25872 9580
rect 23845 9571 23903 9577
rect 23845 9568 23857 9571
rect 23808 9540 23857 9568
rect 23808 9528 23814 9540
rect 23845 9537 23857 9540
rect 23891 9537 23903 9571
rect 23845 9531 23903 9537
rect 24029 9571 24087 9577
rect 24029 9537 24041 9571
rect 24075 9537 24087 9571
rect 24029 9531 24087 9537
rect 24489 9571 24547 9577
rect 24489 9537 24501 9571
rect 24535 9537 24547 9571
rect 24489 9531 24547 9537
rect 24765 9571 24823 9577
rect 24765 9537 24777 9571
rect 24811 9537 24823 9571
rect 25864 9568 25872 9577
rect 25827 9540 25872 9568
rect 24765 9531 24823 9537
rect 25864 9531 25872 9540
rect 20254 9500 20260 9512
rect 17512 9472 20260 9500
rect 17512 9444 17540 9472
rect 20254 9460 20260 9472
rect 20312 9460 20318 9512
rect 20438 9460 20444 9512
rect 20496 9460 20502 9512
rect 22189 9503 22247 9509
rect 22189 9500 22201 9503
rect 20824 9472 22201 9500
rect 17494 9392 17500 9444
rect 17552 9392 17558 9444
rect 17589 9435 17647 9441
rect 17589 9401 17601 9435
rect 17635 9432 17647 9435
rect 18049 9435 18107 9441
rect 18049 9432 18061 9435
rect 17635 9404 18061 9432
rect 17635 9401 17647 9404
rect 17589 9395 17647 9401
rect 18049 9401 18061 9404
rect 18095 9401 18107 9435
rect 18049 9395 18107 9401
rect 20824 9376 20852 9472
rect 22189 9469 22201 9472
rect 22235 9469 22247 9503
rect 22189 9463 22247 9469
rect 22557 9503 22615 9509
rect 22557 9469 22569 9503
rect 22603 9500 22615 9503
rect 23584 9500 23612 9528
rect 22603 9472 23612 9500
rect 22603 9469 22615 9472
rect 22557 9463 22615 9469
rect 22922 9392 22928 9444
rect 22980 9392 22986 9444
rect 23492 9376 23520 9472
rect 24044 9444 24072 9531
rect 24670 9460 24676 9512
rect 24728 9500 24734 9512
rect 24780 9500 24808 9531
rect 25866 9528 25872 9531
rect 25924 9528 25930 9580
rect 25961 9571 26019 9577
rect 25961 9537 25973 9571
rect 26007 9537 26019 9571
rect 25961 9531 26019 9537
rect 26053 9571 26111 9577
rect 26053 9537 26065 9571
rect 26099 9568 26111 9571
rect 26142 9568 26148 9580
rect 26099 9540 26148 9568
rect 26099 9537 26111 9540
rect 26053 9531 26111 9537
rect 24728 9472 24808 9500
rect 25976 9500 26004 9531
rect 26142 9528 26148 9540
rect 26200 9528 26206 9580
rect 26234 9528 26240 9580
rect 26292 9528 26298 9580
rect 26329 9571 26387 9577
rect 26329 9537 26341 9571
rect 26375 9568 26387 9571
rect 26602 9568 26608 9580
rect 26375 9540 26608 9568
rect 26375 9537 26387 9540
rect 26329 9531 26387 9537
rect 26602 9528 26608 9540
rect 26660 9568 26666 9580
rect 26970 9568 26976 9580
rect 26660 9540 26976 9568
rect 26660 9528 26666 9540
rect 26970 9528 26976 9540
rect 27028 9528 27034 9580
rect 27154 9528 27160 9580
rect 27212 9528 27218 9580
rect 27249 9571 27307 9577
rect 27249 9537 27261 9571
rect 27295 9537 27307 9571
rect 27448 9568 27476 9676
rect 28166 9664 28172 9676
rect 28224 9664 28230 9716
rect 28442 9704 28448 9716
rect 28276 9676 28448 9704
rect 28074 9596 28080 9648
rect 28132 9636 28138 9648
rect 28276 9636 28304 9676
rect 28442 9664 28448 9676
rect 28500 9704 28506 9716
rect 28810 9704 28816 9716
rect 28500 9676 28816 9704
rect 28500 9664 28506 9676
rect 28810 9664 28816 9676
rect 28868 9664 28874 9716
rect 33318 9664 33324 9716
rect 33376 9664 33382 9716
rect 28132 9608 28304 9636
rect 28132 9596 28138 9608
rect 29362 9596 29368 9648
rect 29420 9636 29426 9648
rect 29825 9639 29883 9645
rect 29825 9636 29837 9639
rect 29420 9608 29837 9636
rect 29420 9596 29426 9608
rect 29825 9605 29837 9608
rect 29871 9605 29883 9639
rect 29825 9599 29883 9605
rect 30098 9596 30104 9648
rect 30156 9636 30162 9648
rect 33502 9636 33508 9648
rect 30156 9608 33508 9636
rect 30156 9596 30162 9608
rect 33502 9596 33508 9608
rect 33560 9596 33566 9648
rect 34514 9596 34520 9648
rect 34572 9636 34578 9648
rect 34793 9639 34851 9645
rect 34793 9636 34805 9639
rect 34572 9608 34805 9636
rect 34572 9596 34578 9608
rect 34793 9605 34805 9608
rect 34839 9605 34851 9639
rect 34793 9599 34851 9605
rect 27525 9571 27583 9577
rect 27525 9568 27537 9571
rect 27448 9540 27537 9568
rect 27249 9531 27307 9537
rect 27525 9537 27537 9540
rect 27571 9537 27583 9571
rect 27525 9531 27583 9537
rect 27264 9500 27292 9531
rect 29454 9528 29460 9580
rect 29512 9528 29518 9580
rect 29641 9571 29699 9577
rect 29641 9537 29653 9571
rect 29687 9537 29699 9571
rect 29641 9531 29699 9537
rect 28350 9500 28356 9512
rect 25976 9472 28356 9500
rect 24728 9460 24734 9472
rect 28350 9460 28356 9472
rect 28408 9500 28414 9512
rect 29472 9500 29500 9528
rect 28408 9472 29500 9500
rect 29656 9500 29684 9531
rect 29914 9528 29920 9580
rect 29972 9528 29978 9580
rect 30009 9571 30067 9577
rect 30009 9537 30021 9571
rect 30055 9568 30067 9571
rect 30282 9568 30288 9580
rect 30055 9540 30288 9568
rect 30055 9537 30067 9540
rect 30009 9531 30067 9537
rect 30282 9528 30288 9540
rect 30340 9528 30346 9580
rect 32766 9528 32772 9580
rect 32824 9568 32830 9580
rect 32824 9540 33456 9568
rect 32824 9528 32830 9540
rect 30837 9503 30895 9509
rect 30837 9500 30849 9503
rect 29656 9472 30849 9500
rect 28408 9460 28414 9472
rect 30837 9469 30849 9472
rect 30883 9469 30895 9503
rect 30837 9463 30895 9469
rect 31294 9460 31300 9512
rect 31352 9500 31358 9512
rect 31481 9503 31539 9509
rect 31481 9500 31493 9503
rect 31352 9472 31493 9500
rect 31352 9460 31358 9472
rect 31481 9469 31493 9472
rect 31527 9500 31539 9503
rect 31938 9500 31944 9512
rect 31527 9472 31944 9500
rect 31527 9469 31539 9472
rect 31481 9463 31539 9469
rect 31938 9460 31944 9472
rect 31996 9460 32002 9512
rect 32861 9503 32919 9509
rect 32861 9469 32873 9503
rect 32907 9469 32919 9503
rect 32861 9463 32919 9469
rect 32953 9503 33011 9509
rect 32953 9469 32965 9503
rect 32999 9500 33011 9503
rect 33318 9500 33324 9512
rect 32999 9472 33324 9500
rect 32999 9469 33011 9472
rect 32953 9463 33011 9469
rect 24026 9392 24032 9444
rect 24084 9432 24090 9444
rect 24578 9432 24584 9444
rect 24084 9404 24584 9432
rect 24084 9392 24090 9404
rect 24578 9392 24584 9404
rect 24636 9432 24642 9444
rect 25314 9432 25320 9444
rect 24636 9404 25320 9432
rect 24636 9392 24642 9404
rect 25314 9392 25320 9404
rect 25372 9392 25378 9444
rect 25685 9435 25743 9441
rect 25685 9401 25697 9435
rect 25731 9432 25743 9435
rect 25774 9432 25780 9444
rect 25731 9404 25780 9432
rect 25731 9401 25743 9404
rect 25685 9395 25743 9401
rect 25774 9392 25780 9404
rect 25832 9392 25838 9444
rect 26510 9392 26516 9444
rect 26568 9432 26574 9444
rect 26973 9435 27031 9441
rect 26973 9432 26985 9435
rect 26568 9404 26985 9432
rect 26568 9392 26574 9404
rect 26973 9401 26985 9404
rect 27019 9401 27031 9435
rect 26973 9395 27031 9401
rect 27246 9392 27252 9444
rect 27304 9392 27310 9444
rect 29914 9392 29920 9444
rect 29972 9432 29978 9444
rect 32582 9432 32588 9444
rect 29972 9404 32588 9432
rect 29972 9392 29978 9404
rect 32582 9392 32588 9404
rect 32640 9432 32646 9444
rect 32876 9432 32904 9463
rect 32640 9404 32904 9432
rect 32640 9392 32646 9404
rect 17862 9364 17868 9376
rect 17000 9336 17868 9364
rect 17000 9324 17006 9336
rect 17862 9324 17868 9336
rect 17920 9324 17926 9376
rect 17954 9324 17960 9376
rect 18012 9364 18018 9376
rect 18141 9367 18199 9373
rect 18141 9364 18153 9367
rect 18012 9336 18153 9364
rect 18012 9324 18018 9336
rect 18141 9333 18153 9336
rect 18187 9364 18199 9367
rect 19794 9364 19800 9376
rect 18187 9336 19800 9364
rect 18187 9333 18199 9336
rect 18141 9327 18199 9333
rect 19794 9324 19800 9336
rect 19852 9324 19858 9376
rect 20622 9324 20628 9376
rect 20680 9324 20686 9376
rect 20806 9324 20812 9376
rect 20864 9324 20870 9376
rect 22189 9367 22247 9373
rect 22189 9333 22201 9367
rect 22235 9364 22247 9367
rect 22278 9364 22284 9376
rect 22235 9336 22284 9364
rect 22235 9333 22247 9336
rect 22189 9327 22247 9333
rect 22278 9324 22284 9336
rect 22336 9324 22342 9376
rect 22462 9324 22468 9376
rect 22520 9324 22526 9376
rect 23474 9324 23480 9376
rect 23532 9324 23538 9376
rect 24213 9367 24271 9373
rect 24213 9333 24225 9367
rect 24259 9364 24271 9367
rect 27264 9364 27292 9392
rect 24259 9336 27292 9364
rect 30193 9367 30251 9373
rect 24259 9333 24271 9336
rect 24213 9327 24271 9333
rect 30193 9333 30205 9367
rect 30239 9364 30251 9367
rect 30466 9364 30472 9376
rect 30239 9336 30472 9364
rect 30239 9333 30251 9336
rect 30193 9327 30251 9333
rect 30466 9324 30472 9336
rect 30524 9324 30530 9376
rect 32398 9324 32404 9376
rect 32456 9324 32462 9376
rect 32766 9324 32772 9376
rect 32824 9364 32830 9376
rect 32968 9364 32996 9463
rect 33318 9460 33324 9472
rect 33376 9460 33382 9512
rect 33428 9500 33456 9540
rect 33686 9528 33692 9580
rect 33744 9528 33750 9580
rect 34422 9500 34428 9512
rect 33428 9472 34428 9500
rect 34422 9460 34428 9472
rect 34480 9460 34486 9512
rect 35066 9460 35072 9512
rect 35124 9460 35130 9512
rect 32824 9336 32996 9364
rect 32824 9324 32830 9336
rect 1104 9274 38272 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38272 9274
rect 1104 9200 38272 9222
rect 9858 9120 9864 9172
rect 9916 9160 9922 9172
rect 10505 9163 10563 9169
rect 10505 9160 10517 9163
rect 9916 9132 10517 9160
rect 9916 9120 9922 9132
rect 10505 9129 10517 9132
rect 10551 9129 10563 9163
rect 10505 9123 10563 9129
rect 11146 9120 11152 9172
rect 11204 9160 11210 9172
rect 11425 9163 11483 9169
rect 11425 9160 11437 9163
rect 11204 9132 11437 9160
rect 11204 9120 11210 9132
rect 11425 9129 11437 9132
rect 11471 9129 11483 9163
rect 11425 9123 11483 9129
rect 12342 9120 12348 9172
rect 12400 9160 12406 9172
rect 13081 9163 13139 9169
rect 13081 9160 13093 9163
rect 12400 9132 13093 9160
rect 12400 9120 12406 9132
rect 13081 9129 13093 9132
rect 13127 9129 13139 9163
rect 13081 9123 13139 9129
rect 13188 9132 15424 9160
rect 10962 9052 10968 9104
rect 11020 9092 11026 9104
rect 12894 9092 12900 9104
rect 11020 9064 12900 9092
rect 11020 9052 11026 9064
rect 12894 9052 12900 9064
rect 12952 9052 12958 9104
rect 12986 9052 12992 9104
rect 13044 9092 13050 9104
rect 13188 9092 13216 9132
rect 15396 9104 15424 9132
rect 15930 9120 15936 9172
rect 15988 9160 15994 9172
rect 16209 9163 16267 9169
rect 16209 9160 16221 9163
rect 15988 9132 16221 9160
rect 15988 9120 15994 9132
rect 16209 9129 16221 9132
rect 16255 9129 16267 9163
rect 20438 9160 20444 9172
rect 16209 9123 16267 9129
rect 18064 9132 20444 9160
rect 13044 9064 13216 9092
rect 14461 9095 14519 9101
rect 13044 9052 13050 9064
rect 14461 9061 14473 9095
rect 14507 9061 14519 9095
rect 14461 9055 14519 9061
rect 11330 9024 11336 9036
rect 11072 8996 11336 9024
rect 4614 8916 4620 8968
rect 4672 8916 4678 8968
rect 10689 8959 10747 8965
rect 10689 8925 10701 8959
rect 10735 8925 10747 8959
rect 10689 8919 10747 8925
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8956 10839 8959
rect 10870 8956 10876 8968
rect 10827 8928 10876 8956
rect 10827 8925 10839 8928
rect 10781 8919 10839 8925
rect 4632 8888 4660 8916
rect 4632 8860 6960 8888
rect 6932 8832 6960 8860
rect 4522 8780 4528 8832
rect 4580 8780 4586 8832
rect 6914 8780 6920 8832
rect 6972 8780 6978 8832
rect 10704 8820 10732 8919
rect 10870 8916 10876 8928
rect 10928 8916 10934 8968
rect 11072 8965 11100 8996
rect 11330 8984 11336 8996
rect 11388 8984 11394 9036
rect 12066 8984 12072 9036
rect 12124 8984 12130 9036
rect 14476 9024 14504 9055
rect 14918 9052 14924 9104
rect 14976 9092 14982 9104
rect 14976 9064 15148 9092
rect 14976 9052 14982 9064
rect 15120 9033 15148 9064
rect 15378 9052 15384 9104
rect 15436 9052 15442 9104
rect 17310 9092 17316 9104
rect 15580 9064 17316 9092
rect 12820 8996 13216 9024
rect 10965 8959 11023 8965
rect 10965 8925 10977 8959
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 11057 8959 11115 8965
rect 11057 8925 11069 8959
rect 11103 8925 11115 8959
rect 11057 8919 11115 8925
rect 10980 8888 11008 8919
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 11977 8959 12035 8965
rect 11204 8928 11836 8956
rect 11204 8916 11210 8928
rect 11330 8888 11336 8900
rect 10980 8860 11336 8888
rect 11330 8848 11336 8860
rect 11388 8848 11394 8900
rect 11808 8888 11836 8928
rect 11977 8925 11989 8959
rect 12023 8956 12035 8959
rect 12820 8956 12848 8996
rect 12023 8928 12848 8956
rect 12023 8925 12035 8928
rect 11977 8919 12035 8925
rect 12986 8916 12992 8968
rect 13044 8916 13050 8968
rect 13004 8888 13032 8916
rect 11808 8860 13032 8888
rect 13188 8888 13216 8996
rect 13280 8996 14504 9024
rect 15105 9027 15163 9033
rect 13280 8965 13308 8996
rect 15105 8993 15117 9027
rect 15151 8993 15163 9027
rect 15105 8987 15163 8993
rect 13265 8959 13323 8965
rect 13265 8925 13277 8959
rect 13311 8925 13323 8959
rect 13265 8919 13323 8925
rect 13538 8916 13544 8968
rect 13596 8916 13602 8968
rect 13630 8916 13636 8968
rect 13688 8916 13694 8968
rect 13722 8916 13728 8968
rect 13780 8916 13786 8968
rect 13906 8916 13912 8968
rect 13964 8916 13970 8968
rect 14274 8916 14280 8968
rect 14332 8956 14338 8968
rect 14921 8959 14979 8965
rect 14921 8956 14933 8959
rect 14332 8928 14933 8956
rect 14332 8916 14338 8928
rect 14921 8925 14933 8928
rect 14967 8925 14979 8959
rect 14921 8919 14979 8925
rect 15194 8916 15200 8968
rect 15252 8916 15258 8968
rect 15580 8965 15608 9064
rect 17310 9052 17316 9064
rect 17368 9052 17374 9104
rect 15654 8984 15660 9036
rect 15712 9024 15718 9036
rect 15712 8996 16574 9024
rect 15712 8984 15718 8996
rect 15565 8959 15623 8965
rect 15565 8925 15577 8959
rect 15611 8925 15623 8959
rect 15565 8919 15623 8925
rect 15746 8916 15752 8968
rect 15804 8916 15810 8968
rect 15856 8965 15884 8996
rect 15841 8959 15899 8965
rect 15841 8925 15853 8959
rect 15887 8925 15899 8959
rect 15841 8919 15899 8925
rect 15933 8959 15991 8965
rect 15933 8925 15945 8959
rect 15979 8925 15991 8959
rect 15933 8919 15991 8925
rect 13814 8888 13820 8900
rect 13188 8860 13820 8888
rect 13814 8848 13820 8860
rect 13872 8888 13878 8900
rect 14829 8891 14887 8897
rect 14829 8888 14841 8891
rect 13872 8860 14841 8888
rect 13872 8848 13878 8860
rect 14829 8857 14841 8860
rect 14875 8857 14887 8891
rect 15212 8888 15240 8916
rect 15948 8888 15976 8919
rect 15212 8860 15976 8888
rect 16546 8888 16574 8996
rect 17862 8916 17868 8968
rect 17920 8916 17926 8968
rect 18064 8965 18092 9132
rect 20438 9120 20444 9132
rect 20496 9160 20502 9172
rect 20496 9132 20944 9160
rect 20496 9120 20502 9132
rect 18156 9064 18373 9092
rect 18156 8965 18184 9064
rect 18345 9024 18373 9064
rect 18506 9052 18512 9104
rect 18564 9052 18570 9104
rect 18690 9092 18696 9104
rect 18616 9064 18696 9092
rect 18616 9024 18644 9064
rect 18690 9052 18696 9064
rect 18748 9052 18754 9104
rect 19610 9052 19616 9104
rect 19668 9052 19674 9104
rect 19794 9052 19800 9104
rect 19852 9092 19858 9104
rect 19852 9064 20116 9092
rect 19852 9052 19858 9064
rect 18345 8996 20005 9024
rect 18267 8969 18325 8975
rect 18049 8959 18107 8965
rect 18049 8925 18061 8959
rect 18095 8925 18107 8959
rect 18049 8919 18107 8925
rect 18141 8959 18199 8965
rect 18141 8925 18153 8959
rect 18187 8925 18199 8959
rect 18267 8935 18279 8969
rect 18313 8968 18325 8969
rect 18313 8935 18328 8968
rect 18267 8929 18328 8935
rect 18306 8928 18328 8929
rect 18141 8919 18199 8925
rect 18322 8916 18328 8928
rect 18380 8916 18386 8968
rect 19610 8916 19616 8968
rect 19668 8956 19674 8968
rect 19786 8965 19912 8966
rect 19977 8965 20005 8996
rect 20088 8965 20116 9064
rect 20162 9052 20168 9104
rect 20220 9092 20226 9104
rect 20220 9064 20484 9092
rect 20220 9052 20226 9064
rect 19786 8959 19927 8965
rect 19786 8956 19881 8959
rect 19668 8938 19881 8956
rect 19668 8928 19814 8938
rect 19668 8916 19674 8928
rect 19869 8925 19881 8938
rect 19915 8925 19927 8959
rect 19977 8959 20036 8965
rect 19977 8928 19990 8959
rect 19869 8919 19927 8925
rect 19978 8925 19990 8928
rect 20024 8925 20036 8959
rect 19978 8919 20036 8925
rect 20078 8959 20136 8965
rect 20078 8925 20090 8959
rect 20124 8925 20136 8959
rect 20078 8919 20136 8925
rect 20257 8959 20315 8965
rect 20257 8925 20269 8959
rect 20303 8925 20315 8959
rect 20257 8919 20315 8925
rect 20349 8959 20407 8965
rect 20349 8925 20361 8959
rect 20395 8950 20407 8959
rect 20456 8956 20484 9064
rect 20530 9052 20536 9104
rect 20588 9052 20594 9104
rect 20916 9092 20944 9132
rect 20990 9120 20996 9172
rect 21048 9120 21054 9172
rect 21634 9120 21640 9172
rect 21692 9160 21698 9172
rect 22465 9163 22523 9169
rect 22465 9160 22477 9163
rect 21692 9132 22477 9160
rect 21692 9120 21698 9132
rect 22465 9129 22477 9132
rect 22511 9129 22523 9163
rect 22465 9123 22523 9129
rect 23106 9120 23112 9172
rect 23164 9160 23170 9172
rect 23658 9160 23664 9172
rect 23164 9132 23664 9160
rect 23164 9120 23170 9132
rect 23658 9120 23664 9132
rect 23716 9160 23722 9172
rect 25222 9160 25228 9172
rect 23716 9132 25228 9160
rect 23716 9120 23722 9132
rect 25222 9120 25228 9132
rect 25280 9120 25286 9172
rect 25314 9120 25320 9172
rect 25372 9160 25378 9172
rect 28258 9160 28264 9172
rect 25372 9132 28264 9160
rect 25372 9120 25378 9132
rect 28258 9120 28264 9132
rect 28316 9120 28322 9172
rect 28810 9120 28816 9172
rect 28868 9120 28874 9172
rect 28994 9120 29000 9172
rect 29052 9120 29058 9172
rect 30098 9120 30104 9172
rect 30156 9120 30162 9172
rect 30834 9160 30840 9172
rect 30300 9132 30840 9160
rect 22097 9095 22155 9101
rect 20916 9064 21956 9092
rect 20548 9024 20576 9052
rect 21818 9024 21824 9036
rect 20548 8996 21824 9024
rect 20451 8950 20484 8956
rect 20395 8928 20484 8950
rect 20395 8925 20479 8928
rect 20349 8922 20479 8925
rect 20349 8919 20407 8922
rect 19242 8888 19248 8900
rect 16546 8860 19248 8888
rect 14829 8851 14887 8857
rect 19242 8848 19248 8860
rect 19300 8848 19306 8900
rect 20272 8888 20300 8919
rect 20530 8916 20536 8968
rect 20588 8916 20594 8968
rect 20640 8965 20668 8996
rect 21818 8984 21824 8996
rect 21876 8984 21882 9036
rect 21928 9024 21956 9064
rect 22097 9061 22109 9095
rect 22143 9092 22155 9095
rect 22143 9064 22600 9092
rect 22143 9061 22155 9064
rect 22097 9055 22155 9061
rect 22572 9033 22600 9064
rect 22830 9052 22836 9104
rect 22888 9092 22894 9104
rect 28718 9092 28724 9104
rect 22888 9064 28724 9092
rect 22888 9052 22894 9064
rect 28718 9052 28724 9064
rect 28776 9052 28782 9104
rect 30300 9092 30328 9132
rect 30834 9120 30840 9132
rect 30892 9120 30898 9172
rect 31938 9120 31944 9172
rect 31996 9120 32002 9172
rect 32398 9120 32404 9172
rect 32456 9120 32462 9172
rect 34422 9120 34428 9172
rect 34480 9120 34486 9172
rect 29840 9064 30328 9092
rect 22557 9027 22615 9033
rect 21928 8996 22048 9024
rect 20625 8959 20683 8965
rect 20625 8925 20637 8959
rect 20671 8925 20683 8959
rect 20625 8919 20683 8925
rect 20717 8959 20775 8965
rect 20717 8925 20729 8959
rect 20763 8925 20775 8959
rect 20717 8919 20775 8925
rect 21085 8959 21143 8965
rect 21085 8925 21097 8959
rect 21131 8956 21143 8959
rect 21174 8956 21180 8968
rect 21131 8928 21180 8956
rect 21131 8925 21143 8928
rect 21085 8919 21143 8925
rect 20732 8888 20760 8919
rect 21174 8916 21180 8928
rect 21232 8916 21238 8968
rect 21542 8916 21548 8968
rect 21600 8916 21606 8968
rect 21910 8916 21916 8968
rect 21968 8916 21974 8968
rect 22020 8956 22048 8996
rect 22557 8993 22569 9027
rect 22603 8993 22615 9027
rect 22557 8987 22615 8993
rect 24394 8984 24400 9036
rect 24452 8984 24458 9036
rect 25038 8984 25044 9036
rect 25096 9024 25102 9036
rect 26053 9027 26111 9033
rect 26053 9024 26065 9027
rect 25096 8996 26065 9024
rect 25096 8984 25102 8996
rect 22741 8959 22799 8965
rect 22020 8928 22692 8956
rect 20806 8888 20812 8900
rect 20272 8860 20484 8888
rect 20732 8860 20812 8888
rect 20456 8832 20484 8860
rect 20806 8848 20812 8860
rect 20864 8888 20870 8900
rect 21269 8891 21327 8897
rect 20864 8860 21220 8888
rect 20864 8848 20870 8860
rect 21192 8832 21220 8860
rect 21269 8857 21281 8891
rect 21315 8857 21327 8891
rect 21269 8851 21327 8857
rect 21453 8891 21511 8897
rect 21453 8857 21465 8891
rect 21499 8888 21511 8891
rect 21729 8891 21787 8897
rect 21729 8888 21741 8891
rect 21499 8860 21741 8888
rect 21499 8857 21511 8860
rect 21453 8851 21511 8857
rect 21729 8857 21741 8860
rect 21775 8857 21787 8891
rect 21729 8851 21787 8857
rect 11517 8823 11575 8829
rect 11517 8820 11529 8823
rect 10704 8792 11529 8820
rect 11517 8789 11529 8792
rect 11563 8789 11575 8823
rect 11517 8783 11575 8789
rect 11885 8823 11943 8829
rect 11885 8789 11897 8823
rect 11931 8820 11943 8823
rect 12342 8820 12348 8832
rect 11931 8792 12348 8820
rect 11931 8789 11943 8792
rect 11885 8783 11943 8789
rect 12342 8780 12348 8792
rect 12400 8780 12406 8832
rect 12894 8780 12900 8832
rect 12952 8820 12958 8832
rect 13357 8823 13415 8829
rect 13357 8820 13369 8823
rect 12952 8792 13369 8820
rect 12952 8780 12958 8792
rect 13357 8789 13369 8792
rect 13403 8789 13415 8823
rect 13357 8783 13415 8789
rect 15378 8780 15384 8832
rect 15436 8820 15442 8832
rect 18322 8820 18328 8832
rect 15436 8792 18328 8820
rect 15436 8780 15442 8792
rect 18322 8780 18328 8792
rect 18380 8780 18386 8832
rect 20438 8780 20444 8832
rect 20496 8780 20502 8832
rect 21174 8780 21180 8832
rect 21232 8780 21238 8832
rect 21284 8820 21312 8851
rect 21818 8848 21824 8900
rect 21876 8848 21882 8900
rect 22462 8848 22468 8900
rect 22520 8848 22526 8900
rect 22554 8848 22560 8900
rect 22612 8848 22618 8900
rect 22664 8888 22692 8928
rect 22741 8925 22753 8959
rect 22787 8956 22799 8959
rect 22922 8956 22928 8968
rect 22787 8928 22928 8956
rect 22787 8925 22799 8928
rect 22741 8919 22799 8925
rect 22922 8916 22928 8928
rect 22980 8916 22986 8968
rect 24578 8916 24584 8968
rect 24636 8956 24642 8968
rect 25516 8965 25544 8996
rect 26053 8993 26065 8996
rect 26099 8993 26111 9027
rect 26053 8987 26111 8993
rect 26234 8984 26240 9036
rect 26292 9024 26298 9036
rect 26418 9024 26424 9036
rect 26292 8996 26424 9024
rect 26292 8984 26298 8996
rect 26418 8984 26424 8996
rect 26476 8984 26482 9036
rect 28902 8984 28908 9036
rect 28960 8984 28966 9036
rect 24673 8959 24731 8965
rect 24673 8956 24685 8959
rect 24636 8928 24685 8956
rect 24636 8916 24642 8928
rect 24673 8925 24685 8928
rect 24719 8925 24731 8959
rect 24673 8919 24731 8925
rect 24949 8959 25007 8965
rect 24949 8925 24961 8959
rect 24995 8925 25007 8959
rect 24949 8919 25007 8925
rect 25501 8959 25559 8965
rect 25501 8925 25513 8959
rect 25547 8925 25559 8959
rect 25501 8919 25559 8925
rect 24964 8888 24992 8919
rect 25774 8916 25780 8968
rect 25832 8916 25838 8968
rect 25866 8916 25872 8968
rect 25924 8956 25930 8968
rect 25961 8959 26019 8965
rect 25961 8956 25973 8959
rect 25924 8928 25973 8956
rect 25924 8916 25930 8928
rect 25961 8925 25973 8928
rect 26007 8925 26019 8959
rect 25961 8919 26019 8925
rect 27430 8916 27436 8968
rect 27488 8956 27494 8968
rect 27801 8959 27859 8965
rect 27801 8956 27813 8959
rect 27488 8928 27813 8956
rect 27488 8916 27494 8928
rect 27801 8925 27813 8928
rect 27847 8925 27859 8959
rect 27801 8919 27859 8925
rect 27985 8959 28043 8965
rect 27985 8925 27997 8959
rect 28031 8956 28043 8959
rect 28166 8956 28172 8968
rect 28031 8928 28172 8956
rect 28031 8925 28043 8928
rect 27985 8919 28043 8925
rect 28166 8916 28172 8928
rect 28224 8916 28230 8968
rect 22664 8860 24992 8888
rect 27890 8848 27896 8900
rect 27948 8888 27954 8900
rect 28445 8891 28503 8897
rect 28445 8888 28457 8891
rect 27948 8860 28457 8888
rect 27948 8848 27954 8860
rect 28445 8857 28457 8860
rect 28491 8857 28503 8891
rect 28445 8851 28503 8857
rect 28822 8891 28880 8897
rect 28822 8857 28834 8891
rect 28868 8888 28880 8891
rect 28920 8888 28948 8984
rect 29546 8916 29552 8968
rect 29604 8916 29610 8968
rect 29840 8965 29868 9064
rect 31570 9052 31576 9104
rect 31628 9092 31634 9104
rect 31628 9064 31754 9092
rect 31628 9052 31634 9064
rect 30466 8984 30472 9036
rect 30524 8984 30530 9036
rect 31726 9024 31754 9064
rect 31588 8996 32076 9024
rect 29641 8959 29699 8965
rect 29641 8925 29653 8959
rect 29687 8925 29699 8959
rect 29641 8919 29699 8925
rect 29825 8959 29883 8965
rect 29825 8925 29837 8959
rect 29871 8925 29883 8959
rect 29825 8919 29883 8925
rect 28868 8860 28948 8888
rect 29656 8888 29684 8919
rect 29914 8916 29920 8968
rect 29972 8916 29978 8968
rect 30190 8916 30196 8968
rect 30248 8916 30254 8968
rect 31588 8942 31616 8996
rect 30558 8888 30564 8900
rect 29656 8860 30564 8888
rect 28868 8857 28880 8860
rect 28822 8851 28880 8857
rect 30558 8848 30564 8860
rect 30616 8848 30622 8900
rect 32048 8888 32076 8996
rect 32416 8965 32444 9120
rect 33686 9024 33692 9036
rect 32508 8996 33692 9024
rect 32401 8959 32459 8965
rect 32401 8925 32413 8959
rect 32447 8925 32459 8959
rect 32401 8919 32459 8925
rect 32508 8888 32536 8996
rect 33686 8984 33692 8996
rect 33744 8984 33750 9036
rect 32674 8916 32680 8968
rect 32732 8916 32738 8968
rect 32953 8891 33011 8897
rect 32953 8888 32965 8891
rect 32048 8860 32536 8888
rect 32600 8860 32965 8888
rect 22278 8820 22284 8832
rect 21284 8792 22284 8820
rect 22278 8780 22284 8792
rect 22336 8780 22342 8832
rect 22572 8820 22600 8848
rect 22925 8823 22983 8829
rect 22925 8820 22937 8823
rect 22572 8792 22937 8820
rect 22925 8789 22937 8792
rect 22971 8789 22983 8823
rect 22925 8783 22983 8789
rect 26142 8780 26148 8832
rect 26200 8820 26206 8832
rect 32600 8829 32628 8860
rect 32953 8857 32965 8860
rect 32999 8857 33011 8891
rect 32953 8851 33011 8857
rect 33686 8848 33692 8900
rect 33744 8848 33750 8900
rect 26237 8823 26295 8829
rect 26237 8820 26249 8823
rect 26200 8792 26249 8820
rect 26200 8780 26206 8792
rect 26237 8789 26249 8792
rect 26283 8789 26295 8823
rect 26237 8783 26295 8789
rect 32585 8823 32643 8829
rect 32585 8789 32597 8823
rect 32631 8789 32643 8823
rect 32585 8783 32643 8789
rect 1104 8730 38272 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 38272 8730
rect 1104 8656 38272 8678
rect 4522 8576 4528 8628
rect 4580 8576 4586 8628
rect 10410 8576 10416 8628
rect 10468 8616 10474 8628
rect 12342 8616 12348 8628
rect 10468 8588 12348 8616
rect 10468 8576 10474 8588
rect 12342 8576 12348 8588
rect 12400 8616 12406 8628
rect 14090 8616 14096 8628
rect 12400 8588 14096 8616
rect 12400 8576 12406 8588
rect 14090 8576 14096 8588
rect 14148 8576 14154 8628
rect 16114 8616 16120 8628
rect 14568 8588 16120 8616
rect 4540 8548 4568 8576
rect 6086 8548 6092 8560
rect 4172 8520 4568 8548
rect 5658 8520 6092 8548
rect 4172 8489 4200 8520
rect 6086 8508 6092 8520
rect 6144 8508 6150 8560
rect 6178 8508 6184 8560
rect 6236 8548 6242 8560
rect 11146 8548 11152 8560
rect 6236 8520 11152 8548
rect 6236 8508 6242 8520
rect 11146 8508 11152 8520
rect 11204 8508 11210 8560
rect 12066 8508 12072 8560
rect 12124 8548 12130 8560
rect 14274 8548 14280 8560
rect 12124 8520 14280 8548
rect 12124 8508 12130 8520
rect 14274 8508 14280 8520
rect 14332 8508 14338 8560
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8449 4215 8483
rect 4157 8443 4215 8449
rect 6914 8440 6920 8492
rect 6972 8480 6978 8492
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 6972 8452 7849 8480
rect 6972 8440 6978 8452
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 9585 8483 9643 8489
rect 9585 8449 9597 8483
rect 9631 8480 9643 8483
rect 14458 8480 14464 8492
rect 9631 8452 14464 8480
rect 9631 8449 9643 8452
rect 9585 8443 9643 8449
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8412 4491 8415
rect 4890 8412 4896 8424
rect 4479 8384 4896 8412
rect 4479 8381 4491 8384
rect 4433 8375 4491 8381
rect 4890 8372 4896 8384
rect 4948 8372 4954 8424
rect 10502 8372 10508 8424
rect 10560 8412 10566 8424
rect 14568 8412 14596 8588
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 17681 8619 17739 8625
rect 17681 8585 17693 8619
rect 17727 8616 17739 8619
rect 17862 8616 17868 8628
rect 17727 8588 17868 8616
rect 17727 8585 17739 8588
rect 17681 8579 17739 8585
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 18049 8619 18107 8625
rect 18049 8585 18061 8619
rect 18095 8616 18107 8619
rect 18414 8616 18420 8628
rect 18095 8588 18420 8616
rect 18095 8585 18107 8588
rect 18049 8579 18107 8585
rect 18414 8576 18420 8588
rect 18472 8576 18478 8628
rect 19794 8576 19800 8628
rect 19852 8616 19858 8628
rect 20533 8619 20591 8625
rect 20533 8616 20545 8619
rect 19852 8588 20545 8616
rect 19852 8576 19858 8588
rect 20533 8585 20545 8588
rect 20579 8585 20591 8619
rect 20533 8579 20591 8585
rect 20806 8576 20812 8628
rect 20864 8616 20870 8628
rect 20901 8619 20959 8625
rect 20901 8616 20913 8619
rect 20864 8588 20913 8616
rect 20864 8576 20870 8588
rect 20901 8585 20913 8588
rect 20947 8585 20959 8619
rect 20901 8579 20959 8585
rect 21082 8576 21088 8628
rect 21140 8616 21146 8628
rect 21140 8588 21220 8616
rect 21140 8576 21146 8588
rect 14737 8551 14795 8557
rect 14737 8517 14749 8551
rect 14783 8548 14795 8551
rect 19150 8548 19156 8560
rect 14783 8520 19156 8548
rect 14783 8517 14795 8520
rect 14737 8511 14795 8517
rect 19150 8508 19156 8520
rect 19208 8508 19214 8560
rect 20070 8508 20076 8560
rect 20128 8508 20134 8560
rect 20165 8551 20223 8557
rect 20165 8517 20177 8551
rect 20211 8548 20223 8551
rect 20346 8548 20352 8560
rect 20211 8520 20352 8548
rect 20211 8517 20223 8520
rect 20165 8511 20223 8517
rect 20346 8508 20352 8520
rect 20404 8508 20410 8560
rect 15010 8440 15016 8492
rect 15068 8440 15074 8492
rect 15102 8440 15108 8492
rect 15160 8440 15166 8492
rect 15197 8483 15255 8489
rect 15197 8449 15209 8483
rect 15243 8480 15255 8483
rect 16482 8480 16488 8492
rect 15243 8452 16488 8480
rect 15243 8449 15255 8452
rect 15197 8443 15255 8449
rect 16482 8440 16488 8452
rect 16540 8480 16546 8492
rect 17034 8480 17040 8492
rect 16540 8452 17040 8480
rect 16540 8440 16546 8452
rect 17034 8440 17040 8452
rect 17092 8440 17098 8492
rect 17865 8483 17923 8489
rect 17865 8449 17877 8483
rect 17911 8480 17923 8483
rect 17954 8480 17960 8492
rect 17911 8452 17960 8480
rect 17911 8449 17923 8452
rect 17865 8443 17923 8449
rect 17954 8440 17960 8452
rect 18012 8440 18018 8492
rect 18141 8483 18199 8489
rect 18141 8449 18153 8483
rect 18187 8480 18199 8483
rect 19610 8480 19616 8492
rect 18187 8452 19616 8480
rect 18187 8449 18199 8452
rect 18141 8443 18199 8449
rect 10560 8384 14596 8412
rect 10560 8372 10566 8384
rect 16206 8372 16212 8424
rect 16264 8372 16270 8424
rect 17586 8372 17592 8424
rect 17644 8412 17650 8424
rect 18156 8412 18184 8443
rect 19610 8440 19616 8452
rect 19668 8440 19674 8492
rect 19797 8483 19855 8489
rect 19797 8449 19809 8483
rect 19843 8449 19855 8483
rect 19797 8443 19855 8449
rect 19890 8483 19948 8489
rect 19890 8449 19902 8483
rect 19936 8470 19948 8483
rect 19936 8449 20024 8470
rect 19890 8443 20024 8449
rect 17644 8384 18184 8412
rect 19812 8412 19840 8443
rect 19905 8442 20024 8443
rect 19996 8412 20024 8442
rect 20254 8440 20260 8492
rect 20312 8489 20318 8492
rect 20312 8480 20320 8489
rect 20717 8483 20775 8489
rect 20312 8452 20357 8480
rect 20312 8443 20320 8452
rect 20717 8449 20729 8483
rect 20763 8449 20775 8483
rect 20717 8443 20775 8449
rect 20312 8440 20318 8443
rect 19812 8384 19932 8412
rect 19996 8384 20208 8412
rect 17644 8372 17650 8384
rect 12158 8304 12164 8356
rect 12216 8344 12222 8356
rect 13078 8344 13084 8356
rect 12216 8316 13084 8344
rect 12216 8304 12222 8316
rect 13078 8304 13084 8316
rect 13136 8304 13142 8356
rect 13446 8304 13452 8356
rect 13504 8344 13510 8356
rect 13814 8344 13820 8356
rect 13504 8316 13820 8344
rect 13504 8304 13510 8316
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 14829 8347 14887 8353
rect 14829 8313 14841 8347
rect 14875 8313 14887 8347
rect 16224 8344 16252 8372
rect 19904 8356 19932 8384
rect 20180 8356 20208 8384
rect 16224 8316 19840 8344
rect 14829 8307 14887 8313
rect 7190 8236 7196 8288
rect 7248 8276 7254 8288
rect 11606 8276 11612 8288
rect 7248 8248 11612 8276
rect 7248 8236 7254 8248
rect 11606 8236 11612 8248
rect 11664 8276 11670 8288
rect 14844 8276 14872 8307
rect 15010 8276 15016 8288
rect 11664 8248 15016 8276
rect 11664 8236 11670 8248
rect 15010 8236 15016 8248
rect 15068 8236 15074 8288
rect 15378 8236 15384 8288
rect 15436 8236 15442 8288
rect 15654 8236 15660 8288
rect 15712 8276 15718 8288
rect 16298 8276 16304 8288
rect 15712 8248 16304 8276
rect 15712 8236 15718 8248
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 16850 8236 16856 8288
rect 16908 8276 16914 8288
rect 19610 8276 19616 8288
rect 16908 8248 19616 8276
rect 16908 8236 16914 8248
rect 19610 8236 19616 8248
rect 19668 8236 19674 8288
rect 19812 8276 19840 8316
rect 19886 8304 19892 8356
rect 19944 8304 19950 8356
rect 20162 8304 20168 8356
rect 20220 8304 20226 8356
rect 20441 8347 20499 8353
rect 20441 8313 20453 8347
rect 20487 8344 20499 8347
rect 20732 8344 20760 8443
rect 20898 8440 20904 8492
rect 20956 8486 20962 8492
rect 20993 8486 21051 8489
rect 20956 8483 21051 8486
rect 20956 8458 21005 8483
rect 20956 8440 20962 8458
rect 20993 8449 21005 8458
rect 21039 8449 21051 8483
rect 20993 8443 21051 8449
rect 21082 8440 21088 8492
rect 21140 8440 21146 8492
rect 21192 8412 21220 8588
rect 21450 8576 21456 8628
rect 21508 8616 21514 8628
rect 22373 8619 22431 8625
rect 21508 8588 22048 8616
rect 21508 8576 21514 8588
rect 21266 8508 21272 8560
rect 21324 8508 21330 8560
rect 21910 8548 21916 8560
rect 21376 8520 21916 8548
rect 21376 8489 21404 8520
rect 21910 8508 21916 8520
rect 21968 8508 21974 8560
rect 22020 8557 22048 8588
rect 22373 8585 22385 8619
rect 22419 8616 22431 8619
rect 22462 8616 22468 8628
rect 22419 8588 22468 8616
rect 22419 8585 22431 8588
rect 22373 8579 22431 8585
rect 22462 8576 22468 8588
rect 22520 8576 22526 8628
rect 22557 8619 22615 8625
rect 22557 8585 22569 8619
rect 22603 8616 22615 8619
rect 22646 8616 22652 8628
rect 22603 8588 22652 8616
rect 22603 8585 22615 8588
rect 22557 8579 22615 8585
rect 22646 8576 22652 8588
rect 22704 8576 22710 8628
rect 23201 8619 23259 8625
rect 23201 8585 23213 8619
rect 23247 8585 23259 8619
rect 26050 8616 26056 8628
rect 23201 8579 23259 8585
rect 25240 8588 26056 8616
rect 22005 8551 22063 8557
rect 22005 8517 22017 8551
rect 22051 8517 22063 8551
rect 22005 8511 22063 8517
rect 22278 8508 22284 8560
rect 22336 8548 22342 8560
rect 23216 8548 23244 8579
rect 22336 8520 22876 8548
rect 22336 8508 22342 8520
rect 22848 8492 22876 8520
rect 23032 8520 23244 8548
rect 21361 8483 21419 8489
rect 21361 8449 21373 8483
rect 21407 8449 21419 8483
rect 21361 8443 21419 8449
rect 21450 8440 21456 8492
rect 21508 8440 21514 8492
rect 21634 8440 21640 8492
rect 21692 8440 21698 8492
rect 21821 8483 21879 8489
rect 21821 8449 21833 8483
rect 21867 8449 21879 8483
rect 22097 8483 22155 8489
rect 22097 8480 22109 8483
rect 21821 8443 21879 8449
rect 21928 8452 22109 8480
rect 21468 8412 21496 8440
rect 21192 8384 21496 8412
rect 21376 8344 21404 8384
rect 21652 8353 21680 8440
rect 20487 8316 20760 8344
rect 20916 8316 21404 8344
rect 21637 8347 21695 8353
rect 20487 8313 20499 8316
rect 20441 8307 20499 8313
rect 20916 8276 20944 8316
rect 21637 8313 21649 8347
rect 21683 8313 21695 8347
rect 21836 8344 21864 8443
rect 21928 8424 21956 8452
rect 22097 8449 22109 8452
rect 22143 8449 22155 8483
rect 22097 8443 22155 8449
rect 22189 8483 22247 8489
rect 22189 8449 22201 8483
rect 22235 8449 22247 8483
rect 22189 8443 22247 8449
rect 21910 8372 21916 8424
rect 21968 8372 21974 8424
rect 22204 8412 22232 8443
rect 22738 8440 22744 8492
rect 22796 8440 22802 8492
rect 22830 8440 22836 8492
rect 22888 8440 22894 8492
rect 23032 8489 23060 8520
rect 23474 8508 23480 8560
rect 23532 8508 23538 8560
rect 23767 8520 23980 8548
rect 23017 8483 23075 8489
rect 23017 8449 23029 8483
rect 23063 8449 23075 8483
rect 23017 8443 23075 8449
rect 23106 8440 23112 8492
rect 23164 8440 23170 8492
rect 23290 8440 23296 8492
rect 23348 8489 23354 8492
rect 23348 8483 23397 8489
rect 23348 8449 23351 8483
rect 23385 8449 23397 8483
rect 23348 8443 23397 8449
rect 23348 8440 23354 8443
rect 23566 8440 23572 8492
rect 23624 8440 23630 8492
rect 23767 8489 23795 8520
rect 23952 8492 23980 8520
rect 23752 8483 23810 8489
rect 23752 8449 23764 8483
rect 23798 8449 23810 8483
rect 23752 8443 23810 8449
rect 23842 8440 23848 8492
rect 23900 8440 23906 8492
rect 23934 8440 23940 8492
rect 23992 8440 23998 8492
rect 24026 8440 24032 8492
rect 24084 8440 24090 8492
rect 25240 8489 25268 8588
rect 26050 8576 26056 8588
rect 26108 8576 26114 8628
rect 26142 8576 26148 8628
rect 26200 8576 26206 8628
rect 28353 8619 28411 8625
rect 28353 8585 28365 8619
rect 28399 8616 28411 8619
rect 29914 8616 29920 8628
rect 28399 8588 29920 8616
rect 28399 8585 28411 8588
rect 28353 8579 28411 8585
rect 29914 8576 29920 8588
rect 29972 8576 29978 8628
rect 30190 8576 30196 8628
rect 30248 8616 30254 8628
rect 30377 8619 30435 8625
rect 30377 8616 30389 8619
rect 30248 8588 30389 8616
rect 30248 8576 30254 8588
rect 30377 8585 30389 8588
rect 30423 8585 30435 8619
rect 30377 8579 30435 8585
rect 31662 8576 31668 8628
rect 31720 8576 31726 8628
rect 32674 8576 32680 8628
rect 32732 8616 32738 8628
rect 32861 8619 32919 8625
rect 32861 8616 32873 8619
rect 32732 8588 32873 8616
rect 32732 8576 32738 8588
rect 32861 8585 32873 8588
rect 32907 8585 32919 8619
rect 32861 8579 32919 8585
rect 25774 8508 25780 8560
rect 25832 8548 25838 8560
rect 25832 8520 25907 8548
rect 25832 8508 25838 8520
rect 25225 8483 25283 8489
rect 25225 8480 25237 8483
rect 24504 8452 25237 8480
rect 24044 8412 24072 8440
rect 22204 8384 24072 8412
rect 22554 8344 22560 8356
rect 21836 8316 22560 8344
rect 21637 8307 21695 8313
rect 22554 8304 22560 8316
rect 22612 8304 22618 8356
rect 22646 8304 22652 8356
rect 22704 8344 22710 8356
rect 24504 8344 24532 8452
rect 25225 8449 25237 8452
rect 25271 8449 25283 8483
rect 25225 8443 25283 8449
rect 25409 8483 25467 8489
rect 25409 8449 25421 8483
rect 25455 8449 25467 8483
rect 25409 8443 25467 8449
rect 25685 8483 25743 8489
rect 25685 8449 25697 8483
rect 25731 8449 25743 8483
rect 25685 8443 25743 8449
rect 25038 8372 25044 8424
rect 25096 8412 25102 8424
rect 25424 8412 25452 8443
rect 25096 8384 25452 8412
rect 25096 8372 25102 8384
rect 22704 8316 24532 8344
rect 25700 8344 25728 8443
rect 25879 8412 25907 8520
rect 25958 8440 25964 8492
rect 26016 8440 26022 8492
rect 26160 8489 26188 8576
rect 26786 8508 26792 8560
rect 26844 8508 26850 8560
rect 27890 8557 27896 8560
rect 27867 8551 27896 8557
rect 27867 8517 27879 8551
rect 27867 8511 27896 8517
rect 27890 8508 27896 8511
rect 27948 8508 27954 8560
rect 28718 8508 28724 8560
rect 28776 8508 28782 8560
rect 28902 8548 28908 8560
rect 28863 8520 28908 8548
rect 28902 8508 28908 8520
rect 28960 8548 28966 8560
rect 30926 8548 30932 8560
rect 28960 8520 30932 8548
rect 28960 8508 28966 8520
rect 30926 8508 30932 8520
rect 30984 8508 30990 8560
rect 31680 8548 31708 8576
rect 31680 8520 32996 8548
rect 26154 8483 26212 8489
rect 26154 8449 26166 8483
rect 26200 8449 26212 8483
rect 26154 8443 26212 8449
rect 26326 8440 26332 8492
rect 26384 8480 26390 8492
rect 26973 8483 27031 8489
rect 26973 8480 26985 8483
rect 26384 8452 26985 8480
rect 26384 8440 26390 8452
rect 26973 8449 26985 8452
rect 27019 8449 27031 8483
rect 26973 8443 27031 8449
rect 27157 8483 27215 8489
rect 27157 8449 27169 8483
rect 27203 8480 27215 8483
rect 27430 8480 27436 8492
rect 27203 8452 27436 8480
rect 27203 8449 27215 8452
rect 27157 8443 27215 8449
rect 27172 8412 27200 8443
rect 27430 8440 27436 8452
rect 27488 8440 27494 8492
rect 27706 8440 27712 8492
rect 27764 8440 27770 8492
rect 27982 8440 27988 8492
rect 28040 8440 28046 8492
rect 28077 8483 28135 8489
rect 28077 8449 28089 8483
rect 28123 8449 28135 8483
rect 28077 8443 28135 8449
rect 25879 8384 27200 8412
rect 26973 8347 27031 8353
rect 26973 8344 26985 8347
rect 25700 8316 26985 8344
rect 22704 8304 22710 8316
rect 26973 8313 26985 8316
rect 27019 8313 27031 8347
rect 27724 8344 27752 8440
rect 28092 8412 28120 8443
rect 28166 8440 28172 8492
rect 28224 8440 28230 8492
rect 28258 8440 28264 8492
rect 28316 8480 28322 8492
rect 28501 8483 28559 8489
rect 28501 8480 28513 8483
rect 28316 8452 28513 8480
rect 28316 8440 28322 8452
rect 28501 8449 28513 8452
rect 28547 8449 28559 8483
rect 28501 8443 28559 8449
rect 28626 8440 28632 8492
rect 28684 8440 28690 8492
rect 30469 8483 30527 8489
rect 30469 8449 30481 8483
rect 30515 8480 30527 8483
rect 31846 8480 31852 8492
rect 30515 8452 31852 8480
rect 30515 8449 30527 8452
rect 30469 8443 30527 8449
rect 31846 8440 31852 8452
rect 31904 8440 31910 8492
rect 32968 8489 32996 8520
rect 32953 8483 33011 8489
rect 32953 8449 32965 8483
rect 32999 8449 33011 8483
rect 32953 8443 33011 8449
rect 28813 8415 28871 8421
rect 28813 8412 28825 8415
rect 28092 8384 28825 8412
rect 28813 8381 28825 8384
rect 28859 8381 28871 8415
rect 28813 8375 28871 8381
rect 28350 8344 28356 8356
rect 27724 8316 28356 8344
rect 26973 8307 27031 8313
rect 28350 8304 28356 8316
rect 28408 8304 28414 8356
rect 19812 8248 20944 8276
rect 21174 8236 21180 8288
rect 21232 8276 21238 8288
rect 23566 8276 23572 8288
rect 21232 8248 23572 8276
rect 21232 8236 21238 8248
rect 23566 8236 23572 8248
rect 23624 8236 23630 8288
rect 23750 8236 23756 8288
rect 23808 8276 23814 8288
rect 31662 8276 31668 8288
rect 23808 8248 31668 8276
rect 23808 8236 23814 8248
rect 31662 8236 31668 8248
rect 31720 8236 31726 8288
rect 1104 8186 38272 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38272 8186
rect 1104 8112 38272 8134
rect 4890 8032 4896 8084
rect 4948 8032 4954 8084
rect 6822 8032 6828 8084
rect 6880 8032 6886 8084
rect 7926 8032 7932 8084
rect 7984 8072 7990 8084
rect 10962 8072 10968 8084
rect 7984 8044 10968 8072
rect 7984 8032 7990 8044
rect 5353 8007 5411 8013
rect 5353 7973 5365 8007
rect 5399 7973 5411 8007
rect 6840 8004 6868 8032
rect 5353 7967 5411 7973
rect 6012 7976 6868 8004
rect 5077 7871 5135 7877
rect 5077 7837 5089 7871
rect 5123 7868 5135 7871
rect 5368 7868 5396 7967
rect 6012 7945 6040 7976
rect 5997 7939 6055 7945
rect 5997 7905 6009 7939
rect 6043 7905 6055 7939
rect 5997 7899 6055 7905
rect 5123 7840 5396 7868
rect 5123 7837 5135 7840
rect 5077 7831 5135 7837
rect 5718 7828 5724 7880
rect 5776 7868 5782 7880
rect 6178 7868 6184 7880
rect 5776 7840 6184 7868
rect 5776 7828 5782 7840
rect 6178 7828 6184 7840
rect 6236 7828 6242 7880
rect 6730 7828 6736 7880
rect 6788 7828 6794 7880
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 6871 7840 7021 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 7009 7837 7021 7840
rect 7055 7837 7067 7871
rect 8404 7854 8432 8044
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 11422 8032 11428 8084
rect 11480 8072 11486 8084
rect 11517 8075 11575 8081
rect 11517 8072 11529 8075
rect 11480 8044 11529 8072
rect 11480 8032 11486 8044
rect 11517 8041 11529 8044
rect 11563 8041 11575 8075
rect 11517 8035 11575 8041
rect 13906 8032 13912 8084
rect 13964 8072 13970 8084
rect 14093 8075 14151 8081
rect 14093 8072 14105 8075
rect 13964 8044 14105 8072
rect 13964 8032 13970 8044
rect 14093 8041 14105 8044
rect 14139 8041 14151 8075
rect 14093 8035 14151 8041
rect 14826 8032 14832 8084
rect 14884 8072 14890 8084
rect 15102 8072 15108 8084
rect 14884 8044 15108 8072
rect 14884 8032 14890 8044
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 15657 8075 15715 8081
rect 15657 8041 15669 8075
rect 15703 8072 15715 8075
rect 16393 8075 16451 8081
rect 16393 8072 16405 8075
rect 15703 8044 16405 8072
rect 15703 8041 15715 8044
rect 15657 8035 15715 8041
rect 16393 8041 16405 8044
rect 16439 8041 16451 8075
rect 16393 8035 16451 8041
rect 16758 8032 16764 8084
rect 16816 8032 16822 8084
rect 17310 8032 17316 8084
rect 17368 8072 17374 8084
rect 17368 8044 17724 8072
rect 17368 8032 17374 8044
rect 9950 7964 9956 8016
rect 10008 8004 10014 8016
rect 10226 8004 10232 8016
rect 10008 7976 10232 8004
rect 10008 7964 10014 7976
rect 10226 7964 10232 7976
rect 10284 8004 10290 8016
rect 10284 7976 10456 8004
rect 10284 7964 10290 7976
rect 8662 7896 8668 7948
rect 8720 7936 8726 7948
rect 8757 7939 8815 7945
rect 8757 7936 8769 7939
rect 8720 7908 8769 7936
rect 8720 7896 8726 7908
rect 8757 7905 8769 7908
rect 8803 7936 8815 7939
rect 10318 7936 10324 7948
rect 8803 7908 10324 7936
rect 8803 7905 8815 7908
rect 8757 7899 8815 7905
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 10428 7945 10456 7976
rect 15010 7964 15016 8016
rect 15068 8004 15074 8016
rect 17034 8004 17040 8016
rect 15068 7976 17040 8004
rect 15068 7964 15074 7976
rect 17034 7964 17040 7976
rect 17092 8004 17098 8016
rect 17092 7976 17632 8004
rect 17092 7964 17098 7976
rect 10413 7939 10471 7945
rect 10413 7905 10425 7939
rect 10459 7905 10471 7939
rect 12437 7939 12495 7945
rect 10413 7899 10471 7905
rect 11624 7908 11836 7936
rect 11624 7880 11652 7908
rect 9401 7871 9459 7877
rect 9401 7868 9413 7871
rect 7009 7831 7067 7837
rect 8956 7840 9413 7868
rect 7282 7760 7288 7812
rect 7340 7760 7346 7812
rect 8956 7744 8984 7840
rect 9401 7837 9413 7840
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7868 9735 7871
rect 9723 7840 9812 7868
rect 9723 7837 9735 7840
rect 9677 7831 9735 7837
rect 5813 7735 5871 7741
rect 5813 7701 5825 7735
rect 5859 7732 5871 7735
rect 6546 7732 6552 7744
rect 5859 7704 6552 7732
rect 5859 7701 5871 7704
rect 5813 7695 5871 7701
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 8938 7692 8944 7744
rect 8996 7692 9002 7744
rect 9306 7692 9312 7744
rect 9364 7692 9370 7744
rect 9490 7692 9496 7744
rect 9548 7692 9554 7744
rect 9784 7741 9812 7840
rect 11606 7828 11612 7880
rect 11664 7828 11670 7880
rect 11698 7828 11704 7880
rect 11756 7828 11762 7880
rect 11808 7877 11836 7908
rect 12437 7905 12449 7939
rect 12483 7936 12495 7939
rect 12894 7936 12900 7948
rect 12483 7908 12900 7936
rect 12483 7905 12495 7908
rect 12437 7899 12495 7905
rect 12894 7896 12900 7908
rect 12952 7896 12958 7948
rect 16574 7936 16580 7948
rect 13832 7908 16580 7936
rect 11793 7871 11851 7877
rect 11793 7837 11805 7871
rect 11839 7837 11851 7871
rect 11793 7831 11851 7837
rect 11974 7828 11980 7880
rect 12032 7828 12038 7880
rect 12069 7871 12127 7877
rect 12069 7837 12081 7871
rect 12115 7837 12127 7871
rect 12069 7831 12127 7837
rect 10134 7760 10140 7812
rect 10192 7760 10198 7812
rect 12084 7800 12112 7831
rect 12158 7828 12164 7880
rect 12216 7828 12222 7880
rect 13538 7828 13544 7880
rect 13596 7828 13602 7880
rect 12342 7800 12348 7812
rect 12084 7772 12348 7800
rect 12342 7760 12348 7772
rect 12400 7760 12406 7812
rect 9769 7735 9827 7741
rect 9769 7701 9781 7735
rect 9815 7701 9827 7735
rect 9769 7695 9827 7701
rect 10229 7735 10287 7741
rect 10229 7701 10241 7735
rect 10275 7732 10287 7735
rect 10870 7732 10876 7744
rect 10275 7704 10876 7732
rect 10275 7701 10287 7704
rect 10229 7695 10287 7701
rect 10870 7692 10876 7704
rect 10928 7692 10934 7744
rect 11698 7692 11704 7744
rect 11756 7732 11762 7744
rect 13832 7732 13860 7908
rect 14737 7871 14795 7877
rect 14737 7837 14749 7871
rect 14783 7837 14795 7871
rect 14737 7831 14795 7837
rect 14752 7800 14780 7831
rect 14826 7828 14832 7880
rect 14884 7868 14890 7880
rect 15105 7871 15163 7877
rect 15105 7868 15117 7871
rect 14884 7840 15117 7868
rect 14884 7828 14890 7840
rect 15105 7837 15117 7840
rect 15151 7837 15163 7871
rect 15105 7831 15163 7837
rect 15194 7828 15200 7880
rect 15252 7828 15258 7880
rect 15470 7828 15476 7880
rect 15528 7828 15534 7880
rect 15764 7877 15792 7908
rect 16574 7896 16580 7908
rect 16632 7896 16638 7948
rect 15749 7871 15807 7877
rect 15749 7837 15761 7871
rect 15795 7837 15807 7871
rect 15749 7831 15807 7837
rect 15838 7828 15844 7880
rect 15896 7868 15902 7880
rect 15933 7871 15991 7877
rect 15933 7868 15945 7871
rect 15896 7840 15945 7868
rect 15896 7828 15902 7840
rect 15933 7837 15945 7840
rect 15979 7837 15991 7871
rect 15933 7831 15991 7837
rect 16117 7871 16175 7877
rect 16117 7837 16129 7871
rect 16163 7868 16175 7871
rect 16206 7868 16212 7880
rect 16163 7840 16212 7868
rect 16163 7837 16175 7840
rect 16117 7831 16175 7837
rect 16206 7828 16212 7840
rect 16264 7828 16270 7880
rect 16298 7828 16304 7880
rect 16356 7868 16362 7880
rect 16393 7871 16451 7877
rect 16393 7868 16405 7871
rect 16356 7840 16405 7868
rect 16356 7828 16362 7840
rect 16393 7837 16405 7840
rect 16439 7837 16451 7871
rect 16393 7831 16451 7837
rect 16482 7828 16488 7880
rect 16540 7828 16546 7880
rect 16850 7828 16856 7880
rect 16908 7828 16914 7880
rect 17126 7828 17132 7880
rect 17184 7868 17190 7880
rect 17313 7871 17371 7877
rect 17184 7862 17264 7868
rect 17313 7862 17325 7871
rect 17184 7840 17325 7862
rect 17184 7828 17190 7840
rect 17236 7837 17325 7840
rect 17359 7837 17371 7871
rect 17236 7834 17371 7837
rect 17313 7831 17371 7834
rect 17406 7871 17464 7877
rect 17406 7837 17418 7871
rect 17452 7864 17464 7871
rect 17604 7868 17632 7976
rect 17696 7877 17724 8044
rect 17954 8032 17960 8084
rect 18012 8032 18018 8084
rect 18230 8032 18236 8084
rect 18288 8032 18294 8084
rect 18690 8032 18696 8084
rect 18748 8032 18754 8084
rect 20349 8075 20407 8081
rect 19904 8044 20300 8072
rect 18248 8004 18276 8032
rect 18156 7976 18276 8004
rect 17862 7877 17868 7880
rect 17512 7864 17632 7868
rect 17452 7840 17632 7864
rect 17681 7871 17739 7877
rect 17452 7837 17540 7840
rect 17406 7836 17540 7837
rect 17681 7837 17693 7871
rect 17727 7837 17739 7871
rect 17406 7831 17464 7836
rect 17681 7831 17739 7837
rect 17819 7871 17868 7877
rect 17819 7837 17831 7871
rect 17865 7837 17868 7871
rect 17819 7831 17868 7837
rect 17862 7828 17868 7831
rect 17920 7828 17926 7880
rect 18156 7877 18184 7976
rect 18230 7896 18236 7948
rect 18288 7896 18294 7948
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7837 18199 7871
rect 18141 7831 18199 7837
rect 18417 7871 18475 7877
rect 18417 7837 18429 7871
rect 18463 7837 18475 7871
rect 18417 7831 18475 7837
rect 15212 7800 15240 7828
rect 13924 7772 15240 7800
rect 13924 7741 13952 7772
rect 15286 7760 15292 7812
rect 15344 7760 15350 7812
rect 15381 7803 15439 7809
rect 15381 7769 15393 7803
rect 15427 7769 15439 7803
rect 15381 7763 15439 7769
rect 11756 7704 13860 7732
rect 13909 7735 13967 7741
rect 11756 7692 11762 7704
rect 13909 7701 13921 7735
rect 13955 7701 13967 7735
rect 13909 7695 13967 7701
rect 14090 7692 14096 7744
rect 14148 7732 14154 7744
rect 15396 7732 15424 7763
rect 15562 7760 15568 7812
rect 15620 7800 15626 7812
rect 16025 7803 16083 7809
rect 16025 7800 16037 7803
rect 15620 7772 16037 7800
rect 15620 7760 15626 7772
rect 16025 7769 16037 7772
rect 16071 7769 16083 7803
rect 16868 7800 16896 7828
rect 17589 7803 17647 7809
rect 17589 7800 17601 7803
rect 16025 7763 16083 7769
rect 16132 7772 16436 7800
rect 16868 7772 17601 7800
rect 16132 7732 16160 7772
rect 14148 7704 16160 7732
rect 14148 7692 14154 7704
rect 16298 7692 16304 7744
rect 16356 7692 16362 7744
rect 16408 7732 16436 7772
rect 17589 7769 17601 7772
rect 17635 7769 17647 7803
rect 17589 7763 17647 7769
rect 17954 7760 17960 7812
rect 18012 7800 18018 7812
rect 18432 7800 18460 7831
rect 18506 7828 18512 7880
rect 18564 7828 18570 7880
rect 19904 7877 19932 8044
rect 20162 7964 20168 8016
rect 20220 7964 20226 8016
rect 20272 8004 20300 8044
rect 20349 8041 20361 8075
rect 20395 8072 20407 8075
rect 20530 8072 20536 8084
rect 20395 8044 20536 8072
rect 20395 8041 20407 8044
rect 20349 8035 20407 8041
rect 20530 8032 20536 8044
rect 20588 8032 20594 8084
rect 21818 8072 21824 8084
rect 20824 8044 21824 8072
rect 20441 8007 20499 8013
rect 20441 8004 20453 8007
rect 20272 7976 20453 8004
rect 20441 7973 20453 7976
rect 20487 7973 20499 8007
rect 20441 7967 20499 7973
rect 20180 7936 20208 7964
rect 20824 7936 20852 8044
rect 21818 8032 21824 8044
rect 21876 8032 21882 8084
rect 22925 8075 22983 8081
rect 22925 8041 22937 8075
rect 22971 8041 22983 8075
rect 22925 8035 22983 8041
rect 23109 8075 23167 8081
rect 23109 8041 23121 8075
rect 23155 8072 23167 8075
rect 23842 8072 23848 8084
rect 23155 8044 23848 8072
rect 23155 8041 23167 8044
rect 23109 8035 23167 8041
rect 22738 8004 22744 8016
rect 20088 7908 20852 7936
rect 20916 7976 22744 8004
rect 20088 7877 20116 7908
rect 19797 7871 19855 7877
rect 19797 7868 19809 7871
rect 19306 7840 19809 7868
rect 18012 7772 18460 7800
rect 18012 7760 18018 7772
rect 18690 7760 18696 7812
rect 18748 7800 18754 7812
rect 19306 7800 19334 7840
rect 19797 7837 19809 7840
rect 19843 7837 19855 7871
rect 19797 7831 19855 7837
rect 19889 7871 19947 7877
rect 19889 7837 19901 7871
rect 19935 7837 19947 7871
rect 19889 7831 19947 7837
rect 20073 7871 20131 7877
rect 20073 7837 20085 7871
rect 20119 7837 20131 7871
rect 20073 7831 20131 7837
rect 20165 7871 20223 7877
rect 20165 7837 20177 7871
rect 20211 7868 20223 7871
rect 20438 7868 20444 7880
rect 20211 7840 20444 7868
rect 20211 7837 20223 7840
rect 20165 7831 20223 7837
rect 20438 7828 20444 7840
rect 20496 7828 20502 7880
rect 20530 7828 20536 7880
rect 20588 7878 20594 7880
rect 20588 7877 20668 7878
rect 20588 7871 20683 7877
rect 20588 7850 20637 7871
rect 20588 7828 20594 7850
rect 20625 7837 20637 7850
rect 20671 7837 20683 7871
rect 20625 7831 20683 7837
rect 20809 7871 20867 7877
rect 20809 7837 20821 7871
rect 20855 7868 20867 7871
rect 20916 7868 20944 7976
rect 22738 7964 22744 7976
rect 22796 7964 22802 8016
rect 22940 8004 22968 8035
rect 23842 8032 23848 8044
rect 23900 8032 23906 8084
rect 24578 8032 24584 8084
rect 24636 8072 24642 8084
rect 24765 8075 24823 8081
rect 24765 8072 24777 8075
rect 24636 8044 24777 8072
rect 24636 8032 24642 8044
rect 24765 8041 24777 8044
rect 24811 8041 24823 8075
rect 24765 8035 24823 8041
rect 27893 8075 27951 8081
rect 27893 8041 27905 8075
rect 27939 8072 27951 8075
rect 27982 8072 27988 8084
rect 27939 8044 27988 8072
rect 27939 8041 27951 8044
rect 27893 8035 27951 8041
rect 27982 8032 27988 8044
rect 28040 8032 28046 8084
rect 28810 8032 28816 8084
rect 28868 8072 28874 8084
rect 29549 8075 29607 8081
rect 29549 8072 29561 8075
rect 28868 8044 29561 8072
rect 28868 8032 28874 8044
rect 29549 8041 29561 8044
rect 29595 8041 29607 8075
rect 29549 8035 29607 8041
rect 29730 8032 29736 8084
rect 29788 8032 29794 8084
rect 30558 8032 30564 8084
rect 30616 8032 30622 8084
rect 30926 8032 30932 8084
rect 30984 8032 30990 8084
rect 23382 8004 23388 8016
rect 22940 7976 23388 8004
rect 23382 7964 23388 7976
rect 23440 8004 23446 8016
rect 27246 8004 27252 8016
rect 23440 7976 27252 8004
rect 23440 7964 23446 7976
rect 27246 7964 27252 7976
rect 27304 7964 27310 8016
rect 21358 7896 21364 7948
rect 21416 7936 21422 7948
rect 23106 7936 23112 7948
rect 21416 7908 23112 7936
rect 21416 7896 21422 7908
rect 23106 7896 23112 7908
rect 23164 7936 23170 7948
rect 23164 7908 25268 7936
rect 23164 7896 23170 7908
rect 20855 7840 20944 7868
rect 20993 7871 21051 7877
rect 20855 7837 20867 7840
rect 20809 7831 20867 7837
rect 20993 7837 21005 7871
rect 21039 7868 21051 7871
rect 21082 7868 21088 7880
rect 21039 7840 21088 7868
rect 21039 7837 21051 7840
rect 20993 7831 21051 7837
rect 21082 7828 21088 7840
rect 21140 7828 21146 7880
rect 24946 7828 24952 7880
rect 25004 7828 25010 7880
rect 25240 7877 25268 7908
rect 25774 7896 25780 7948
rect 25832 7936 25838 7948
rect 28902 7936 28908 7948
rect 25832 7908 28908 7936
rect 25832 7896 25838 7908
rect 28902 7896 28908 7908
rect 28960 7896 28966 7948
rect 29748 7936 29776 8032
rect 30944 8004 30972 8032
rect 30392 7976 30972 8004
rect 29748 7908 30144 7936
rect 25225 7871 25283 7877
rect 25225 7837 25237 7871
rect 25271 7868 25283 7871
rect 25406 7868 25412 7880
rect 25271 7840 25412 7868
rect 25271 7837 25283 7840
rect 25225 7831 25283 7837
rect 25406 7828 25412 7840
rect 25464 7828 25470 7880
rect 27798 7828 27804 7880
rect 27856 7828 27862 7880
rect 27985 7871 28043 7877
rect 27985 7868 27997 7871
rect 27908 7840 27997 7868
rect 18748 7772 19334 7800
rect 20717 7803 20775 7809
rect 18748 7760 18754 7772
rect 20717 7769 20729 7803
rect 20763 7800 20775 7803
rect 20898 7800 20904 7812
rect 20763 7772 20904 7800
rect 20763 7769 20775 7772
rect 20717 7763 20775 7769
rect 20898 7760 20904 7772
rect 20956 7800 20962 7812
rect 21910 7800 21916 7812
rect 20956 7772 21916 7800
rect 20956 7760 20962 7772
rect 21910 7760 21916 7772
rect 21968 7760 21974 7812
rect 22462 7760 22468 7812
rect 22520 7800 22526 7812
rect 22741 7803 22799 7809
rect 22741 7800 22753 7803
rect 22520 7772 22753 7800
rect 22520 7760 22526 7772
rect 22741 7769 22753 7772
rect 22787 7769 22799 7803
rect 22741 7763 22799 7769
rect 22957 7803 23015 7809
rect 22957 7769 22969 7803
rect 23003 7800 23015 7803
rect 23003 7772 27844 7800
rect 23003 7769 23015 7772
rect 22957 7763 23015 7769
rect 18414 7732 18420 7744
rect 16408 7704 18420 7732
rect 18414 7692 18420 7704
rect 18472 7692 18478 7744
rect 19058 7692 19064 7744
rect 19116 7732 19122 7744
rect 21266 7732 21272 7744
rect 19116 7704 21272 7732
rect 19116 7692 19122 7704
rect 21266 7692 21272 7704
rect 21324 7732 21330 7744
rect 22972 7732 23000 7763
rect 27816 7744 27844 7772
rect 27908 7744 27936 7840
rect 27985 7837 27997 7840
rect 28031 7837 28043 7871
rect 27985 7831 28043 7837
rect 29638 7828 29644 7880
rect 29696 7868 29702 7880
rect 29733 7871 29791 7877
rect 29733 7868 29745 7871
rect 29696 7840 29745 7868
rect 29696 7828 29702 7840
rect 29733 7837 29745 7840
rect 29779 7837 29791 7871
rect 29733 7831 29791 7837
rect 29825 7871 29883 7877
rect 29825 7837 29837 7871
rect 29871 7837 29883 7871
rect 29825 7831 29883 7837
rect 29840 7800 29868 7831
rect 30006 7828 30012 7880
rect 30064 7828 30070 7880
rect 30116 7877 30144 7908
rect 30392 7877 30420 7976
rect 30561 7939 30619 7945
rect 30561 7905 30573 7939
rect 30607 7936 30619 7939
rect 30834 7936 30840 7948
rect 30607 7908 30840 7936
rect 30607 7905 30619 7908
rect 30561 7899 30619 7905
rect 30834 7896 30840 7908
rect 30892 7896 30898 7948
rect 30101 7871 30159 7877
rect 30101 7837 30113 7871
rect 30147 7868 30159 7871
rect 30193 7871 30251 7877
rect 30193 7868 30205 7871
rect 30147 7840 30205 7868
rect 30147 7837 30159 7840
rect 30101 7831 30159 7837
rect 30193 7837 30205 7840
rect 30239 7837 30251 7871
rect 30193 7831 30251 7837
rect 30377 7871 30435 7877
rect 30377 7837 30389 7871
rect 30423 7837 30435 7871
rect 30377 7831 30435 7837
rect 30466 7828 30472 7880
rect 30524 7828 30530 7880
rect 31846 7828 31852 7880
rect 31904 7868 31910 7880
rect 32401 7871 32459 7877
rect 32401 7868 32413 7871
rect 31904 7840 32413 7868
rect 31904 7828 31910 7840
rect 32401 7837 32413 7840
rect 32447 7837 32459 7871
rect 32401 7831 32459 7837
rect 29748 7772 29868 7800
rect 29748 7744 29776 7772
rect 31662 7760 31668 7812
rect 31720 7800 31726 7812
rect 33226 7800 33232 7812
rect 31720 7772 33232 7800
rect 31720 7760 31726 7772
rect 33226 7760 33232 7772
rect 33284 7760 33290 7812
rect 21324 7704 23000 7732
rect 25133 7735 25191 7741
rect 21324 7692 21330 7704
rect 25133 7701 25145 7735
rect 25179 7732 25191 7735
rect 26142 7732 26148 7744
rect 25179 7704 26148 7732
rect 25179 7701 25191 7704
rect 25133 7695 25191 7701
rect 26142 7692 26148 7704
rect 26200 7692 26206 7744
rect 27798 7692 27804 7744
rect 27856 7692 27862 7744
rect 27890 7692 27896 7744
rect 27948 7692 27954 7744
rect 29730 7692 29736 7744
rect 29788 7692 29794 7744
rect 32306 7692 32312 7744
rect 32364 7692 32370 7744
rect 1104 7642 38272 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 38272 7642
rect 1104 7568 38272 7590
rect 6365 7531 6423 7537
rect 6365 7497 6377 7531
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 6825 7531 6883 7537
rect 6825 7497 6837 7531
rect 6871 7528 6883 7531
rect 7190 7528 7196 7540
rect 6871 7500 7196 7528
rect 6871 7497 6883 7500
rect 6825 7491 6883 7497
rect 6089 7395 6147 7401
rect 6089 7361 6101 7395
rect 6135 7392 6147 7395
rect 6380 7392 6408 7491
rect 7190 7488 7196 7500
rect 7248 7488 7254 7540
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 7653 7531 7711 7537
rect 7653 7528 7665 7531
rect 7340 7500 7665 7528
rect 7340 7488 7346 7500
rect 7653 7497 7665 7500
rect 7699 7497 7711 7531
rect 7653 7491 7711 7497
rect 8389 7531 8447 7537
rect 8389 7497 8401 7531
rect 8435 7528 8447 7531
rect 8662 7528 8668 7540
rect 8435 7500 8668 7528
rect 8435 7497 8447 7500
rect 8389 7491 8447 7497
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 9306 7488 9312 7540
rect 9364 7488 9370 7540
rect 9490 7488 9496 7540
rect 9548 7488 9554 7540
rect 10318 7488 10324 7540
rect 10376 7528 10382 7540
rect 11698 7528 11704 7540
rect 10376 7500 11704 7528
rect 10376 7488 10382 7500
rect 6546 7420 6552 7472
rect 6604 7460 6610 7472
rect 6733 7463 6791 7469
rect 6733 7460 6745 7463
rect 6604 7432 6745 7460
rect 6604 7420 6610 7432
rect 6733 7429 6745 7432
rect 6779 7460 6791 7463
rect 9324 7460 9352 7488
rect 6779 7432 8524 7460
rect 6779 7429 6791 7432
rect 6733 7423 6791 7429
rect 8496 7401 8524 7432
rect 9140 7432 9352 7460
rect 9401 7463 9459 7469
rect 9140 7401 9168 7432
rect 9401 7429 9413 7463
rect 9447 7460 9459 7463
rect 9508 7460 9536 7488
rect 10962 7460 10968 7472
rect 9447 7432 9536 7460
rect 10626 7432 10968 7460
rect 9447 7429 9459 7432
rect 9401 7423 9459 7429
rect 10962 7420 10968 7432
rect 11020 7420 11026 7472
rect 6135 7364 6408 7392
rect 7837 7395 7895 7401
rect 6135 7361 6147 7364
rect 6089 7355 6147 7361
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 8481 7395 8539 7401
rect 7883 7364 8064 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 6917 7327 6975 7333
rect 6917 7293 6929 7327
rect 6963 7293 6975 7327
rect 6917 7287 6975 7293
rect 6638 7216 6644 7268
rect 6696 7256 6702 7268
rect 6932 7256 6960 7287
rect 8036 7265 8064 7364
rect 8481 7361 8493 7395
rect 8527 7392 8539 7395
rect 9125 7395 9183 7401
rect 8527 7364 8708 7392
rect 8527 7361 8539 7364
rect 8481 7355 8539 7361
rect 8294 7284 8300 7336
rect 8352 7324 8358 7336
rect 8573 7327 8631 7333
rect 8573 7324 8585 7327
rect 8352 7296 8585 7324
rect 8352 7284 8358 7296
rect 8573 7293 8585 7296
rect 8619 7293 8631 7327
rect 8680 7324 8708 7364
rect 9125 7361 9137 7395
rect 9171 7361 9183 7395
rect 11532 7392 11560 7500
rect 11698 7488 11704 7500
rect 11756 7488 11762 7540
rect 12158 7488 12164 7540
rect 12216 7528 12222 7540
rect 12345 7531 12403 7537
rect 12345 7528 12357 7531
rect 12216 7500 12357 7528
rect 12216 7488 12222 7500
rect 12345 7497 12357 7500
rect 12391 7497 12403 7531
rect 12345 7491 12403 7497
rect 12526 7488 12532 7540
rect 12584 7528 12590 7540
rect 16025 7531 16083 7537
rect 12584 7500 13032 7528
rect 12584 7488 12590 7500
rect 11790 7420 11796 7472
rect 11848 7420 11854 7472
rect 12618 7420 12624 7472
rect 12676 7420 12682 7472
rect 13004 7469 13032 7500
rect 16025 7497 16037 7531
rect 16071 7528 16083 7531
rect 16482 7528 16488 7540
rect 16071 7500 16488 7528
rect 16071 7497 16083 7500
rect 16025 7491 16083 7497
rect 16482 7488 16488 7500
rect 16540 7488 16546 7540
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 17310 7528 17316 7540
rect 16632 7500 17316 7528
rect 16632 7488 16638 7500
rect 17310 7488 17316 7500
rect 17368 7488 17374 7540
rect 18325 7531 18383 7537
rect 18064 7500 18276 7528
rect 12989 7463 13047 7469
rect 12989 7429 13001 7463
rect 13035 7429 13047 7463
rect 12989 7423 13047 7429
rect 14737 7463 14795 7469
rect 14737 7429 14749 7463
rect 14783 7460 14795 7463
rect 16758 7460 16764 7472
rect 14783 7432 16764 7460
rect 14783 7429 14795 7432
rect 14737 7423 14795 7429
rect 16758 7420 16764 7432
rect 16816 7420 16822 7472
rect 11609 7395 11667 7401
rect 11609 7392 11621 7395
rect 11532 7364 11621 7392
rect 9125 7355 9183 7361
rect 11609 7361 11621 7364
rect 11655 7361 11667 7395
rect 11609 7355 11667 7361
rect 11885 7395 11943 7401
rect 11885 7361 11897 7395
rect 11931 7361 11943 7395
rect 11885 7355 11943 7361
rect 11977 7395 12035 7401
rect 11977 7361 11989 7395
rect 12023 7361 12035 7395
rect 11977 7355 12035 7361
rect 12437 7395 12495 7401
rect 12437 7361 12449 7395
rect 12483 7392 12495 7395
rect 12636 7392 12664 7420
rect 12483 7364 12664 7392
rect 12483 7361 12495 7364
rect 12437 7355 12495 7361
rect 10134 7324 10140 7336
rect 8680 7296 10140 7324
rect 8573 7287 8631 7293
rect 10134 7284 10140 7296
rect 10192 7284 10198 7336
rect 10870 7284 10876 7336
rect 10928 7324 10934 7336
rect 11900 7324 11928 7355
rect 10928 7296 11928 7324
rect 11992 7324 12020 7355
rect 15378 7352 15384 7404
rect 15436 7352 15442 7404
rect 15470 7352 15476 7404
rect 15528 7392 15534 7404
rect 15528 7364 15573 7392
rect 15528 7352 15534 7364
rect 15654 7352 15660 7404
rect 15712 7352 15718 7404
rect 15749 7395 15807 7401
rect 15749 7361 15761 7395
rect 15795 7361 15807 7395
rect 15749 7355 15807 7361
rect 15887 7395 15945 7401
rect 15887 7361 15899 7395
rect 15933 7392 15945 7395
rect 16022 7392 16028 7404
rect 15933 7364 16028 7392
rect 15933 7361 15945 7364
rect 15887 7355 15945 7361
rect 12802 7324 12808 7336
rect 11992 7296 12808 7324
rect 10928 7284 10934 7296
rect 6696 7228 6960 7256
rect 8021 7259 8079 7265
rect 6696 7216 6702 7228
rect 8021 7225 8033 7259
rect 8067 7225 8079 7259
rect 8021 7219 8079 7225
rect 5902 7148 5908 7200
rect 5960 7148 5966 7200
rect 11900 7188 11928 7296
rect 12802 7284 12808 7296
rect 12860 7324 12866 7336
rect 14826 7324 14832 7336
rect 12860 7296 14832 7324
rect 12860 7284 12866 7296
rect 14826 7284 14832 7296
rect 14884 7284 14890 7336
rect 15194 7284 15200 7336
rect 15252 7324 15258 7336
rect 15764 7324 15792 7355
rect 16022 7352 16028 7364
rect 16080 7352 16086 7404
rect 16301 7395 16359 7401
rect 16301 7361 16313 7395
rect 16347 7361 16359 7395
rect 16301 7355 16359 7361
rect 15252 7296 16252 7324
rect 15252 7284 15258 7296
rect 11974 7216 11980 7268
rect 12032 7256 12038 7268
rect 12161 7259 12219 7265
rect 12161 7256 12173 7259
rect 12032 7228 12173 7256
rect 12032 7216 12038 7228
rect 12161 7225 12173 7228
rect 12207 7225 12219 7259
rect 12161 7219 12219 7225
rect 12342 7216 12348 7268
rect 12400 7256 12406 7268
rect 14734 7256 14740 7268
rect 12400 7228 14740 7256
rect 12400 7216 12406 7228
rect 14734 7216 14740 7228
rect 14792 7216 14798 7268
rect 15286 7216 15292 7268
rect 15344 7216 15350 7268
rect 16117 7259 16175 7265
rect 16117 7225 16129 7259
rect 16163 7225 16175 7259
rect 16117 7219 16175 7225
rect 14090 7188 14096 7200
rect 11900 7160 14096 7188
rect 14090 7148 14096 7160
rect 14148 7148 14154 7200
rect 15304 7188 15332 7216
rect 16132 7188 16160 7219
rect 15304 7160 16160 7188
rect 16224 7188 16252 7296
rect 16316 7256 16344 7355
rect 16390 7352 16396 7404
rect 16448 7392 16454 7404
rect 16485 7395 16543 7401
rect 16485 7392 16497 7395
rect 16448 7364 16497 7392
rect 16448 7352 16454 7364
rect 16485 7361 16497 7364
rect 16531 7361 16543 7395
rect 16485 7355 16543 7361
rect 17034 7352 17040 7404
rect 17092 7352 17098 7404
rect 17126 7352 17132 7404
rect 17184 7352 17190 7404
rect 17218 7352 17224 7404
rect 17276 7352 17282 7404
rect 17328 7401 17356 7488
rect 18064 7469 18092 7500
rect 18049 7463 18107 7469
rect 18049 7429 18061 7463
rect 18095 7429 18107 7463
rect 18248 7460 18276 7500
rect 18325 7497 18337 7531
rect 18371 7528 18383 7531
rect 18506 7528 18512 7540
rect 18371 7500 18512 7528
rect 18371 7497 18383 7500
rect 18325 7491 18383 7497
rect 18506 7488 18512 7500
rect 18564 7488 18570 7540
rect 19794 7528 19800 7540
rect 18616 7500 19800 7528
rect 18616 7460 18644 7500
rect 19794 7488 19800 7500
rect 19852 7488 19858 7540
rect 19978 7488 19984 7540
rect 20036 7528 20042 7540
rect 20165 7531 20223 7537
rect 20165 7528 20177 7531
rect 20036 7500 20177 7528
rect 20036 7488 20042 7500
rect 20165 7497 20177 7500
rect 20211 7528 20223 7531
rect 20530 7528 20536 7540
rect 20211 7500 20536 7528
rect 20211 7497 20223 7500
rect 20165 7491 20223 7497
rect 20530 7488 20536 7500
rect 20588 7528 20594 7540
rect 21174 7528 21180 7540
rect 20588 7500 21180 7528
rect 20588 7488 20594 7500
rect 21174 7488 21180 7500
rect 21232 7488 21238 7540
rect 22370 7488 22376 7540
rect 22428 7488 22434 7540
rect 22554 7488 22560 7540
rect 22612 7528 22618 7540
rect 23014 7528 23020 7540
rect 22612 7500 23020 7528
rect 22612 7488 22618 7500
rect 23014 7488 23020 7500
rect 23072 7488 23078 7540
rect 23198 7488 23204 7540
rect 23256 7528 23262 7540
rect 23293 7531 23351 7537
rect 23293 7528 23305 7531
rect 23256 7500 23305 7528
rect 23256 7488 23262 7500
rect 23293 7497 23305 7500
rect 23339 7497 23351 7531
rect 23293 7491 23351 7497
rect 24946 7488 24952 7540
rect 25004 7528 25010 7540
rect 25317 7531 25375 7537
rect 25317 7528 25329 7531
rect 25004 7500 25329 7528
rect 25004 7488 25010 7500
rect 25317 7497 25329 7500
rect 25363 7497 25375 7531
rect 25317 7491 25375 7497
rect 25406 7488 25412 7540
rect 25464 7488 25470 7540
rect 26237 7531 26295 7537
rect 26237 7497 26249 7531
rect 26283 7528 26295 7531
rect 26326 7528 26332 7540
rect 26283 7500 26332 7528
rect 26283 7497 26295 7500
rect 26237 7491 26295 7497
rect 26326 7488 26332 7500
rect 26384 7528 26390 7540
rect 28718 7528 28724 7540
rect 26384 7500 28724 7528
rect 26384 7488 26390 7500
rect 28718 7488 28724 7500
rect 28776 7488 28782 7540
rect 29365 7531 29423 7537
rect 29365 7497 29377 7531
rect 29411 7528 29423 7531
rect 30006 7528 30012 7540
rect 29411 7500 30012 7528
rect 29411 7497 29423 7500
rect 29365 7491 29423 7497
rect 30006 7488 30012 7500
rect 30064 7488 30070 7540
rect 30377 7531 30435 7537
rect 30377 7497 30389 7531
rect 30423 7528 30435 7531
rect 30466 7528 30472 7540
rect 30423 7500 30472 7528
rect 30423 7497 30435 7500
rect 30377 7491 30435 7497
rect 30466 7488 30472 7500
rect 30524 7488 30530 7540
rect 31386 7488 31392 7540
rect 31444 7528 31450 7540
rect 31570 7528 31576 7540
rect 31444 7500 31576 7528
rect 31444 7488 31450 7500
rect 31570 7488 31576 7500
rect 31628 7488 31634 7540
rect 32306 7488 32312 7540
rect 32364 7488 32370 7540
rect 18248 7432 18368 7460
rect 18049 7423 18107 7429
rect 17313 7395 17371 7401
rect 17313 7361 17325 7395
rect 17359 7361 17371 7395
rect 17313 7355 17371 7361
rect 17405 7395 17463 7401
rect 17405 7361 17417 7395
rect 17451 7392 17463 7395
rect 17494 7392 17500 7404
rect 17451 7364 17500 7392
rect 17451 7361 17463 7364
rect 17405 7355 17463 7361
rect 17494 7352 17500 7364
rect 17552 7352 17558 7404
rect 17678 7352 17684 7404
rect 17736 7352 17742 7404
rect 17770 7352 17776 7404
rect 17828 7352 17834 7404
rect 17862 7352 17868 7404
rect 17920 7392 17926 7404
rect 17957 7395 18015 7401
rect 17957 7392 17969 7395
rect 17920 7364 17969 7392
rect 17920 7352 17926 7364
rect 17957 7361 17969 7364
rect 18003 7361 18015 7395
rect 17957 7355 18015 7361
rect 18146 7395 18204 7401
rect 18146 7361 18158 7395
rect 18192 7361 18204 7395
rect 18146 7355 18204 7361
rect 17144 7324 17172 7352
rect 18156 7324 18184 7355
rect 17144 7296 18184 7324
rect 18340 7324 18368 7432
rect 18524 7432 18644 7460
rect 18414 7352 18420 7404
rect 18472 7401 18478 7404
rect 18472 7395 18495 7401
rect 18483 7361 18495 7395
rect 18524 7392 18552 7432
rect 19150 7420 19156 7472
rect 19208 7460 19214 7472
rect 20714 7460 20720 7472
rect 19208 7432 20720 7460
rect 19208 7420 19214 7432
rect 20714 7420 20720 7432
rect 20772 7420 20778 7472
rect 23385 7463 23443 7469
rect 23385 7460 23397 7463
rect 20916 7432 23397 7460
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 18524 7364 18613 7392
rect 18472 7355 18495 7361
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 18601 7355 18659 7361
rect 18693 7395 18751 7401
rect 18693 7361 18705 7395
rect 18739 7361 18751 7395
rect 18693 7355 18751 7361
rect 18785 7395 18843 7401
rect 18785 7361 18797 7395
rect 18831 7390 18843 7395
rect 18831 7361 18852 7390
rect 18785 7355 18852 7361
rect 18472 7352 18478 7355
rect 18708 7324 18736 7355
rect 18340 7296 18736 7324
rect 16574 7256 16580 7268
rect 16316 7228 16580 7256
rect 16574 7216 16580 7228
rect 16632 7216 16638 7268
rect 18340 7256 18368 7296
rect 16684 7228 18368 7256
rect 18824 7256 18852 7355
rect 18966 7352 18972 7404
rect 19024 7392 19030 7404
rect 19886 7392 19892 7404
rect 19024 7364 19892 7392
rect 19024 7352 19030 7364
rect 19886 7352 19892 7364
rect 19944 7392 19950 7404
rect 20530 7392 20536 7404
rect 19944 7364 20536 7392
rect 19944 7352 19950 7364
rect 20530 7352 20536 7364
rect 20588 7352 20594 7404
rect 20625 7395 20683 7401
rect 20625 7361 20637 7395
rect 20671 7361 20683 7395
rect 20732 7392 20760 7420
rect 20916 7392 20944 7432
rect 23385 7429 23397 7432
rect 23431 7429 23443 7463
rect 25424 7460 25452 7488
rect 25424 7432 26372 7460
rect 23385 7423 23443 7429
rect 20732 7364 20944 7392
rect 20625 7355 20683 7361
rect 19426 7324 19432 7336
rect 19306 7296 19432 7324
rect 19306 7256 19334 7296
rect 19426 7284 19432 7296
rect 19484 7284 19490 7336
rect 20640 7324 20668 7355
rect 21266 7352 21272 7404
rect 21324 7352 21330 7404
rect 21450 7352 21456 7404
rect 21508 7352 21514 7404
rect 21818 7352 21824 7404
rect 21876 7352 21882 7404
rect 21910 7352 21916 7404
rect 21968 7392 21974 7404
rect 22005 7395 22063 7401
rect 22005 7392 22017 7395
rect 21968 7364 22017 7392
rect 21968 7352 21974 7364
rect 22005 7361 22017 7364
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 22097 7395 22155 7401
rect 22097 7361 22109 7395
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 21468 7324 21496 7352
rect 20640 7296 21496 7324
rect 22112 7324 22140 7355
rect 22186 7352 22192 7404
rect 22244 7352 22250 7404
rect 22462 7352 22468 7404
rect 22520 7392 22526 7404
rect 22741 7395 22799 7401
rect 22741 7392 22753 7395
rect 22520 7364 22753 7392
rect 22520 7352 22526 7364
rect 22741 7361 22753 7364
rect 22787 7361 22799 7395
rect 22741 7355 22799 7361
rect 22925 7395 22983 7401
rect 22925 7361 22937 7395
rect 22971 7361 22983 7395
rect 22925 7355 22983 7361
rect 22278 7324 22284 7336
rect 22112 7296 22284 7324
rect 22278 7284 22284 7296
rect 22336 7284 22342 7336
rect 22940 7324 22968 7355
rect 23014 7352 23020 7404
rect 23072 7352 23078 7404
rect 23106 7352 23112 7404
rect 23164 7352 23170 7404
rect 24210 7352 24216 7404
rect 24268 7392 24274 7404
rect 24670 7392 24676 7404
rect 24268 7364 24676 7392
rect 24268 7352 24274 7364
rect 24670 7352 24676 7364
rect 24728 7352 24734 7404
rect 25498 7401 25504 7404
rect 25496 7392 25504 7401
rect 25459 7364 25504 7392
rect 25496 7355 25504 7364
rect 25498 7352 25504 7355
rect 25556 7352 25562 7404
rect 25590 7352 25596 7404
rect 25648 7352 25654 7404
rect 25685 7395 25743 7401
rect 25685 7361 25697 7395
rect 25731 7361 25743 7395
rect 25866 7392 25872 7404
rect 25827 7364 25872 7392
rect 25685 7355 25743 7361
rect 25700 7324 25728 7355
rect 25866 7352 25872 7364
rect 25924 7352 25930 7404
rect 25961 7395 26019 7401
rect 25961 7361 25973 7395
rect 26007 7361 26019 7395
rect 25961 7355 26019 7361
rect 22940 7296 25728 7324
rect 25976 7324 26004 7355
rect 26050 7352 26056 7404
rect 26108 7352 26114 7404
rect 26344 7401 26372 7432
rect 28994 7420 29000 7472
rect 29052 7420 29058 7472
rect 29914 7460 29920 7472
rect 29196 7432 29920 7460
rect 26329 7395 26387 7401
rect 26329 7361 26341 7395
rect 26375 7361 26387 7395
rect 26329 7355 26387 7361
rect 26510 7352 26516 7404
rect 26568 7352 26574 7404
rect 26602 7352 26608 7404
rect 26660 7392 26666 7404
rect 29196 7401 29224 7432
rect 29914 7420 29920 7432
rect 29972 7460 29978 7472
rect 32030 7460 32036 7472
rect 29972 7432 30052 7460
rect 29972 7420 29978 7432
rect 28813 7395 28871 7401
rect 28813 7392 28825 7395
rect 26660 7364 28825 7392
rect 26660 7352 26666 7364
rect 28813 7361 28825 7364
rect 28859 7361 28871 7395
rect 28813 7355 28871 7361
rect 29089 7395 29147 7401
rect 29089 7361 29101 7395
rect 29135 7361 29147 7395
rect 29089 7355 29147 7361
rect 29181 7395 29239 7401
rect 29181 7361 29193 7395
rect 29227 7361 29239 7395
rect 29181 7355 29239 7361
rect 26528 7324 26556 7352
rect 25976 7296 26556 7324
rect 18824 7228 19334 7256
rect 16684 7188 16712 7228
rect 19610 7216 19616 7268
rect 19668 7256 19674 7268
rect 20070 7256 20076 7268
rect 19668 7228 20076 7256
rect 19668 7216 19674 7228
rect 20070 7216 20076 7228
rect 20128 7256 20134 7268
rect 22940 7256 22968 7296
rect 20128 7228 22968 7256
rect 20128 7216 20134 7228
rect 16224 7160 16712 7188
rect 17589 7191 17647 7197
rect 17589 7157 17601 7191
rect 17635 7188 17647 7191
rect 18414 7188 18420 7200
rect 17635 7160 18420 7188
rect 17635 7157 17647 7160
rect 17589 7151 17647 7157
rect 18414 7148 18420 7160
rect 18472 7148 18478 7200
rect 18966 7148 18972 7200
rect 19024 7148 19030 7200
rect 19058 7148 19064 7200
rect 19116 7188 19122 7200
rect 20254 7188 20260 7200
rect 19116 7160 20260 7188
rect 19116 7148 19122 7160
rect 20254 7148 20260 7160
rect 20312 7148 20318 7200
rect 20346 7148 20352 7200
rect 20404 7188 20410 7200
rect 21082 7188 21088 7200
rect 20404 7160 21088 7188
rect 20404 7148 20410 7160
rect 21082 7148 21088 7160
rect 21140 7148 21146 7200
rect 22186 7148 22192 7200
rect 22244 7188 22250 7200
rect 24302 7188 24308 7200
rect 22244 7160 24308 7188
rect 22244 7148 22250 7160
rect 24302 7148 24308 7160
rect 24360 7148 24366 7200
rect 24670 7148 24676 7200
rect 24728 7148 24734 7200
rect 25700 7188 25728 7296
rect 29104 7268 29132 7355
rect 29546 7352 29552 7404
rect 29604 7392 29610 7404
rect 29733 7395 29791 7401
rect 29733 7392 29745 7395
rect 29604 7364 29745 7392
rect 29604 7352 29610 7364
rect 29733 7361 29745 7364
rect 29779 7361 29791 7395
rect 29733 7355 29791 7361
rect 29822 7352 29828 7404
rect 29880 7392 29886 7404
rect 30024 7401 30052 7432
rect 30116 7432 32036 7460
rect 30116 7404 30144 7432
rect 32030 7420 32036 7432
rect 32088 7420 32094 7472
rect 32324 7460 32352 7488
rect 33686 7460 33692 7472
rect 32140 7432 32352 7460
rect 33626 7432 33692 7460
rect 30009 7395 30067 7401
rect 29880 7364 29925 7392
rect 29880 7352 29886 7364
rect 30009 7361 30021 7395
rect 30055 7361 30067 7395
rect 30009 7355 30067 7361
rect 30098 7352 30104 7404
rect 30156 7352 30162 7404
rect 30198 7395 30256 7401
rect 30198 7361 30210 7395
rect 30244 7361 30256 7395
rect 31662 7392 31668 7404
rect 30198 7355 30256 7361
rect 31404 7364 31668 7392
rect 29638 7284 29644 7336
rect 29696 7324 29702 7336
rect 30208 7324 30236 7355
rect 31404 7333 31432 7364
rect 31662 7352 31668 7364
rect 31720 7352 31726 7404
rect 32140 7401 32168 7432
rect 33686 7420 33692 7432
rect 33744 7420 33750 7472
rect 32125 7395 32183 7401
rect 32125 7361 32137 7395
rect 32171 7361 32183 7395
rect 32125 7355 32183 7361
rect 29696 7296 30236 7324
rect 31389 7327 31447 7333
rect 29696 7284 29702 7296
rect 31389 7293 31401 7327
rect 31435 7293 31447 7327
rect 31389 7287 31447 7293
rect 31481 7327 31539 7333
rect 31481 7293 31493 7327
rect 31527 7324 31539 7327
rect 31527 7296 32260 7324
rect 31527 7293 31539 7296
rect 31481 7287 31539 7293
rect 25958 7216 25964 7268
rect 26016 7256 26022 7268
rect 26053 7259 26111 7265
rect 26053 7256 26065 7259
rect 26016 7228 26065 7256
rect 26016 7216 26022 7228
rect 26053 7225 26065 7228
rect 26099 7225 26111 7259
rect 26053 7219 26111 7225
rect 26142 7216 26148 7268
rect 26200 7256 26206 7268
rect 28626 7256 28632 7268
rect 26200 7228 28632 7256
rect 26200 7216 26206 7228
rect 28626 7216 28632 7228
rect 28684 7256 28690 7268
rect 29086 7256 29092 7268
rect 28684 7228 29092 7256
rect 28684 7216 28690 7228
rect 29086 7216 29092 7228
rect 29144 7216 29150 7268
rect 29822 7216 29828 7268
rect 29880 7256 29886 7268
rect 31496 7256 31524 7287
rect 29880 7228 31524 7256
rect 29880 7216 29886 7228
rect 26234 7188 26240 7200
rect 25700 7160 26240 7188
rect 26234 7148 26240 7160
rect 26292 7148 26298 7200
rect 27890 7148 27896 7200
rect 27948 7188 27954 7200
rect 30098 7188 30104 7200
rect 27948 7160 30104 7188
rect 27948 7148 27954 7160
rect 30098 7148 30104 7160
rect 30156 7148 30162 7200
rect 31938 7148 31944 7200
rect 31996 7148 32002 7200
rect 32232 7188 32260 7296
rect 32398 7284 32404 7336
rect 32456 7284 32462 7336
rect 33873 7191 33931 7197
rect 33873 7188 33885 7191
rect 32232 7160 33885 7188
rect 33873 7157 33885 7160
rect 33919 7157 33931 7191
rect 33873 7151 33931 7157
rect 1104 7098 38272 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38272 7098
rect 1104 7024 38272 7046
rect 5708 6987 5766 6993
rect 5708 6953 5720 6987
rect 5754 6984 5766 6987
rect 5902 6984 5908 6996
rect 5754 6956 5908 6984
rect 5754 6953 5766 6956
rect 5708 6947 5766 6953
rect 5902 6944 5908 6956
rect 5960 6944 5966 6996
rect 7190 6944 7196 6996
rect 7248 6944 7254 6996
rect 14734 6944 14740 6996
rect 14792 6984 14798 6996
rect 18141 6987 18199 6993
rect 14792 6956 18092 6984
rect 14792 6944 14798 6956
rect 16574 6916 16580 6928
rect 14936 6888 16580 6916
rect 14090 6808 14096 6860
rect 14148 6848 14154 6860
rect 14936 6848 14964 6888
rect 16574 6876 16580 6888
rect 16632 6916 16638 6928
rect 17770 6916 17776 6928
rect 16632 6888 17776 6916
rect 16632 6876 16638 6888
rect 17770 6876 17776 6888
rect 17828 6876 17834 6928
rect 18064 6916 18092 6956
rect 18141 6953 18153 6987
rect 18187 6984 18199 6987
rect 18230 6984 18236 6996
rect 18187 6956 18236 6984
rect 18187 6953 18199 6956
rect 18141 6947 18199 6953
rect 18230 6944 18236 6956
rect 18288 6944 18294 6996
rect 18690 6984 18696 6996
rect 18340 6956 18696 6984
rect 18340 6916 18368 6956
rect 18690 6944 18696 6956
rect 18748 6944 18754 6996
rect 20530 6944 20536 6996
rect 20588 6984 20594 6996
rect 20588 6956 21956 6984
rect 20588 6944 20594 6956
rect 18064 6888 18368 6916
rect 18414 6876 18420 6928
rect 18472 6876 18478 6928
rect 18708 6916 18736 6944
rect 21542 6916 21548 6928
rect 18708 6888 21548 6916
rect 21542 6876 21548 6888
rect 21600 6876 21606 6928
rect 21634 6876 21640 6928
rect 21692 6916 21698 6928
rect 21928 6916 21956 6956
rect 22278 6944 22284 6996
rect 22336 6984 22342 6996
rect 22830 6984 22836 6996
rect 22336 6956 22836 6984
rect 22336 6944 22342 6956
rect 22830 6944 22836 6956
rect 22888 6984 22894 6996
rect 25869 6987 25927 6993
rect 22888 6956 23520 6984
rect 22888 6944 22894 6956
rect 21692 6888 21864 6916
rect 21928 6888 23336 6916
rect 21692 6876 21698 6888
rect 15470 6848 15476 6860
rect 14148 6820 14964 6848
rect 15028 6820 15476 6848
rect 14148 6808 14154 6820
rect 5169 6783 5227 6789
rect 5169 6749 5181 6783
rect 5215 6749 5227 6783
rect 5169 6743 5227 6749
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6780 5319 6783
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 5307 6752 5457 6780
rect 5307 6749 5319 6752
rect 5261 6743 5319 6749
rect 5445 6749 5457 6752
rect 5491 6749 5503 6783
rect 7742 6780 7748 6792
rect 6854 6752 7748 6780
rect 5445 6743 5503 6749
rect 5184 6712 5212 6743
rect 7742 6740 7748 6752
rect 7800 6780 7806 6792
rect 7926 6780 7932 6792
rect 7800 6752 7932 6780
rect 7800 6740 7806 6752
rect 7926 6740 7932 6752
rect 7984 6740 7990 6792
rect 8938 6740 8944 6792
rect 8996 6780 9002 6792
rect 11885 6783 11943 6789
rect 11885 6780 11897 6783
rect 8996 6752 11897 6780
rect 8996 6740 9002 6752
rect 11885 6749 11897 6752
rect 11931 6780 11943 6783
rect 11931 6752 12434 6780
rect 11931 6749 11943 6752
rect 11885 6743 11943 6749
rect 5994 6712 6000 6724
rect 5184 6684 6000 6712
rect 5994 6672 6000 6684
rect 6052 6672 6058 6724
rect 12406 6656 12434 6752
rect 14182 6740 14188 6792
rect 14240 6740 14246 6792
rect 14366 6740 14372 6792
rect 14424 6740 14430 6792
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 14645 6783 14703 6789
rect 14645 6780 14657 6783
rect 14599 6752 14657 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 14645 6749 14657 6752
rect 14691 6749 14703 6783
rect 14645 6743 14703 6749
rect 14738 6783 14796 6789
rect 14738 6749 14750 6783
rect 14784 6780 14796 6783
rect 15028 6780 15056 6820
rect 15470 6808 15476 6820
rect 15528 6848 15534 6860
rect 15528 6820 17172 6848
rect 15528 6808 15534 6820
rect 14784 6752 15056 6780
rect 14784 6749 14796 6752
rect 14738 6743 14796 6749
rect 14752 6712 14780 6743
rect 15102 6740 15108 6792
rect 15160 6789 15166 6792
rect 15160 6780 15168 6789
rect 15160 6752 15205 6780
rect 15160 6743 15168 6752
rect 15160 6740 15166 6743
rect 15654 6740 15660 6792
rect 15712 6780 15718 6792
rect 17144 6789 17172 6820
rect 18230 6808 18236 6860
rect 18288 6848 18294 6860
rect 18509 6851 18567 6857
rect 18288 6820 18460 6848
rect 18288 6808 18294 6820
rect 16853 6783 16911 6789
rect 16853 6780 16865 6783
rect 15712 6752 16865 6780
rect 15712 6740 15718 6752
rect 16853 6749 16865 6752
rect 16899 6749 16911 6783
rect 16853 6743 16911 6749
rect 17129 6783 17187 6789
rect 17129 6749 17141 6783
rect 17175 6749 17187 6783
rect 17129 6743 17187 6749
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6780 17279 6783
rect 17586 6780 17592 6792
rect 17267 6752 17592 6780
rect 17267 6749 17279 6752
rect 17221 6743 17279 6749
rect 17586 6740 17592 6752
rect 17644 6740 17650 6792
rect 18046 6740 18052 6792
rect 18104 6740 18110 6792
rect 18322 6740 18328 6792
rect 18380 6740 18386 6792
rect 18432 6780 18460 6820
rect 18509 6817 18521 6851
rect 18555 6848 18567 6851
rect 18966 6848 18972 6860
rect 18555 6820 18972 6848
rect 18555 6817 18567 6820
rect 18509 6811 18567 6817
rect 18966 6808 18972 6820
rect 19024 6808 19030 6860
rect 20254 6808 20260 6860
rect 20312 6808 20318 6860
rect 21082 6808 21088 6860
rect 21140 6848 21146 6860
rect 21140 6820 21772 6848
rect 21140 6808 21146 6820
rect 18601 6783 18659 6789
rect 18601 6780 18613 6783
rect 18432 6752 18613 6780
rect 18601 6749 18613 6752
rect 18647 6749 18659 6783
rect 18601 6743 18659 6749
rect 18690 6740 18696 6792
rect 18748 6780 18754 6792
rect 18785 6783 18843 6789
rect 18785 6780 18797 6783
rect 18748 6752 18797 6780
rect 18748 6740 18754 6752
rect 18785 6749 18797 6752
rect 18831 6749 18843 6783
rect 18785 6743 18843 6749
rect 20070 6740 20076 6792
rect 20128 6740 20134 6792
rect 21545 6783 21603 6789
rect 21545 6780 21557 6783
rect 20180 6752 21557 6780
rect 14568 6684 14780 6712
rect 14568 6656 14596 6684
rect 14826 6672 14832 6724
rect 14884 6712 14890 6724
rect 14921 6715 14979 6721
rect 14921 6712 14933 6715
rect 14884 6684 14933 6712
rect 14884 6672 14890 6684
rect 14921 6681 14933 6684
rect 14967 6681 14979 6715
rect 14921 6675 14979 6681
rect 15013 6715 15071 6721
rect 15013 6681 15025 6715
rect 15059 6712 15071 6715
rect 15672 6712 15700 6740
rect 17037 6715 17095 6721
rect 17037 6712 17049 6715
rect 15059 6684 15700 6712
rect 16868 6684 17049 6712
rect 15059 6681 15071 6684
rect 15013 6675 15071 6681
rect 16868 6656 16896 6684
rect 17037 6681 17049 6684
rect 17083 6681 17095 6715
rect 17037 6675 17095 6681
rect 17954 6672 17960 6724
rect 18012 6672 18018 6724
rect 18064 6712 18092 6740
rect 20180 6712 20208 6752
rect 21545 6749 21557 6752
rect 21591 6749 21603 6783
rect 21545 6743 21603 6749
rect 21638 6783 21696 6789
rect 21638 6749 21650 6783
rect 21684 6749 21696 6783
rect 21638 6743 21696 6749
rect 18064 6684 20208 6712
rect 20622 6672 20628 6724
rect 20680 6712 20686 6724
rect 20898 6712 20904 6724
rect 20680 6684 20904 6712
rect 20680 6672 20686 6684
rect 20898 6672 20904 6684
rect 20956 6712 20962 6724
rect 21653 6712 21681 6743
rect 20956 6684 21681 6712
rect 21744 6712 21772 6820
rect 21836 6789 21864 6888
rect 23308 6860 23336 6888
rect 21928 6820 23060 6848
rect 21928 6789 21956 6820
rect 23032 6792 23060 6820
rect 23290 6808 23296 6860
rect 23348 6808 23354 6860
rect 21821 6783 21879 6789
rect 21821 6749 21833 6783
rect 21867 6749 21879 6783
rect 21821 6743 21879 6749
rect 21913 6783 21971 6789
rect 21913 6749 21925 6783
rect 21959 6749 21971 6783
rect 21913 6743 21971 6749
rect 22002 6740 22008 6792
rect 22060 6789 22066 6792
rect 22060 6783 22109 6789
rect 22060 6749 22063 6783
rect 22097 6749 22109 6783
rect 22060 6743 22109 6749
rect 22060 6740 22066 6743
rect 22186 6740 22192 6792
rect 22244 6780 22250 6792
rect 22281 6783 22339 6789
rect 22281 6780 22293 6783
rect 22244 6752 22293 6780
rect 22244 6740 22250 6752
rect 22281 6749 22293 6752
rect 22327 6749 22339 6783
rect 22281 6743 22339 6749
rect 22374 6783 22432 6789
rect 22374 6749 22386 6783
rect 22420 6749 22432 6783
rect 22374 6743 22432 6749
rect 22787 6783 22845 6789
rect 22787 6749 22799 6783
rect 22833 6780 22845 6783
rect 22922 6780 22928 6792
rect 22833 6752 22928 6780
rect 22833 6749 22845 6752
rect 22787 6743 22845 6749
rect 22389 6712 22417 6743
rect 22922 6740 22928 6752
rect 22980 6740 22986 6792
rect 23014 6740 23020 6792
rect 23072 6740 23078 6792
rect 23196 6783 23254 6789
rect 23196 6749 23208 6783
rect 23242 6780 23254 6783
rect 23308 6780 23336 6808
rect 23242 6752 23336 6780
rect 23492 6780 23520 6956
rect 25869 6953 25881 6987
rect 25915 6984 25927 6987
rect 26050 6984 26056 6996
rect 25915 6956 26056 6984
rect 25915 6953 25927 6956
rect 25869 6947 25927 6953
rect 26050 6944 26056 6956
rect 26108 6944 26114 6996
rect 28534 6984 28540 6996
rect 27724 6956 28540 6984
rect 25682 6916 25688 6928
rect 24872 6888 25688 6916
rect 23566 6780 23572 6792
rect 23492 6752 23572 6780
rect 23242 6749 23254 6752
rect 23196 6743 23254 6749
rect 23566 6740 23572 6752
rect 23624 6740 23630 6792
rect 23658 6740 23664 6792
rect 23716 6740 23722 6792
rect 24872 6780 24900 6888
rect 25682 6876 25688 6888
rect 25740 6876 25746 6928
rect 26142 6876 26148 6928
rect 26200 6876 26206 6928
rect 25222 6808 25228 6860
rect 25280 6848 25286 6860
rect 26160 6848 26188 6876
rect 25280 6820 25360 6848
rect 25280 6808 25286 6820
rect 25332 6789 25360 6820
rect 25700 6820 26188 6848
rect 25700 6789 25728 6820
rect 24689 6752 24900 6780
rect 24949 6783 25007 6789
rect 21744 6684 22417 6712
rect 20956 6672 20962 6684
rect 22554 6672 22560 6724
rect 22612 6672 22618 6724
rect 22649 6715 22707 6721
rect 22649 6681 22661 6715
rect 22695 6712 22707 6715
rect 23290 6712 23296 6724
rect 22695 6684 23296 6712
rect 22695 6681 22707 6684
rect 22649 6675 22707 6681
rect 23290 6672 23296 6684
rect 23348 6672 23354 6724
rect 23385 6715 23443 6721
rect 23385 6681 23397 6715
rect 23431 6712 23443 6715
rect 24689 6712 24717 6752
rect 24949 6749 24961 6783
rect 24995 6749 25007 6783
rect 24949 6743 25007 6749
rect 25041 6783 25099 6789
rect 25041 6749 25053 6783
rect 25087 6780 25099 6783
rect 25317 6783 25375 6789
rect 25087 6752 25268 6780
rect 25087 6749 25099 6752
rect 25041 6743 25099 6749
rect 23431 6684 24717 6712
rect 24765 6715 24823 6721
rect 23431 6681 23443 6684
rect 23385 6675 23443 6681
rect 24765 6681 24777 6715
rect 24811 6712 24823 6715
rect 24854 6712 24860 6724
rect 24811 6684 24860 6712
rect 24811 6681 24823 6684
rect 24765 6675 24823 6681
rect 24854 6672 24860 6684
rect 24912 6672 24918 6724
rect 24964 6712 24992 6743
rect 24964 6684 25176 6712
rect 11790 6604 11796 6656
rect 11848 6604 11854 6656
rect 12342 6604 12348 6656
rect 12400 6644 12434 6656
rect 12526 6644 12532 6656
rect 12400 6616 12532 6644
rect 12400 6604 12406 6616
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 14550 6604 14556 6656
rect 14608 6604 14614 6656
rect 15289 6647 15347 6653
rect 15289 6613 15301 6647
rect 15335 6644 15347 6647
rect 15746 6644 15752 6656
rect 15335 6616 15752 6644
rect 15335 6613 15347 6616
rect 15289 6607 15347 6613
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 16850 6604 16856 6656
rect 16908 6604 16914 6656
rect 17405 6647 17463 6653
rect 17405 6613 17417 6647
rect 17451 6644 17463 6647
rect 17972 6644 18000 6672
rect 17451 6616 18000 6644
rect 17451 6613 17463 6616
rect 17405 6607 17463 6613
rect 19794 6604 19800 6656
rect 19852 6644 19858 6656
rect 21634 6644 21640 6656
rect 19852 6616 21640 6644
rect 19852 6604 19858 6616
rect 21634 6604 21640 6616
rect 21692 6604 21698 6656
rect 22186 6604 22192 6656
rect 22244 6604 22250 6656
rect 22278 6604 22284 6656
rect 22336 6644 22342 6656
rect 22925 6647 22983 6653
rect 22925 6644 22937 6647
rect 22336 6616 22937 6644
rect 22336 6604 22342 6616
rect 22925 6613 22937 6616
rect 22971 6613 22983 6647
rect 22925 6607 22983 6613
rect 23014 6604 23020 6656
rect 23072 6604 23078 6656
rect 23106 6604 23112 6656
rect 23164 6644 23170 6656
rect 23934 6644 23940 6656
rect 23164 6616 23940 6644
rect 23164 6604 23170 6616
rect 23934 6604 23940 6616
rect 23992 6604 23998 6656
rect 25038 6604 25044 6656
rect 25096 6604 25102 6656
rect 25148 6653 25176 6684
rect 25133 6647 25191 6653
rect 25133 6613 25145 6647
rect 25179 6613 25191 6647
rect 25240 6644 25268 6752
rect 25317 6749 25329 6783
rect 25363 6749 25375 6783
rect 25317 6743 25375 6749
rect 25685 6783 25743 6789
rect 25685 6749 25697 6783
rect 25731 6749 25743 6783
rect 25685 6743 25743 6749
rect 25774 6740 25780 6792
rect 25832 6780 25838 6792
rect 26007 6783 26065 6789
rect 26007 6780 26019 6783
rect 25832 6752 26019 6780
rect 25832 6740 25838 6752
rect 26007 6749 26019 6752
rect 26053 6749 26065 6783
rect 26007 6743 26065 6749
rect 26142 6740 26148 6792
rect 26200 6740 26206 6792
rect 26234 6740 26240 6792
rect 26292 6740 26298 6792
rect 26418 6780 26424 6792
rect 26379 6752 26424 6780
rect 26418 6740 26424 6752
rect 26476 6740 26482 6792
rect 26510 6740 26516 6792
rect 26568 6740 26574 6792
rect 27246 6740 27252 6792
rect 27304 6740 27310 6792
rect 27617 6783 27675 6789
rect 27617 6780 27629 6783
rect 27448 6752 27629 6780
rect 25406 6672 25412 6724
rect 25464 6672 25470 6724
rect 25498 6672 25504 6724
rect 25556 6672 25562 6724
rect 25590 6672 25596 6724
rect 25648 6712 25654 6724
rect 26602 6712 26608 6724
rect 25648 6684 26608 6712
rect 25648 6672 25654 6684
rect 26602 6672 26608 6684
rect 26660 6712 26666 6724
rect 26973 6715 27031 6721
rect 26973 6712 26985 6715
rect 26660 6684 26985 6712
rect 26660 6672 26666 6684
rect 26973 6681 26985 6684
rect 27019 6681 27031 6715
rect 26973 6675 27031 6681
rect 25314 6644 25320 6656
rect 25240 6616 25320 6644
rect 25133 6607 25191 6613
rect 25314 6604 25320 6616
rect 25372 6604 25378 6656
rect 25424 6644 25452 6672
rect 26786 6644 26792 6656
rect 25424 6616 26792 6644
rect 26786 6604 26792 6616
rect 26844 6604 26850 6656
rect 27154 6604 27160 6656
rect 27212 6604 27218 6656
rect 27341 6647 27399 6653
rect 27341 6613 27353 6647
rect 27387 6644 27399 6647
rect 27448 6644 27476 6752
rect 27617 6749 27629 6752
rect 27663 6749 27675 6783
rect 27724 6780 27752 6956
rect 28534 6944 28540 6956
rect 28592 6984 28598 6996
rect 29733 6987 29791 6993
rect 29733 6984 29745 6987
rect 28592 6956 29745 6984
rect 28592 6944 28598 6956
rect 29733 6953 29745 6956
rect 29779 6953 29791 6987
rect 29733 6947 29791 6953
rect 31757 6987 31815 6993
rect 31757 6953 31769 6987
rect 31803 6984 31815 6987
rect 32398 6984 32404 6996
rect 31803 6956 32404 6984
rect 31803 6953 31815 6956
rect 31757 6947 31815 6953
rect 32398 6944 32404 6956
rect 32456 6944 32462 6996
rect 28350 6916 28356 6928
rect 28000 6888 28356 6916
rect 28000 6848 28028 6888
rect 28350 6876 28356 6888
rect 28408 6876 28414 6928
rect 28718 6876 28724 6928
rect 28776 6916 28782 6928
rect 29822 6916 29828 6928
rect 28776 6888 29828 6916
rect 28776 6876 28782 6888
rect 29822 6876 29828 6888
rect 29880 6876 29886 6928
rect 27908 6820 28028 6848
rect 28261 6851 28319 6857
rect 27908 6789 27936 6820
rect 28261 6817 28273 6851
rect 28307 6848 28319 6851
rect 28537 6851 28595 6857
rect 28537 6848 28549 6851
rect 28307 6820 28549 6848
rect 28307 6817 28319 6820
rect 28261 6811 28319 6817
rect 28537 6817 28549 6820
rect 28583 6817 28595 6851
rect 28736 6848 28764 6876
rect 28736 6820 28856 6848
rect 28537 6811 28595 6817
rect 27801 6783 27859 6789
rect 27801 6780 27813 6783
rect 27724 6752 27813 6780
rect 27617 6743 27675 6749
rect 27801 6749 27813 6752
rect 27847 6749 27859 6783
rect 27801 6743 27859 6749
rect 27893 6783 27951 6789
rect 27893 6749 27905 6783
rect 27939 6749 27951 6783
rect 27893 6743 27951 6749
rect 27985 6783 28043 6789
rect 27985 6749 27997 6783
rect 28031 6780 28043 6783
rect 28074 6780 28080 6792
rect 28031 6752 28080 6780
rect 28031 6749 28043 6752
rect 27985 6743 28043 6749
rect 28074 6740 28080 6752
rect 28132 6740 28138 6792
rect 28166 6740 28172 6792
rect 28224 6780 28230 6792
rect 28353 6783 28411 6789
rect 28353 6780 28365 6783
rect 28224 6752 28365 6780
rect 28224 6740 28230 6752
rect 28353 6749 28365 6752
rect 28399 6749 28411 6783
rect 28353 6743 28411 6749
rect 28629 6783 28687 6789
rect 28629 6749 28641 6783
rect 28675 6749 28687 6783
rect 28629 6743 28687 6749
rect 27525 6715 27583 6721
rect 27525 6681 27537 6715
rect 27571 6712 27583 6715
rect 28644 6712 28672 6743
rect 28718 6740 28724 6792
rect 28776 6740 28782 6792
rect 28828 6789 28856 6820
rect 28813 6783 28871 6789
rect 28813 6749 28825 6783
rect 28859 6749 28871 6783
rect 28813 6743 28871 6749
rect 28997 6783 29055 6789
rect 28997 6749 29009 6783
rect 29043 6780 29055 6783
rect 29178 6780 29184 6792
rect 29043 6752 29184 6780
rect 29043 6749 29055 6752
rect 28997 6743 29055 6749
rect 29178 6740 29184 6752
rect 29236 6740 29242 6792
rect 31573 6783 31631 6789
rect 31573 6749 31585 6783
rect 31619 6780 31631 6783
rect 31938 6780 31944 6792
rect 31619 6752 31944 6780
rect 31619 6749 31631 6752
rect 31573 6743 31631 6749
rect 31938 6740 31944 6752
rect 31996 6740 32002 6792
rect 29917 6715 29975 6721
rect 29917 6712 29929 6715
rect 27571 6684 28672 6712
rect 28966 6684 29929 6712
rect 27571 6681 27583 6684
rect 27525 6675 27583 6681
rect 27982 6644 27988 6656
rect 27387 6616 27988 6644
rect 27387 6613 27399 6616
rect 27341 6607 27399 6613
rect 27982 6604 27988 6616
rect 28040 6604 28046 6656
rect 28074 6604 28080 6656
rect 28132 6644 28138 6656
rect 28966 6644 28994 6684
rect 29917 6681 29929 6684
rect 29963 6712 29975 6715
rect 30466 6712 30472 6724
rect 29963 6684 30472 6712
rect 29963 6681 29975 6684
rect 29917 6675 29975 6681
rect 30466 6672 30472 6684
rect 30524 6672 30530 6724
rect 28132 6616 28994 6644
rect 28132 6604 28138 6616
rect 29546 6604 29552 6656
rect 29604 6604 29610 6656
rect 29707 6647 29765 6653
rect 29707 6613 29719 6647
rect 29753 6644 29765 6647
rect 29822 6644 29828 6656
rect 29753 6616 29828 6644
rect 29753 6613 29765 6616
rect 29707 6607 29765 6613
rect 29822 6604 29828 6616
rect 29880 6604 29886 6656
rect 1104 6554 38272 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 38272 6554
rect 1104 6480 38272 6502
rect 5994 6400 6000 6452
rect 6052 6400 6058 6452
rect 11790 6400 11796 6452
rect 11848 6400 11854 6452
rect 13357 6443 13415 6449
rect 13357 6409 13369 6443
rect 13403 6440 13415 6443
rect 13817 6443 13875 6449
rect 13817 6440 13829 6443
rect 13403 6412 13829 6440
rect 13403 6409 13415 6412
rect 13357 6403 13415 6409
rect 13817 6409 13829 6412
rect 13863 6440 13875 6443
rect 14090 6440 14096 6452
rect 13863 6412 14096 6440
rect 13863 6409 13875 6412
rect 13817 6403 13875 6409
rect 14090 6400 14096 6412
rect 14148 6400 14154 6452
rect 14274 6400 14280 6452
rect 14332 6440 14338 6452
rect 15562 6440 15568 6452
rect 14332 6412 15568 6440
rect 14332 6400 14338 6412
rect 15562 6400 15568 6412
rect 15620 6400 15626 6452
rect 16942 6400 16948 6452
rect 17000 6440 17006 6452
rect 17037 6443 17095 6449
rect 17037 6440 17049 6443
rect 17000 6412 17049 6440
rect 17000 6400 17006 6412
rect 17037 6409 17049 6412
rect 17083 6409 17095 6443
rect 17037 6403 17095 6409
rect 17221 6443 17279 6449
rect 17221 6409 17233 6443
rect 17267 6440 17279 6443
rect 17402 6440 17408 6452
rect 17267 6412 17408 6440
rect 17267 6409 17279 6412
rect 17221 6403 17279 6409
rect 17402 6400 17408 6412
rect 17460 6400 17466 6452
rect 17589 6443 17647 6449
rect 17589 6409 17601 6443
rect 17635 6440 17647 6443
rect 17770 6440 17776 6452
rect 17635 6412 17776 6440
rect 17635 6409 17647 6412
rect 17589 6403 17647 6409
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 18233 6443 18291 6449
rect 18233 6409 18245 6443
rect 18279 6440 18291 6443
rect 18322 6440 18328 6452
rect 18279 6412 18328 6440
rect 18279 6409 18291 6412
rect 18233 6403 18291 6409
rect 18322 6400 18328 6412
rect 18380 6400 18386 6452
rect 20070 6400 20076 6452
rect 20128 6440 20134 6452
rect 20165 6443 20223 6449
rect 20165 6440 20177 6443
rect 20128 6412 20177 6440
rect 20128 6400 20134 6412
rect 20165 6409 20177 6412
rect 20211 6409 20223 6443
rect 20165 6403 20223 6409
rect 21269 6443 21327 6449
rect 21269 6409 21281 6443
rect 21315 6440 21327 6443
rect 21637 6443 21695 6449
rect 21315 6412 21588 6440
rect 21315 6409 21327 6412
rect 21269 6403 21327 6409
rect 6012 6372 6040 6400
rect 11808 6372 11836 6400
rect 6012 6344 10548 6372
rect 6730 6264 6736 6316
rect 6788 6304 6794 6316
rect 8938 6304 8944 6316
rect 6788 6276 8944 6304
rect 6788 6264 6794 6276
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 10520 6313 10548 6344
rect 11624 6344 11836 6372
rect 11624 6313 11652 6344
rect 13630 6332 13636 6384
rect 13688 6372 13694 6384
rect 13906 6372 13912 6384
rect 13688 6344 13912 6372
rect 13688 6332 13694 6344
rect 13906 6332 13912 6344
rect 13964 6332 13970 6384
rect 21450 6372 21456 6384
rect 17604 6344 21456 6372
rect 17604 6316 17632 6344
rect 21450 6332 21456 6344
rect 21508 6332 21514 6384
rect 21560 6372 21588 6412
rect 21637 6409 21649 6443
rect 21683 6440 21695 6443
rect 22094 6440 22100 6452
rect 21683 6412 22100 6440
rect 21683 6409 21695 6412
rect 21637 6403 21695 6409
rect 22094 6400 22100 6412
rect 22152 6400 22158 6452
rect 22186 6400 22192 6452
rect 22244 6400 22250 6452
rect 22278 6400 22284 6452
rect 22336 6400 22342 6452
rect 22370 6400 22376 6452
rect 22428 6440 22434 6452
rect 22428 6412 22508 6440
rect 22428 6400 22434 6412
rect 21560 6344 22048 6372
rect 10505 6307 10563 6313
rect 10505 6273 10517 6307
rect 10551 6273 10563 6307
rect 10505 6267 10563 6273
rect 11609 6307 11667 6313
rect 11609 6273 11621 6307
rect 11655 6273 11667 6307
rect 13538 6304 13544 6316
rect 13018 6276 13544 6304
rect 11609 6267 11667 6273
rect 10520 6236 10548 6267
rect 13538 6264 13544 6276
rect 13596 6264 13602 6316
rect 15013 6307 15071 6313
rect 15013 6273 15025 6307
rect 15059 6273 15071 6307
rect 15013 6267 15071 6273
rect 10520 6208 11468 6236
rect 5442 6128 5448 6180
rect 5500 6168 5506 6180
rect 11330 6168 11336 6180
rect 5500 6140 11336 6168
rect 5500 6128 5506 6140
rect 11330 6128 11336 6140
rect 11388 6128 11394 6180
rect 8662 6060 8668 6112
rect 8720 6100 8726 6112
rect 8849 6103 8907 6109
rect 8849 6100 8861 6103
rect 8720 6072 8861 6100
rect 8720 6060 8726 6072
rect 8849 6069 8861 6072
rect 8895 6069 8907 6103
rect 8849 6063 8907 6069
rect 10318 6060 10324 6112
rect 10376 6100 10382 6112
rect 10413 6103 10471 6109
rect 10413 6100 10425 6103
rect 10376 6072 10425 6100
rect 10376 6060 10382 6072
rect 10413 6069 10425 6072
rect 10459 6069 10471 6103
rect 11440 6100 11468 6208
rect 11882 6196 11888 6248
rect 11940 6196 11946 6248
rect 13998 6196 14004 6248
rect 14056 6196 14062 6248
rect 15028 6236 15056 6267
rect 16666 6264 16672 6316
rect 16724 6304 16730 6316
rect 17129 6307 17187 6313
rect 17129 6304 17141 6307
rect 16724 6276 17141 6304
rect 16724 6264 16730 6276
rect 17129 6273 17141 6276
rect 17175 6304 17187 6307
rect 17402 6304 17408 6316
rect 17175 6276 17408 6304
rect 17175 6273 17187 6276
rect 17129 6267 17187 6273
rect 17402 6264 17408 6276
rect 17460 6264 17466 6316
rect 17497 6307 17555 6313
rect 17497 6273 17509 6307
rect 17543 6273 17555 6307
rect 17497 6267 17555 6273
rect 17034 6236 17040 6248
rect 15028 6208 17040 6236
rect 13814 6168 13820 6180
rect 13372 6140 13820 6168
rect 13372 6100 13400 6140
rect 13814 6128 13820 6140
rect 13872 6168 13878 6180
rect 15028 6168 15056 6208
rect 17034 6196 17040 6208
rect 17092 6196 17098 6248
rect 17512 6236 17540 6267
rect 17586 6264 17592 6316
rect 17644 6264 17650 6316
rect 17770 6264 17776 6316
rect 17828 6264 17834 6316
rect 17957 6307 18015 6313
rect 17957 6273 17969 6307
rect 18003 6304 18015 6307
rect 18046 6304 18052 6316
rect 18003 6276 18052 6304
rect 18003 6273 18015 6276
rect 17957 6267 18015 6273
rect 18046 6264 18052 6276
rect 18104 6264 18110 6316
rect 19981 6307 20039 6313
rect 19981 6304 19993 6307
rect 19260 6276 19993 6304
rect 18138 6236 18144 6248
rect 17512 6208 18144 6236
rect 18138 6196 18144 6208
rect 18196 6196 18202 6248
rect 13872 6140 15056 6168
rect 13872 6128 13878 6140
rect 15470 6128 15476 6180
rect 15528 6168 15534 6180
rect 16853 6171 16911 6177
rect 16853 6168 16865 6171
rect 15528 6140 16865 6168
rect 15528 6128 15534 6140
rect 16853 6137 16865 6140
rect 16899 6137 16911 6171
rect 16853 6131 16911 6137
rect 16942 6128 16948 6180
rect 17000 6128 17006 6180
rect 17405 6171 17463 6177
rect 17405 6137 17417 6171
rect 17451 6168 17463 6171
rect 17865 6171 17923 6177
rect 17865 6168 17877 6171
rect 17451 6140 17877 6168
rect 17451 6137 17463 6140
rect 17405 6131 17463 6137
rect 17865 6137 17877 6140
rect 17911 6137 17923 6171
rect 17865 6131 17923 6137
rect 17954 6128 17960 6180
rect 18012 6168 18018 6180
rect 19260 6168 19288 6276
rect 19981 6273 19993 6276
rect 20027 6304 20039 6307
rect 21358 6304 21364 6316
rect 20027 6276 21364 6304
rect 20027 6273 20039 6276
rect 19981 6267 20039 6273
rect 21358 6264 21364 6276
rect 21416 6264 21422 6316
rect 21560 6304 21588 6344
rect 22020 6316 22048 6344
rect 21468 6276 21588 6304
rect 19797 6239 19855 6245
rect 19797 6205 19809 6239
rect 19843 6236 19855 6239
rect 21468 6236 21496 6276
rect 21910 6264 21916 6316
rect 21968 6264 21974 6316
rect 22002 6264 22008 6316
rect 22060 6264 22066 6316
rect 22204 6313 22232 6400
rect 22296 6313 22324 6400
rect 22097 6307 22155 6313
rect 22097 6273 22109 6307
rect 22143 6273 22155 6307
rect 22097 6267 22155 6273
rect 22189 6307 22247 6313
rect 22189 6273 22201 6307
rect 22235 6273 22247 6307
rect 22189 6267 22247 6273
rect 22281 6307 22339 6313
rect 22281 6273 22293 6307
rect 22327 6273 22339 6307
rect 22281 6267 22339 6273
rect 22373 6307 22431 6313
rect 22373 6273 22385 6307
rect 22419 6304 22431 6307
rect 22480 6304 22508 6412
rect 23014 6400 23020 6452
rect 23072 6400 23078 6452
rect 23474 6400 23480 6452
rect 23532 6400 23538 6452
rect 23842 6400 23848 6452
rect 23900 6440 23906 6452
rect 24397 6443 24455 6449
rect 24397 6440 24409 6443
rect 23900 6412 24409 6440
rect 23900 6400 23906 6412
rect 24397 6409 24409 6412
rect 24443 6409 24455 6443
rect 24397 6403 24455 6409
rect 24486 6400 24492 6452
rect 24544 6400 24550 6452
rect 24854 6400 24860 6452
rect 24912 6400 24918 6452
rect 25501 6443 25559 6449
rect 25501 6409 25513 6443
rect 25547 6440 25559 6443
rect 25590 6440 25596 6452
rect 25547 6412 25596 6440
rect 25547 6409 25559 6412
rect 25501 6403 25559 6409
rect 25590 6400 25596 6412
rect 25648 6400 25654 6452
rect 26418 6400 26424 6452
rect 26476 6440 26482 6452
rect 27890 6440 27896 6452
rect 26476 6412 27896 6440
rect 26476 6400 26482 6412
rect 27890 6400 27896 6412
rect 27948 6400 27954 6452
rect 28077 6443 28135 6449
rect 28077 6409 28089 6443
rect 28123 6440 28135 6443
rect 28718 6440 28724 6452
rect 28123 6412 28724 6440
rect 28123 6409 28135 6412
rect 28077 6403 28135 6409
rect 28718 6400 28724 6412
rect 28776 6400 28782 6452
rect 29822 6400 29828 6452
rect 29880 6400 29886 6452
rect 23032 6372 23060 6400
rect 23032 6344 23336 6372
rect 22419 6276 22508 6304
rect 22419 6273 22431 6276
rect 22373 6267 22431 6273
rect 19843 6208 21496 6236
rect 19843 6205 19855 6208
rect 19797 6199 19855 6205
rect 18012 6140 19288 6168
rect 18012 6128 18018 6140
rect 11440 6072 13400 6100
rect 10413 6063 10471 6069
rect 13446 6060 13452 6112
rect 13504 6060 13510 6112
rect 14734 6060 14740 6112
rect 14792 6100 14798 6112
rect 14921 6103 14979 6109
rect 14921 6100 14933 6103
rect 14792 6072 14933 6100
rect 14792 6060 14798 6072
rect 14921 6069 14933 6072
rect 14967 6069 14979 6103
rect 16960 6100 16988 6128
rect 19812 6100 19840 6199
rect 21542 6196 21548 6248
rect 21600 6236 21606 6248
rect 22112 6236 22140 6267
rect 23198 6264 23204 6316
rect 23256 6264 23262 6316
rect 23308 6313 23336 6344
rect 24302 6332 24308 6384
rect 24360 6372 24366 6384
rect 26053 6375 26111 6381
rect 26053 6372 26065 6375
rect 24360 6344 26065 6372
rect 24360 6332 24366 6344
rect 26053 6341 26065 6344
rect 26099 6372 26111 6375
rect 26878 6372 26884 6384
rect 26099 6344 26884 6372
rect 26099 6341 26111 6344
rect 26053 6335 26111 6341
rect 26878 6332 26884 6344
rect 26936 6332 26942 6384
rect 27154 6332 27160 6384
rect 27212 6372 27218 6384
rect 27709 6375 27767 6381
rect 27709 6372 27721 6375
rect 27212 6344 27721 6372
rect 27212 6332 27218 6344
rect 27709 6341 27721 6344
rect 27755 6341 27767 6375
rect 27709 6335 27767 6341
rect 23293 6307 23351 6313
rect 23293 6273 23305 6307
rect 23339 6273 23351 6307
rect 23293 6267 23351 6273
rect 24578 6264 24584 6316
rect 24636 6264 24642 6316
rect 25133 6307 25191 6313
rect 25133 6273 25145 6307
rect 25179 6304 25191 6307
rect 25179 6276 25452 6304
rect 25179 6273 25191 6276
rect 25133 6267 25191 6273
rect 21600 6208 22140 6236
rect 21600 6196 21606 6208
rect 22830 6196 22836 6248
rect 22888 6236 22894 6248
rect 22925 6239 22983 6245
rect 22925 6236 22937 6239
rect 22888 6208 22937 6236
rect 22888 6196 22894 6208
rect 22925 6205 22937 6208
rect 22971 6205 22983 6239
rect 22925 6199 22983 6205
rect 24213 6239 24271 6245
rect 24213 6205 24225 6239
rect 24259 6236 24271 6239
rect 25317 6239 25375 6245
rect 25317 6236 25329 6239
rect 24259 6208 25329 6236
rect 24259 6205 24271 6208
rect 24213 6199 24271 6205
rect 25317 6205 25329 6208
rect 25363 6205 25375 6239
rect 25424 6236 25452 6276
rect 25590 6264 25596 6316
rect 25648 6264 25654 6316
rect 25866 6264 25872 6316
rect 25924 6264 25930 6316
rect 25958 6264 25964 6316
rect 26016 6264 26022 6316
rect 26142 6264 26148 6316
rect 26200 6304 26206 6316
rect 26237 6307 26295 6313
rect 26237 6304 26249 6307
rect 26200 6276 26249 6304
rect 26200 6264 26206 6276
rect 26237 6273 26249 6276
rect 26283 6304 26295 6307
rect 26283 6276 26832 6304
rect 26283 6273 26295 6276
rect 26237 6267 26295 6273
rect 26694 6236 26700 6248
rect 25424 6208 26700 6236
rect 25317 6199 25375 6205
rect 26694 6196 26700 6208
rect 26752 6196 26758 6248
rect 26804 6236 26832 6276
rect 27246 6264 27252 6316
rect 27304 6304 27310 6316
rect 27801 6307 27859 6313
rect 27801 6304 27813 6307
rect 27304 6276 27813 6304
rect 27304 6264 27310 6276
rect 27801 6273 27813 6276
rect 27847 6273 27859 6307
rect 27801 6267 27859 6273
rect 27890 6264 27896 6316
rect 27948 6304 27954 6316
rect 29840 6304 29868 6400
rect 27948 6276 29868 6304
rect 27948 6264 27954 6276
rect 30190 6264 30196 6316
rect 30248 6264 30254 6316
rect 28074 6236 28080 6248
rect 26804 6208 28080 6236
rect 28074 6196 28080 6208
rect 28132 6196 28138 6248
rect 21085 6171 21143 6177
rect 21085 6137 21097 6171
rect 21131 6168 21143 6171
rect 22278 6168 22284 6180
rect 21131 6140 22284 6168
rect 21131 6137 21143 6140
rect 21085 6131 21143 6137
rect 22278 6128 22284 6140
rect 22336 6128 22342 6180
rect 24765 6171 24823 6177
rect 24765 6137 24777 6171
rect 24811 6168 24823 6171
rect 26326 6168 26332 6180
rect 24811 6140 26332 6168
rect 24811 6137 24823 6140
rect 24765 6131 24823 6137
rect 26326 6128 26332 6140
rect 26384 6128 26390 6180
rect 26786 6128 26792 6180
rect 26844 6168 26850 6180
rect 27062 6168 27068 6180
rect 26844 6140 27068 6168
rect 26844 6128 26850 6140
rect 27062 6128 27068 6140
rect 27120 6168 27126 6180
rect 27525 6171 27583 6177
rect 27525 6168 27537 6171
rect 27120 6140 27537 6168
rect 27120 6128 27126 6140
rect 27525 6137 27537 6140
rect 27571 6137 27583 6171
rect 27525 6131 27583 6137
rect 16960 6072 19840 6100
rect 22557 6103 22615 6109
rect 14921 6063 14979 6069
rect 22557 6069 22569 6103
rect 22603 6100 22615 6103
rect 23017 6103 23075 6109
rect 23017 6100 23029 6103
rect 22603 6072 23029 6100
rect 22603 6069 22615 6072
rect 22557 6063 22615 6069
rect 23017 6069 23029 6072
rect 23063 6069 23075 6103
rect 23017 6063 23075 6069
rect 24946 6060 24952 6112
rect 25004 6100 25010 6112
rect 25225 6103 25283 6109
rect 25225 6100 25237 6103
rect 25004 6072 25237 6100
rect 25004 6060 25010 6072
rect 25225 6069 25237 6072
rect 25271 6069 25283 6103
rect 25225 6063 25283 6069
rect 25314 6060 25320 6112
rect 25372 6100 25378 6112
rect 25685 6103 25743 6109
rect 25685 6100 25697 6103
rect 25372 6072 25697 6100
rect 25372 6060 25378 6072
rect 25685 6069 25697 6072
rect 25731 6069 25743 6103
rect 25685 6063 25743 6069
rect 30006 6060 30012 6112
rect 30064 6060 30070 6112
rect 1104 6010 38272 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38272 6010
rect 1104 5936 38272 5958
rect 10318 5856 10324 5908
rect 10376 5856 10382 5908
rect 11882 5856 11888 5908
rect 11940 5896 11946 5908
rect 12345 5899 12403 5905
rect 12345 5896 12357 5899
rect 11940 5868 12357 5896
rect 11940 5856 11946 5868
rect 12345 5865 12357 5868
rect 12391 5865 12403 5899
rect 12345 5859 12403 5865
rect 14642 5856 14648 5908
rect 14700 5856 14706 5908
rect 23658 5896 23664 5908
rect 15488 5868 23664 5896
rect 9309 5831 9367 5837
rect 9309 5797 9321 5831
rect 9355 5797 9367 5831
rect 9309 5791 9367 5797
rect 5537 5763 5595 5769
rect 5537 5729 5549 5763
rect 5583 5760 5595 5763
rect 5718 5760 5724 5772
rect 5583 5732 5724 5760
rect 5583 5729 5595 5732
rect 5537 5723 5595 5729
rect 5718 5720 5724 5732
rect 5776 5720 5782 5772
rect 6549 5763 6607 5769
rect 6549 5729 6561 5763
rect 6595 5760 6607 5763
rect 6733 5763 6791 5769
rect 6733 5760 6745 5763
rect 6595 5732 6745 5760
rect 6595 5729 6607 5732
rect 6549 5723 6607 5729
rect 6733 5729 6745 5732
rect 6779 5729 6791 5763
rect 6733 5723 6791 5729
rect 8570 5720 8576 5772
rect 8628 5760 8634 5772
rect 8757 5763 8815 5769
rect 8757 5760 8769 5763
rect 8628 5732 8769 5760
rect 8628 5720 8634 5732
rect 8757 5729 8769 5732
rect 8803 5760 8815 5763
rect 9122 5760 9128 5772
rect 8803 5732 9128 5760
rect 8803 5729 8815 5732
rect 8757 5723 8815 5729
rect 9122 5720 9128 5732
rect 9180 5720 9186 5772
rect 5353 5695 5411 5701
rect 5353 5661 5365 5695
rect 5399 5692 5411 5695
rect 5442 5692 5448 5704
rect 5399 5664 5448 5692
rect 5399 5661 5411 5664
rect 5353 5655 5411 5661
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5692 6699 5695
rect 9217 5695 9275 5701
rect 6687 5664 6776 5692
rect 6687 5661 6699 5664
rect 6641 5655 6699 5661
rect 6748 5636 6776 5664
rect 9217 5661 9229 5695
rect 9263 5692 9275 5695
rect 9324 5692 9352 5791
rect 9766 5720 9772 5772
rect 9824 5720 9830 5772
rect 9950 5720 9956 5772
rect 10008 5720 10014 5772
rect 10229 5763 10287 5769
rect 10229 5729 10241 5763
rect 10275 5760 10287 5763
rect 10336 5760 10364 5856
rect 14660 5828 14688 5856
rect 14826 5828 14832 5840
rect 12406 5800 14832 5828
rect 10275 5732 10364 5760
rect 10275 5729 10287 5732
rect 10229 5723 10287 5729
rect 10594 5720 10600 5772
rect 10652 5760 10658 5772
rect 11514 5760 11520 5772
rect 10652 5732 11520 5760
rect 10652 5720 10658 5732
rect 11514 5720 11520 5732
rect 11572 5720 11578 5772
rect 12250 5720 12256 5772
rect 12308 5720 12314 5772
rect 9263 5664 9352 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 6730 5584 6736 5636
rect 6788 5584 6794 5636
rect 7006 5584 7012 5636
rect 7064 5584 7070 5636
rect 7742 5584 7748 5636
rect 7800 5584 7806 5636
rect 9677 5627 9735 5633
rect 9677 5624 9689 5627
rect 8312 5596 9689 5624
rect 4154 5516 4160 5568
rect 4212 5556 4218 5568
rect 5169 5559 5227 5565
rect 5169 5556 5181 5559
rect 4212 5528 5181 5556
rect 4212 5516 4218 5528
rect 5169 5525 5181 5528
rect 5215 5525 5227 5559
rect 5169 5519 5227 5525
rect 8018 5516 8024 5568
rect 8076 5556 8082 5568
rect 8312 5556 8340 5596
rect 9677 5593 9689 5596
rect 9723 5593 9735 5627
rect 9784 5624 9812 5720
rect 12406 5692 12434 5800
rect 14826 5788 14832 5800
rect 14884 5788 14890 5840
rect 13446 5760 13452 5772
rect 12544 5732 13452 5760
rect 12544 5701 12572 5732
rect 13446 5720 13452 5732
rect 13504 5720 13510 5772
rect 14737 5763 14795 5769
rect 14737 5729 14749 5763
rect 14783 5760 14795 5763
rect 14918 5760 14924 5772
rect 14783 5732 14924 5760
rect 14783 5729 14795 5732
rect 14737 5723 14795 5729
rect 14918 5720 14924 5732
rect 14976 5760 14982 5772
rect 15488 5760 15516 5868
rect 23658 5856 23664 5868
rect 23716 5856 23722 5908
rect 24765 5899 24823 5905
rect 24765 5865 24777 5899
rect 24811 5896 24823 5899
rect 24946 5896 24952 5908
rect 24811 5868 24952 5896
rect 24811 5865 24823 5868
rect 24765 5859 24823 5865
rect 24946 5856 24952 5868
rect 25004 5856 25010 5908
rect 31478 5856 31484 5908
rect 31536 5856 31542 5908
rect 17402 5788 17408 5840
rect 17460 5828 17466 5840
rect 17862 5828 17868 5840
rect 17460 5800 17868 5828
rect 17460 5788 17466 5800
rect 17862 5788 17868 5800
rect 17920 5788 17926 5840
rect 18506 5788 18512 5840
rect 18564 5828 18570 5840
rect 23382 5828 23388 5840
rect 18564 5800 23388 5828
rect 18564 5788 18570 5800
rect 23382 5788 23388 5800
rect 23440 5788 23446 5840
rect 25317 5831 25375 5837
rect 25317 5797 25329 5831
rect 25363 5828 25375 5831
rect 26418 5828 26424 5840
rect 25363 5800 26424 5828
rect 25363 5797 25375 5800
rect 25317 5791 25375 5797
rect 26418 5788 26424 5800
rect 26476 5788 26482 5840
rect 14976 5732 15516 5760
rect 14976 5720 14982 5732
rect 15562 5720 15568 5772
rect 15620 5760 15626 5772
rect 22554 5760 22560 5772
rect 15620 5732 22560 5760
rect 15620 5720 15626 5732
rect 22554 5720 22560 5732
rect 22612 5720 22618 5772
rect 25130 5720 25136 5772
rect 25188 5720 25194 5772
rect 29917 5763 29975 5769
rect 29917 5729 29929 5763
rect 29963 5760 29975 5763
rect 30006 5760 30012 5772
rect 29963 5732 30012 5760
rect 29963 5729 29975 5732
rect 29917 5723 29975 5729
rect 30006 5720 30012 5732
rect 30064 5720 30070 5772
rect 31496 5760 31524 5856
rect 31036 5732 32904 5760
rect 11638 5664 12434 5692
rect 12529 5695 12587 5701
rect 12529 5661 12541 5695
rect 12575 5661 12587 5695
rect 12529 5655 12587 5661
rect 12618 5652 12624 5704
rect 12676 5692 12682 5704
rect 13081 5695 13139 5701
rect 13081 5692 13093 5695
rect 12676 5664 13093 5692
rect 12676 5652 12682 5664
rect 13081 5661 13093 5664
rect 13127 5661 13139 5695
rect 13081 5655 13139 5661
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 14461 5695 14519 5701
rect 14461 5692 14473 5695
rect 13964 5664 14473 5692
rect 13964 5652 13970 5664
rect 14461 5661 14473 5664
rect 14507 5692 14519 5695
rect 15289 5695 15347 5701
rect 14507 5664 15240 5692
rect 14507 5661 14519 5664
rect 14461 5655 14519 5661
rect 10226 5624 10232 5636
rect 9784 5596 10232 5624
rect 9677 5587 9735 5593
rect 10226 5584 10232 5596
rect 10284 5584 10290 5636
rect 10505 5627 10563 5633
rect 10505 5593 10517 5627
rect 10551 5624 10563 5627
rect 10594 5624 10600 5636
rect 10551 5596 10600 5624
rect 10551 5593 10563 5596
rect 10505 5587 10563 5593
rect 10594 5584 10600 5596
rect 10652 5584 10658 5636
rect 15212 5624 15240 5664
rect 15289 5661 15301 5695
rect 15335 5692 15347 5695
rect 15654 5692 15660 5704
rect 15335 5664 15660 5692
rect 15335 5661 15347 5664
rect 15289 5655 15347 5661
rect 15654 5652 15660 5664
rect 15712 5692 15718 5704
rect 17221 5695 17279 5701
rect 17221 5692 17233 5695
rect 15712 5664 17233 5692
rect 15712 5652 15718 5664
rect 17221 5661 17233 5664
rect 17267 5661 17279 5695
rect 17221 5655 17279 5661
rect 17402 5652 17408 5704
rect 17460 5692 17466 5704
rect 17497 5695 17555 5701
rect 17497 5692 17509 5695
rect 17460 5664 17509 5692
rect 17460 5652 17466 5664
rect 17497 5661 17509 5664
rect 17543 5661 17555 5695
rect 17497 5655 17555 5661
rect 17586 5652 17592 5704
rect 17644 5652 17650 5704
rect 19426 5652 19432 5704
rect 19484 5652 19490 5704
rect 19521 5695 19579 5701
rect 19521 5661 19533 5695
rect 19567 5661 19579 5695
rect 19521 5655 19579 5661
rect 15212 5596 15424 5624
rect 8076 5528 8340 5556
rect 8076 5516 8082 5528
rect 9030 5516 9036 5568
rect 9088 5516 9094 5568
rect 12802 5516 12808 5568
rect 12860 5556 12866 5568
rect 12989 5559 13047 5565
rect 12989 5556 13001 5559
rect 12860 5528 13001 5556
rect 12860 5516 12866 5528
rect 12989 5525 13001 5528
rect 13035 5525 13047 5559
rect 12989 5519 13047 5525
rect 14090 5516 14096 5568
rect 14148 5516 14154 5568
rect 14550 5516 14556 5568
rect 14608 5516 14614 5568
rect 14921 5559 14979 5565
rect 14921 5525 14933 5559
rect 14967 5556 14979 5559
rect 15194 5556 15200 5568
rect 14967 5528 15200 5556
rect 14967 5525 14979 5528
rect 14921 5519 14979 5525
rect 15194 5516 15200 5528
rect 15252 5516 15258 5568
rect 15396 5565 15424 5596
rect 16942 5584 16948 5636
rect 17000 5584 17006 5636
rect 17034 5584 17040 5636
rect 17092 5624 17098 5636
rect 19536 5624 19564 5655
rect 21450 5652 21456 5704
rect 21508 5692 21514 5704
rect 24949 5695 25007 5701
rect 24949 5692 24961 5695
rect 21508 5664 24961 5692
rect 21508 5652 21514 5664
rect 24949 5661 24961 5664
rect 24995 5692 25007 5695
rect 25148 5692 25176 5720
rect 31036 5704 31064 5732
rect 24995 5664 25176 5692
rect 24995 5661 25007 5664
rect 24949 5655 25007 5661
rect 29638 5652 29644 5704
rect 29696 5652 29702 5704
rect 31018 5652 31024 5704
rect 31076 5652 31082 5704
rect 31478 5652 31484 5704
rect 31536 5652 31542 5704
rect 32876 5678 32904 5732
rect 17092 5596 19564 5624
rect 17092 5584 17098 5596
rect 22002 5584 22008 5636
rect 22060 5624 22066 5636
rect 24578 5624 24584 5636
rect 22060 5596 24584 5624
rect 22060 5584 22066 5596
rect 24578 5584 24584 5596
rect 24636 5624 24642 5636
rect 25133 5627 25191 5633
rect 25133 5624 25145 5627
rect 24636 5596 25145 5624
rect 24636 5584 24642 5596
rect 25133 5593 25145 5596
rect 25179 5593 25191 5627
rect 25133 5587 25191 5593
rect 31754 5584 31760 5636
rect 31812 5584 31818 5636
rect 32030 5584 32036 5636
rect 32088 5584 32094 5636
rect 15381 5559 15439 5565
rect 15381 5525 15393 5559
rect 15427 5525 15439 5559
rect 16960 5556 16988 5584
rect 17405 5559 17463 5565
rect 17405 5556 17417 5559
rect 16960 5528 17417 5556
rect 15381 5519 15439 5525
rect 17405 5525 17417 5528
rect 17451 5525 17463 5559
rect 17405 5519 17463 5525
rect 17770 5516 17776 5568
rect 17828 5516 17834 5568
rect 19242 5516 19248 5568
rect 19300 5516 19306 5568
rect 19610 5516 19616 5568
rect 19668 5516 19674 5568
rect 21358 5516 21364 5568
rect 21416 5556 21422 5568
rect 24486 5556 24492 5568
rect 21416 5528 24492 5556
rect 21416 5516 21422 5528
rect 24486 5516 24492 5528
rect 24544 5556 24550 5568
rect 25041 5559 25099 5565
rect 25041 5556 25053 5559
rect 24544 5528 25053 5556
rect 24544 5516 24550 5528
rect 25041 5525 25053 5528
rect 25087 5525 25099 5559
rect 25041 5519 25099 5525
rect 31386 5516 31392 5568
rect 31444 5516 31450 5568
rect 32048 5556 32076 5584
rect 33229 5559 33287 5565
rect 33229 5556 33241 5559
rect 32048 5528 33241 5556
rect 33229 5525 33241 5528
rect 33275 5525 33287 5559
rect 33229 5519 33287 5525
rect 1104 5466 38272 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 38272 5466
rect 1104 5392 38272 5414
rect 5537 5355 5595 5361
rect 5537 5321 5549 5355
rect 5583 5352 5595 5355
rect 18874 5352 18880 5364
rect 5583 5324 18880 5352
rect 5583 5321 5595 5324
rect 5537 5315 5595 5321
rect 18874 5312 18880 5324
rect 18932 5312 18938 5364
rect 19610 5312 19616 5364
rect 19668 5312 19674 5364
rect 22554 5312 22560 5364
rect 22612 5352 22618 5364
rect 27338 5352 27344 5364
rect 22612 5324 27344 5352
rect 22612 5312 22618 5324
rect 27338 5312 27344 5324
rect 27396 5312 27402 5364
rect 27433 5355 27491 5361
rect 27433 5321 27445 5355
rect 27479 5352 27491 5355
rect 28074 5352 28080 5364
rect 27479 5324 28080 5352
rect 27479 5321 27491 5324
rect 27433 5315 27491 5321
rect 28074 5312 28080 5324
rect 28132 5312 28138 5364
rect 29638 5312 29644 5364
rect 29696 5352 29702 5364
rect 29825 5355 29883 5361
rect 29825 5352 29837 5355
rect 29696 5324 29837 5352
rect 29696 5312 29702 5324
rect 29825 5321 29837 5324
rect 29871 5321 29883 5355
rect 29825 5315 29883 5321
rect 30009 5355 30067 5361
rect 30009 5321 30021 5355
rect 30055 5352 30067 5355
rect 30190 5352 30196 5364
rect 30055 5324 30196 5352
rect 30055 5321 30067 5324
rect 30009 5315 30067 5321
rect 30190 5312 30196 5324
rect 30248 5312 30254 5364
rect 30377 5355 30435 5361
rect 30377 5321 30389 5355
rect 30423 5352 30435 5355
rect 30466 5352 30472 5364
rect 30423 5324 30472 5352
rect 30423 5321 30435 5324
rect 30377 5315 30435 5321
rect 30466 5312 30472 5324
rect 30524 5352 30530 5364
rect 31386 5352 31392 5364
rect 30524 5324 31392 5352
rect 30524 5312 30530 5324
rect 31386 5312 31392 5324
rect 31444 5312 31450 5364
rect 31478 5312 31484 5364
rect 31536 5352 31542 5364
rect 31665 5355 31723 5361
rect 31665 5352 31677 5355
rect 31536 5324 31677 5352
rect 31536 5312 31542 5324
rect 31665 5321 31677 5324
rect 31711 5321 31723 5355
rect 31665 5315 31723 5321
rect 32030 5312 32036 5364
rect 32088 5352 32094 5364
rect 32493 5355 32551 5361
rect 32493 5352 32505 5355
rect 32088 5324 32505 5352
rect 32088 5312 32094 5324
rect 32493 5321 32505 5324
rect 32539 5321 32551 5355
rect 32493 5315 32551 5321
rect 8021 5287 8079 5293
rect 8021 5253 8033 5287
rect 8067 5284 8079 5287
rect 8570 5284 8576 5296
rect 8067 5256 8576 5284
rect 8067 5253 8079 5256
rect 8021 5247 8079 5253
rect 8570 5244 8576 5256
rect 8628 5244 8634 5296
rect 8941 5287 8999 5293
rect 8941 5253 8953 5287
rect 8987 5284 8999 5287
rect 9030 5284 9036 5296
rect 8987 5256 9036 5284
rect 8987 5253 8999 5256
rect 8941 5247 8999 5253
rect 9030 5244 9036 5256
rect 9088 5244 9094 5296
rect 10226 5244 10232 5296
rect 10284 5284 10290 5296
rect 10689 5287 10747 5293
rect 10689 5284 10701 5287
rect 10284 5256 10701 5284
rect 10284 5244 10290 5256
rect 10689 5253 10701 5256
rect 10735 5253 10747 5287
rect 10689 5247 10747 5253
rect 11054 5244 11060 5296
rect 11112 5284 11118 5296
rect 11977 5287 12035 5293
rect 11112 5256 11836 5284
rect 11112 5244 11118 5256
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5216 2007 5219
rect 4154 5216 4160 5228
rect 1995 5188 4160 5216
rect 1995 5185 2007 5188
rect 1949 5179 2007 5185
rect 4154 5176 4160 5188
rect 4212 5176 4218 5228
rect 5353 5219 5411 5225
rect 5353 5185 5365 5219
rect 5399 5185 5411 5219
rect 5353 5179 5411 5185
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5216 7527 5219
rect 10965 5219 11023 5225
rect 7515 5188 7696 5216
rect 10074 5188 10916 5216
rect 7515 5185 7527 5188
rect 7469 5179 7527 5185
rect 5368 5148 5396 5179
rect 6914 5148 6920 5160
rect 5368 5120 6920 5148
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7006 5040 7012 5092
rect 7064 5080 7070 5092
rect 7668 5089 7696 5188
rect 8018 5108 8024 5160
rect 8076 5148 8082 5160
rect 8113 5151 8171 5157
rect 8113 5148 8125 5151
rect 8076 5120 8125 5148
rect 8076 5108 8082 5120
rect 8113 5117 8125 5120
rect 8159 5117 8171 5151
rect 8113 5111 8171 5117
rect 8205 5151 8263 5157
rect 8205 5117 8217 5151
rect 8251 5148 8263 5151
rect 8294 5148 8300 5160
rect 8251 5120 8300 5148
rect 8251 5117 8263 5120
rect 8205 5111 8263 5117
rect 8294 5108 8300 5120
rect 8352 5108 8358 5160
rect 8662 5108 8668 5160
rect 8720 5108 8726 5160
rect 10594 5108 10600 5160
rect 10652 5108 10658 5160
rect 10888 5148 10916 5188
rect 10965 5185 10977 5219
rect 11011 5216 11023 5219
rect 11011 5188 11560 5216
rect 11011 5185 11023 5188
rect 10965 5179 11023 5185
rect 11422 5148 11428 5160
rect 10888 5120 11428 5148
rect 11422 5108 11428 5120
rect 11480 5108 11486 5160
rect 7285 5083 7343 5089
rect 7285 5080 7297 5083
rect 7064 5052 7297 5080
rect 7064 5040 7070 5052
rect 7285 5049 7297 5052
rect 7331 5049 7343 5083
rect 7285 5043 7343 5049
rect 7653 5083 7711 5089
rect 7653 5049 7665 5083
rect 7699 5049 7711 5083
rect 7653 5043 7711 5049
rect 1762 4972 1768 5024
rect 1820 4972 1826 5024
rect 8312 5012 8340 5108
rect 10612 5080 10640 5108
rect 11532 5089 11560 5188
rect 11808 5148 11836 5256
rect 11977 5253 11989 5287
rect 12023 5284 12035 5287
rect 12250 5284 12256 5296
rect 12023 5256 12256 5284
rect 12023 5253 12035 5256
rect 11977 5247 12035 5253
rect 12250 5244 12256 5256
rect 12308 5244 12314 5296
rect 13170 5284 13176 5296
rect 12728 5256 13176 5284
rect 11882 5176 11888 5228
rect 11940 5216 11946 5228
rect 12728 5216 12756 5256
rect 13170 5244 13176 5256
rect 13228 5244 13234 5296
rect 13538 5244 13544 5296
rect 13596 5244 13602 5296
rect 19628 5284 19656 5312
rect 22186 5284 22192 5296
rect 18984 5256 19656 5284
rect 20470 5256 22192 5284
rect 17678 5216 17684 5228
rect 11940 5188 12756 5216
rect 16146 5188 17684 5216
rect 11940 5176 11946 5188
rect 12069 5151 12127 5157
rect 12069 5148 12081 5151
rect 11808 5120 12081 5148
rect 12069 5117 12081 5120
rect 12115 5148 12127 5151
rect 12618 5148 12624 5160
rect 12115 5120 12624 5148
rect 12115 5117 12127 5120
rect 12069 5111 12127 5117
rect 12618 5108 12624 5120
rect 12676 5108 12682 5160
rect 12802 5108 12808 5160
rect 12860 5108 12866 5160
rect 13078 5108 13084 5160
rect 13136 5108 13142 5160
rect 14550 5108 14556 5160
rect 14608 5108 14614 5160
rect 14734 5108 14740 5160
rect 14792 5108 14798 5160
rect 15010 5108 15016 5160
rect 15068 5108 15074 5160
rect 15654 5108 15660 5160
rect 15712 5148 15718 5160
rect 16485 5151 16543 5157
rect 16485 5148 16497 5151
rect 15712 5120 16497 5148
rect 15712 5108 15718 5120
rect 16485 5117 16497 5120
rect 16531 5117 16543 5151
rect 16485 5111 16543 5117
rect 10781 5083 10839 5089
rect 10781 5080 10793 5083
rect 10612 5052 10793 5080
rect 10781 5049 10793 5052
rect 10827 5049 10839 5083
rect 10781 5043 10839 5049
rect 11517 5083 11575 5089
rect 11517 5049 11529 5083
rect 11563 5049 11575 5083
rect 11517 5043 11575 5049
rect 11054 5012 11060 5024
rect 8312 4984 11060 5012
rect 11054 4972 11060 4984
rect 11112 4972 11118 5024
rect 14826 4972 14832 5024
rect 14884 5012 14890 5024
rect 16592 5012 16620 5188
rect 17678 5176 17684 5188
rect 17736 5176 17742 5228
rect 18984 5225 19012 5256
rect 22186 5244 22192 5256
rect 22244 5244 22250 5296
rect 22373 5287 22431 5293
rect 22373 5253 22385 5287
rect 22419 5284 22431 5287
rect 23290 5284 23296 5296
rect 22419 5256 23296 5284
rect 22419 5253 22431 5256
rect 22373 5247 22431 5253
rect 23290 5244 23296 5256
rect 23348 5244 23354 5296
rect 23382 5244 23388 5296
rect 23440 5284 23446 5296
rect 23440 5256 27823 5284
rect 23440 5244 23446 5256
rect 18969 5219 19027 5225
rect 18969 5185 18981 5219
rect 19015 5185 19027 5219
rect 18969 5179 19027 5185
rect 22278 5176 22284 5228
rect 22336 5216 22342 5228
rect 22830 5216 22836 5228
rect 22336 5188 22836 5216
rect 22336 5176 22342 5188
rect 22830 5176 22836 5188
rect 22888 5176 22894 5228
rect 23308 5216 23336 5244
rect 23845 5219 23903 5225
rect 23845 5216 23857 5219
rect 23308 5188 23857 5216
rect 23845 5185 23857 5188
rect 23891 5185 23903 5219
rect 23845 5179 23903 5185
rect 23934 5176 23940 5228
rect 23992 5176 23998 5228
rect 24044 5188 26556 5216
rect 19242 5108 19248 5160
rect 19300 5108 19306 5160
rect 22554 5108 22560 5160
rect 22612 5108 22618 5160
rect 23658 5108 23664 5160
rect 23716 5108 23722 5160
rect 23753 5151 23811 5157
rect 23753 5117 23765 5151
rect 23799 5148 23811 5151
rect 23952 5148 23980 5176
rect 23799 5120 23980 5148
rect 23799 5117 23811 5120
rect 23753 5111 23811 5117
rect 24044 5080 24072 5188
rect 26528 5160 26556 5188
rect 26970 5176 26976 5228
rect 27028 5176 27034 5228
rect 27246 5176 27252 5228
rect 27304 5176 27310 5228
rect 27709 5219 27767 5225
rect 27709 5216 27721 5219
rect 27632 5188 27721 5216
rect 27632 5160 27660 5188
rect 27709 5185 27721 5188
rect 27755 5185 27767 5219
rect 27709 5179 27767 5185
rect 26510 5108 26516 5160
rect 26568 5108 26574 5160
rect 27614 5108 27620 5160
rect 27672 5108 27678 5160
rect 27795 5148 27823 5256
rect 28092 5256 31800 5284
rect 27890 5176 27896 5228
rect 27948 5216 27954 5228
rect 28092 5225 28120 5256
rect 28077 5219 28135 5225
rect 28077 5216 28089 5219
rect 27948 5188 28089 5216
rect 27948 5176 27954 5188
rect 28077 5185 28089 5188
rect 28123 5185 28135 5219
rect 28077 5179 28135 5185
rect 28258 5176 28264 5228
rect 28316 5216 28322 5228
rect 29917 5219 29975 5225
rect 29917 5216 29929 5219
rect 28316 5188 29929 5216
rect 28316 5176 28322 5188
rect 29917 5185 29929 5188
rect 29963 5216 29975 5219
rect 30282 5216 30288 5228
rect 29963 5188 30288 5216
rect 29963 5185 29975 5188
rect 29917 5179 29975 5185
rect 30282 5176 30288 5188
rect 30340 5176 30346 5228
rect 31772 5225 31800 5256
rect 30469 5219 30527 5225
rect 30469 5185 30481 5219
rect 30515 5216 30527 5219
rect 31297 5219 31355 5225
rect 30515 5188 31248 5216
rect 30515 5185 30527 5188
rect 30469 5179 30527 5185
rect 30561 5151 30619 5157
rect 30561 5148 30573 5151
rect 27795 5120 30573 5148
rect 30561 5117 30573 5120
rect 30607 5117 30619 5151
rect 30561 5111 30619 5117
rect 24762 5080 24768 5092
rect 20272 5052 24072 5080
rect 24136 5052 24768 5080
rect 14884 4984 16620 5012
rect 14884 4972 14890 4984
rect 19886 4972 19892 5024
rect 19944 5012 19950 5024
rect 20272 5012 20300 5052
rect 19944 4984 20300 5012
rect 19944 4972 19950 4984
rect 20714 4972 20720 5024
rect 20772 4972 20778 5024
rect 21910 4972 21916 5024
rect 21968 4972 21974 5024
rect 22738 4972 22744 5024
rect 22796 5012 22802 5024
rect 24136 5012 24164 5052
rect 24762 5040 24768 5052
rect 24820 5080 24826 5092
rect 27890 5080 27896 5092
rect 24820 5052 27896 5080
rect 24820 5040 24826 5052
rect 27890 5040 27896 5052
rect 27948 5040 27954 5092
rect 22796 4984 24164 5012
rect 22796 4972 22802 4984
rect 24210 4972 24216 5024
rect 24268 4972 24274 5024
rect 27154 4972 27160 5024
rect 27212 4972 27218 5024
rect 27522 4972 27528 5024
rect 27580 5012 27586 5024
rect 27617 5015 27675 5021
rect 27617 5012 27629 5015
rect 27580 4984 27629 5012
rect 27580 4972 27586 4984
rect 27617 4981 27629 4984
rect 27663 4981 27675 5015
rect 27617 4975 27675 4981
rect 27798 4972 27804 5024
rect 27856 5012 27862 5024
rect 27985 5015 28043 5021
rect 27985 5012 27997 5015
rect 27856 4984 27997 5012
rect 27856 4972 27862 4984
rect 27985 4981 27997 4984
rect 28031 4981 28043 5015
rect 31220 5012 31248 5188
rect 31297 5185 31309 5219
rect 31343 5185 31355 5219
rect 31297 5179 31355 5185
rect 31757 5219 31815 5225
rect 31757 5185 31769 5219
rect 31803 5185 31815 5219
rect 31757 5179 31815 5185
rect 31312 5148 31340 5179
rect 32585 5151 32643 5157
rect 31312 5120 32168 5148
rect 31481 5083 31539 5089
rect 31481 5049 31493 5083
rect 31527 5080 31539 5083
rect 31754 5080 31760 5092
rect 31527 5052 31760 5080
rect 31527 5049 31539 5052
rect 31481 5043 31539 5049
rect 31754 5040 31760 5052
rect 31812 5040 31818 5092
rect 32140 5089 32168 5120
rect 32585 5117 32597 5151
rect 32631 5117 32643 5151
rect 32585 5111 32643 5117
rect 32125 5083 32183 5089
rect 32125 5049 32137 5083
rect 32171 5049 32183 5083
rect 32125 5043 32183 5049
rect 31570 5012 31576 5024
rect 31220 4984 31576 5012
rect 27985 4975 28043 4981
rect 31570 4972 31576 4984
rect 31628 5012 31634 5024
rect 32600 5012 32628 5111
rect 32674 5108 32680 5160
rect 32732 5108 32738 5160
rect 31628 4984 32628 5012
rect 31628 4972 31634 4984
rect 1104 4922 38272 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38272 4922
rect 1104 4848 38272 4870
rect 1581 4811 1639 4817
rect 1581 4777 1593 4811
rect 1627 4808 1639 4811
rect 6270 4808 6276 4820
rect 1627 4780 6276 4808
rect 1627 4777 1639 4780
rect 1581 4771 1639 4777
rect 6270 4768 6276 4780
rect 6328 4768 6334 4820
rect 9766 4768 9772 4820
rect 9824 4808 9830 4820
rect 19334 4808 19340 4820
rect 9824 4780 19340 4808
rect 9824 4768 9830 4780
rect 19334 4768 19340 4780
rect 19392 4768 19398 4820
rect 22830 4768 22836 4820
rect 22888 4768 22894 4820
rect 24210 4808 24216 4820
rect 23768 4780 24216 4808
rect 12618 4700 12624 4752
rect 12676 4700 12682 4752
rect 13078 4700 13084 4752
rect 13136 4740 13142 4752
rect 13357 4743 13415 4749
rect 13357 4740 13369 4743
rect 13136 4712 13369 4740
rect 13136 4700 13142 4712
rect 13357 4709 13369 4712
rect 13403 4709 13415 4743
rect 13357 4703 13415 4709
rect 14090 4700 14096 4752
rect 14148 4700 14154 4752
rect 15010 4700 15016 4752
rect 15068 4700 15074 4752
rect 15194 4700 15200 4752
rect 15252 4700 15258 4752
rect 17034 4700 17040 4752
rect 17092 4700 17098 4752
rect 8941 4607 8999 4613
rect 8941 4573 8953 4607
rect 8987 4604 8999 4607
rect 8987 4576 9076 4604
rect 8987 4573 8999 4576
rect 8941 4567 8999 4573
rect 934 4496 940 4548
rect 992 4536 998 4548
rect 1489 4539 1547 4545
rect 1489 4536 1501 4539
rect 992 4508 1501 4536
rect 992 4496 998 4508
rect 1489 4505 1501 4508
rect 1535 4505 1547 4539
rect 1489 4499 1547 4505
rect 9048 4480 9076 4576
rect 12636 4536 12664 4700
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4604 13599 4607
rect 14108 4604 14136 4700
rect 15212 4613 15240 4700
rect 13587 4576 14136 4604
rect 15197 4607 15255 4613
rect 13587 4573 13599 4576
rect 13541 4567 13599 4573
rect 15197 4573 15209 4607
rect 15243 4573 15255 4607
rect 15197 4567 15255 4573
rect 16945 4607 17003 4613
rect 16945 4573 16957 4607
rect 16991 4604 17003 4607
rect 17052 4604 17080 4700
rect 19886 4672 19892 4684
rect 16991 4576 17080 4604
rect 18156 4644 19892 4672
rect 16991 4573 17003 4576
rect 16945 4567 17003 4573
rect 18156 4536 18184 4644
rect 19886 4632 19892 4644
rect 19944 4632 19950 4684
rect 20901 4675 20959 4681
rect 20901 4641 20913 4675
rect 20947 4672 20959 4675
rect 21085 4675 21143 4681
rect 21085 4672 21097 4675
rect 20947 4644 21097 4672
rect 20947 4641 20959 4644
rect 20901 4635 20959 4641
rect 21085 4641 21097 4644
rect 21131 4641 21143 4675
rect 21085 4635 21143 4641
rect 23382 4632 23388 4684
rect 23440 4672 23446 4684
rect 23477 4675 23535 4681
rect 23477 4672 23489 4675
rect 23440 4644 23489 4672
rect 23440 4632 23446 4644
rect 23477 4641 23489 4644
rect 23523 4641 23535 4675
rect 23477 4635 23535 4641
rect 19426 4564 19432 4616
rect 19484 4564 19490 4616
rect 19797 4607 19855 4613
rect 19797 4573 19809 4607
rect 19843 4604 19855 4607
rect 20162 4604 20168 4616
rect 19843 4576 20168 4604
rect 19843 4573 19855 4576
rect 19797 4567 19855 4573
rect 20162 4564 20168 4576
rect 20220 4604 20226 4616
rect 20714 4604 20720 4616
rect 20220 4576 20720 4604
rect 20220 4564 20226 4576
rect 20714 4564 20720 4576
rect 20772 4564 20778 4616
rect 20993 4607 21051 4613
rect 20993 4573 21005 4607
rect 21039 4573 21051 4607
rect 20993 4567 21051 4573
rect 23293 4607 23351 4613
rect 23293 4573 23305 4607
rect 23339 4604 23351 4607
rect 23566 4604 23572 4616
rect 23339 4576 23572 4604
rect 23339 4573 23351 4576
rect 23293 4567 23351 4573
rect 12636 4508 18184 4536
rect 9030 4428 9036 4480
rect 9088 4428 9094 4480
rect 9122 4428 9128 4480
rect 9180 4428 9186 4480
rect 9950 4428 9956 4480
rect 10008 4468 10014 4480
rect 15838 4468 15844 4480
rect 10008 4440 15844 4468
rect 10008 4428 10014 4440
rect 15838 4428 15844 4440
rect 15896 4428 15902 4480
rect 16666 4428 16672 4480
rect 16724 4468 16730 4480
rect 16853 4471 16911 4477
rect 16853 4468 16865 4471
rect 16724 4440 16865 4468
rect 16724 4428 16730 4440
rect 16853 4437 16865 4440
rect 16899 4437 16911 4471
rect 16853 4431 16911 4437
rect 19337 4471 19395 4477
rect 19337 4437 19349 4471
rect 19383 4468 19395 4471
rect 19444 4468 19472 4564
rect 19383 4440 19472 4468
rect 19383 4437 19395 4440
rect 19337 4431 19395 4437
rect 19702 4428 19708 4480
rect 19760 4428 19766 4480
rect 21008 4468 21036 4567
rect 23566 4564 23572 4576
rect 23624 4564 23630 4616
rect 23768 4613 23796 4780
rect 24210 4768 24216 4780
rect 24268 4768 24274 4820
rect 24302 4768 24308 4820
rect 24360 4808 24366 4820
rect 26145 4811 26203 4817
rect 26145 4808 26157 4811
rect 24360 4780 26157 4808
rect 24360 4768 24366 4780
rect 26145 4777 26157 4780
rect 26191 4777 26203 4811
rect 26145 4771 26203 4777
rect 27157 4811 27215 4817
rect 27157 4777 27169 4811
rect 27203 4808 27215 4811
rect 27246 4808 27252 4820
rect 27203 4780 27252 4808
rect 27203 4777 27215 4780
rect 27157 4771 27215 4777
rect 27246 4768 27252 4780
rect 27304 4768 27310 4820
rect 27338 4768 27344 4820
rect 27396 4808 27402 4820
rect 27396 4780 31754 4808
rect 27396 4768 27402 4780
rect 23937 4743 23995 4749
rect 23937 4709 23949 4743
rect 23983 4740 23995 4743
rect 23983 4712 24532 4740
rect 23983 4709 23995 4712
rect 23937 4703 23995 4709
rect 24121 4675 24179 4681
rect 24121 4641 24133 4675
rect 24167 4672 24179 4675
rect 24397 4675 24455 4681
rect 24397 4672 24409 4675
rect 24167 4644 24409 4672
rect 24167 4641 24179 4644
rect 24121 4635 24179 4641
rect 24397 4641 24409 4644
rect 24443 4641 24455 4675
rect 24504 4672 24532 4712
rect 29086 4700 29092 4752
rect 29144 4740 29150 4752
rect 29181 4743 29239 4749
rect 29181 4740 29193 4743
rect 29144 4712 29193 4740
rect 29144 4700 29150 4712
rect 29181 4709 29193 4712
rect 29227 4709 29239 4743
rect 31726 4740 31754 4780
rect 32674 4740 32680 4752
rect 31726 4712 32680 4740
rect 29181 4703 29239 4709
rect 32674 4700 32680 4712
rect 32732 4700 32738 4752
rect 24673 4675 24731 4681
rect 24673 4672 24685 4675
rect 24504 4644 24685 4672
rect 24397 4635 24455 4641
rect 24673 4641 24685 4644
rect 24719 4641 24731 4675
rect 24673 4635 24731 4641
rect 26510 4632 26516 4684
rect 26568 4632 26574 4684
rect 26620 4644 28948 4672
rect 23753 4607 23811 4613
rect 23753 4573 23765 4607
rect 23799 4573 23811 4607
rect 23753 4567 23811 4573
rect 24213 4607 24271 4613
rect 24213 4573 24225 4607
rect 24259 4573 24271 4607
rect 24213 4567 24271 4573
rect 21358 4496 21364 4548
rect 21416 4496 21422 4548
rect 22646 4536 22652 4548
rect 22586 4508 22652 4536
rect 22646 4496 22652 4508
rect 22704 4496 22710 4548
rect 22738 4468 22744 4480
rect 21008 4440 22744 4468
rect 22738 4428 22744 4440
rect 22796 4428 22802 4480
rect 22922 4428 22928 4480
rect 22980 4428 22986 4480
rect 23290 4428 23296 4480
rect 23348 4468 23354 4480
rect 23385 4471 23443 4477
rect 23385 4468 23397 4471
rect 23348 4440 23397 4468
rect 23348 4428 23354 4440
rect 23385 4437 23397 4440
rect 23431 4437 23443 4471
rect 24228 4468 24256 4567
rect 25774 4564 25780 4616
rect 25832 4604 25838 4616
rect 26620 4604 26648 4644
rect 25832 4576 26648 4604
rect 26697 4607 26755 4613
rect 25832 4564 25838 4576
rect 26697 4573 26709 4607
rect 26743 4604 26755 4607
rect 27062 4604 27068 4616
rect 26743 4576 27068 4604
rect 26743 4573 26755 4576
rect 26697 4567 26755 4573
rect 27062 4564 27068 4576
rect 27120 4564 27126 4616
rect 27430 4564 27436 4616
rect 27488 4564 27494 4616
rect 27614 4536 27620 4548
rect 26068 4508 27620 4536
rect 26068 4468 26096 4508
rect 27614 4496 27620 4508
rect 27672 4496 27678 4548
rect 27709 4539 27767 4545
rect 27709 4505 27721 4539
rect 27755 4505 27767 4539
rect 28920 4536 28948 4644
rect 28920 4522 29500 4536
rect 28934 4508 29500 4522
rect 27709 4499 27767 4505
rect 24228 4440 26096 4468
rect 23385 4431 23443 4437
rect 26786 4428 26792 4480
rect 26844 4428 26850 4480
rect 27154 4428 27160 4480
rect 27212 4468 27218 4480
rect 27724 4468 27752 4499
rect 27212 4440 27752 4468
rect 27212 4428 27218 4440
rect 28534 4428 28540 4480
rect 28592 4468 28598 4480
rect 29012 4468 29040 4508
rect 29472 4480 29500 4508
rect 28592 4440 29040 4468
rect 28592 4428 28598 4440
rect 29454 4428 29460 4480
rect 29512 4428 29518 4480
rect 1104 4378 38272 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 38272 4378
rect 1104 4304 38272 4326
rect 11790 4224 11796 4276
rect 11848 4264 11854 4276
rect 12710 4264 12716 4276
rect 11848 4236 12716 4264
rect 11848 4224 11854 4236
rect 12710 4224 12716 4236
rect 12768 4264 12774 4276
rect 16206 4264 16212 4276
rect 12768 4236 16212 4264
rect 12768 4224 12774 4236
rect 16206 4224 16212 4236
rect 16264 4224 16270 4276
rect 21358 4224 21364 4276
rect 21416 4264 21422 4276
rect 21821 4267 21879 4273
rect 21821 4264 21833 4267
rect 21416 4236 21833 4264
rect 21416 4224 21422 4236
rect 21821 4233 21833 4236
rect 21867 4233 21879 4267
rect 21821 4227 21879 4233
rect 22186 4224 22192 4276
rect 22244 4264 22250 4276
rect 22646 4264 22652 4276
rect 22244 4236 22652 4264
rect 22244 4224 22250 4236
rect 22646 4224 22652 4236
rect 22704 4264 22710 4276
rect 23382 4264 23388 4276
rect 22704 4236 23388 4264
rect 22704 4224 22710 4236
rect 23382 4224 23388 4236
rect 23440 4264 23446 4276
rect 25774 4264 25780 4276
rect 23440 4236 25780 4264
rect 23440 4224 23446 4236
rect 25774 4224 25780 4236
rect 25832 4224 25838 4276
rect 26786 4224 26792 4276
rect 26844 4224 26850 4276
rect 26970 4224 26976 4276
rect 27028 4224 27034 4276
rect 27062 4224 27068 4276
rect 27120 4264 27126 4276
rect 29549 4267 29607 4273
rect 29549 4264 29561 4267
rect 27120 4236 29561 4264
rect 27120 4224 27126 4236
rect 29549 4233 29561 4236
rect 29595 4264 29607 4267
rect 29730 4264 29736 4276
rect 29595 4236 29736 4264
rect 29595 4233 29607 4236
rect 29549 4227 29607 4233
rect 29730 4224 29736 4236
rect 29788 4224 29794 4276
rect 11422 4156 11428 4208
rect 11480 4196 11486 4208
rect 13446 4196 13452 4208
rect 11480 4168 13452 4196
rect 11480 4156 11486 4168
rect 13446 4156 13452 4168
rect 13504 4196 13510 4208
rect 16114 4196 16120 4208
rect 13504 4168 16120 4196
rect 13504 4156 13510 4168
rect 16114 4156 16120 4168
rect 16172 4196 16178 4208
rect 16172 4168 17434 4196
rect 16172 4156 16178 4168
rect 20990 4156 20996 4208
rect 21048 4196 21054 4208
rect 25314 4196 25320 4208
rect 21048 4168 25320 4196
rect 21048 4156 21054 4168
rect 25314 4156 25320 4168
rect 25372 4156 25378 4208
rect 26804 4196 26832 4224
rect 27341 4199 27399 4205
rect 27341 4196 27353 4199
rect 26804 4168 27353 4196
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4128 12311 4131
rect 12342 4128 12348 4140
rect 12299 4100 12348 4128
rect 12299 4097 12311 4100
rect 12253 4091 12311 4097
rect 12342 4088 12348 4100
rect 12400 4128 12406 4140
rect 12529 4131 12587 4137
rect 12400 4088 12434 4128
rect 12529 4097 12541 4131
rect 12575 4128 12587 4131
rect 12802 4128 12808 4140
rect 12575 4100 12808 4128
rect 12575 4097 12587 4100
rect 12529 4091 12587 4097
rect 12802 4088 12808 4100
rect 12860 4088 12866 4140
rect 16298 4088 16304 4140
rect 16356 4088 16362 4140
rect 19334 4088 19340 4140
rect 19392 4128 19398 4140
rect 21542 4128 21548 4140
rect 19392 4100 21548 4128
rect 19392 4088 19398 4100
rect 21542 4088 21548 4100
rect 21600 4088 21606 4140
rect 21910 4088 21916 4140
rect 21968 4128 21974 4140
rect 22005 4131 22063 4137
rect 22005 4128 22017 4131
rect 21968 4100 22017 4128
rect 21968 4088 21974 4100
rect 22005 4097 22017 4100
rect 22051 4097 22063 4131
rect 22005 4091 22063 4097
rect 24762 4088 24768 4140
rect 24820 4128 24826 4140
rect 26804 4128 26832 4168
rect 27341 4165 27353 4168
rect 27387 4165 27399 4199
rect 29454 4196 29460 4208
rect 29302 4168 29460 4196
rect 27341 4159 27399 4165
rect 29454 4156 29460 4168
rect 29512 4196 29518 4208
rect 31018 4196 31024 4208
rect 29512 4168 31024 4196
rect 29512 4156 29518 4168
rect 31018 4156 31024 4168
rect 31076 4156 31082 4208
rect 24820 4100 26832 4128
rect 27433 4131 27491 4137
rect 24820 4088 24826 4100
rect 27433 4097 27445 4131
rect 27479 4128 27491 4131
rect 27479 4100 27660 4128
rect 27479 4097 27491 4100
rect 27433 4091 27491 4097
rect 12406 4060 12434 4088
rect 12406 4032 14688 4060
rect 11054 3952 11060 4004
rect 11112 3992 11118 4004
rect 11974 3992 11980 4004
rect 11112 3964 11980 3992
rect 11112 3952 11118 3964
rect 11974 3952 11980 3964
rect 12032 3992 12038 4004
rect 14550 3992 14556 4004
rect 12032 3964 14556 3992
rect 12032 3952 12038 3964
rect 14550 3952 14556 3964
rect 14608 3952 14614 4004
rect 14660 3936 14688 4032
rect 16666 4020 16672 4072
rect 16724 4020 16730 4072
rect 16945 4063 17003 4069
rect 16945 4060 16957 4063
rect 16776 4032 16957 4060
rect 16485 3995 16543 4001
rect 16485 3961 16497 3995
rect 16531 3992 16543 3995
rect 16776 3992 16804 4032
rect 16945 4029 16957 4032
rect 16991 4029 17003 4063
rect 16945 4023 17003 4029
rect 27525 4063 27583 4069
rect 27525 4029 27537 4063
rect 27571 4029 27583 4063
rect 27525 4023 27583 4029
rect 20346 3992 20352 4004
rect 16531 3964 16804 3992
rect 18432 3964 20352 3992
rect 16531 3961 16543 3964
rect 16485 3955 16543 3961
rect 12158 3884 12164 3936
rect 12216 3884 12222 3936
rect 12250 3884 12256 3936
rect 12308 3924 12314 3936
rect 12345 3927 12403 3933
rect 12345 3924 12357 3927
rect 12308 3896 12357 3924
rect 12308 3884 12314 3896
rect 12345 3893 12357 3896
rect 12391 3893 12403 3927
rect 12345 3887 12403 3893
rect 14642 3884 14648 3936
rect 14700 3884 14706 3936
rect 17494 3884 17500 3936
rect 17552 3924 17558 3936
rect 18432 3933 18460 3964
rect 20346 3952 20352 3964
rect 20404 3952 20410 4004
rect 18417 3927 18475 3933
rect 18417 3924 18429 3927
rect 17552 3896 18429 3924
rect 17552 3884 17558 3896
rect 18417 3893 18429 3896
rect 18463 3893 18475 3927
rect 18417 3887 18475 3893
rect 19794 3884 19800 3936
rect 19852 3924 19858 3936
rect 27540 3924 27568 4023
rect 19852 3896 27568 3924
rect 27632 3924 27660 4100
rect 27798 4020 27804 4072
rect 27856 4020 27862 4072
rect 28074 4020 28080 4072
rect 28132 4020 28138 4072
rect 29086 3924 29092 3936
rect 27632 3896 29092 3924
rect 19852 3884 19858 3896
rect 29086 3884 29092 3896
rect 29144 3884 29150 3936
rect 1104 3834 38272 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38272 3834
rect 1104 3760 38272 3782
rect 7101 3723 7159 3729
rect 7101 3689 7113 3723
rect 7147 3720 7159 3723
rect 9766 3720 9772 3732
rect 7147 3692 9772 3720
rect 7147 3689 7159 3692
rect 7101 3683 7159 3689
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 12158 3720 12164 3732
rect 11900 3692 12164 3720
rect 11900 3593 11928 3692
rect 12158 3680 12164 3692
rect 12216 3680 12222 3732
rect 14550 3680 14556 3732
rect 14608 3720 14614 3732
rect 14608 3692 16252 3720
rect 14608 3680 14614 3692
rect 15197 3655 15255 3661
rect 15197 3621 15209 3655
rect 15243 3621 15255 3655
rect 15197 3615 15255 3621
rect 11885 3587 11943 3593
rect 11885 3553 11897 3587
rect 11931 3553 11943 3587
rect 11885 3547 11943 3553
rect 12161 3587 12219 3593
rect 12161 3553 12173 3587
rect 12207 3584 12219 3587
rect 12250 3584 12256 3596
rect 12207 3556 12256 3584
rect 12207 3553 12219 3556
rect 12161 3547 12219 3553
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 14366 3544 14372 3596
rect 14424 3584 14430 3596
rect 14461 3587 14519 3593
rect 14461 3584 14473 3587
rect 14424 3556 14473 3584
rect 14424 3544 14430 3556
rect 14461 3553 14473 3556
rect 14507 3553 14519 3587
rect 14461 3547 14519 3553
rect 6914 3476 6920 3528
rect 6972 3476 6978 3528
rect 9030 3476 9036 3528
rect 9088 3476 9094 3528
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3516 9183 3519
rect 9309 3519 9367 3525
rect 9309 3516 9321 3519
rect 9171 3488 9321 3516
rect 9171 3485 9183 3488
rect 9125 3479 9183 3485
rect 9309 3485 9321 3488
rect 9355 3485 9367 3519
rect 11422 3516 11428 3528
rect 10718 3488 11428 3516
rect 9309 3479 9367 3485
rect 11422 3476 11428 3488
rect 11480 3476 11486 3528
rect 11606 3476 11612 3528
rect 11664 3476 11670 3528
rect 11698 3476 11704 3528
rect 11756 3476 11762 3528
rect 13446 3516 13452 3528
rect 13294 3488 13452 3516
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 14274 3476 14280 3528
rect 14332 3476 14338 3528
rect 14642 3476 14648 3528
rect 14700 3476 14706 3528
rect 15105 3519 15163 3525
rect 15105 3485 15117 3519
rect 15151 3516 15163 3519
rect 15212 3516 15240 3615
rect 15838 3544 15844 3596
rect 15896 3544 15902 3596
rect 16224 3584 16252 3692
rect 16298 3680 16304 3732
rect 16356 3720 16362 3732
rect 17129 3723 17187 3729
rect 17129 3720 17141 3723
rect 16356 3692 17141 3720
rect 16356 3680 16362 3692
rect 17129 3689 17141 3692
rect 17175 3689 17187 3723
rect 17129 3683 17187 3689
rect 17696 3692 26096 3720
rect 17696 3593 17724 3692
rect 17954 3612 17960 3664
rect 18012 3612 18018 3664
rect 18233 3655 18291 3661
rect 18233 3652 18245 3655
rect 18156 3624 18245 3652
rect 17681 3587 17739 3593
rect 17681 3584 17693 3587
rect 16224 3556 17693 3584
rect 17681 3553 17693 3556
rect 17727 3553 17739 3587
rect 17681 3547 17739 3553
rect 18156 3525 18184 3624
rect 18233 3621 18245 3624
rect 18279 3621 18291 3655
rect 18233 3615 18291 3621
rect 20441 3655 20499 3661
rect 20441 3621 20453 3655
rect 20487 3652 20499 3655
rect 20487 3624 20760 3652
rect 20487 3621 20499 3624
rect 20441 3615 20499 3621
rect 18782 3544 18788 3596
rect 18840 3544 18846 3596
rect 19794 3544 19800 3596
rect 19852 3544 19858 3596
rect 16853 3519 16911 3525
rect 16853 3516 16865 3519
rect 15151 3488 15240 3516
rect 15304 3488 16865 3516
rect 15151 3485 15163 3488
rect 15105 3479 15163 3485
rect 9048 3448 9076 3476
rect 9490 3448 9496 3460
rect 9048 3420 9496 3448
rect 9490 3408 9496 3420
rect 9548 3408 9554 3460
rect 9582 3408 9588 3460
rect 9640 3408 9646 3460
rect 11238 3408 11244 3460
rect 11296 3448 11302 3460
rect 11333 3451 11391 3457
rect 11333 3448 11345 3451
rect 11296 3420 11345 3448
rect 11296 3408 11302 3420
rect 11333 3417 11345 3420
rect 11379 3448 11391 3451
rect 11379 3420 12388 3448
rect 11379 3417 11391 3420
rect 11333 3411 11391 3417
rect 12360 3392 12388 3420
rect 13906 3408 13912 3460
rect 13964 3408 13970 3460
rect 15304 3448 15332 3488
rect 16853 3485 16865 3488
rect 16899 3516 16911 3519
rect 18141 3519 18199 3525
rect 16899 3488 16988 3516
rect 16899 3485 16911 3488
rect 16853 3479 16911 3485
rect 14660 3420 15332 3448
rect 16960 3448 16988 3488
rect 18141 3485 18153 3519
rect 18187 3485 18199 3519
rect 18141 3479 18199 3485
rect 18598 3476 18604 3528
rect 18656 3476 18662 3528
rect 18874 3476 18880 3528
rect 18932 3516 18938 3528
rect 19812 3516 19840 3544
rect 18932 3488 19840 3516
rect 19981 3519 20039 3525
rect 18932 3476 18938 3488
rect 19981 3485 19993 3519
rect 20027 3516 20039 3519
rect 20622 3516 20628 3528
rect 20027 3488 20628 3516
rect 20027 3485 20039 3488
rect 19981 3479 20039 3485
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 20732 3525 20760 3624
rect 22296 3556 24072 3584
rect 20717 3519 20775 3525
rect 20717 3485 20729 3519
rect 20763 3485 20775 3519
rect 20717 3479 20775 3485
rect 20993 3519 21051 3525
rect 20993 3485 21005 3519
rect 21039 3516 21051 3519
rect 22097 3519 22155 3525
rect 22097 3516 22109 3519
rect 21039 3488 22109 3516
rect 21039 3485 21051 3488
rect 20993 3479 21051 3485
rect 22097 3485 22109 3488
rect 22143 3516 22155 3519
rect 22296 3516 22324 3556
rect 22143 3488 22324 3516
rect 22373 3519 22431 3525
rect 22143 3485 22155 3488
rect 22097 3479 22155 3485
rect 22373 3485 22385 3519
rect 22419 3516 22431 3519
rect 22922 3516 22928 3528
rect 22419 3488 22928 3516
rect 22419 3485 22431 3488
rect 22373 3479 22431 3485
rect 22922 3476 22928 3488
rect 22980 3476 22986 3528
rect 23937 3519 23995 3525
rect 23937 3485 23949 3519
rect 23983 3485 23995 3519
rect 23937 3479 23995 3485
rect 23952 3448 23980 3479
rect 16960 3420 23980 3448
rect 24044 3448 24072 3556
rect 24578 3544 24584 3596
rect 24636 3544 24642 3596
rect 24762 3544 24768 3596
rect 24820 3544 24826 3596
rect 25222 3544 25228 3596
rect 25280 3544 25286 3596
rect 25314 3544 25320 3596
rect 25372 3544 25378 3596
rect 26068 3593 26096 3692
rect 29362 3680 29368 3732
rect 29420 3720 29426 3732
rect 37645 3723 37703 3729
rect 37645 3720 37657 3723
rect 29420 3692 37657 3720
rect 29420 3680 29426 3692
rect 37645 3689 37657 3692
rect 37691 3689 37703 3723
rect 37645 3683 37703 3689
rect 26326 3612 26332 3664
rect 26384 3652 26390 3664
rect 26384 3624 31248 3652
rect 26384 3612 26390 3624
rect 31220 3596 31248 3624
rect 26053 3587 26111 3593
rect 26053 3553 26065 3587
rect 26099 3553 26111 3587
rect 26053 3547 26111 3553
rect 26237 3587 26295 3593
rect 26237 3553 26249 3587
rect 26283 3584 26295 3587
rect 26786 3584 26792 3596
rect 26283 3556 26792 3584
rect 26283 3553 26295 3556
rect 26237 3547 26295 3553
rect 26786 3544 26792 3556
rect 26844 3544 26850 3596
rect 27172 3556 28396 3584
rect 25240 3516 25268 3544
rect 25501 3519 25559 3525
rect 25501 3516 25513 3519
rect 25240 3488 25513 3516
rect 25501 3485 25513 3488
rect 25547 3516 25559 3519
rect 27172 3516 27200 3556
rect 25547 3488 27200 3516
rect 27249 3519 27307 3525
rect 25547 3485 25559 3488
rect 25501 3479 25559 3485
rect 27249 3485 27261 3519
rect 27295 3485 27307 3519
rect 27249 3479 27307 3485
rect 24670 3448 24676 3460
rect 24044 3420 24676 3448
rect 14660 3392 14688 3420
rect 24670 3408 24676 3420
rect 24728 3448 24734 3460
rect 27264 3448 27292 3479
rect 27706 3476 27712 3528
rect 27764 3516 27770 3528
rect 28169 3519 28227 3525
rect 28169 3516 28181 3519
rect 27764 3488 28181 3516
rect 27764 3476 27770 3488
rect 28169 3485 28181 3488
rect 28215 3485 28227 3519
rect 28169 3479 28227 3485
rect 28258 3476 28264 3528
rect 28316 3476 28322 3528
rect 28368 3525 28396 3556
rect 31202 3544 31208 3596
rect 31260 3544 31266 3596
rect 28353 3519 28411 3525
rect 28353 3485 28365 3519
rect 28399 3485 28411 3519
rect 28353 3479 28411 3485
rect 37458 3476 37464 3528
rect 37516 3476 37522 3528
rect 28276 3448 28304 3476
rect 24728 3420 28304 3448
rect 24728 3408 24734 3420
rect 9214 3340 9220 3392
rect 9272 3380 9278 3392
rect 11425 3383 11483 3389
rect 11425 3380 11437 3383
rect 9272 3352 11437 3380
rect 9272 3340 9278 3352
rect 11425 3349 11437 3352
rect 11471 3349 11483 3383
rect 11425 3343 11483 3349
rect 12342 3340 12348 3392
rect 12400 3340 12406 3392
rect 12434 3340 12440 3392
rect 12492 3380 12498 3392
rect 14093 3383 14151 3389
rect 14093 3380 14105 3383
rect 12492 3352 14105 3380
rect 12492 3340 12498 3352
rect 14093 3349 14105 3352
rect 14139 3349 14151 3383
rect 14093 3343 14151 3349
rect 14642 3340 14648 3392
rect 14700 3340 14706 3392
rect 14734 3340 14740 3392
rect 14792 3340 14798 3392
rect 14918 3340 14924 3392
rect 14976 3340 14982 3392
rect 15562 3340 15568 3392
rect 15620 3340 15626 3392
rect 15657 3383 15715 3389
rect 15657 3349 15669 3383
rect 15703 3380 15715 3383
rect 16298 3380 16304 3392
rect 15703 3352 16304 3380
rect 15703 3349 15715 3352
rect 15657 3343 15715 3349
rect 16298 3340 16304 3352
rect 16356 3340 16362 3392
rect 16942 3340 16948 3392
rect 17000 3340 17006 3392
rect 17494 3340 17500 3392
rect 17552 3340 17558 3392
rect 17586 3340 17592 3392
rect 17644 3380 17650 3392
rect 18693 3383 18751 3389
rect 18693 3380 18705 3383
rect 17644 3352 18705 3380
rect 17644 3340 17650 3352
rect 18693 3349 18705 3352
rect 18739 3380 18751 3383
rect 19702 3380 19708 3392
rect 18739 3352 19708 3380
rect 18739 3349 18751 3352
rect 18693 3343 18751 3349
rect 19702 3340 19708 3352
rect 19760 3380 19766 3392
rect 20073 3383 20131 3389
rect 20073 3380 20085 3383
rect 19760 3352 20085 3380
rect 19760 3340 19766 3352
rect 20073 3349 20085 3352
rect 20119 3349 20131 3383
rect 20073 3343 20131 3349
rect 20346 3340 20352 3392
rect 20404 3380 20410 3392
rect 20533 3383 20591 3389
rect 20533 3380 20545 3383
rect 20404 3352 20545 3380
rect 20404 3340 20410 3352
rect 20533 3349 20545 3352
rect 20579 3349 20591 3383
rect 20533 3343 20591 3349
rect 20898 3340 20904 3392
rect 20956 3340 20962 3392
rect 22002 3340 22008 3392
rect 22060 3340 22066 3392
rect 22186 3340 22192 3392
rect 22244 3340 22250 3392
rect 24026 3340 24032 3392
rect 24084 3340 24090 3392
rect 24854 3340 24860 3392
rect 24912 3340 24918 3392
rect 25222 3340 25228 3392
rect 25280 3340 25286 3392
rect 25682 3340 25688 3392
rect 25740 3340 25746 3392
rect 26329 3383 26387 3389
rect 26329 3349 26341 3383
rect 26375 3380 26387 3383
rect 26510 3380 26516 3392
rect 26375 3352 26516 3380
rect 26375 3349 26387 3352
rect 26329 3343 26387 3349
rect 26510 3340 26516 3352
rect 26568 3340 26574 3392
rect 26694 3340 26700 3392
rect 26752 3340 26758 3392
rect 27154 3340 27160 3392
rect 27212 3340 27218 3392
rect 28537 3383 28595 3389
rect 28537 3349 28549 3383
rect 28583 3380 28595 3383
rect 36906 3380 36912 3392
rect 28583 3352 36912 3380
rect 28583 3349 28595 3352
rect 28537 3343 28595 3349
rect 36906 3340 36912 3352
rect 36964 3340 36970 3392
rect 1104 3290 38272 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 38272 3290
rect 1104 3216 38272 3238
rect 9214 3136 9220 3188
rect 9272 3136 9278 3188
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 14642 3176 14648 3188
rect 9548 3148 14648 3176
rect 9548 3136 9554 3148
rect 1762 3068 1768 3120
rect 1820 3068 1826 3120
rect 2133 3043 2191 3049
rect 2133 3009 2145 3043
rect 2179 3040 2191 3043
rect 7009 3043 7067 3049
rect 2179 3012 2774 3040
rect 2179 3009 2191 3012
rect 2133 3003 2191 3009
rect 2746 2972 2774 3012
rect 7009 3009 7021 3043
rect 7055 3040 7067 3043
rect 9232 3040 9260 3136
rect 9582 3068 9588 3120
rect 9640 3068 9646 3120
rect 12434 3108 12440 3120
rect 9968 3080 12440 3108
rect 7055 3012 9260 3040
rect 7055 3009 7067 3012
rect 7009 3003 7067 3009
rect 2746 2944 7052 2972
rect 1486 2796 1492 2848
rect 1544 2796 1550 2848
rect 1946 2796 1952 2848
rect 2004 2796 2010 2848
rect 6825 2839 6883 2845
rect 6825 2805 6837 2839
rect 6871 2836 6883 2839
rect 6914 2836 6920 2848
rect 6871 2808 6920 2836
rect 6871 2805 6883 2808
rect 6825 2799 6883 2805
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 7024 2836 7052 2944
rect 9600 2904 9628 3068
rect 9861 2907 9919 2913
rect 9861 2904 9873 2907
rect 9600 2876 9873 2904
rect 9861 2873 9873 2876
rect 9907 2873 9919 2907
rect 9861 2867 9919 2873
rect 9968 2836 9996 3080
rect 12434 3068 12440 3080
rect 12492 3068 12498 3120
rect 12728 3117 12756 3148
rect 14642 3136 14648 3148
rect 14700 3136 14706 3188
rect 14734 3136 14740 3188
rect 14792 3136 14798 3188
rect 14918 3176 14924 3188
rect 14844 3148 14924 3176
rect 12713 3111 12771 3117
rect 12713 3077 12725 3111
rect 12759 3077 12771 3111
rect 12713 3071 12771 3077
rect 14458 3068 14464 3120
rect 14516 3068 14522 3120
rect 14752 3108 14780 3136
rect 14844 3117 14872 3148
rect 14918 3136 14924 3148
rect 14976 3136 14982 3188
rect 16942 3136 16948 3188
rect 17000 3136 17006 3188
rect 17954 3176 17960 3188
rect 17604 3148 17960 3176
rect 14568 3080 14780 3108
rect 14829 3111 14887 3117
rect 10045 3043 10103 3049
rect 10045 3009 10057 3043
rect 10091 3040 10103 3043
rect 10781 3043 10839 3049
rect 10091 3012 10456 3040
rect 10091 3009 10103 3012
rect 10045 3003 10103 3009
rect 10428 2913 10456 3012
rect 10781 3009 10793 3043
rect 10827 3009 10839 3043
rect 10781 3003 10839 3009
rect 10873 3043 10931 3049
rect 10873 3009 10885 3043
rect 10919 3040 10931 3043
rect 10919 3012 11468 3040
rect 10919 3009 10931 3012
rect 10873 3003 10931 3009
rect 10796 2972 10824 3003
rect 10796 2944 10916 2972
rect 10413 2907 10471 2913
rect 10413 2873 10425 2907
rect 10459 2873 10471 2907
rect 10888 2904 10916 2944
rect 10962 2932 10968 2984
rect 11020 2932 11026 2984
rect 11238 2932 11244 2984
rect 11296 2932 11302 2984
rect 11440 2972 11468 3012
rect 11514 3000 11520 3052
rect 11572 3000 11578 3052
rect 11606 3000 11612 3052
rect 11664 3000 11670 3052
rect 11790 3000 11796 3052
rect 11848 3000 11854 3052
rect 11882 3000 11888 3052
rect 11940 3040 11946 3052
rect 12161 3043 12219 3049
rect 12161 3040 12173 3043
rect 11940 3012 12173 3040
rect 11940 3000 11946 3012
rect 12161 3009 12173 3012
rect 12207 3009 12219 3043
rect 12161 3003 12219 3009
rect 12253 3043 12311 3049
rect 12253 3009 12265 3043
rect 12299 3040 12311 3043
rect 13906 3040 13912 3052
rect 12299 3012 13912 3040
rect 12299 3009 12311 3012
rect 12253 3003 12311 3009
rect 11900 2972 11928 3000
rect 11440 2944 11928 2972
rect 11974 2932 11980 2984
rect 12032 2932 12038 2984
rect 12176 2972 12204 3003
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 14568 3049 14596 3080
rect 14829 3077 14841 3111
rect 14875 3077 14887 3111
rect 16114 3108 16120 3120
rect 16054 3080 16120 3108
rect 14829 3071 14887 3077
rect 16114 3068 16120 3080
rect 16172 3068 16178 3120
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3009 14611 3043
rect 16960 3040 16988 3136
rect 17604 3117 17632 3148
rect 17954 3136 17960 3148
rect 18012 3136 18018 3188
rect 18230 3136 18236 3188
rect 18288 3176 18294 3188
rect 19518 3176 19524 3188
rect 18288 3148 19524 3176
rect 18288 3136 18294 3148
rect 19518 3136 19524 3148
rect 19576 3136 19582 3188
rect 20898 3176 20904 3188
rect 19812 3148 20904 3176
rect 17589 3111 17647 3117
rect 17589 3077 17601 3111
rect 17635 3077 17647 3111
rect 17589 3071 17647 3077
rect 17678 3068 17684 3120
rect 17736 3108 17742 3120
rect 17736 3080 18078 3108
rect 17736 3068 17742 3080
rect 19812 3049 19840 3148
rect 20898 3136 20904 3148
rect 20956 3136 20962 3188
rect 22002 3136 22008 3188
rect 22060 3136 22066 3188
rect 22186 3136 22192 3188
rect 22244 3136 22250 3188
rect 23566 3136 23572 3188
rect 23624 3136 23630 3188
rect 24026 3136 24032 3188
rect 24084 3136 24090 3188
rect 24854 3136 24860 3188
rect 24912 3176 24918 3188
rect 27338 3176 27344 3188
rect 24912 3148 27344 3176
rect 24912 3136 24918 3148
rect 20073 3111 20131 3117
rect 20073 3077 20085 3111
rect 20119 3108 20131 3111
rect 20346 3108 20352 3120
rect 20119 3080 20352 3108
rect 20119 3077 20131 3080
rect 20073 3071 20131 3077
rect 20346 3068 20352 3080
rect 20404 3068 20410 3120
rect 22020 3108 22048 3136
rect 21836 3080 22048 3108
rect 22097 3111 22155 3117
rect 21836 3049 21864 3080
rect 22097 3077 22109 3111
rect 22143 3108 22155 3111
rect 22204 3108 22232 3136
rect 23382 3108 23388 3120
rect 22143 3080 22232 3108
rect 23322 3094 23388 3108
rect 23308 3080 23388 3094
rect 22143 3077 22155 3080
rect 22097 3071 22155 3077
rect 17313 3043 17371 3049
rect 17313 3040 17325 3043
rect 16960 3012 17325 3040
rect 14553 3003 14611 3009
rect 17313 3009 17325 3012
rect 17359 3009 17371 3043
rect 17313 3003 17371 3009
rect 19541 3043 19599 3049
rect 19541 3009 19553 3043
rect 19587 3040 19599 3043
rect 19797 3043 19855 3049
rect 19587 3012 19748 3040
rect 19587 3009 19599 3012
rect 19541 3003 19599 3009
rect 15562 2972 15568 2984
rect 12176 2944 15568 2972
rect 15562 2932 15568 2944
rect 15620 2932 15626 2984
rect 18230 2972 18236 2984
rect 16224 2944 18236 2972
rect 11256 2904 11284 2932
rect 10888 2876 11284 2904
rect 12621 2907 12679 2913
rect 10413 2867 10471 2873
rect 12621 2873 12633 2907
rect 12667 2904 12679 2907
rect 12802 2904 12808 2916
rect 12667 2876 12808 2904
rect 12667 2873 12679 2876
rect 12621 2867 12679 2873
rect 12802 2864 12808 2876
rect 12860 2864 12866 2916
rect 13906 2864 13912 2916
rect 13964 2864 13970 2916
rect 7024 2808 9996 2836
rect 11701 2839 11759 2845
rect 11701 2805 11713 2839
rect 11747 2836 11759 2839
rect 12526 2836 12532 2848
rect 11747 2808 12532 2836
rect 11747 2805 11759 2808
rect 11701 2799 11759 2805
rect 12526 2796 12532 2808
rect 12584 2796 12590 2848
rect 13924 2836 13952 2864
rect 16224 2836 16252 2944
rect 18230 2932 18236 2944
rect 18288 2932 18294 2984
rect 18598 2932 18604 2984
rect 18656 2972 18662 2984
rect 19061 2975 19119 2981
rect 19061 2972 19073 2975
rect 18656 2944 19073 2972
rect 18656 2932 18662 2944
rect 19061 2941 19073 2944
rect 19107 2972 19119 2975
rect 19334 2972 19340 2984
rect 19107 2944 19340 2972
rect 19107 2941 19119 2944
rect 19061 2935 19119 2941
rect 19334 2932 19340 2944
rect 19392 2932 19398 2984
rect 19720 2972 19748 3012
rect 19797 3009 19809 3043
rect 19843 3009 19855 3043
rect 21821 3043 21879 3049
rect 19797 3003 19855 3009
rect 19720 2944 19840 2972
rect 18690 2864 18696 2916
rect 18748 2864 18754 2916
rect 13924 2808 16252 2836
rect 16298 2796 16304 2848
rect 16356 2836 16362 2848
rect 18708 2836 18736 2864
rect 19812 2848 19840 2944
rect 20622 2932 20628 2984
rect 20680 2972 20686 2984
rect 21192 2972 21220 3026
rect 21821 3009 21833 3043
rect 21867 3009 21879 3043
rect 21821 3003 21879 3009
rect 23308 2972 23336 3080
rect 23382 3068 23388 3080
rect 23440 3068 23446 3120
rect 24044 3108 24072 3136
rect 25884 3117 25912 3148
rect 27338 3136 27344 3148
rect 27396 3176 27402 3188
rect 31849 3179 31907 3185
rect 27396 3148 30880 3176
rect 27396 3136 27402 3148
rect 23860 3080 24072 3108
rect 25869 3111 25927 3117
rect 23860 3049 23888 3080
rect 25869 3077 25881 3111
rect 25915 3077 25927 3111
rect 27154 3108 27160 3120
rect 25869 3071 25927 3077
rect 26988 3080 27160 3108
rect 23845 3043 23903 3049
rect 23845 3009 23857 3043
rect 23891 3009 23903 3043
rect 23845 3003 23903 3009
rect 20680 2944 21128 2972
rect 21192 2944 23336 2972
rect 24121 2975 24179 2981
rect 20680 2932 20686 2944
rect 21100 2904 21128 2944
rect 24121 2941 24133 2975
rect 24167 2972 24179 2975
rect 25130 2972 25136 2984
rect 24167 2944 25136 2972
rect 24167 2941 24179 2944
rect 24121 2935 24179 2941
rect 25130 2932 25136 2944
rect 25188 2932 25194 2984
rect 25240 2972 25268 3026
rect 25682 3000 25688 3052
rect 25740 3040 25746 3052
rect 25961 3043 26019 3049
rect 25961 3040 25973 3043
rect 25740 3012 25973 3040
rect 25740 3000 25746 3012
rect 25961 3009 25973 3012
rect 26007 3009 26019 3043
rect 25961 3003 26019 3009
rect 26421 3043 26479 3049
rect 26421 3009 26433 3043
rect 26467 3040 26479 3043
rect 26694 3040 26700 3052
rect 26467 3012 26700 3040
rect 26467 3009 26479 3012
rect 26421 3003 26479 3009
rect 26694 3000 26700 3012
rect 26752 3000 26758 3052
rect 26988 3049 27016 3080
rect 27154 3068 27160 3080
rect 27212 3068 27218 3120
rect 28534 3108 28540 3120
rect 28474 3080 28540 3108
rect 28534 3068 28540 3080
rect 28592 3068 28598 3120
rect 30852 3049 30880 3148
rect 31849 3145 31861 3179
rect 31895 3145 31907 3179
rect 31849 3139 31907 3145
rect 31864 3108 31892 3139
rect 37553 3111 37611 3117
rect 37553 3108 37565 3111
rect 31864 3080 37565 3108
rect 37553 3077 37565 3080
rect 37599 3077 37611 3111
rect 37553 3071 37611 3077
rect 26973 3043 27031 3049
rect 26973 3009 26985 3043
rect 27019 3009 27031 3043
rect 26973 3003 27031 3009
rect 30837 3043 30895 3049
rect 30837 3009 30849 3043
rect 30883 3009 30895 3043
rect 30837 3003 30895 3009
rect 31018 3000 31024 3052
rect 31076 3040 31082 3052
rect 31205 3043 31263 3049
rect 31076 3012 31156 3040
rect 31076 3000 31082 3012
rect 25774 2972 25780 2984
rect 25240 2944 25780 2972
rect 25774 2932 25780 2944
rect 25832 2932 25838 2984
rect 27249 2975 27307 2981
rect 27249 2972 27261 2975
rect 26620 2944 27261 2972
rect 21545 2907 21603 2913
rect 21545 2904 21557 2907
rect 21100 2876 21557 2904
rect 21545 2873 21557 2876
rect 21591 2873 21603 2907
rect 26326 2904 26332 2916
rect 21545 2867 21603 2873
rect 25148 2876 26332 2904
rect 16356 2808 18736 2836
rect 16356 2796 16362 2808
rect 19702 2796 19708 2848
rect 19760 2796 19766 2848
rect 19794 2796 19800 2848
rect 19852 2836 19858 2848
rect 25148 2836 25176 2876
rect 26326 2864 26332 2876
rect 26384 2864 26390 2916
rect 26510 2864 26516 2916
rect 26568 2864 26574 2916
rect 26620 2913 26648 2944
rect 27249 2941 27261 2944
rect 27295 2941 27307 2975
rect 31128 2972 31156 3012
rect 31205 3009 31217 3043
rect 31251 3040 31263 3043
rect 31665 3043 31723 3049
rect 31665 3040 31677 3043
rect 31251 3012 31677 3040
rect 31251 3009 31263 3012
rect 31205 3003 31263 3009
rect 31665 3009 31677 3012
rect 31711 3009 31723 3043
rect 31665 3003 31723 3009
rect 32122 3000 32128 3052
rect 32180 3000 32186 3052
rect 36906 3000 36912 3052
rect 36964 3000 36970 3052
rect 32140 2972 32168 3000
rect 31128 2944 32168 2972
rect 27249 2935 27307 2941
rect 26605 2907 26663 2913
rect 26605 2873 26617 2907
rect 26651 2873 26663 2907
rect 26605 2867 26663 2873
rect 19852 2808 25176 2836
rect 26145 2839 26203 2845
rect 19852 2796 19858 2808
rect 26145 2805 26157 2839
rect 26191 2836 26203 2839
rect 26418 2836 26424 2848
rect 26191 2808 26424 2836
rect 26191 2805 26203 2808
rect 26145 2799 26203 2805
rect 26418 2796 26424 2808
rect 26476 2796 26482 2848
rect 26528 2836 26556 2864
rect 28721 2839 28779 2845
rect 28721 2836 28733 2839
rect 26528 2808 28733 2836
rect 28721 2805 28733 2808
rect 28767 2805 28779 2839
rect 28721 2799 28779 2805
rect 37093 2839 37151 2845
rect 37093 2805 37105 2839
rect 37139 2836 37151 2839
rect 37274 2836 37280 2848
rect 37139 2808 37280 2836
rect 37139 2805 37151 2808
rect 37093 2799 37151 2805
rect 37274 2796 37280 2808
rect 37332 2796 37338 2848
rect 37826 2796 37832 2848
rect 37884 2796 37890 2848
rect 1104 2746 38272 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38272 2746
rect 1104 2672 38272 2694
rect 9122 2632 9128 2644
rect 2424 2604 9128 2632
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2428 1823 2431
rect 1946 2428 1952 2440
rect 1811 2400 1952 2428
rect 1811 2397 1823 2400
rect 1765 2391 1823 2397
rect 1946 2388 1952 2400
rect 2004 2388 2010 2440
rect 2424 2437 2452 2604
rect 9122 2592 9128 2604
rect 9180 2592 9186 2644
rect 11606 2592 11612 2644
rect 11664 2632 11670 2644
rect 13219 2635 13277 2641
rect 13219 2632 13231 2635
rect 11664 2604 13231 2632
rect 11664 2592 11670 2604
rect 13219 2601 13231 2604
rect 13265 2601 13277 2635
rect 19794 2632 19800 2644
rect 13219 2595 13277 2601
rect 15125 2604 19800 2632
rect 11514 2524 11520 2576
rect 11572 2564 11578 2576
rect 15125 2564 15153 2604
rect 19794 2592 19800 2604
rect 19852 2592 19858 2644
rect 25130 2592 25136 2644
rect 25188 2592 25194 2644
rect 31018 2564 31024 2576
rect 11572 2536 15153 2564
rect 11572 2524 11578 2536
rect 8938 2496 8944 2508
rect 4356 2468 8944 2496
rect 4356 2437 4384 2468
rect 8938 2456 8944 2468
rect 8996 2456 9002 2508
rect 2409 2431 2467 2437
rect 2409 2397 2421 2431
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2397 4399 2431
rect 4341 2391 4399 2397
rect 6914 2388 6920 2440
rect 6972 2388 6978 2440
rect 12268 2437 12296 2536
rect 12618 2456 12624 2508
rect 12676 2456 12682 2508
rect 13354 2456 13360 2508
rect 13412 2456 13418 2508
rect 14366 2456 14372 2508
rect 14424 2456 14430 2508
rect 10873 2431 10931 2437
rect 10873 2397 10885 2431
rect 10919 2428 10931 2431
rect 12069 2431 12127 2437
rect 12069 2428 12081 2431
rect 10919 2400 12081 2428
rect 10919 2397 10931 2400
rect 10873 2391 10931 2397
rect 12069 2397 12081 2400
rect 12115 2397 12127 2431
rect 12069 2391 12127 2397
rect 12253 2431 12311 2437
rect 12253 2397 12265 2431
rect 12299 2397 12311 2431
rect 12253 2391 12311 2397
rect 12434 2388 12440 2440
rect 12492 2388 12498 2440
rect 12526 2388 12532 2440
rect 12584 2388 12590 2440
rect 12986 2388 12992 2440
rect 13044 2388 13050 2440
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 72 2332 1409 2360
rect 72 2320 78 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 2038 2320 2044 2372
rect 2096 2320 2102 2372
rect 3970 2320 3976 2372
rect 4028 2320 4034 2372
rect 6546 2320 6552 2372
rect 6604 2320 6610 2372
rect 11609 2363 11667 2369
rect 11609 2360 11621 2363
rect 11072 2332 11621 2360
rect 11072 2301 11100 2332
rect 11609 2329 11621 2332
rect 11655 2329 11667 2363
rect 12452 2360 12480 2388
rect 13372 2360 13400 2456
rect 15125 2437 15153 2536
rect 16132 2536 31024 2564
rect 16132 2505 16160 2536
rect 31018 2524 31024 2536
rect 31076 2524 31082 2576
rect 16117 2499 16175 2505
rect 16117 2496 16129 2499
rect 15489 2468 16129 2496
rect 15105 2431 15163 2437
rect 15105 2397 15117 2431
rect 15151 2397 15163 2431
rect 15105 2391 15163 2397
rect 12452 2332 13400 2360
rect 11609 2323 11667 2329
rect 14366 2320 14372 2372
rect 14424 2360 14430 2372
rect 15489 2360 15517 2468
rect 16117 2465 16129 2468
rect 16163 2465 16175 2499
rect 16117 2459 16175 2465
rect 16206 2456 16212 2508
rect 16264 2456 16270 2508
rect 19702 2456 19708 2508
rect 19760 2456 19766 2508
rect 25222 2456 25228 2508
rect 25280 2456 25286 2508
rect 31110 2456 31116 2508
rect 31168 2496 31174 2508
rect 31205 2499 31263 2505
rect 31205 2496 31217 2499
rect 31168 2468 31217 2496
rect 31168 2456 31174 2468
rect 31205 2465 31217 2468
rect 31251 2465 31263 2499
rect 31205 2459 31263 2465
rect 16224 2428 16252 2456
rect 16301 2431 16359 2437
rect 16301 2428 16313 2431
rect 16224 2400 16313 2428
rect 16301 2397 16313 2400
rect 16347 2397 16359 2431
rect 16301 2391 16359 2397
rect 16485 2431 16543 2437
rect 16485 2397 16497 2431
rect 16531 2428 16543 2431
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16531 2400 16865 2428
rect 16531 2397 16543 2400
rect 16485 2391 16543 2397
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 19720 2428 19748 2456
rect 19797 2431 19855 2437
rect 19797 2428 19809 2431
rect 19720 2400 19809 2428
rect 16853 2391 16911 2397
rect 19797 2397 19809 2400
rect 19843 2397 19855 2431
rect 19797 2391 19855 2397
rect 24670 2388 24676 2440
rect 24728 2388 24734 2440
rect 25240 2428 25268 2456
rect 25317 2431 25375 2437
rect 25317 2428 25329 2431
rect 25240 2400 25329 2428
rect 25317 2397 25329 2400
rect 25363 2397 25375 2431
rect 25317 2391 25375 2397
rect 26694 2388 26700 2440
rect 26752 2428 26758 2440
rect 27065 2431 27123 2437
rect 27065 2428 27077 2431
rect 26752 2400 27077 2428
rect 26752 2388 26758 2400
rect 27065 2397 27077 2400
rect 27111 2397 27123 2431
rect 27065 2391 27123 2397
rect 31018 2388 31024 2440
rect 31076 2388 31082 2440
rect 35526 2388 35532 2440
rect 35584 2388 35590 2440
rect 37274 2388 37280 2440
rect 37332 2428 37338 2440
rect 37369 2431 37427 2437
rect 37369 2428 37381 2431
rect 37332 2400 37381 2428
rect 37332 2388 37338 2400
rect 37369 2397 37381 2400
rect 37415 2397 37427 2431
rect 37369 2391 37427 2397
rect 14424 2332 15517 2360
rect 14424 2320 14430 2332
rect 15562 2320 15568 2372
rect 15620 2320 15626 2372
rect 15933 2363 15991 2369
rect 15933 2329 15945 2363
rect 15979 2360 15991 2363
rect 20165 2363 20223 2369
rect 20165 2360 20177 2363
rect 15979 2332 16574 2360
rect 15979 2329 15991 2332
rect 15933 2323 15991 2329
rect 11057 2295 11115 2301
rect 11057 2261 11069 2295
rect 11103 2261 11115 2295
rect 11057 2255 11115 2261
rect 11146 2252 11152 2304
rect 11204 2292 11210 2304
rect 11701 2295 11759 2301
rect 11701 2292 11713 2295
rect 11204 2264 11713 2292
rect 11204 2252 11210 2264
rect 11701 2261 11713 2264
rect 11747 2261 11759 2295
rect 16546 2292 16574 2332
rect 19996 2332 20177 2360
rect 19996 2301 20024 2332
rect 20165 2329 20177 2332
rect 20211 2329 20223 2363
rect 20165 2323 20223 2329
rect 16669 2295 16727 2301
rect 16669 2292 16681 2295
rect 16546 2264 16681 2292
rect 11701 2255 11759 2261
rect 16669 2261 16681 2264
rect 16715 2261 16727 2295
rect 16669 2255 16727 2261
rect 19981 2295 20039 2301
rect 19981 2261 19993 2295
rect 20027 2261 20039 2295
rect 19981 2255 20039 2261
rect 20254 2252 20260 2304
rect 20312 2252 20318 2304
rect 24578 2252 24584 2304
rect 24636 2292 24642 2304
rect 24949 2295 25007 2301
rect 24949 2292 24961 2295
rect 24636 2264 24961 2292
rect 24636 2252 24642 2264
rect 24949 2261 24961 2264
rect 24995 2261 25007 2295
rect 24949 2255 25007 2261
rect 26418 2252 26424 2304
rect 26476 2292 26482 2304
rect 27157 2295 27215 2301
rect 27157 2292 27169 2295
rect 26476 2264 27169 2292
rect 26476 2252 26482 2264
rect 27157 2261 27169 2264
rect 27203 2261 27215 2295
rect 27157 2255 27215 2261
rect 35710 2252 35716 2304
rect 35768 2252 35774 2304
rect 37645 2295 37703 2301
rect 37645 2261 37657 2295
rect 37691 2292 37703 2295
rect 37734 2292 37740 2304
rect 37691 2264 37740 2292
rect 37691 2261 37703 2264
rect 37645 2255 37703 2261
rect 37734 2252 37740 2264
rect 37792 2252 37798 2304
rect 1104 2202 38272 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 38272 2202
rect 1104 2128 38272 2150
<< via1 >>
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 35594 39142 35646 39194
rect 35658 39142 35710 39194
rect 35722 39142 35774 39194
rect 35786 39142 35838 39194
rect 35850 39142 35902 39194
rect 664 39040 716 39092
rect 1124 38972 1176 39024
rect 5264 39040 5316 39092
rect 9772 39040 9824 39092
rect 14188 39040 14240 39092
rect 17592 39083 17644 39092
rect 17592 39049 17601 39083
rect 17601 39049 17635 39083
rect 17635 39049 17644 39083
rect 17592 39040 17644 39049
rect 23204 39040 23256 39092
rect 25136 39040 25188 39092
rect 27344 39083 27396 39092
rect 27344 39049 27353 39083
rect 27353 39049 27387 39083
rect 27387 39049 27396 39083
rect 27344 39040 27396 39049
rect 31852 39040 31904 39092
rect 34152 39040 34204 39092
rect 36360 39083 36412 39092
rect 36360 39049 36369 39083
rect 36369 39049 36403 39083
rect 36403 39049 36412 39083
rect 36360 39040 36412 39049
rect 20720 38972 20772 39024
rect 23940 38972 23992 39024
rect 1768 38947 1820 38956
rect 1768 38913 1777 38947
rect 1777 38913 1811 38947
rect 1811 38913 1820 38947
rect 1768 38904 1820 38913
rect 2044 38947 2096 38956
rect 2044 38913 2053 38947
rect 2053 38913 2087 38947
rect 2087 38913 2096 38947
rect 2044 38904 2096 38913
rect 9680 38904 9732 38956
rect 10140 38947 10192 38956
rect 10140 38913 10149 38947
rect 10149 38913 10183 38947
rect 10183 38913 10192 38947
rect 10140 38904 10192 38913
rect 14740 38947 14792 38956
rect 14740 38913 14749 38947
rect 14749 38913 14783 38947
rect 14783 38913 14792 38947
rect 14740 38904 14792 38913
rect 17776 38947 17828 38956
rect 17776 38913 17785 38947
rect 17785 38913 17819 38947
rect 17819 38913 17828 38947
rect 17776 38904 17828 38913
rect 23388 38947 23440 38956
rect 23388 38913 23397 38947
rect 23397 38913 23431 38947
rect 23431 38913 23440 38947
rect 23388 38904 23440 38913
rect 25228 38947 25280 38956
rect 25228 38913 25237 38947
rect 25237 38913 25271 38947
rect 25271 38913 25280 38947
rect 25228 38904 25280 38913
rect 27252 38947 27304 38956
rect 27252 38913 27261 38947
rect 27261 38913 27295 38947
rect 27295 38913 27304 38947
rect 27252 38904 27304 38913
rect 14832 38836 14884 38888
rect 33600 38904 33652 38956
rect 37188 38972 37240 39024
rect 13912 38768 13964 38820
rect 14648 38700 14700 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 2044 38496 2096 38548
rect 9680 38496 9732 38548
rect 19432 38496 19484 38548
rect 21088 38496 21140 38548
rect 11612 38335 11664 38344
rect 11612 38301 11621 38335
rect 11621 38301 11655 38335
rect 11655 38301 11664 38335
rect 11612 38292 11664 38301
rect 14188 38292 14240 38344
rect 17960 38360 18012 38412
rect 23204 38428 23256 38480
rect 23480 38428 23532 38480
rect 21088 38292 21140 38344
rect 23204 38292 23256 38344
rect 24032 38335 24084 38344
rect 24032 38301 24041 38335
rect 24041 38301 24075 38335
rect 24075 38301 24084 38335
rect 24032 38292 24084 38301
rect 15292 38267 15344 38276
rect 15292 38233 15301 38267
rect 15301 38233 15335 38267
rect 15335 38233 15344 38267
rect 15292 38224 15344 38233
rect 15844 38224 15896 38276
rect 17592 38267 17644 38276
rect 17592 38233 17601 38267
rect 17601 38233 17635 38267
rect 17635 38233 17644 38267
rect 17592 38224 17644 38233
rect 19432 38224 19484 38276
rect 19984 38267 20036 38276
rect 19984 38233 19993 38267
rect 19993 38233 20027 38267
rect 20027 38233 20036 38267
rect 19984 38224 20036 38233
rect 22100 38267 22152 38276
rect 22100 38233 22109 38267
rect 22109 38233 22143 38267
rect 22143 38233 22152 38267
rect 22100 38224 22152 38233
rect 23480 38224 23532 38276
rect 24124 38224 24176 38276
rect 10324 38156 10376 38208
rect 16764 38199 16816 38208
rect 16764 38165 16773 38199
rect 16773 38165 16807 38199
rect 16807 38165 16816 38199
rect 16764 38156 16816 38165
rect 19064 38199 19116 38208
rect 19064 38165 19073 38199
rect 19073 38165 19107 38199
rect 19107 38165 19116 38199
rect 19064 38156 19116 38165
rect 20720 38156 20772 38208
rect 21456 38199 21508 38208
rect 21456 38165 21465 38199
rect 21465 38165 21499 38199
rect 21499 38165 21508 38199
rect 21456 38156 21508 38165
rect 22928 38156 22980 38208
rect 25044 38156 25096 38208
rect 26056 38156 26108 38208
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 35594 38054 35646 38106
rect 35658 38054 35710 38106
rect 35722 38054 35774 38106
rect 35786 38054 35838 38106
rect 35850 38054 35902 38106
rect 10140 37952 10192 38004
rect 10324 37952 10376 38004
rect 15292 37952 15344 38004
rect 14004 37884 14056 37936
rect 16396 37952 16448 38004
rect 16764 37952 16816 38004
rect 17776 37952 17828 38004
rect 12072 37816 12124 37868
rect 12992 37859 13044 37868
rect 12992 37825 13001 37859
rect 13001 37825 13035 37859
rect 13035 37825 13044 37859
rect 12992 37816 13044 37825
rect 17684 37884 17736 37936
rect 19064 37952 19116 38004
rect 19984 37952 20036 38004
rect 20720 37995 20772 38004
rect 20720 37961 20729 37995
rect 20729 37961 20763 37995
rect 20763 37961 20772 37995
rect 20720 37952 20772 37961
rect 22100 37952 22152 38004
rect 14004 37748 14056 37800
rect 16120 37859 16172 37868
rect 16120 37825 16129 37859
rect 16129 37825 16163 37859
rect 16163 37825 16172 37859
rect 16120 37816 16172 37825
rect 16212 37859 16264 37868
rect 16212 37825 16221 37859
rect 16221 37825 16255 37859
rect 16255 37825 16264 37859
rect 16212 37816 16264 37825
rect 16304 37859 16356 37868
rect 16304 37825 16313 37859
rect 16313 37825 16347 37859
rect 16347 37825 16356 37859
rect 16304 37816 16356 37825
rect 16396 37816 16448 37868
rect 17132 37791 17184 37800
rect 17132 37757 17141 37791
rect 17141 37757 17175 37791
rect 17175 37757 17184 37791
rect 17132 37748 17184 37757
rect 17316 37791 17368 37800
rect 17316 37757 17325 37791
rect 17325 37757 17359 37791
rect 17359 37757 17368 37791
rect 17316 37748 17368 37757
rect 18052 37791 18104 37800
rect 18052 37757 18061 37791
rect 18061 37757 18095 37791
rect 18095 37757 18104 37791
rect 18052 37748 18104 37757
rect 19800 37748 19852 37800
rect 940 37612 992 37664
rect 1768 37612 1820 37664
rect 19984 37680 20036 37732
rect 20812 37791 20864 37800
rect 20812 37757 20821 37791
rect 20821 37757 20855 37791
rect 20855 37757 20864 37791
rect 20812 37748 20864 37757
rect 22928 37995 22980 38004
rect 22928 37961 22937 37995
rect 22937 37961 22971 37995
rect 22971 37961 22980 37995
rect 22928 37952 22980 37961
rect 24032 37952 24084 38004
rect 25044 37952 25096 38004
rect 25228 37995 25280 38004
rect 25228 37961 25237 37995
rect 25237 37961 25271 37995
rect 25271 37961 25280 37995
rect 25228 37952 25280 37961
rect 27252 37952 27304 38004
rect 23020 37791 23072 37800
rect 23020 37757 23029 37791
rect 23029 37757 23063 37791
rect 23063 37757 23072 37791
rect 23020 37748 23072 37757
rect 23756 37748 23808 37800
rect 24860 37791 24912 37800
rect 24860 37757 24869 37791
rect 24869 37757 24903 37791
rect 24903 37757 24912 37791
rect 24860 37748 24912 37757
rect 25596 37859 25648 37868
rect 25596 37825 25605 37859
rect 25605 37825 25639 37859
rect 25639 37825 25648 37859
rect 25596 37816 25648 37825
rect 25688 37859 25740 37868
rect 25688 37825 25697 37859
rect 25697 37825 25731 37859
rect 25731 37825 25740 37859
rect 25688 37816 25740 37825
rect 25780 37748 25832 37800
rect 24952 37612 25004 37664
rect 26148 37859 26200 37868
rect 26148 37825 26157 37859
rect 26157 37825 26191 37859
rect 26191 37825 26200 37859
rect 26148 37816 26200 37825
rect 27252 37816 27304 37868
rect 37648 37859 37700 37868
rect 37648 37825 37657 37859
rect 37657 37825 37691 37859
rect 37691 37825 37700 37859
rect 37648 37816 37700 37825
rect 37832 37655 37884 37664
rect 37832 37621 37841 37655
rect 37841 37621 37875 37655
rect 37875 37621 37884 37655
rect 37832 37612 37884 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 11612 37451 11664 37460
rect 11612 37417 11621 37451
rect 11621 37417 11655 37451
rect 11655 37417 11664 37451
rect 11612 37408 11664 37417
rect 12072 37451 12124 37460
rect 12072 37417 12081 37451
rect 12081 37417 12115 37451
rect 12115 37417 12124 37451
rect 12072 37408 12124 37417
rect 16120 37408 16172 37460
rect 16304 37408 16356 37460
rect 19984 37451 20036 37460
rect 19984 37417 19993 37451
rect 19993 37417 20027 37451
rect 20027 37417 20036 37451
rect 19984 37408 20036 37417
rect 20352 37408 20404 37460
rect 21088 37408 21140 37460
rect 22836 37408 22888 37460
rect 25688 37408 25740 37460
rect 26148 37408 26200 37460
rect 24676 37340 24728 37392
rect 2596 37272 2648 37324
rect 8484 37272 8536 37324
rect 11980 37315 12032 37324
rect 11980 37281 11989 37315
rect 11989 37281 12023 37315
rect 12023 37281 12032 37315
rect 11980 37272 12032 37281
rect 14464 37272 14516 37324
rect 16120 37272 16172 37324
rect 12440 37247 12492 37256
rect 12440 37213 12449 37247
rect 12449 37213 12483 37247
rect 12483 37213 12492 37247
rect 12440 37204 12492 37213
rect 12716 37247 12768 37256
rect 12716 37213 12725 37247
rect 12725 37213 12759 37247
rect 12759 37213 12768 37247
rect 12716 37204 12768 37213
rect 16304 37204 16356 37256
rect 16764 37204 16816 37256
rect 20168 37272 20220 37324
rect 21548 37272 21600 37324
rect 13544 37136 13596 37188
rect 19892 37204 19944 37256
rect 19340 37136 19392 37188
rect 20536 37204 20588 37256
rect 20996 37204 21048 37256
rect 22928 37204 22980 37256
rect 21088 37179 21140 37188
rect 21088 37145 21097 37179
rect 21097 37145 21131 37179
rect 21131 37145 21140 37179
rect 21088 37136 21140 37145
rect 22836 37136 22888 37188
rect 25136 37136 25188 37188
rect 11612 37068 11664 37120
rect 12900 37111 12952 37120
rect 12900 37077 12909 37111
rect 12909 37077 12943 37111
rect 12943 37077 12952 37111
rect 12900 37068 12952 37077
rect 19064 37068 19116 37120
rect 21548 37068 21600 37120
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 12716 36907 12768 36916
rect 12716 36873 12725 36907
rect 12725 36873 12759 36907
rect 12759 36873 12768 36907
rect 12716 36864 12768 36873
rect 12900 36864 12952 36916
rect 10692 36660 10744 36712
rect 12992 36796 13044 36848
rect 20812 36864 20864 36916
rect 21272 36864 21324 36916
rect 21732 36864 21784 36916
rect 19432 36796 19484 36848
rect 21456 36796 21508 36848
rect 21916 36796 21968 36848
rect 23020 36864 23072 36916
rect 33600 36907 33652 36916
rect 33600 36873 33609 36907
rect 33609 36873 33643 36907
rect 33643 36873 33652 36907
rect 33600 36864 33652 36873
rect 37648 36864 37700 36916
rect 12348 36771 12400 36780
rect 12348 36737 12357 36771
rect 12357 36737 12391 36771
rect 12391 36737 12400 36771
rect 12348 36728 12400 36737
rect 14096 36728 14148 36780
rect 15844 36728 15896 36780
rect 17960 36728 18012 36780
rect 21364 36728 21416 36780
rect 22928 36728 22980 36780
rect 23664 36771 23716 36780
rect 23664 36737 23673 36771
rect 23673 36737 23707 36771
rect 23707 36737 23716 36771
rect 23664 36728 23716 36737
rect 12716 36660 12768 36712
rect 18420 36703 18472 36712
rect 18420 36669 18429 36703
rect 18429 36669 18463 36703
rect 18463 36669 18472 36703
rect 18420 36660 18472 36669
rect 21180 36703 21232 36712
rect 21180 36669 21189 36703
rect 21189 36669 21223 36703
rect 21223 36669 21232 36703
rect 21180 36660 21232 36669
rect 21272 36703 21324 36712
rect 21272 36669 21281 36703
rect 21281 36669 21315 36703
rect 21315 36669 21324 36703
rect 21272 36660 21324 36669
rect 25136 36771 25188 36780
rect 25136 36737 25145 36771
rect 25145 36737 25179 36771
rect 25179 36737 25188 36771
rect 25136 36728 25188 36737
rect 25412 36660 25464 36712
rect 14188 36524 14240 36576
rect 14556 36567 14608 36576
rect 14556 36533 14565 36567
rect 14565 36533 14599 36567
rect 14599 36533 14608 36567
rect 14556 36524 14608 36533
rect 21272 36524 21324 36576
rect 22008 36567 22060 36576
rect 22008 36533 22017 36567
rect 22017 36533 22051 36567
rect 22051 36533 22060 36567
rect 22008 36524 22060 36533
rect 28448 36728 28500 36780
rect 37372 36771 37424 36780
rect 37372 36737 37381 36771
rect 37381 36737 37415 36771
rect 37415 36737 37424 36771
rect 37372 36728 37424 36737
rect 25320 36567 25372 36576
rect 25320 36533 25329 36567
rect 25329 36533 25363 36567
rect 25363 36533 25372 36567
rect 25320 36524 25372 36533
rect 25964 36524 26016 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 9864 36184 9916 36236
rect 14096 36320 14148 36372
rect 14832 36363 14884 36372
rect 14832 36329 14841 36363
rect 14841 36329 14875 36363
rect 14875 36329 14884 36363
rect 14832 36320 14884 36329
rect 17132 36320 17184 36372
rect 18420 36320 18472 36372
rect 21180 36320 21232 36372
rect 24860 36363 24912 36372
rect 24860 36329 24869 36363
rect 24869 36329 24903 36363
rect 24903 36329 24912 36363
rect 24860 36320 24912 36329
rect 25320 36320 25372 36372
rect 25964 36363 26016 36372
rect 25964 36329 25973 36363
rect 25973 36329 26007 36363
rect 26007 36329 26016 36363
rect 25964 36320 26016 36329
rect 28448 36363 28500 36372
rect 28448 36329 28457 36363
rect 28457 36329 28491 36363
rect 28491 36329 28500 36363
rect 28448 36320 28500 36329
rect 37372 36320 37424 36372
rect 12992 36252 13044 36304
rect 8300 36116 8352 36168
rect 9220 36116 9272 36168
rect 9772 36091 9824 36100
rect 9772 36057 9781 36091
rect 9781 36057 9815 36091
rect 9815 36057 9824 36091
rect 9772 36048 9824 36057
rect 11612 36048 11664 36100
rect 13544 36091 13596 36100
rect 13544 36057 13553 36091
rect 13553 36057 13587 36091
rect 13587 36057 13596 36091
rect 13544 36048 13596 36057
rect 14096 36116 14148 36168
rect 15384 36227 15436 36236
rect 15384 36193 15393 36227
rect 15393 36193 15427 36227
rect 15427 36193 15436 36227
rect 15384 36184 15436 36193
rect 17316 36252 17368 36304
rect 16580 36184 16632 36236
rect 14464 36159 14516 36168
rect 14464 36125 14473 36159
rect 14473 36125 14507 36159
rect 14507 36125 14516 36159
rect 14464 36116 14516 36125
rect 15200 36116 15252 36168
rect 15752 36116 15804 36168
rect 16304 36159 16356 36168
rect 16304 36125 16313 36159
rect 16313 36125 16347 36159
rect 16347 36125 16356 36159
rect 16304 36116 16356 36125
rect 16764 36116 16816 36168
rect 18788 36184 18840 36236
rect 21272 36252 21324 36304
rect 19800 36227 19852 36236
rect 19800 36193 19809 36227
rect 19809 36193 19843 36227
rect 19843 36193 19852 36227
rect 19800 36184 19852 36193
rect 19616 36159 19668 36168
rect 19616 36125 19625 36159
rect 19625 36125 19659 36159
rect 19659 36125 19668 36159
rect 19616 36116 19668 36125
rect 11244 36023 11296 36032
rect 11244 35989 11253 36023
rect 11253 35989 11287 36023
rect 11287 35989 11296 36023
rect 11244 35980 11296 35989
rect 12624 35980 12676 36032
rect 14924 36023 14976 36032
rect 14924 35989 14933 36023
rect 14933 35989 14967 36023
rect 14967 35989 14976 36023
rect 14924 35980 14976 35989
rect 17132 36023 17184 36032
rect 17132 35989 17141 36023
rect 17141 35989 17175 36023
rect 17175 35989 17184 36023
rect 17132 35980 17184 35989
rect 19708 36023 19760 36032
rect 19708 35989 19717 36023
rect 19717 35989 19751 36023
rect 19751 35989 19760 36023
rect 19708 35980 19760 35989
rect 20996 36048 21048 36100
rect 21916 36184 21968 36236
rect 22100 36116 22152 36168
rect 25412 36227 25464 36236
rect 25412 36193 25421 36227
rect 25421 36193 25455 36227
rect 25455 36193 25464 36227
rect 25412 36184 25464 36193
rect 25688 36159 25740 36168
rect 25688 36125 25697 36159
rect 25697 36125 25731 36159
rect 25731 36125 25740 36159
rect 25688 36116 25740 36125
rect 22836 36048 22888 36100
rect 26056 36116 26108 36168
rect 27804 36116 27856 36168
rect 28632 36159 28684 36168
rect 28632 36125 28641 36159
rect 28641 36125 28675 36159
rect 28675 36125 28684 36159
rect 28632 36116 28684 36125
rect 23112 36023 23164 36032
rect 23112 35989 23121 36023
rect 23121 35989 23155 36023
rect 23155 35989 23164 36023
rect 23112 35980 23164 35989
rect 25228 36023 25280 36032
rect 25228 35989 25237 36023
rect 25237 35989 25271 36023
rect 25271 35989 25280 36023
rect 25228 35980 25280 35989
rect 25872 35980 25924 36032
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 9772 35776 9824 35828
rect 9864 35708 9916 35760
rect 8208 35683 8260 35692
rect 8208 35649 8217 35683
rect 8217 35649 8251 35683
rect 8251 35649 8260 35683
rect 8208 35640 8260 35649
rect 11244 35776 11296 35828
rect 12624 35776 12676 35828
rect 12716 35776 12768 35828
rect 13360 35776 13412 35828
rect 8944 35572 8996 35624
rect 9956 35615 10008 35624
rect 9956 35581 9965 35615
rect 9965 35581 9999 35615
rect 9999 35581 10008 35615
rect 9956 35572 10008 35581
rect 11060 35615 11112 35624
rect 11060 35581 11069 35615
rect 11069 35581 11103 35615
rect 11103 35581 11112 35615
rect 11060 35572 11112 35581
rect 11244 35572 11296 35624
rect 12440 35683 12492 35692
rect 12440 35649 12449 35683
rect 12449 35649 12483 35683
rect 12483 35649 12492 35683
rect 12440 35640 12492 35649
rect 13452 35708 13504 35760
rect 15844 35708 15896 35760
rect 16580 35776 16632 35828
rect 16396 35708 16448 35760
rect 18052 35776 18104 35828
rect 19616 35776 19668 35828
rect 12532 35615 12584 35624
rect 12532 35581 12541 35615
rect 12541 35581 12575 35615
rect 12575 35581 12584 35615
rect 12532 35572 12584 35581
rect 12992 35572 13044 35624
rect 11796 35504 11848 35556
rect 10692 35436 10744 35488
rect 11888 35479 11940 35488
rect 11888 35445 11897 35479
rect 11897 35445 11931 35479
rect 11931 35445 11940 35479
rect 11888 35436 11940 35445
rect 12348 35436 12400 35488
rect 14188 35615 14240 35624
rect 14188 35581 14197 35615
rect 14197 35581 14231 35615
rect 14231 35581 14240 35615
rect 14188 35572 14240 35581
rect 14464 35615 14516 35624
rect 14464 35581 14473 35615
rect 14473 35581 14507 35615
rect 14507 35581 14516 35615
rect 14464 35572 14516 35581
rect 16856 35615 16908 35624
rect 16856 35581 16865 35615
rect 16865 35581 16899 35615
rect 16899 35581 16908 35615
rect 16856 35572 16908 35581
rect 13636 35504 13688 35556
rect 17684 35615 17736 35624
rect 17684 35581 17693 35615
rect 17693 35581 17727 35615
rect 17727 35581 17736 35615
rect 17684 35572 17736 35581
rect 18052 35683 18104 35692
rect 18052 35649 18061 35683
rect 18061 35649 18095 35683
rect 18095 35649 18104 35683
rect 18052 35640 18104 35649
rect 18880 35640 18932 35692
rect 18788 35615 18840 35624
rect 18788 35581 18797 35615
rect 18797 35581 18831 35615
rect 18831 35581 18840 35615
rect 18788 35572 18840 35581
rect 13176 35479 13228 35488
rect 13176 35445 13185 35479
rect 13185 35445 13219 35479
rect 13219 35445 13228 35479
rect 13176 35436 13228 35445
rect 15752 35436 15804 35488
rect 16120 35479 16172 35488
rect 16120 35445 16129 35479
rect 16129 35445 16163 35479
rect 16163 35445 16172 35479
rect 16120 35436 16172 35445
rect 17868 35504 17920 35556
rect 25136 35776 25188 35828
rect 22100 35708 22152 35760
rect 22744 35640 22796 35692
rect 22468 35615 22520 35624
rect 22468 35581 22477 35615
rect 22477 35581 22511 35615
rect 22511 35581 22520 35615
rect 22468 35572 22520 35581
rect 25688 35708 25740 35760
rect 25872 35708 25924 35760
rect 25136 35683 25188 35692
rect 25136 35649 25145 35683
rect 25145 35649 25179 35683
rect 25179 35649 25188 35683
rect 25136 35640 25188 35649
rect 37648 35683 37700 35692
rect 37648 35649 37657 35683
rect 37657 35649 37691 35683
rect 37691 35649 37700 35683
rect 37648 35640 37700 35649
rect 16488 35436 16540 35488
rect 17684 35436 17736 35488
rect 18144 35436 18196 35488
rect 19616 35479 19668 35488
rect 19616 35445 19625 35479
rect 19625 35445 19659 35479
rect 19659 35445 19668 35479
rect 19616 35436 19668 35445
rect 22652 35436 22704 35488
rect 25504 35479 25556 35488
rect 25504 35445 25513 35479
rect 25513 35445 25547 35479
rect 25547 35445 25556 35479
rect 25504 35436 25556 35445
rect 26056 35436 26108 35488
rect 37832 35479 37884 35488
rect 37832 35445 37841 35479
rect 37841 35445 37875 35479
rect 37875 35445 37884 35479
rect 37832 35436 37884 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 8944 35275 8996 35284
rect 8944 35241 8953 35275
rect 8953 35241 8987 35275
rect 8987 35241 8996 35275
rect 8944 35232 8996 35241
rect 9956 35232 10008 35284
rect 11060 35232 11112 35284
rect 11796 35232 11848 35284
rect 11888 35232 11940 35284
rect 12440 35232 12492 35284
rect 12624 35232 12676 35284
rect 13360 35275 13412 35284
rect 13360 35241 13369 35275
rect 13369 35241 13403 35275
rect 13403 35241 13412 35275
rect 13360 35232 13412 35241
rect 14464 35232 14516 35284
rect 15384 35232 15436 35284
rect 16856 35232 16908 35284
rect 17868 35232 17920 35284
rect 18052 35232 18104 35284
rect 19708 35232 19760 35284
rect 23388 35232 23440 35284
rect 25504 35232 25556 35284
rect 37648 35232 37700 35284
rect 10692 35096 10744 35148
rect 940 34960 992 35012
rect 6000 34960 6052 35012
rect 12900 35096 12952 35148
rect 16764 35164 16816 35216
rect 18788 35164 18840 35216
rect 11980 35071 12032 35080
rect 11980 35037 11989 35071
rect 11989 35037 12023 35071
rect 12023 35037 12032 35071
rect 11980 35028 12032 35037
rect 12348 35071 12400 35080
rect 12348 35037 12357 35071
rect 12357 35037 12391 35071
rect 12391 35037 12400 35071
rect 12348 35028 12400 35037
rect 12440 35071 12492 35080
rect 12440 35037 12449 35071
rect 12449 35037 12483 35071
rect 12483 35037 12492 35071
rect 12440 35028 12492 35037
rect 11704 35003 11756 35012
rect 11704 34969 11713 35003
rect 11713 34969 11747 35003
rect 11747 34969 11756 35003
rect 11704 34960 11756 34969
rect 9864 34935 9916 34944
rect 9864 34901 9873 34935
rect 9873 34901 9907 34935
rect 9907 34901 9916 34935
rect 9864 34892 9916 34901
rect 11612 34892 11664 34944
rect 12532 34960 12584 35012
rect 12992 35071 13044 35080
rect 12992 35037 13001 35071
rect 13001 35037 13035 35071
rect 13035 35037 13044 35071
rect 12992 35028 13044 35037
rect 13268 35096 13320 35148
rect 15844 35096 15896 35148
rect 13452 35071 13504 35080
rect 13452 35037 13461 35071
rect 13461 35037 13495 35071
rect 13495 35037 13504 35071
rect 13452 35028 13504 35037
rect 14924 35028 14976 35080
rect 12716 34892 12768 34944
rect 13636 35003 13688 35012
rect 13636 34969 13645 35003
rect 13645 34969 13679 35003
rect 13679 34969 13688 35003
rect 13636 34960 13688 34969
rect 14556 34960 14608 35012
rect 16580 35071 16632 35080
rect 16580 35037 16589 35071
rect 16589 35037 16623 35071
rect 16623 35037 16632 35071
rect 16580 35028 16632 35037
rect 16764 35071 16816 35080
rect 16764 35037 16773 35071
rect 16773 35037 16807 35071
rect 16807 35037 16816 35071
rect 16764 35028 16816 35037
rect 15292 34960 15344 35012
rect 16672 35003 16724 35012
rect 16672 34969 16681 35003
rect 16681 34969 16715 35003
rect 16715 34969 16724 35003
rect 16672 34960 16724 34969
rect 16856 35003 16908 35012
rect 16856 34969 16891 35003
rect 16891 34969 16908 35003
rect 17868 35028 17920 35080
rect 18144 35071 18196 35080
rect 18144 35037 18153 35071
rect 18153 35037 18187 35071
rect 18187 35037 18196 35071
rect 18144 35028 18196 35037
rect 18236 35028 18288 35080
rect 19340 35096 19392 35148
rect 22468 35164 22520 35216
rect 19616 35096 19668 35148
rect 20536 35096 20588 35148
rect 21732 35139 21784 35148
rect 21732 35105 21741 35139
rect 21741 35105 21775 35139
rect 21775 35105 21784 35139
rect 21732 35096 21784 35105
rect 20260 35071 20312 35080
rect 20260 35037 20269 35071
rect 20269 35037 20303 35071
rect 20303 35037 20312 35071
rect 20260 35028 20312 35037
rect 20352 35071 20404 35080
rect 20352 35037 20361 35071
rect 20361 35037 20395 35071
rect 20395 35037 20404 35071
rect 20352 35028 20404 35037
rect 21180 35071 21232 35080
rect 21180 35037 21189 35071
rect 21189 35037 21223 35071
rect 21223 35037 21232 35071
rect 21180 35028 21232 35037
rect 22652 35071 22704 35080
rect 22652 35037 22661 35071
rect 22661 35037 22695 35071
rect 22695 35037 22704 35071
rect 22652 35028 22704 35037
rect 22744 35071 22796 35080
rect 22744 35037 22753 35071
rect 22753 35037 22787 35071
rect 22787 35037 22796 35071
rect 22744 35028 22796 35037
rect 23756 35096 23808 35148
rect 25412 35096 25464 35148
rect 25136 35028 25188 35080
rect 37372 35071 37424 35080
rect 37372 35037 37381 35071
rect 37381 35037 37415 35071
rect 37415 35037 37424 35071
rect 37372 35028 37424 35037
rect 16856 34960 16908 34969
rect 17868 34892 17920 34944
rect 19064 34935 19116 34944
rect 19064 34901 19073 34935
rect 19073 34901 19107 34935
rect 19107 34901 19116 34935
rect 19064 34892 19116 34901
rect 20168 34892 20220 34944
rect 20996 34935 21048 34944
rect 20996 34901 21005 34935
rect 21005 34901 21039 34935
rect 21039 34901 21048 34935
rect 20996 34892 21048 34901
rect 21272 34892 21324 34944
rect 22376 34935 22428 34944
rect 22376 34901 22385 34935
rect 22385 34901 22419 34935
rect 22419 34901 22428 34935
rect 22376 34892 22428 34901
rect 24400 34935 24452 34944
rect 24400 34901 24409 34935
rect 24409 34901 24443 34935
rect 24443 34901 24452 34935
rect 24400 34892 24452 34901
rect 25596 34935 25648 34944
rect 25596 34901 25605 34935
rect 25605 34901 25639 34935
rect 25639 34901 25648 34935
rect 25596 34892 25648 34901
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 9864 34688 9916 34740
rect 11704 34688 11756 34740
rect 11612 34552 11664 34604
rect 12348 34620 12400 34672
rect 13452 34688 13504 34740
rect 14372 34688 14424 34740
rect 16672 34688 16724 34740
rect 20260 34688 20312 34740
rect 20352 34688 20404 34740
rect 21180 34688 21232 34740
rect 22376 34688 22428 34740
rect 22468 34688 22520 34740
rect 25136 34688 25188 34740
rect 26608 34688 26660 34740
rect 27528 34688 27580 34740
rect 13636 34620 13688 34672
rect 18236 34620 18288 34672
rect 12256 34552 12308 34604
rect 12992 34552 13044 34604
rect 15292 34552 15344 34604
rect 16120 34595 16172 34604
rect 16120 34561 16129 34595
rect 16129 34561 16163 34595
rect 16163 34561 16172 34595
rect 16120 34552 16172 34561
rect 24124 34620 24176 34672
rect 19984 34552 20036 34604
rect 29368 34595 29420 34604
rect 29368 34561 29377 34595
rect 29377 34561 29411 34595
rect 29411 34561 29420 34595
rect 29368 34552 29420 34561
rect 19432 34484 19484 34536
rect 21456 34484 21508 34536
rect 11980 34416 12032 34468
rect 12716 34416 12768 34468
rect 16856 34416 16908 34468
rect 12624 34348 12676 34400
rect 12900 34348 12952 34400
rect 15200 34348 15252 34400
rect 18236 34348 18288 34400
rect 23296 34527 23348 34536
rect 23296 34493 23305 34527
rect 23305 34493 23339 34527
rect 23339 34493 23348 34527
rect 23296 34484 23348 34493
rect 23572 34527 23624 34536
rect 23572 34493 23581 34527
rect 23581 34493 23615 34527
rect 23615 34493 23624 34527
rect 23572 34484 23624 34493
rect 28908 34484 28960 34536
rect 29828 34595 29880 34604
rect 29828 34561 29837 34595
rect 29837 34561 29871 34595
rect 29871 34561 29880 34595
rect 29828 34552 29880 34561
rect 23756 34348 23808 34400
rect 30104 34391 30156 34400
rect 30104 34357 30113 34391
rect 30113 34357 30147 34391
rect 30147 34357 30156 34391
rect 30104 34348 30156 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 14740 34187 14792 34196
rect 14740 34153 14749 34187
rect 14749 34153 14783 34187
rect 14783 34153 14792 34187
rect 14740 34144 14792 34153
rect 17868 34144 17920 34196
rect 22468 34187 22520 34196
rect 22468 34153 22477 34187
rect 22477 34153 22511 34187
rect 22511 34153 22520 34187
rect 22468 34144 22520 34153
rect 23572 34144 23624 34196
rect 26792 34144 26844 34196
rect 6920 34119 6972 34128
rect 6920 34085 6929 34119
rect 6929 34085 6963 34119
rect 6963 34085 6972 34119
rect 6920 34076 6972 34085
rect 23020 34076 23072 34128
rect 12440 34008 12492 34060
rect 12992 34008 13044 34060
rect 14188 34008 14240 34060
rect 23296 34008 23348 34060
rect 4068 33940 4120 33992
rect 14096 33983 14148 33992
rect 14096 33949 14105 33983
rect 14105 33949 14139 33983
rect 14139 33949 14148 33983
rect 14096 33940 14148 33949
rect 5724 33872 5776 33924
rect 5356 33804 5408 33856
rect 12900 33872 12952 33924
rect 14372 33983 14424 33992
rect 14372 33949 14381 33983
rect 14381 33949 14415 33983
rect 14415 33949 14424 33983
rect 14372 33940 14424 33949
rect 15384 33983 15436 33992
rect 15384 33949 15393 33983
rect 15393 33949 15427 33983
rect 15427 33949 15436 33983
rect 15384 33940 15436 33949
rect 15476 33940 15528 33992
rect 15108 33872 15160 33924
rect 15660 33872 15712 33924
rect 15936 33872 15988 33924
rect 18144 33940 18196 33992
rect 22468 33940 22520 33992
rect 24400 33940 24452 33992
rect 25136 33940 25188 33992
rect 27344 34076 27396 34128
rect 27528 34187 27580 34196
rect 27528 34153 27537 34187
rect 27537 34153 27571 34187
rect 27571 34153 27580 34187
rect 27528 34144 27580 34153
rect 26424 34008 26476 34060
rect 26608 33983 26660 33992
rect 26608 33949 26617 33983
rect 26617 33949 26651 33983
rect 26651 33949 26660 33983
rect 26608 33940 26660 33949
rect 30104 34008 30156 34060
rect 27528 33983 27580 33992
rect 27528 33949 27537 33983
rect 27537 33949 27571 33983
rect 27571 33949 27580 33983
rect 27528 33940 27580 33949
rect 29736 33940 29788 33992
rect 31392 34008 31444 34060
rect 20996 33915 21048 33924
rect 20996 33881 21005 33915
rect 21005 33881 21039 33915
rect 21039 33881 21048 33915
rect 20996 33872 21048 33881
rect 21456 33872 21508 33924
rect 23020 33872 23072 33924
rect 17408 33804 17460 33856
rect 17776 33847 17828 33856
rect 17776 33813 17785 33847
rect 17785 33813 17819 33847
rect 17819 33813 17828 33847
rect 17776 33804 17828 33813
rect 17868 33804 17920 33856
rect 23296 33847 23348 33856
rect 23296 33813 23305 33847
rect 23305 33813 23339 33847
rect 23339 33813 23348 33847
rect 23296 33804 23348 33813
rect 24124 33804 24176 33856
rect 25044 33847 25096 33856
rect 25044 33813 25053 33847
rect 25053 33813 25087 33847
rect 25087 33813 25096 33847
rect 25044 33804 25096 33813
rect 26332 33847 26384 33856
rect 26332 33813 26341 33847
rect 26341 33813 26375 33847
rect 26375 33813 26384 33847
rect 26332 33804 26384 33813
rect 27068 33847 27120 33856
rect 27068 33813 27077 33847
rect 27077 33813 27111 33847
rect 27111 33813 27120 33847
rect 27068 33804 27120 33813
rect 29092 33872 29144 33924
rect 31760 33940 31812 33992
rect 27252 33804 27304 33856
rect 27896 33804 27948 33856
rect 30472 33804 30524 33856
rect 30564 33847 30616 33856
rect 30564 33813 30573 33847
rect 30573 33813 30607 33847
rect 30607 33813 30616 33847
rect 30564 33804 30616 33813
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 5724 33600 5776 33652
rect 4620 33532 4672 33584
rect 5356 33532 5408 33584
rect 8300 33600 8352 33652
rect 11796 33600 11848 33652
rect 9772 33532 9824 33584
rect 9956 33532 10008 33584
rect 12256 33600 12308 33652
rect 12900 33643 12952 33652
rect 12900 33609 12909 33643
rect 12909 33609 12943 33643
rect 12943 33609 12952 33643
rect 12900 33600 12952 33609
rect 14188 33600 14240 33652
rect 11980 33575 12032 33584
rect 11980 33541 12015 33575
rect 12015 33541 12032 33575
rect 11980 33532 12032 33541
rect 13544 33532 13596 33584
rect 6092 33507 6144 33516
rect 6092 33473 6101 33507
rect 6101 33473 6135 33507
rect 6135 33473 6144 33507
rect 6092 33464 6144 33473
rect 6736 33507 6788 33516
rect 6736 33473 6745 33507
rect 6745 33473 6779 33507
rect 6779 33473 6788 33507
rect 6736 33464 6788 33473
rect 8944 33464 8996 33516
rect 4068 33439 4120 33448
rect 4068 33405 4077 33439
rect 4077 33405 4111 33439
rect 4111 33405 4120 33439
rect 4068 33396 4120 33405
rect 7012 33439 7064 33448
rect 7012 33405 7021 33439
rect 7021 33405 7055 33439
rect 7055 33405 7064 33439
rect 7012 33396 7064 33405
rect 11704 33507 11756 33516
rect 11704 33473 11713 33507
rect 11713 33473 11747 33507
rect 11747 33473 11756 33507
rect 11704 33464 11756 33473
rect 11796 33507 11848 33516
rect 11796 33473 11805 33507
rect 11805 33473 11839 33507
rect 11839 33473 11848 33507
rect 11796 33464 11848 33473
rect 11888 33507 11940 33516
rect 11888 33473 11897 33507
rect 11897 33473 11931 33507
rect 11931 33473 11940 33507
rect 11888 33464 11940 33473
rect 12716 33507 12768 33516
rect 12716 33473 12725 33507
rect 12725 33473 12759 33507
rect 12759 33473 12768 33507
rect 12716 33464 12768 33473
rect 9220 33439 9272 33448
rect 9220 33405 9229 33439
rect 9229 33405 9263 33439
rect 9263 33405 9272 33439
rect 9220 33396 9272 33405
rect 9956 33396 10008 33448
rect 11612 33396 11664 33448
rect 12440 33396 12492 33448
rect 13176 33464 13228 33516
rect 14832 33507 14884 33516
rect 14832 33473 14841 33507
rect 14841 33473 14875 33507
rect 14875 33473 14884 33507
rect 14832 33464 14884 33473
rect 15016 33507 15068 33516
rect 15016 33473 15025 33507
rect 15025 33473 15059 33507
rect 15059 33473 15068 33507
rect 15016 33464 15068 33473
rect 15384 33600 15436 33652
rect 15660 33643 15712 33652
rect 15660 33609 15669 33643
rect 15669 33609 15703 33643
rect 15703 33609 15712 33643
rect 15660 33600 15712 33609
rect 17132 33600 17184 33652
rect 21640 33600 21692 33652
rect 24676 33600 24728 33652
rect 26424 33600 26476 33652
rect 27068 33600 27120 33652
rect 15936 33507 15988 33516
rect 15936 33473 15945 33507
rect 15945 33473 15979 33507
rect 15979 33473 15988 33507
rect 15936 33464 15988 33473
rect 16028 33507 16080 33516
rect 16028 33473 16037 33507
rect 16037 33473 16071 33507
rect 16071 33473 16080 33507
rect 16028 33464 16080 33473
rect 17684 33464 17736 33516
rect 18328 33464 18380 33516
rect 17408 33439 17460 33448
rect 17408 33405 17417 33439
rect 17417 33405 17451 33439
rect 17451 33405 17460 33439
rect 17408 33396 17460 33405
rect 18052 33439 18104 33448
rect 18052 33405 18061 33439
rect 18061 33405 18095 33439
rect 18095 33405 18104 33439
rect 19340 33464 19392 33516
rect 19616 33464 19668 33516
rect 18052 33396 18104 33405
rect 20076 33464 20128 33516
rect 25872 33507 25924 33516
rect 25872 33473 25881 33507
rect 25881 33473 25915 33507
rect 25915 33473 25924 33507
rect 25872 33464 25924 33473
rect 26332 33464 26384 33516
rect 26516 33507 26568 33516
rect 26516 33473 26525 33507
rect 26525 33473 26559 33507
rect 26559 33473 26568 33507
rect 26516 33464 26568 33473
rect 27528 33507 27580 33516
rect 27528 33473 27537 33507
rect 27537 33473 27571 33507
rect 27571 33473 27580 33507
rect 27528 33464 27580 33473
rect 26608 33396 26660 33448
rect 27896 33439 27948 33448
rect 27896 33405 27905 33439
rect 27905 33405 27939 33439
rect 27939 33405 27948 33439
rect 27896 33396 27948 33405
rect 28172 33507 28224 33516
rect 28172 33473 28181 33507
rect 28181 33473 28215 33507
rect 28215 33473 28224 33507
rect 28172 33464 28224 33473
rect 29092 33643 29144 33652
rect 29092 33609 29101 33643
rect 29101 33609 29135 33643
rect 29135 33609 29144 33643
rect 29092 33600 29144 33609
rect 29736 33600 29788 33652
rect 30564 33600 30616 33652
rect 31760 33643 31812 33652
rect 31760 33609 31769 33643
rect 31769 33609 31803 33643
rect 31803 33609 31812 33643
rect 31760 33600 31812 33609
rect 29184 33464 29236 33516
rect 29276 33507 29328 33516
rect 29276 33473 29285 33507
rect 29285 33473 29319 33507
rect 29319 33473 29328 33507
rect 29276 33464 29328 33473
rect 5816 33303 5868 33312
rect 5816 33269 5825 33303
rect 5825 33269 5859 33303
rect 5859 33269 5868 33303
rect 20812 33328 20864 33380
rect 5816 33260 5868 33269
rect 10968 33303 11020 33312
rect 10968 33269 10977 33303
rect 10977 33269 11011 33303
rect 11011 33269 11020 33303
rect 10968 33260 11020 33269
rect 11520 33303 11572 33312
rect 11520 33269 11529 33303
rect 11529 33269 11563 33303
rect 11563 33269 11572 33303
rect 11520 33260 11572 33269
rect 12348 33260 12400 33312
rect 15200 33303 15252 33312
rect 15200 33269 15209 33303
rect 15209 33269 15243 33303
rect 15243 33269 15252 33303
rect 15200 33260 15252 33269
rect 15384 33260 15436 33312
rect 18512 33303 18564 33312
rect 18512 33269 18521 33303
rect 18521 33269 18555 33303
rect 18555 33269 18564 33303
rect 18512 33260 18564 33269
rect 19800 33303 19852 33312
rect 19800 33269 19809 33303
rect 19809 33269 19843 33303
rect 19843 33269 19852 33303
rect 19800 33260 19852 33269
rect 25688 33303 25740 33312
rect 25688 33269 25697 33303
rect 25697 33269 25731 33303
rect 25731 33269 25740 33303
rect 25688 33260 25740 33269
rect 27252 33328 27304 33380
rect 27436 33371 27488 33380
rect 27436 33337 27445 33371
rect 27445 33337 27479 33371
rect 27479 33337 27488 33371
rect 27436 33328 27488 33337
rect 28080 33371 28132 33380
rect 28080 33337 28089 33371
rect 28089 33337 28123 33371
rect 28123 33337 28132 33371
rect 28080 33328 28132 33337
rect 30104 33328 30156 33380
rect 29644 33303 29696 33312
rect 29644 33269 29653 33303
rect 29653 33269 29687 33303
rect 29687 33269 29696 33303
rect 29644 33260 29696 33269
rect 30288 33439 30340 33448
rect 30288 33405 30297 33439
rect 30297 33405 30331 33439
rect 30331 33405 30340 33439
rect 30288 33396 30340 33405
rect 30472 33396 30524 33448
rect 31208 33396 31260 33448
rect 31484 33507 31536 33516
rect 31484 33473 31493 33507
rect 31493 33473 31527 33507
rect 31527 33473 31536 33507
rect 31484 33464 31536 33473
rect 31852 33464 31904 33516
rect 32312 33464 32364 33516
rect 32036 33396 32088 33448
rect 31392 33328 31444 33380
rect 31484 33328 31536 33380
rect 33140 33328 33192 33380
rect 34152 33328 34204 33380
rect 31760 33260 31812 33312
rect 34060 33260 34112 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 4620 33056 4672 33108
rect 6092 33056 6144 33108
rect 6736 33056 6788 33108
rect 9772 33099 9824 33108
rect 9772 33065 9781 33099
rect 9781 33065 9815 33099
rect 9815 33065 9824 33099
rect 9772 33056 9824 33065
rect 11704 33056 11756 33108
rect 11796 33099 11848 33108
rect 11796 33065 11805 33099
rect 11805 33065 11839 33099
rect 11839 33065 11848 33099
rect 11796 33056 11848 33065
rect 16028 33099 16080 33108
rect 16028 33065 16037 33099
rect 16037 33065 16071 33099
rect 16071 33065 16080 33099
rect 16028 33056 16080 33065
rect 7472 32963 7524 32972
rect 7472 32929 7481 32963
rect 7481 32929 7515 32963
rect 7515 32929 7524 32963
rect 7472 32920 7524 32929
rect 5356 32852 5408 32904
rect 5816 32852 5868 32904
rect 6920 32852 6972 32904
rect 7104 32852 7156 32904
rect 7932 32827 7984 32836
rect 7932 32793 7941 32827
rect 7941 32793 7975 32827
rect 7975 32793 7984 32827
rect 7932 32784 7984 32793
rect 5724 32716 5776 32768
rect 6736 32716 6788 32768
rect 8300 32852 8352 32904
rect 10692 32920 10744 32972
rect 11520 32920 11572 32972
rect 11612 32920 11664 32972
rect 14832 32988 14884 33040
rect 15016 32988 15068 33040
rect 17500 33056 17552 33108
rect 18144 33056 18196 33108
rect 19064 33056 19116 33108
rect 19708 33056 19760 33108
rect 19984 33056 20036 33108
rect 20076 33099 20128 33108
rect 20076 33065 20085 33099
rect 20085 33065 20119 33099
rect 20119 33065 20128 33099
rect 20076 33056 20128 33065
rect 21732 33056 21784 33108
rect 23848 33056 23900 33108
rect 26516 33099 26568 33108
rect 26516 33065 26525 33099
rect 26525 33065 26559 33099
rect 26559 33065 26568 33099
rect 26516 33056 26568 33065
rect 26608 33056 26660 33108
rect 29184 33056 29236 33108
rect 29276 33056 29328 33108
rect 30012 33099 30064 33108
rect 30012 33065 30021 33099
rect 30021 33065 30055 33099
rect 30055 33065 30064 33099
rect 30012 33056 30064 33065
rect 8208 32716 8260 32768
rect 11704 32895 11756 32904
rect 11704 32861 11713 32895
rect 11713 32861 11747 32895
rect 11747 32861 11756 32895
rect 11704 32852 11756 32861
rect 10784 32716 10836 32768
rect 12716 32852 12768 32904
rect 12256 32784 12308 32836
rect 12624 32827 12676 32836
rect 12624 32793 12633 32827
rect 12633 32793 12667 32827
rect 12667 32793 12676 32827
rect 12624 32784 12676 32793
rect 10968 32716 11020 32768
rect 11980 32716 12032 32768
rect 13544 32895 13596 32904
rect 13544 32861 13553 32895
rect 13553 32861 13587 32895
rect 13587 32861 13596 32895
rect 13544 32852 13596 32861
rect 13268 32784 13320 32836
rect 15200 32852 15252 32904
rect 15476 32895 15528 32904
rect 15476 32861 15485 32895
rect 15485 32861 15519 32895
rect 15519 32861 15528 32895
rect 15476 32852 15528 32861
rect 16304 32920 16356 32972
rect 17040 32920 17092 32972
rect 14372 32716 14424 32768
rect 14464 32716 14516 32768
rect 14556 32759 14608 32768
rect 14556 32725 14565 32759
rect 14565 32725 14599 32759
rect 14599 32725 14608 32759
rect 14556 32716 14608 32725
rect 17684 32852 17736 32904
rect 17776 32895 17828 32904
rect 17776 32861 17785 32895
rect 17785 32861 17819 32895
rect 17819 32861 17828 32895
rect 17776 32852 17828 32861
rect 18144 32920 18196 32972
rect 18236 32963 18288 32972
rect 18236 32929 18245 32963
rect 18245 32929 18279 32963
rect 18279 32929 18288 32963
rect 18236 32920 18288 32929
rect 17960 32895 18012 32904
rect 17960 32861 17970 32895
rect 17970 32861 18004 32895
rect 18004 32861 18012 32895
rect 17960 32852 18012 32861
rect 18512 32852 18564 32904
rect 15936 32759 15988 32768
rect 15936 32725 15945 32759
rect 15945 32725 15979 32759
rect 15979 32725 15988 32759
rect 15936 32716 15988 32725
rect 16028 32716 16080 32768
rect 16304 32716 16356 32768
rect 16488 32759 16540 32768
rect 16488 32725 16497 32759
rect 16497 32725 16531 32759
rect 16531 32725 16540 32759
rect 16488 32716 16540 32725
rect 17408 32759 17460 32768
rect 17408 32725 17417 32759
rect 17417 32725 17451 32759
rect 17451 32725 17460 32759
rect 17408 32716 17460 32725
rect 17868 32716 17920 32768
rect 17960 32716 18012 32768
rect 18788 32895 18840 32904
rect 18788 32861 18797 32895
rect 18797 32861 18831 32895
rect 18831 32861 18840 32895
rect 18788 32852 18840 32861
rect 19432 33031 19484 33040
rect 19432 32997 19441 33031
rect 19441 32997 19475 33031
rect 19475 32997 19484 33031
rect 19432 32988 19484 32997
rect 22744 32988 22796 33040
rect 19340 32852 19392 32904
rect 19616 32895 19668 32904
rect 19616 32861 19625 32895
rect 19625 32861 19659 32895
rect 19659 32861 19668 32895
rect 19616 32852 19668 32861
rect 19248 32784 19300 32836
rect 19800 32852 19852 32904
rect 19984 32895 20036 32904
rect 19984 32861 19993 32895
rect 19993 32861 20027 32895
rect 20027 32861 20036 32895
rect 19984 32852 20036 32861
rect 21180 32920 21232 32972
rect 21732 32895 21784 32904
rect 21732 32861 21741 32895
rect 21741 32861 21775 32895
rect 21775 32861 21784 32895
rect 21732 32852 21784 32861
rect 22008 32852 22060 32904
rect 23020 32852 23072 32904
rect 26792 32988 26844 33040
rect 28172 32988 28224 33040
rect 25688 32895 25740 32904
rect 25688 32861 25697 32895
rect 25697 32861 25731 32895
rect 25731 32861 25740 32895
rect 25688 32852 25740 32861
rect 27620 32963 27672 32972
rect 27620 32929 27629 32963
rect 27629 32929 27663 32963
rect 27663 32929 27672 32963
rect 27620 32920 27672 32929
rect 29736 32988 29788 33040
rect 33048 33056 33100 33108
rect 33324 33056 33376 33108
rect 29644 32920 29696 32972
rect 31852 32988 31904 33040
rect 27160 32852 27212 32904
rect 21824 32827 21876 32836
rect 21824 32793 21833 32827
rect 21833 32793 21867 32827
rect 21867 32793 21876 32827
rect 21824 32784 21876 32793
rect 22376 32784 22428 32836
rect 26516 32784 26568 32836
rect 30104 32895 30156 32904
rect 30104 32861 30113 32895
rect 30113 32861 30147 32895
rect 30147 32861 30156 32895
rect 30104 32852 30156 32861
rect 30288 32784 30340 32836
rect 31208 32852 31260 32904
rect 31576 32895 31628 32904
rect 31576 32861 31585 32895
rect 31585 32861 31619 32895
rect 31619 32861 31628 32895
rect 31576 32852 31628 32861
rect 31944 32895 31996 32904
rect 31944 32861 31953 32895
rect 31953 32861 31987 32895
rect 31987 32861 31996 32895
rect 34152 33031 34204 33040
rect 34152 32997 34161 33031
rect 34161 32997 34195 33031
rect 34195 32997 34204 33031
rect 34152 32988 34204 32997
rect 35164 32988 35216 33040
rect 31944 32852 31996 32861
rect 33140 32852 33192 32904
rect 34060 32852 34112 32904
rect 20444 32759 20496 32768
rect 20444 32725 20453 32759
rect 20453 32725 20487 32759
rect 20487 32725 20496 32759
rect 20444 32716 20496 32725
rect 20720 32716 20772 32768
rect 21456 32716 21508 32768
rect 22284 32759 22336 32768
rect 22284 32725 22293 32759
rect 22293 32725 22327 32759
rect 22327 32725 22336 32759
rect 22284 32716 22336 32725
rect 23480 32716 23532 32768
rect 24216 32716 24268 32768
rect 24308 32716 24360 32768
rect 28816 32716 28868 32768
rect 29552 32716 29604 32768
rect 31760 32716 31812 32768
rect 32404 32827 32456 32836
rect 32404 32793 32413 32827
rect 32413 32793 32447 32827
rect 32447 32793 32456 32827
rect 32404 32784 32456 32793
rect 33692 32784 33744 32836
rect 34980 32895 35032 32904
rect 34980 32861 34989 32895
rect 34989 32861 35023 32895
rect 35023 32861 35032 32895
rect 34980 32852 35032 32861
rect 36636 32852 36688 32904
rect 38292 32852 38344 32904
rect 33600 32759 33652 32768
rect 33600 32725 33609 32759
rect 33609 32725 33643 32759
rect 33643 32725 33652 32759
rect 33600 32716 33652 32725
rect 34980 32716 35032 32768
rect 35992 32716 36044 32768
rect 37740 32759 37792 32768
rect 37740 32725 37749 32759
rect 37749 32725 37783 32759
rect 37783 32725 37792 32759
rect 37740 32716 37792 32725
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 8208 32512 8260 32564
rect 17316 32512 17368 32564
rect 18236 32512 18288 32564
rect 18788 32512 18840 32564
rect 18972 32512 19024 32564
rect 20352 32512 20404 32564
rect 20444 32555 20496 32564
rect 20444 32521 20453 32555
rect 20453 32521 20487 32555
rect 20487 32521 20496 32555
rect 20444 32512 20496 32521
rect 21824 32555 21876 32564
rect 21824 32521 21833 32555
rect 21833 32521 21867 32555
rect 21867 32521 21876 32555
rect 21824 32512 21876 32521
rect 22284 32512 22336 32564
rect 22376 32512 22428 32564
rect 8944 32444 8996 32496
rect 12348 32444 12400 32496
rect 11336 32376 11388 32428
rect 7656 32351 7708 32360
rect 7656 32317 7665 32351
rect 7665 32317 7699 32351
rect 7699 32317 7708 32351
rect 7656 32308 7708 32317
rect 7932 32308 7984 32360
rect 11612 32308 11664 32360
rect 12808 32376 12860 32428
rect 13544 32376 13596 32428
rect 17868 32376 17920 32428
rect 13268 32308 13320 32360
rect 16028 32308 16080 32360
rect 17960 32308 18012 32360
rect 18052 32308 18104 32360
rect 18604 32308 18656 32360
rect 18788 32419 18840 32428
rect 18788 32385 18797 32419
rect 18797 32385 18831 32419
rect 18831 32385 18840 32419
rect 18788 32376 18840 32385
rect 19340 32376 19392 32428
rect 19064 32308 19116 32360
rect 19156 32351 19208 32360
rect 19156 32317 19165 32351
rect 19165 32317 19199 32351
rect 19199 32317 19208 32351
rect 19156 32308 19208 32317
rect 19248 32308 19300 32360
rect 20444 32376 20496 32428
rect 20628 32419 20680 32428
rect 20628 32385 20637 32419
rect 20637 32385 20671 32419
rect 20671 32385 20680 32419
rect 20628 32376 20680 32385
rect 21456 32419 21508 32428
rect 14372 32240 14424 32292
rect 20076 32351 20128 32360
rect 20076 32317 20085 32351
rect 20085 32317 20119 32351
rect 20119 32317 20128 32351
rect 20076 32308 20128 32317
rect 21456 32385 21465 32419
rect 21465 32385 21499 32419
rect 21499 32385 21508 32419
rect 21456 32376 21508 32385
rect 22652 32487 22704 32496
rect 22652 32453 22661 32487
rect 22661 32453 22695 32487
rect 22695 32453 22704 32487
rect 22652 32444 22704 32453
rect 22284 32351 22336 32360
rect 22284 32317 22293 32351
rect 22293 32317 22327 32351
rect 22327 32317 22336 32351
rect 22284 32308 22336 32317
rect 12624 32172 12676 32224
rect 18052 32172 18104 32224
rect 18512 32172 18564 32224
rect 21180 32240 21232 32292
rect 21456 32240 21508 32292
rect 23848 32444 23900 32496
rect 23020 32376 23072 32428
rect 23204 32419 23256 32428
rect 23204 32385 23213 32419
rect 23213 32385 23247 32419
rect 23247 32385 23256 32419
rect 23204 32376 23256 32385
rect 23572 32419 23624 32428
rect 23572 32385 23581 32419
rect 23581 32385 23615 32419
rect 23615 32385 23624 32419
rect 23572 32376 23624 32385
rect 24124 32487 24176 32496
rect 24124 32453 24133 32487
rect 24133 32453 24167 32487
rect 24167 32453 24176 32487
rect 24124 32444 24176 32453
rect 29552 32512 29604 32564
rect 30012 32555 30064 32564
rect 30012 32521 30021 32555
rect 30021 32521 30055 32555
rect 30055 32521 30064 32555
rect 30012 32512 30064 32521
rect 30196 32512 30248 32564
rect 31484 32512 31536 32564
rect 23388 32308 23440 32360
rect 29184 32444 29236 32496
rect 31576 32444 31628 32496
rect 24400 32419 24452 32428
rect 24400 32385 24409 32419
rect 24409 32385 24443 32419
rect 24443 32385 24452 32419
rect 24400 32376 24452 32385
rect 23756 32240 23808 32292
rect 24584 32376 24636 32428
rect 25136 32376 25188 32428
rect 32128 32419 32180 32428
rect 32128 32385 32137 32419
rect 32137 32385 32171 32419
rect 32171 32385 32180 32419
rect 32128 32376 32180 32385
rect 32404 32376 32456 32428
rect 32864 32376 32916 32428
rect 33600 32444 33652 32496
rect 33692 32419 33744 32428
rect 33692 32385 33701 32419
rect 33701 32385 33735 32419
rect 33735 32385 33744 32419
rect 33692 32376 33744 32385
rect 22008 32172 22060 32224
rect 22468 32215 22520 32224
rect 22468 32181 22477 32215
rect 22477 32181 22511 32215
rect 22511 32181 22520 32215
rect 22468 32172 22520 32181
rect 23020 32172 23072 32224
rect 23480 32172 23532 32224
rect 23572 32172 23624 32224
rect 24124 32172 24176 32224
rect 24216 32172 24268 32224
rect 24860 32215 24912 32224
rect 24860 32181 24869 32215
rect 24869 32181 24903 32215
rect 24903 32181 24912 32215
rect 24860 32172 24912 32181
rect 26056 32240 26108 32292
rect 33416 32351 33468 32360
rect 33416 32317 33425 32351
rect 33425 32317 33459 32351
rect 33459 32317 33468 32351
rect 33416 32308 33468 32317
rect 34336 32308 34388 32360
rect 34612 32351 34664 32360
rect 34612 32317 34621 32351
rect 34621 32317 34655 32351
rect 34655 32317 34664 32351
rect 34612 32308 34664 32317
rect 34704 32351 34756 32360
rect 34704 32317 34713 32351
rect 34713 32317 34747 32351
rect 34747 32317 34756 32351
rect 34704 32308 34756 32317
rect 35348 32308 35400 32360
rect 37740 32308 37792 32360
rect 27804 32172 27856 32224
rect 29736 32172 29788 32224
rect 33324 32172 33376 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 4804 31968 4856 32020
rect 19064 31968 19116 32020
rect 20720 31968 20772 32020
rect 21824 31968 21876 32020
rect 14556 31900 14608 31952
rect 3332 31764 3384 31816
rect 4068 31832 4120 31884
rect 7012 31832 7064 31884
rect 7656 31832 7708 31884
rect 8484 31832 8536 31884
rect 12992 31832 13044 31884
rect 4160 31764 4212 31816
rect 5264 31739 5316 31748
rect 5264 31705 5273 31739
rect 5273 31705 5307 31739
rect 5307 31705 5316 31739
rect 5264 31696 5316 31705
rect 6644 31739 6696 31748
rect 6644 31705 6653 31739
rect 6653 31705 6687 31739
rect 6687 31705 6696 31739
rect 6644 31696 6696 31705
rect 5448 31628 5500 31680
rect 8668 31764 8720 31816
rect 9588 31764 9640 31816
rect 11520 31764 11572 31816
rect 11796 31807 11848 31816
rect 11796 31773 11805 31807
rect 11805 31773 11839 31807
rect 11839 31773 11848 31807
rect 11796 31764 11848 31773
rect 11980 31807 12032 31816
rect 11980 31773 11989 31807
rect 11989 31773 12023 31807
rect 12023 31773 12032 31807
rect 11980 31764 12032 31773
rect 11704 31696 11756 31748
rect 12256 31764 12308 31816
rect 12348 31764 12400 31816
rect 12532 31764 12584 31816
rect 14832 31807 14884 31816
rect 14832 31773 14841 31807
rect 14841 31773 14875 31807
rect 14875 31773 14884 31807
rect 14832 31764 14884 31773
rect 16488 31832 16540 31884
rect 19892 31900 19944 31952
rect 21732 31900 21784 31952
rect 18512 31832 18564 31884
rect 8116 31671 8168 31680
rect 8116 31637 8125 31671
rect 8125 31637 8159 31671
rect 8159 31637 8168 31671
rect 16120 31807 16172 31816
rect 16120 31773 16129 31807
rect 16129 31773 16163 31807
rect 16163 31773 16172 31807
rect 16120 31764 16172 31773
rect 16212 31807 16264 31816
rect 16212 31773 16221 31807
rect 16221 31773 16255 31807
rect 16255 31773 16264 31807
rect 16212 31764 16264 31773
rect 19064 31764 19116 31816
rect 23020 31968 23072 32020
rect 23204 31968 23256 32020
rect 22008 31832 22060 31884
rect 22744 31875 22796 31884
rect 22744 31841 22753 31875
rect 22753 31841 22787 31875
rect 22787 31841 22796 31875
rect 22744 31832 22796 31841
rect 18788 31696 18840 31748
rect 22468 31696 22520 31748
rect 24860 31968 24912 32020
rect 27160 31968 27212 32020
rect 23388 31807 23440 31816
rect 23388 31773 23397 31807
rect 23397 31773 23431 31807
rect 23431 31773 23440 31807
rect 23388 31764 23440 31773
rect 23756 31900 23808 31952
rect 8116 31628 8168 31637
rect 13820 31628 13872 31680
rect 14096 31628 14148 31680
rect 15292 31628 15344 31680
rect 15476 31628 15528 31680
rect 16396 31671 16448 31680
rect 16396 31637 16405 31671
rect 16405 31637 16439 31671
rect 16439 31637 16448 31671
rect 16396 31628 16448 31637
rect 16580 31628 16632 31680
rect 20168 31628 20220 31680
rect 22192 31671 22244 31680
rect 22192 31637 22201 31671
rect 22201 31637 22235 31671
rect 22235 31637 22244 31671
rect 22192 31628 22244 31637
rect 23756 31764 23808 31816
rect 27804 31943 27856 31952
rect 27804 31909 27813 31943
rect 27813 31909 27847 31943
rect 27847 31909 27856 31943
rect 27804 31900 27856 31909
rect 24584 31875 24636 31884
rect 24584 31841 24593 31875
rect 24593 31841 24627 31875
rect 24627 31841 24636 31875
rect 24584 31832 24636 31841
rect 29736 31832 29788 31884
rect 31576 31875 31628 31884
rect 31576 31841 31585 31875
rect 31585 31841 31619 31875
rect 31619 31841 31628 31875
rect 31576 31832 31628 31841
rect 27896 31807 27948 31816
rect 24400 31628 24452 31680
rect 25688 31628 25740 31680
rect 25780 31628 25832 31680
rect 27896 31773 27905 31807
rect 27905 31773 27939 31807
rect 27939 31773 27948 31807
rect 27896 31764 27948 31773
rect 28080 31764 28132 31816
rect 31484 31807 31536 31816
rect 31484 31773 31493 31807
rect 31493 31773 31527 31807
rect 31527 31773 31536 31807
rect 34704 31968 34756 32020
rect 32128 31900 32180 31952
rect 32312 31832 32364 31884
rect 31484 31764 31536 31773
rect 30012 31696 30064 31748
rect 34152 31875 34204 31884
rect 34152 31841 34161 31875
rect 34161 31841 34195 31875
rect 34195 31841 34204 31875
rect 34152 31832 34204 31841
rect 34336 31875 34388 31884
rect 34336 31841 34345 31875
rect 34345 31841 34379 31875
rect 34379 31841 34388 31875
rect 34336 31832 34388 31841
rect 26332 31628 26384 31680
rect 34244 31628 34296 31680
rect 34336 31628 34388 31680
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 5264 31424 5316 31476
rect 6644 31424 6696 31476
rect 7656 31424 7708 31476
rect 9220 31424 9272 31476
rect 6460 31356 6512 31408
rect 7472 31399 7524 31408
rect 7472 31365 7481 31399
rect 7481 31365 7515 31399
rect 7515 31365 7524 31399
rect 12440 31424 12492 31476
rect 7472 31356 7524 31365
rect 9864 31356 9916 31408
rect 11888 31399 11940 31408
rect 11888 31365 11897 31399
rect 11897 31365 11931 31399
rect 11931 31365 11940 31399
rect 11888 31356 11940 31365
rect 12164 31356 12216 31408
rect 3332 31331 3384 31340
rect 3332 31297 3341 31331
rect 3341 31297 3375 31331
rect 3375 31297 3384 31331
rect 3332 31288 3384 31297
rect 4160 31288 4212 31340
rect 4988 31288 5040 31340
rect 3056 31263 3108 31272
rect 3056 31229 3065 31263
rect 3065 31229 3099 31263
rect 3099 31229 3108 31263
rect 3056 31220 3108 31229
rect 3424 31263 3476 31272
rect 3424 31229 3433 31263
rect 3433 31229 3467 31263
rect 3467 31229 3476 31263
rect 3424 31220 3476 31229
rect 4620 31220 4672 31272
rect 5080 31220 5132 31272
rect 8116 31288 8168 31340
rect 9220 31288 9272 31340
rect 11152 31331 11204 31340
rect 11152 31297 11161 31331
rect 11161 31297 11195 31331
rect 11195 31297 11204 31331
rect 11152 31288 11204 31297
rect 11520 31288 11572 31340
rect 12072 31288 12124 31340
rect 12624 31424 12676 31476
rect 13544 31424 13596 31476
rect 14280 31424 14332 31476
rect 15568 31424 15620 31476
rect 12532 31331 12584 31340
rect 12532 31297 12541 31331
rect 12541 31297 12575 31331
rect 12575 31297 12584 31331
rect 12532 31288 12584 31297
rect 6920 31220 6972 31272
rect 7380 31220 7432 31272
rect 9588 31263 9640 31272
rect 9588 31229 9597 31263
rect 9597 31229 9631 31263
rect 9631 31229 9640 31263
rect 9588 31220 9640 31229
rect 4068 31127 4120 31136
rect 4068 31093 4077 31127
rect 4077 31093 4111 31127
rect 4111 31093 4120 31127
rect 4068 31084 4120 31093
rect 5264 31084 5316 31136
rect 9404 31084 9456 31136
rect 12808 31288 12860 31340
rect 12348 31152 12400 31204
rect 12716 31152 12768 31204
rect 11060 31127 11112 31136
rect 11060 31093 11069 31127
rect 11069 31093 11103 31127
rect 11103 31093 11112 31127
rect 11060 31084 11112 31093
rect 11520 31127 11572 31136
rect 11520 31093 11529 31127
rect 11529 31093 11563 31127
rect 11563 31093 11572 31127
rect 11520 31084 11572 31093
rect 13636 31331 13688 31340
rect 13636 31297 13645 31331
rect 13645 31297 13679 31331
rect 13679 31297 13688 31331
rect 13636 31288 13688 31297
rect 13728 31331 13780 31340
rect 13728 31297 13737 31331
rect 13737 31297 13771 31331
rect 13771 31297 13780 31331
rect 13728 31288 13780 31297
rect 13820 31288 13872 31340
rect 14096 31399 14148 31408
rect 14096 31365 14105 31399
rect 14105 31365 14139 31399
rect 14139 31365 14148 31399
rect 14096 31356 14148 31365
rect 13820 31152 13872 31204
rect 14556 31331 14608 31340
rect 14556 31297 14565 31331
rect 14565 31297 14599 31331
rect 14599 31297 14608 31331
rect 14556 31288 14608 31297
rect 14832 31288 14884 31340
rect 15016 31288 15068 31340
rect 14832 31195 14884 31204
rect 14832 31161 14841 31195
rect 14841 31161 14875 31195
rect 14875 31161 14884 31195
rect 14832 31152 14884 31161
rect 15844 31331 15896 31340
rect 15844 31297 15853 31331
rect 15853 31297 15887 31331
rect 15887 31297 15896 31331
rect 16396 31424 16448 31476
rect 15844 31288 15896 31297
rect 16580 31288 16632 31340
rect 16672 31288 16724 31340
rect 17040 31331 17092 31340
rect 17040 31297 17049 31331
rect 17049 31297 17083 31331
rect 17083 31297 17092 31331
rect 17040 31288 17092 31297
rect 18144 31399 18196 31408
rect 18144 31365 18153 31399
rect 18153 31365 18187 31399
rect 18187 31365 18196 31399
rect 18144 31356 18196 31365
rect 18604 31356 18656 31408
rect 19064 31467 19116 31476
rect 19064 31433 19073 31467
rect 19073 31433 19107 31467
rect 19107 31433 19116 31467
rect 19064 31424 19116 31433
rect 19340 31424 19392 31476
rect 20628 31424 20680 31476
rect 20168 31356 20220 31408
rect 16304 31263 16356 31272
rect 15292 31152 15344 31204
rect 15200 31084 15252 31136
rect 16304 31229 16313 31263
rect 16313 31229 16347 31263
rect 16347 31229 16356 31263
rect 16304 31220 16356 31229
rect 16580 31152 16632 31204
rect 15936 31127 15988 31136
rect 15936 31093 15945 31127
rect 15945 31093 15979 31127
rect 15979 31093 15988 31127
rect 15936 31084 15988 31093
rect 16028 31084 16080 31136
rect 18236 31331 18288 31340
rect 18236 31297 18245 31331
rect 18245 31297 18279 31331
rect 18279 31297 18288 31331
rect 18236 31288 18288 31297
rect 18604 31263 18656 31272
rect 18604 31229 18613 31263
rect 18613 31229 18647 31263
rect 18647 31229 18656 31263
rect 18604 31220 18656 31229
rect 19064 31288 19116 31340
rect 22192 31331 22244 31340
rect 22192 31297 22198 31331
rect 22198 31297 22244 31331
rect 19156 31152 19208 31204
rect 22192 31288 22244 31297
rect 22468 31424 22520 31476
rect 24400 31424 24452 31476
rect 26332 31424 26384 31476
rect 27620 31424 27672 31476
rect 30104 31424 30156 31476
rect 25044 31356 25096 31408
rect 24124 31331 24176 31340
rect 24124 31297 24133 31331
rect 24133 31297 24167 31331
rect 24167 31297 24176 31331
rect 24124 31288 24176 31297
rect 24492 31288 24544 31340
rect 24952 31331 25004 31340
rect 24952 31297 24961 31331
rect 24961 31297 24995 31331
rect 24995 31297 25004 31331
rect 24952 31288 25004 31297
rect 25136 31331 25188 31340
rect 25136 31297 25145 31331
rect 25145 31297 25179 31331
rect 25179 31297 25188 31331
rect 25136 31288 25188 31297
rect 25596 31356 25648 31408
rect 32312 31424 32364 31476
rect 21916 31195 21968 31204
rect 21916 31161 21925 31195
rect 21925 31161 21959 31195
rect 21959 31161 21968 31195
rect 21916 31152 21968 31161
rect 17224 31127 17276 31136
rect 17224 31093 17233 31127
rect 17233 31093 17267 31127
rect 17267 31093 17276 31127
rect 17224 31084 17276 31093
rect 17960 31084 18012 31136
rect 18604 31084 18656 31136
rect 21824 31084 21876 31136
rect 27160 31331 27212 31340
rect 27160 31297 27169 31331
rect 27169 31297 27203 31331
rect 27203 31297 27212 31331
rect 27160 31288 27212 31297
rect 28356 31331 28408 31340
rect 28356 31297 28365 31331
rect 28365 31297 28399 31331
rect 28399 31297 28408 31331
rect 28356 31288 28408 31297
rect 28540 31331 28592 31340
rect 28540 31297 28549 31331
rect 28549 31297 28583 31331
rect 28583 31297 28592 31331
rect 28540 31288 28592 31297
rect 28908 31331 28960 31340
rect 28908 31297 28917 31331
rect 28917 31297 28951 31331
rect 28951 31297 28960 31331
rect 28908 31288 28960 31297
rect 29920 31331 29972 31340
rect 29920 31297 29929 31331
rect 29929 31297 29963 31331
rect 29963 31297 29972 31331
rect 29920 31288 29972 31297
rect 30012 31288 30064 31340
rect 30196 31288 30248 31340
rect 26976 31263 27028 31272
rect 26976 31229 26985 31263
rect 26985 31229 27019 31263
rect 27019 31229 27028 31263
rect 26976 31220 27028 31229
rect 27252 31220 27304 31272
rect 28448 31220 28500 31272
rect 31484 31288 31536 31340
rect 33416 31424 33468 31476
rect 33048 31356 33100 31408
rect 31024 31263 31076 31272
rect 29092 31152 29144 31204
rect 28632 31084 28684 31136
rect 28724 31084 28776 31136
rect 31024 31229 31033 31263
rect 31033 31229 31067 31263
rect 31067 31229 31076 31263
rect 31024 31220 31076 31229
rect 31300 31220 31352 31272
rect 30380 31152 30432 31204
rect 32496 31263 32548 31272
rect 32496 31229 32505 31263
rect 32505 31229 32539 31263
rect 32539 31229 32548 31263
rect 32496 31220 32548 31229
rect 32864 31288 32916 31340
rect 33416 31331 33468 31340
rect 33416 31297 33425 31331
rect 33425 31297 33459 31331
rect 33459 31297 33468 31331
rect 33416 31288 33468 31297
rect 33600 31331 33652 31340
rect 33600 31297 33609 31331
rect 33609 31297 33643 31331
rect 33643 31297 33652 31331
rect 33600 31288 33652 31297
rect 34152 31331 34204 31340
rect 34152 31297 34161 31331
rect 34161 31297 34195 31331
rect 34195 31297 34204 31331
rect 34152 31288 34204 31297
rect 34336 31288 34388 31340
rect 35440 31424 35492 31476
rect 35992 31424 36044 31476
rect 34612 31331 34664 31340
rect 34612 31297 34621 31331
rect 34621 31297 34655 31331
rect 34655 31297 34664 31331
rect 34612 31288 34664 31297
rect 35348 31356 35400 31408
rect 34796 31331 34848 31340
rect 34796 31297 34805 31331
rect 34805 31297 34839 31331
rect 34839 31297 34848 31331
rect 34796 31288 34848 31297
rect 35440 31331 35492 31340
rect 35440 31297 35449 31331
rect 35449 31297 35483 31331
rect 35483 31297 35492 31331
rect 35440 31288 35492 31297
rect 35716 31288 35768 31340
rect 36084 31331 36136 31340
rect 36084 31297 36093 31331
rect 36093 31297 36127 31331
rect 36127 31297 36136 31331
rect 36084 31288 36136 31297
rect 36268 31331 36320 31340
rect 36268 31297 36277 31331
rect 36277 31297 36311 31331
rect 36311 31297 36320 31331
rect 36268 31288 36320 31297
rect 36360 31331 36412 31340
rect 36360 31297 36369 31331
rect 36369 31297 36403 31331
rect 36403 31297 36412 31331
rect 36360 31288 36412 31297
rect 36544 31331 36596 31340
rect 36544 31297 36553 31331
rect 36553 31297 36587 31331
rect 36587 31297 36596 31331
rect 36544 31288 36596 31297
rect 34244 31152 34296 31204
rect 32496 31084 32548 31136
rect 32956 31127 33008 31136
rect 32956 31093 32965 31127
rect 32965 31093 32999 31127
rect 32999 31093 33008 31127
rect 32956 31084 33008 31093
rect 33968 31084 34020 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 3056 30880 3108 30932
rect 3332 30719 3384 30728
rect 3332 30685 3341 30719
rect 3341 30685 3375 30719
rect 3375 30685 3384 30719
rect 3332 30676 3384 30685
rect 4068 30880 4120 30932
rect 4620 30880 4672 30932
rect 5080 30923 5132 30932
rect 5080 30889 5089 30923
rect 5089 30889 5123 30923
rect 5123 30889 5132 30923
rect 5080 30880 5132 30889
rect 9588 30880 9640 30932
rect 4528 30855 4580 30864
rect 4528 30821 4537 30855
rect 4537 30821 4571 30855
rect 4571 30821 4580 30855
rect 4528 30812 4580 30821
rect 3976 30719 4028 30728
rect 3976 30685 3983 30719
rect 3983 30685 4028 30719
rect 3976 30676 4028 30685
rect 4068 30651 4120 30660
rect 4068 30617 4077 30651
rect 4077 30617 4111 30651
rect 4111 30617 4120 30651
rect 4068 30608 4120 30617
rect 4344 30676 4396 30728
rect 7012 30787 7064 30796
rect 7012 30753 7021 30787
rect 7021 30753 7055 30787
rect 7055 30753 7064 30787
rect 7012 30744 7064 30753
rect 7380 30744 7432 30796
rect 9404 30787 9456 30796
rect 9404 30753 9413 30787
rect 9413 30753 9447 30787
rect 9447 30753 9456 30787
rect 9404 30744 9456 30753
rect 11520 30880 11572 30932
rect 11152 30812 11204 30864
rect 11796 30880 11848 30932
rect 10876 30787 10928 30796
rect 10876 30753 10885 30787
rect 10885 30753 10919 30787
rect 10919 30753 10928 30787
rect 10876 30744 10928 30753
rect 12532 30812 12584 30864
rect 4804 30676 4856 30728
rect 8668 30676 8720 30728
rect 4712 30651 4764 30660
rect 4712 30617 4721 30651
rect 4721 30617 4755 30651
rect 4755 30617 4764 30651
rect 4712 30608 4764 30617
rect 4988 30608 5040 30660
rect 6552 30651 6604 30660
rect 6552 30617 6561 30651
rect 6561 30617 6595 30651
rect 6595 30617 6604 30651
rect 6552 30608 6604 30617
rect 7288 30651 7340 30660
rect 7288 30617 7297 30651
rect 7297 30617 7331 30651
rect 7331 30617 7340 30651
rect 7288 30608 7340 30617
rect 4436 30540 4488 30592
rect 8944 30583 8996 30592
rect 8944 30549 8953 30583
rect 8953 30549 8987 30583
rect 8987 30549 8996 30583
rect 8944 30540 8996 30549
rect 9312 30583 9364 30592
rect 9312 30549 9321 30583
rect 9321 30549 9355 30583
rect 9355 30549 9364 30583
rect 9312 30540 9364 30549
rect 11060 30676 11112 30728
rect 11704 30608 11756 30660
rect 11980 30608 12032 30660
rect 12716 30719 12768 30728
rect 12716 30685 12725 30719
rect 12725 30685 12759 30719
rect 12759 30685 12768 30719
rect 12716 30676 12768 30685
rect 12808 30719 12860 30728
rect 12808 30685 12817 30719
rect 12817 30685 12851 30719
rect 12851 30685 12860 30719
rect 12808 30676 12860 30685
rect 12532 30608 12584 30660
rect 13176 30812 13228 30864
rect 13728 30880 13780 30932
rect 14280 30880 14332 30932
rect 15936 30880 15988 30932
rect 16212 30880 16264 30932
rect 18604 30923 18656 30932
rect 18604 30889 18613 30923
rect 18613 30889 18647 30923
rect 18647 30889 18656 30923
rect 18604 30880 18656 30889
rect 20076 30880 20128 30932
rect 26976 30880 27028 30932
rect 32956 30880 33008 30932
rect 34612 30880 34664 30932
rect 36360 30880 36412 30932
rect 15016 30744 15068 30796
rect 15936 30787 15988 30796
rect 15936 30753 15945 30787
rect 15945 30753 15979 30787
rect 15979 30753 15988 30787
rect 15936 30744 15988 30753
rect 16028 30744 16080 30796
rect 16120 30787 16172 30796
rect 16120 30753 16129 30787
rect 16129 30753 16163 30787
rect 16163 30753 16172 30787
rect 16120 30744 16172 30753
rect 16304 30787 16356 30796
rect 16304 30753 16313 30787
rect 16313 30753 16347 30787
rect 16347 30753 16356 30787
rect 16304 30744 16356 30753
rect 16580 30719 16632 30728
rect 16580 30685 16589 30719
rect 16589 30685 16623 30719
rect 16623 30685 16632 30719
rect 16580 30676 16632 30685
rect 17592 30812 17644 30864
rect 25228 30812 25280 30864
rect 25688 30812 25740 30864
rect 18236 30676 18288 30728
rect 19064 30744 19116 30796
rect 20076 30744 20128 30796
rect 22376 30744 22428 30796
rect 12716 30540 12768 30592
rect 13452 30583 13504 30592
rect 13452 30549 13461 30583
rect 13461 30549 13495 30583
rect 13495 30549 13504 30583
rect 13452 30540 13504 30549
rect 17960 30608 18012 30660
rect 25780 30608 25832 30660
rect 26700 30608 26752 30660
rect 27712 30719 27764 30728
rect 27712 30685 27721 30719
rect 27721 30685 27755 30719
rect 27755 30685 27764 30719
rect 27712 30676 27764 30685
rect 28172 30744 28224 30796
rect 28724 30744 28776 30796
rect 28264 30676 28316 30728
rect 28816 30676 28868 30728
rect 29092 30676 29144 30728
rect 28448 30608 28500 30660
rect 30380 30744 30432 30796
rect 32772 30744 32824 30796
rect 20168 30540 20220 30592
rect 23572 30540 23624 30592
rect 31944 30676 31996 30728
rect 34612 30744 34664 30796
rect 35716 30744 35768 30796
rect 35992 30787 36044 30796
rect 35992 30753 36001 30787
rect 36001 30753 36035 30787
rect 36035 30753 36044 30787
rect 35992 30744 36044 30753
rect 35440 30676 35492 30728
rect 36084 30676 36136 30728
rect 33508 30608 33560 30660
rect 34060 30608 34112 30660
rect 34336 30608 34388 30660
rect 30932 30540 30984 30592
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 4068 30336 4120 30388
rect 4436 30379 4488 30388
rect 4436 30345 4445 30379
rect 4445 30345 4479 30379
rect 4479 30345 4488 30379
rect 4436 30336 4488 30345
rect 4528 30336 4580 30388
rect 7288 30336 7340 30388
rect 8944 30336 8996 30388
rect 13452 30336 13504 30388
rect 5264 30268 5316 30320
rect 3332 30200 3384 30252
rect 3424 30243 3476 30252
rect 3424 30209 3433 30243
rect 3433 30209 3467 30243
rect 3467 30209 3476 30243
rect 3424 30200 3476 30209
rect 3516 30243 3568 30252
rect 3516 30209 3525 30243
rect 3525 30209 3559 30243
rect 3559 30209 3568 30243
rect 3516 30200 3568 30209
rect 3608 30175 3660 30184
rect 3608 30141 3617 30175
rect 3617 30141 3651 30175
rect 3651 30141 3660 30175
rect 3608 30132 3660 30141
rect 4620 30243 4672 30252
rect 4620 30209 4629 30243
rect 4629 30209 4663 30243
rect 4663 30209 4672 30243
rect 4620 30200 4672 30209
rect 4988 30132 5040 30184
rect 4712 30064 4764 30116
rect 4804 30064 4856 30116
rect 5448 30200 5500 30252
rect 13268 30243 13320 30252
rect 13268 30209 13277 30243
rect 13277 30209 13311 30243
rect 13311 30209 13320 30243
rect 13268 30200 13320 30209
rect 13544 30268 13596 30320
rect 6552 30132 6604 30184
rect 13820 30200 13872 30252
rect 14096 30200 14148 30252
rect 17684 30268 17736 30320
rect 20996 30268 21048 30320
rect 21916 30268 21968 30320
rect 22744 30268 22796 30320
rect 23388 30268 23440 30320
rect 19616 30200 19668 30252
rect 20076 30200 20128 30252
rect 3976 29996 4028 30048
rect 4344 29996 4396 30048
rect 13728 30064 13780 30116
rect 19892 30064 19944 30116
rect 4988 29996 5040 30048
rect 10600 29996 10652 30048
rect 12624 29996 12676 30048
rect 13636 29996 13688 30048
rect 15660 29996 15712 30048
rect 23480 30200 23532 30252
rect 23756 30243 23808 30252
rect 23756 30209 23765 30243
rect 23765 30209 23799 30243
rect 23799 30209 23808 30243
rect 23756 30200 23808 30209
rect 23572 30132 23624 30184
rect 23848 30175 23900 30184
rect 23848 30141 23857 30175
rect 23857 30141 23891 30175
rect 23891 30141 23900 30175
rect 23848 30132 23900 30141
rect 23480 30107 23532 30116
rect 23480 30073 23489 30107
rect 23489 30073 23523 30107
rect 23523 30073 23532 30107
rect 23480 30064 23532 30073
rect 28080 30336 28132 30388
rect 28540 30336 28592 30388
rect 28632 30336 28684 30388
rect 37556 30336 37608 30388
rect 27712 30268 27764 30320
rect 24860 30200 24912 30252
rect 26424 30200 26476 30252
rect 28172 30268 28224 30320
rect 30196 30268 30248 30320
rect 28264 30243 28316 30252
rect 28264 30209 28273 30243
rect 28273 30209 28307 30243
rect 28307 30209 28316 30243
rect 28264 30200 28316 30209
rect 29644 30132 29696 30184
rect 29920 30200 29972 30252
rect 30380 30200 30432 30252
rect 31392 30268 31444 30320
rect 34612 30268 34664 30320
rect 32772 30243 32824 30252
rect 32772 30209 32781 30243
rect 32781 30209 32815 30243
rect 32815 30209 32824 30243
rect 32772 30200 32824 30209
rect 30932 30175 30984 30184
rect 30932 30141 30941 30175
rect 30941 30141 30975 30175
rect 30975 30141 30984 30175
rect 30932 30132 30984 30141
rect 32680 30175 32732 30184
rect 32680 30141 32689 30175
rect 32689 30141 32723 30175
rect 32723 30141 32732 30175
rect 32680 30132 32732 30141
rect 20352 30039 20404 30048
rect 20352 30005 20361 30039
rect 20361 30005 20395 30039
rect 20395 30005 20404 30039
rect 20352 29996 20404 30005
rect 20720 30039 20772 30048
rect 20720 30005 20729 30039
rect 20729 30005 20763 30039
rect 20763 30005 20772 30039
rect 20720 29996 20772 30005
rect 24032 29996 24084 30048
rect 24124 29996 24176 30048
rect 28172 29996 28224 30048
rect 29460 29996 29512 30048
rect 29644 29996 29696 30048
rect 29920 29996 29972 30048
rect 37188 29996 37240 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 1768 29656 1820 29708
rect 12808 29792 12860 29844
rect 3608 29724 3660 29776
rect 4804 29724 4856 29776
rect 4988 29724 5040 29776
rect 2688 29588 2740 29640
rect 2780 29588 2832 29640
rect 4528 29588 4580 29640
rect 8024 29656 8076 29708
rect 12072 29724 12124 29776
rect 12348 29724 12400 29776
rect 12716 29724 12768 29776
rect 15108 29724 15160 29776
rect 10692 29699 10744 29708
rect 10692 29665 10701 29699
rect 10701 29665 10735 29699
rect 10735 29665 10744 29699
rect 10692 29656 10744 29665
rect 10876 29656 10928 29708
rect 1676 29563 1728 29572
rect 1676 29529 1685 29563
rect 1685 29529 1719 29563
rect 1719 29529 1728 29563
rect 1676 29520 1728 29529
rect 4344 29520 4396 29572
rect 4712 29520 4764 29572
rect 11152 29588 11204 29640
rect 7288 29563 7340 29572
rect 7288 29529 7297 29563
rect 7297 29529 7331 29563
rect 7331 29529 7340 29563
rect 7288 29520 7340 29529
rect 10876 29520 10928 29572
rect 12716 29520 12768 29572
rect 13176 29656 13228 29708
rect 13360 29656 13412 29708
rect 13728 29656 13780 29708
rect 15844 29724 15896 29776
rect 18144 29724 18196 29776
rect 15660 29656 15712 29708
rect 15936 29656 15988 29708
rect 16120 29699 16172 29708
rect 16120 29665 16129 29699
rect 16129 29665 16163 29699
rect 16163 29665 16172 29699
rect 16120 29656 16172 29665
rect 20352 29792 20404 29844
rect 12900 29588 12952 29640
rect 13268 29588 13320 29640
rect 14188 29520 14240 29572
rect 8300 29452 8352 29504
rect 8760 29495 8812 29504
rect 8760 29461 8769 29495
rect 8769 29461 8803 29495
rect 8803 29461 8812 29495
rect 8760 29452 8812 29461
rect 9680 29495 9732 29504
rect 9680 29461 9689 29495
rect 9689 29461 9723 29495
rect 9723 29461 9732 29495
rect 9680 29452 9732 29461
rect 11520 29452 11572 29504
rect 11796 29495 11848 29504
rect 11796 29461 11805 29495
rect 11805 29461 11839 29495
rect 11839 29461 11848 29495
rect 11796 29452 11848 29461
rect 12900 29452 12952 29504
rect 13452 29495 13504 29504
rect 13452 29461 13461 29495
rect 13461 29461 13495 29495
rect 13495 29461 13504 29495
rect 13452 29452 13504 29461
rect 15844 29588 15896 29640
rect 17224 29588 17276 29640
rect 20444 29631 20496 29640
rect 20444 29597 20453 29631
rect 20453 29597 20487 29631
rect 20487 29597 20496 29631
rect 20444 29588 20496 29597
rect 20720 29792 20772 29844
rect 23388 29792 23440 29844
rect 24032 29792 24084 29844
rect 26608 29792 26660 29844
rect 27160 29792 27212 29844
rect 20904 29724 20956 29776
rect 22192 29724 22244 29776
rect 26056 29724 26108 29776
rect 28540 29724 28592 29776
rect 28908 29724 28960 29776
rect 31024 29835 31076 29844
rect 31024 29801 31033 29835
rect 31033 29801 31067 29835
rect 31067 29801 31076 29835
rect 31024 29792 31076 29801
rect 34796 29792 34848 29844
rect 15568 29452 15620 29504
rect 16212 29452 16264 29504
rect 20996 29588 21048 29640
rect 21180 29631 21232 29640
rect 21180 29597 21189 29631
rect 21189 29597 21223 29631
rect 21223 29597 21232 29631
rect 21180 29588 21232 29597
rect 21272 29563 21324 29572
rect 21272 29529 21281 29563
rect 21281 29529 21315 29563
rect 21315 29529 21324 29563
rect 21272 29520 21324 29529
rect 23480 29631 23532 29640
rect 23480 29597 23489 29631
rect 23489 29597 23523 29631
rect 23523 29597 23532 29631
rect 23480 29588 23532 29597
rect 23756 29631 23808 29640
rect 23756 29597 23765 29631
rect 23765 29597 23799 29631
rect 23799 29597 23808 29631
rect 23756 29588 23808 29597
rect 24584 29631 24636 29640
rect 24584 29597 24586 29631
rect 24586 29597 24620 29631
rect 24620 29597 24636 29631
rect 24584 29588 24636 29597
rect 26424 29631 26476 29640
rect 26424 29597 26433 29631
rect 26433 29597 26467 29631
rect 26467 29597 26476 29631
rect 26424 29588 26476 29597
rect 26608 29631 26660 29640
rect 26608 29597 26617 29631
rect 26617 29597 26651 29631
rect 26651 29597 26660 29631
rect 26608 29588 26660 29597
rect 26976 29631 27028 29640
rect 26976 29597 26985 29631
rect 26985 29597 27019 29631
rect 27019 29597 27028 29631
rect 26976 29588 27028 29597
rect 28080 29631 28132 29640
rect 28816 29699 28868 29708
rect 28816 29665 28831 29699
rect 28831 29665 28865 29699
rect 28865 29665 28868 29699
rect 28816 29656 28868 29665
rect 31668 29656 31720 29708
rect 28080 29597 28112 29631
rect 28112 29597 28132 29631
rect 28080 29588 28132 29597
rect 28540 29631 28592 29640
rect 28540 29597 28549 29631
rect 28549 29597 28583 29631
rect 28583 29597 28592 29631
rect 28540 29588 28592 29597
rect 28724 29631 28776 29640
rect 28724 29597 28733 29631
rect 28733 29597 28767 29631
rect 28767 29597 28776 29631
rect 28724 29588 28776 29597
rect 28908 29631 28960 29640
rect 28908 29597 28917 29631
rect 28917 29597 28951 29631
rect 28951 29597 28960 29631
rect 28908 29588 28960 29597
rect 30380 29588 30432 29640
rect 30840 29631 30892 29640
rect 30840 29597 30849 29631
rect 30849 29597 30883 29631
rect 30883 29597 30892 29631
rect 30840 29588 30892 29597
rect 20996 29495 21048 29504
rect 20996 29461 21005 29495
rect 21005 29461 21039 29495
rect 21039 29461 21048 29495
rect 20996 29452 21048 29461
rect 21456 29452 21508 29504
rect 23848 29452 23900 29504
rect 24768 29452 24820 29504
rect 26240 29495 26292 29504
rect 26240 29461 26249 29495
rect 26249 29461 26283 29495
rect 26283 29461 26292 29495
rect 26240 29452 26292 29461
rect 27344 29452 27396 29504
rect 28080 29452 28132 29504
rect 30012 29520 30064 29572
rect 32036 29631 32088 29640
rect 32036 29597 32045 29631
rect 32045 29597 32079 29631
rect 32079 29597 32088 29631
rect 32036 29588 32088 29597
rect 33784 29631 33836 29640
rect 33784 29597 33793 29631
rect 33793 29597 33827 29631
rect 33827 29597 33836 29631
rect 33784 29588 33836 29597
rect 33968 29631 34020 29640
rect 33968 29597 33977 29631
rect 33977 29597 34011 29631
rect 34011 29597 34020 29631
rect 33968 29588 34020 29597
rect 34336 29724 34388 29776
rect 36452 29699 36504 29708
rect 36452 29665 36461 29699
rect 36461 29665 36495 29699
rect 36495 29665 36504 29699
rect 36452 29656 36504 29665
rect 31484 29520 31536 29572
rect 34428 29588 34480 29640
rect 36360 29631 36412 29640
rect 36360 29597 36369 29631
rect 36369 29597 36403 29631
rect 36403 29597 36412 29631
rect 36360 29588 36412 29597
rect 37188 29631 37240 29640
rect 37188 29597 37197 29631
rect 37197 29597 37231 29631
rect 37231 29597 37240 29631
rect 37188 29588 37240 29597
rect 31944 29452 31996 29504
rect 32772 29452 32824 29504
rect 34980 29452 35032 29504
rect 36820 29495 36872 29504
rect 36820 29461 36829 29495
rect 36829 29461 36863 29495
rect 36863 29461 36872 29495
rect 36820 29452 36872 29461
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 1676 29248 1728 29300
rect 3976 29248 4028 29300
rect 4528 29248 4580 29300
rect 5080 29248 5132 29300
rect 7288 29248 7340 29300
rect 4344 29087 4396 29096
rect 4344 29053 4353 29087
rect 4353 29053 4387 29087
rect 4387 29053 4396 29087
rect 4344 29044 4396 29053
rect 4804 29155 4856 29164
rect 4804 29121 4837 29155
rect 4837 29121 4856 29155
rect 4804 29112 4856 29121
rect 4988 29155 5040 29164
rect 4988 29121 4997 29155
rect 4997 29121 5031 29155
rect 5031 29121 5040 29155
rect 4988 29112 5040 29121
rect 8760 29180 8812 29232
rect 9680 29180 9732 29232
rect 9864 29180 9916 29232
rect 5264 29155 5316 29164
rect 5264 29121 5273 29155
rect 5273 29121 5307 29155
rect 5307 29121 5316 29155
rect 5264 29112 5316 29121
rect 6828 29112 6880 29164
rect 6920 29044 6972 29096
rect 7288 29087 7340 29096
rect 7288 29053 7297 29087
rect 7297 29053 7331 29087
rect 7331 29053 7340 29087
rect 7288 29044 7340 29053
rect 4620 28976 4672 29028
rect 4988 29019 5040 29028
rect 4988 28985 4997 29019
rect 4997 28985 5031 29019
rect 5031 28985 5040 29019
rect 4988 28976 5040 28985
rect 8024 29044 8076 29096
rect 10876 29291 10928 29300
rect 10876 29257 10885 29291
rect 10885 29257 10919 29291
rect 10919 29257 10928 29291
rect 10876 29248 10928 29257
rect 11520 29291 11572 29300
rect 11520 29257 11529 29291
rect 11529 29257 11563 29291
rect 11563 29257 11572 29291
rect 11520 29248 11572 29257
rect 11796 29248 11848 29300
rect 12164 29248 12216 29300
rect 11152 29155 11204 29164
rect 11152 29121 11161 29155
rect 11161 29121 11195 29155
rect 11195 29121 11204 29155
rect 11152 29112 11204 29121
rect 11888 29223 11940 29232
rect 11888 29189 11897 29223
rect 11897 29189 11931 29223
rect 11931 29189 11940 29223
rect 11888 29180 11940 29189
rect 12256 29180 12308 29232
rect 12348 29180 12400 29232
rect 11796 29155 11848 29164
rect 11796 29121 11805 29155
rect 11805 29121 11839 29155
rect 11839 29121 11848 29155
rect 11796 29112 11848 29121
rect 12808 29248 12860 29300
rect 13452 29248 13504 29300
rect 14188 29248 14240 29300
rect 15936 29248 15988 29300
rect 13360 29180 13412 29232
rect 13360 29044 13412 29096
rect 13820 29044 13872 29096
rect 20904 29180 20956 29232
rect 15936 29155 15988 29164
rect 15936 29121 15945 29155
rect 15945 29121 15979 29155
rect 15979 29121 15988 29155
rect 15936 29112 15988 29121
rect 16120 29155 16172 29164
rect 16120 29121 16129 29155
rect 16129 29121 16163 29155
rect 16163 29121 16172 29155
rect 16120 29112 16172 29121
rect 17868 29155 17920 29164
rect 17868 29121 17877 29155
rect 17877 29121 17911 29155
rect 17911 29121 17920 29155
rect 17868 29112 17920 29121
rect 17960 29155 18012 29164
rect 17960 29121 17969 29155
rect 17969 29121 18003 29155
rect 18003 29121 18012 29155
rect 17960 29112 18012 29121
rect 18144 29155 18196 29164
rect 18144 29121 18153 29155
rect 18153 29121 18187 29155
rect 18187 29121 18196 29155
rect 18144 29112 18196 29121
rect 19524 29112 19576 29164
rect 21272 29223 21324 29232
rect 21272 29189 21281 29223
rect 21281 29189 21315 29223
rect 21315 29189 21324 29223
rect 21272 29180 21324 29189
rect 21456 29223 21508 29232
rect 21456 29189 21481 29223
rect 21481 29189 21508 29223
rect 21456 29180 21508 29189
rect 21732 29112 21784 29164
rect 26056 29248 26108 29300
rect 26792 29248 26844 29300
rect 27528 29248 27580 29300
rect 27896 29248 27948 29300
rect 28264 29291 28316 29300
rect 28264 29257 28273 29291
rect 28273 29257 28307 29291
rect 28307 29257 28316 29291
rect 28264 29248 28316 29257
rect 26424 29180 26476 29232
rect 21916 29087 21968 29096
rect 21916 29053 21925 29087
rect 21925 29053 21959 29087
rect 21959 29053 21968 29087
rect 21916 29044 21968 29053
rect 12256 28976 12308 29028
rect 12808 28976 12860 29028
rect 15108 28976 15160 29028
rect 17132 28976 17184 29028
rect 19432 28976 19484 29028
rect 19892 28976 19944 29028
rect 20812 28976 20864 29028
rect 20996 28976 21048 29028
rect 22100 28976 22152 29028
rect 23388 28976 23440 29028
rect 24124 29044 24176 29096
rect 26148 29112 26200 29164
rect 26240 29044 26292 29096
rect 26884 29112 26936 29164
rect 27528 29155 27580 29164
rect 27528 29121 27537 29155
rect 27537 29121 27571 29155
rect 27571 29121 27580 29155
rect 27528 29112 27580 29121
rect 27620 29112 27672 29164
rect 28632 29112 28684 29164
rect 29000 29155 29052 29164
rect 29000 29121 29009 29155
rect 29009 29121 29043 29155
rect 29043 29121 29052 29155
rect 29000 29112 29052 29121
rect 29644 29112 29696 29164
rect 30012 29155 30064 29164
rect 30012 29121 30021 29155
rect 30021 29121 30055 29155
rect 30055 29121 30064 29155
rect 30012 29112 30064 29121
rect 30104 29155 30156 29164
rect 30104 29121 30113 29155
rect 30113 29121 30147 29155
rect 30147 29121 30156 29155
rect 30104 29112 30156 29121
rect 31944 29112 31996 29164
rect 33048 29248 33100 29300
rect 36360 29248 36412 29300
rect 4712 28951 4764 28960
rect 4712 28917 4721 28951
rect 4721 28917 4755 28951
rect 4755 28917 4764 28951
rect 4712 28908 4764 28917
rect 6184 28908 6236 28960
rect 18512 28951 18564 28960
rect 18512 28917 18521 28951
rect 18521 28917 18555 28951
rect 18555 28917 18564 28951
rect 18512 28908 18564 28917
rect 21272 28908 21324 28960
rect 22284 28951 22336 28960
rect 22284 28917 22293 28951
rect 22293 28917 22327 28951
rect 22327 28917 22336 28951
rect 22284 28908 22336 28917
rect 25412 28908 25464 28960
rect 27528 28976 27580 29028
rect 28264 28976 28316 29028
rect 28540 28976 28592 29028
rect 31668 29044 31720 29096
rect 31024 28976 31076 29028
rect 33140 29155 33192 29164
rect 33140 29121 33149 29155
rect 33149 29121 33183 29155
rect 33183 29121 33192 29155
rect 33140 29112 33192 29121
rect 34980 29223 35032 29232
rect 33508 29155 33560 29164
rect 33508 29121 33517 29155
rect 33517 29121 33551 29155
rect 33551 29121 33560 29155
rect 33508 29112 33560 29121
rect 34152 29155 34204 29164
rect 34152 29121 34161 29155
rect 34161 29121 34195 29155
rect 34195 29121 34204 29155
rect 34152 29112 34204 29121
rect 34980 29189 34989 29223
rect 34989 29189 35023 29223
rect 35023 29189 35032 29223
rect 34980 29180 35032 29189
rect 34428 29112 34480 29164
rect 34796 29112 34848 29164
rect 35164 29155 35216 29164
rect 35164 29121 35173 29155
rect 35173 29121 35207 29155
rect 35207 29121 35216 29155
rect 35164 29112 35216 29121
rect 35532 29112 35584 29164
rect 34336 29087 34388 29096
rect 34336 29053 34345 29087
rect 34345 29053 34379 29087
rect 34379 29053 34388 29087
rect 34336 29044 34388 29053
rect 35992 29112 36044 29164
rect 36176 29155 36228 29164
rect 36176 29121 36185 29155
rect 36185 29121 36219 29155
rect 36219 29121 36228 29155
rect 36176 29112 36228 29121
rect 36360 29155 36412 29164
rect 36360 29121 36369 29155
rect 36369 29121 36403 29155
rect 36403 29121 36412 29155
rect 36360 29112 36412 29121
rect 36728 29044 36780 29096
rect 35440 28976 35492 29028
rect 28080 28908 28132 28960
rect 28816 28908 28868 28960
rect 32036 28908 32088 28960
rect 34428 28908 34480 28960
rect 35808 28908 35860 28960
rect 36728 28908 36780 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 3516 28704 3568 28756
rect 1768 28568 1820 28620
rect 2136 28568 2188 28620
rect 4620 28747 4672 28756
rect 4620 28713 4629 28747
rect 4629 28713 4663 28747
rect 4663 28713 4672 28747
rect 4620 28704 4672 28713
rect 5264 28747 5316 28756
rect 5264 28713 5273 28747
rect 5273 28713 5307 28747
rect 5307 28713 5316 28747
rect 5264 28704 5316 28713
rect 6828 28747 6880 28756
rect 6828 28713 6837 28747
rect 6837 28713 6871 28747
rect 6871 28713 6880 28747
rect 6828 28704 6880 28713
rect 16120 28704 16172 28756
rect 21732 28704 21784 28756
rect 22192 28747 22244 28756
rect 22192 28713 22201 28747
rect 22201 28713 22235 28747
rect 22235 28713 22244 28747
rect 22192 28704 22244 28713
rect 24860 28704 24912 28756
rect 26148 28704 26200 28756
rect 27436 28704 27488 28756
rect 28172 28704 28224 28756
rect 28816 28704 28868 28756
rect 29092 28704 29144 28756
rect 4988 28500 5040 28552
rect 2780 28432 2832 28484
rect 5540 28543 5592 28552
rect 5540 28509 5549 28543
rect 5549 28509 5583 28543
rect 5583 28509 5592 28543
rect 5540 28500 5592 28509
rect 5816 28432 5868 28484
rect 6092 28543 6144 28552
rect 6092 28509 6101 28543
rect 6101 28509 6135 28543
rect 6135 28509 6144 28543
rect 6092 28500 6144 28509
rect 6184 28500 6236 28552
rect 6828 28568 6880 28620
rect 17224 28636 17276 28688
rect 6368 28500 6420 28552
rect 7380 28500 7432 28552
rect 12716 28500 12768 28552
rect 15108 28500 15160 28552
rect 17316 28611 17368 28620
rect 17316 28577 17325 28611
rect 17325 28577 17359 28611
rect 17359 28577 17368 28611
rect 17316 28568 17368 28577
rect 6736 28432 6788 28484
rect 12900 28432 12952 28484
rect 17132 28500 17184 28552
rect 18052 28636 18104 28688
rect 17776 28611 17828 28620
rect 17776 28577 17785 28611
rect 17785 28577 17819 28611
rect 17819 28577 17828 28611
rect 17776 28568 17828 28577
rect 19800 28636 19852 28688
rect 22100 28636 22152 28688
rect 23480 28636 23532 28688
rect 24952 28636 25004 28688
rect 18512 28543 18564 28552
rect 18512 28509 18521 28543
rect 18521 28509 18555 28543
rect 18555 28509 18564 28543
rect 18512 28500 18564 28509
rect 18972 28432 19024 28484
rect 19064 28432 19116 28484
rect 19800 28543 19852 28552
rect 19800 28509 19809 28543
rect 19809 28509 19843 28543
rect 19843 28509 19852 28543
rect 19800 28500 19852 28509
rect 19892 28543 19944 28552
rect 19892 28509 19901 28543
rect 19901 28509 19935 28543
rect 19935 28509 19944 28543
rect 19892 28500 19944 28509
rect 19984 28500 20036 28552
rect 22284 28568 22336 28620
rect 5632 28364 5684 28416
rect 6460 28407 6512 28416
rect 6460 28373 6469 28407
rect 6469 28373 6503 28407
rect 6503 28373 6512 28407
rect 6460 28364 6512 28373
rect 13176 28407 13228 28416
rect 13176 28373 13185 28407
rect 13185 28373 13219 28407
rect 13219 28373 13228 28407
rect 13176 28364 13228 28373
rect 15384 28407 15436 28416
rect 15384 28373 15393 28407
rect 15393 28373 15427 28407
rect 15427 28373 15436 28407
rect 15384 28364 15436 28373
rect 17960 28364 18012 28416
rect 19248 28407 19300 28416
rect 19248 28373 19257 28407
rect 19257 28373 19291 28407
rect 19291 28373 19300 28407
rect 19248 28364 19300 28373
rect 23848 28500 23900 28552
rect 24768 28543 24820 28552
rect 24768 28509 24777 28543
rect 24777 28509 24811 28543
rect 24811 28509 24820 28543
rect 24768 28500 24820 28509
rect 30104 28568 30156 28620
rect 30840 28611 30892 28620
rect 30840 28577 30849 28611
rect 30849 28577 30883 28611
rect 30883 28577 30892 28611
rect 30840 28568 30892 28577
rect 31576 28704 31628 28756
rect 32036 28704 32088 28756
rect 32496 28704 32548 28756
rect 33048 28747 33100 28756
rect 33048 28713 33057 28747
rect 33057 28713 33091 28747
rect 33091 28713 33100 28747
rect 33048 28704 33100 28713
rect 35624 28747 35676 28756
rect 35624 28713 35633 28747
rect 35633 28713 35667 28747
rect 35667 28713 35676 28747
rect 35624 28704 35676 28713
rect 36268 28704 36320 28756
rect 36360 28704 36412 28756
rect 36728 28704 36780 28756
rect 33140 28636 33192 28688
rect 35440 28679 35492 28688
rect 35440 28645 35449 28679
rect 35449 28645 35483 28679
rect 35483 28645 35492 28679
rect 35440 28636 35492 28645
rect 35532 28636 35584 28688
rect 22192 28432 22244 28484
rect 23020 28432 23072 28484
rect 26700 28543 26752 28552
rect 26700 28509 26709 28543
rect 26709 28509 26743 28543
rect 26743 28509 26752 28543
rect 26700 28500 26752 28509
rect 26792 28543 26844 28552
rect 26792 28509 26801 28543
rect 26801 28509 26835 28543
rect 26835 28509 26844 28543
rect 26792 28500 26844 28509
rect 26976 28543 27028 28552
rect 26976 28509 26985 28543
rect 26985 28509 27019 28543
rect 27019 28509 27028 28543
rect 26976 28500 27028 28509
rect 27804 28500 27856 28552
rect 28448 28500 28500 28552
rect 29736 28543 29788 28552
rect 29736 28509 29745 28543
rect 29745 28509 29779 28543
rect 29779 28509 29788 28543
rect 29736 28500 29788 28509
rect 30656 28500 30708 28552
rect 30748 28543 30800 28552
rect 30748 28509 30757 28543
rect 30757 28509 30791 28543
rect 30791 28509 30800 28543
rect 30748 28500 30800 28509
rect 31116 28543 31168 28552
rect 31116 28509 31125 28543
rect 31125 28509 31159 28543
rect 31159 28509 31168 28543
rect 31116 28500 31168 28509
rect 32772 28568 32824 28620
rect 36268 28568 36320 28620
rect 36728 28611 36780 28620
rect 36728 28577 36737 28611
rect 36737 28577 36771 28611
rect 36771 28577 36780 28611
rect 36728 28568 36780 28577
rect 20352 28364 20404 28416
rect 22468 28407 22520 28416
rect 22468 28373 22477 28407
rect 22477 28373 22511 28407
rect 22511 28373 22520 28407
rect 22468 28364 22520 28373
rect 22836 28407 22888 28416
rect 22836 28373 22845 28407
rect 22845 28373 22879 28407
rect 22879 28373 22888 28407
rect 22836 28364 22888 28373
rect 24400 28407 24452 28416
rect 24400 28373 24409 28407
rect 24409 28373 24443 28407
rect 24443 28373 24452 28407
rect 24400 28364 24452 28373
rect 26056 28364 26108 28416
rect 28632 28364 28684 28416
rect 30932 28364 30984 28416
rect 32496 28500 32548 28552
rect 33048 28543 33100 28552
rect 33048 28509 33057 28543
rect 33057 28509 33091 28543
rect 33091 28509 33100 28543
rect 33048 28500 33100 28509
rect 35808 28500 35860 28552
rect 35900 28543 35952 28552
rect 35900 28509 35909 28543
rect 35909 28509 35943 28543
rect 35943 28509 35952 28543
rect 35900 28500 35952 28509
rect 35992 28543 36044 28552
rect 35992 28509 36001 28543
rect 36001 28509 36035 28543
rect 36035 28509 36044 28543
rect 35992 28500 36044 28509
rect 33324 28432 33376 28484
rect 34428 28432 34480 28484
rect 35256 28432 35308 28484
rect 35624 28432 35676 28484
rect 37096 28500 37148 28552
rect 35900 28364 35952 28416
rect 36452 28364 36504 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 5816 28160 5868 28212
rect 9036 28160 9088 28212
rect 12624 28160 12676 28212
rect 13176 28160 13228 28212
rect 15384 28160 15436 28212
rect 15936 28160 15988 28212
rect 17776 28160 17828 28212
rect 17868 28160 17920 28212
rect 4712 28135 4764 28144
rect 4712 28101 4721 28135
rect 4721 28101 4755 28135
rect 4755 28101 4764 28135
rect 4712 28092 4764 28101
rect 8300 28092 8352 28144
rect 8576 28092 8628 28144
rect 2688 28024 2740 28076
rect 1768 27863 1820 27872
rect 1768 27829 1777 27863
rect 1777 27829 1811 27863
rect 1811 27829 1820 27863
rect 1768 27820 1820 27829
rect 5264 27820 5316 27872
rect 6092 27820 6144 27872
rect 7380 28024 7432 28076
rect 11704 28067 11756 28076
rect 11704 28033 11713 28067
rect 11713 28033 11747 28067
rect 11747 28033 11756 28067
rect 11704 28024 11756 28033
rect 8024 27999 8076 28008
rect 8024 27965 8033 27999
rect 8033 27965 8067 27999
rect 8067 27965 8076 27999
rect 8024 27956 8076 27965
rect 8300 27999 8352 28008
rect 8300 27965 8309 27999
rect 8309 27965 8343 27999
rect 8343 27965 8352 27999
rect 8300 27956 8352 27965
rect 8944 27956 8996 28008
rect 6828 27820 6880 27872
rect 9588 27820 9640 27872
rect 9772 27863 9824 27872
rect 9772 27829 9781 27863
rect 9781 27829 9815 27863
rect 9815 27829 9824 27863
rect 9772 27820 9824 27829
rect 11796 27999 11848 28008
rect 11796 27965 11805 27999
rect 11805 27965 11839 27999
rect 11839 27965 11848 27999
rect 11796 27956 11848 27965
rect 13636 28067 13688 28076
rect 13636 28033 13645 28067
rect 13645 28033 13679 28067
rect 13679 28033 13688 28067
rect 13636 28024 13688 28033
rect 13820 28024 13872 28076
rect 14464 28024 14516 28076
rect 19064 28160 19116 28212
rect 19248 28160 19300 28212
rect 19892 28203 19944 28212
rect 19892 28169 19901 28203
rect 19901 28169 19935 28203
rect 19935 28169 19944 28203
rect 19892 28160 19944 28169
rect 16120 28024 16172 28076
rect 17960 28024 18012 28076
rect 18512 28024 18564 28076
rect 24308 28160 24360 28212
rect 24400 28160 24452 28212
rect 27344 28160 27396 28212
rect 30748 28160 30800 28212
rect 31116 28160 31168 28212
rect 33784 28160 33836 28212
rect 34152 28160 34204 28212
rect 35992 28160 36044 28212
rect 15016 27956 15068 28008
rect 17132 27999 17184 28008
rect 17132 27965 17141 27999
rect 17141 27965 17175 27999
rect 17175 27965 17184 27999
rect 17132 27956 17184 27965
rect 18972 27956 19024 28008
rect 12532 27888 12584 27940
rect 18144 27888 18196 27940
rect 19340 27931 19392 27940
rect 19340 27897 19349 27931
rect 19349 27897 19383 27931
rect 19383 27897 19392 27931
rect 19340 27888 19392 27897
rect 19892 28024 19944 28076
rect 22284 28024 22336 28076
rect 22836 28067 22888 28076
rect 22836 28033 22848 28067
rect 22848 28033 22882 28067
rect 22882 28033 22888 28067
rect 22836 28024 22888 28033
rect 19984 27956 20036 28008
rect 22468 27956 22520 28008
rect 27252 28092 27304 28144
rect 24860 28067 24912 28076
rect 24860 28033 24869 28067
rect 24869 28033 24903 28067
rect 24903 28033 24912 28067
rect 24860 28024 24912 28033
rect 24952 28024 25004 28076
rect 25596 28067 25648 28076
rect 25596 28033 25605 28067
rect 25605 28033 25639 28067
rect 25639 28033 25648 28067
rect 25596 28024 25648 28033
rect 25872 28067 25924 28076
rect 25872 28033 25881 28067
rect 25881 28033 25915 28067
rect 25915 28033 25924 28067
rect 25872 28024 25924 28033
rect 26608 28024 26660 28076
rect 26792 28024 26844 28076
rect 27160 28067 27212 28076
rect 27160 28033 27169 28067
rect 27169 28033 27203 28067
rect 27203 28033 27212 28067
rect 27160 28024 27212 28033
rect 28540 28024 28592 28076
rect 32128 28067 32180 28076
rect 32128 28033 32137 28067
rect 32137 28033 32171 28067
rect 32171 28033 32180 28067
rect 32128 28024 32180 28033
rect 32404 28067 32456 28076
rect 32404 28033 32413 28067
rect 32413 28033 32447 28067
rect 32447 28033 32456 28067
rect 32404 28024 32456 28033
rect 32772 28024 32824 28076
rect 32956 28024 33008 28076
rect 33324 28024 33376 28076
rect 25412 27888 25464 27940
rect 22376 27820 22428 27872
rect 22468 27820 22520 27872
rect 22744 27863 22796 27872
rect 22744 27829 22753 27863
rect 22753 27829 22787 27863
rect 22787 27829 22796 27863
rect 22744 27820 22796 27829
rect 23112 27863 23164 27872
rect 23112 27829 23121 27863
rect 23121 27829 23155 27863
rect 23155 27829 23164 27863
rect 23112 27820 23164 27829
rect 23940 27863 23992 27872
rect 23940 27829 23949 27863
rect 23949 27829 23983 27863
rect 23983 27829 23992 27863
rect 23940 27820 23992 27829
rect 25136 27820 25188 27872
rect 25780 27931 25832 27940
rect 25780 27897 25789 27931
rect 25789 27897 25823 27931
rect 25823 27897 25832 27931
rect 25780 27888 25832 27897
rect 32588 27956 32640 28008
rect 33600 28024 33652 28076
rect 33876 28067 33928 28076
rect 33876 28033 33885 28067
rect 33885 28033 33919 28067
rect 33919 28033 33928 28067
rect 33876 28024 33928 28033
rect 34428 28067 34480 28076
rect 34428 28033 34437 28067
rect 34437 28033 34471 28067
rect 34471 28033 34480 28067
rect 34428 28024 34480 28033
rect 34704 28024 34756 28076
rect 35256 28024 35308 28076
rect 36728 28160 36780 28212
rect 35440 27999 35492 28008
rect 35440 27965 35449 27999
rect 35449 27965 35483 27999
rect 35483 27965 35492 27999
rect 35440 27956 35492 27965
rect 36728 27888 36780 27940
rect 26792 27820 26844 27872
rect 32496 27820 32548 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 4804 27616 4856 27668
rect 5540 27616 5592 27668
rect 4160 27548 4212 27600
rect 6920 27616 6972 27668
rect 7012 27616 7064 27668
rect 8300 27659 8352 27668
rect 8300 27625 8309 27659
rect 8309 27625 8343 27659
rect 8343 27625 8352 27659
rect 8300 27616 8352 27625
rect 8576 27616 8628 27668
rect 9864 27616 9916 27668
rect 7104 27548 7156 27600
rect 7288 27548 7340 27600
rect 9772 27548 9824 27600
rect 4620 27276 4672 27328
rect 4712 27319 4764 27328
rect 4712 27285 4721 27319
rect 4721 27285 4755 27319
rect 4755 27285 4764 27319
rect 4712 27276 4764 27285
rect 5264 27276 5316 27328
rect 6920 27412 6972 27464
rect 7656 27412 7708 27464
rect 9680 27480 9732 27532
rect 10692 27480 10744 27532
rect 12716 27548 12768 27600
rect 13084 27548 13136 27600
rect 8208 27344 8260 27396
rect 7288 27276 7340 27328
rect 7564 27319 7616 27328
rect 7564 27285 7573 27319
rect 7573 27285 7607 27319
rect 7607 27285 7616 27319
rect 7564 27276 7616 27285
rect 9588 27276 9640 27328
rect 11244 27319 11296 27328
rect 11244 27285 11253 27319
rect 11253 27285 11287 27319
rect 11287 27285 11296 27319
rect 11244 27276 11296 27285
rect 12348 27455 12400 27464
rect 12348 27421 12357 27455
rect 12357 27421 12391 27455
rect 12391 27421 12400 27455
rect 12348 27412 12400 27421
rect 12532 27455 12584 27464
rect 12532 27421 12541 27455
rect 12541 27421 12575 27455
rect 12575 27421 12584 27455
rect 12532 27412 12584 27421
rect 14832 27548 14884 27600
rect 11704 27387 11756 27396
rect 11704 27353 11713 27387
rect 11713 27353 11747 27387
rect 11747 27353 11756 27387
rect 15016 27616 15068 27668
rect 19340 27616 19392 27668
rect 19984 27659 20036 27668
rect 19984 27625 19993 27659
rect 19993 27625 20027 27659
rect 20027 27625 20036 27659
rect 19984 27616 20036 27625
rect 20352 27659 20404 27668
rect 20352 27625 20361 27659
rect 20361 27625 20395 27659
rect 20395 27625 20404 27659
rect 20352 27616 20404 27625
rect 22376 27616 22428 27668
rect 25412 27616 25464 27668
rect 16396 27548 16448 27600
rect 19524 27548 19576 27600
rect 11704 27344 11756 27353
rect 13268 27344 13320 27396
rect 14096 27344 14148 27396
rect 14372 27455 14424 27464
rect 14372 27421 14381 27455
rect 14381 27421 14415 27455
rect 14415 27421 14424 27455
rect 14372 27412 14424 27421
rect 14832 27455 14884 27464
rect 14832 27421 14841 27455
rect 14841 27421 14875 27455
rect 14875 27421 14884 27455
rect 14832 27412 14884 27421
rect 15660 27412 15712 27464
rect 17684 27412 17736 27464
rect 17500 27344 17552 27396
rect 13176 27319 13228 27328
rect 13176 27285 13185 27319
rect 13185 27285 13219 27319
rect 13219 27285 13228 27319
rect 13176 27276 13228 27285
rect 14188 27319 14240 27328
rect 14188 27285 14197 27319
rect 14197 27285 14231 27319
rect 14231 27285 14240 27319
rect 14188 27276 14240 27285
rect 15384 27276 15436 27328
rect 18696 27344 18748 27396
rect 19248 27344 19300 27396
rect 19524 27412 19576 27464
rect 19892 27455 19944 27464
rect 19892 27421 19901 27455
rect 19901 27421 19935 27455
rect 19935 27421 19944 27455
rect 19892 27412 19944 27421
rect 22192 27412 22244 27464
rect 23020 27548 23072 27600
rect 23112 27548 23164 27600
rect 24400 27548 24452 27600
rect 25964 27548 26016 27600
rect 27528 27548 27580 27600
rect 27804 27548 27856 27600
rect 29460 27548 29512 27600
rect 22744 27455 22796 27464
rect 22744 27421 22753 27455
rect 22753 27421 22787 27455
rect 22787 27421 22796 27455
rect 22744 27412 22796 27421
rect 22836 27412 22888 27464
rect 25136 27412 25188 27464
rect 27160 27412 27212 27464
rect 27436 27455 27488 27464
rect 27436 27421 27445 27455
rect 27445 27421 27479 27455
rect 27479 27421 27488 27455
rect 27436 27412 27488 27421
rect 17684 27276 17736 27328
rect 23112 27344 23164 27396
rect 25228 27344 25280 27396
rect 29736 27480 29788 27532
rect 32864 27480 32916 27532
rect 28724 27412 28776 27464
rect 29368 27455 29420 27464
rect 29368 27421 29377 27455
rect 29377 27421 29411 27455
rect 29411 27421 29420 27455
rect 29368 27412 29420 27421
rect 29644 27387 29696 27396
rect 29644 27353 29653 27387
rect 29653 27353 29687 27387
rect 29687 27353 29696 27387
rect 29644 27344 29696 27353
rect 22284 27276 22336 27328
rect 24584 27276 24636 27328
rect 28908 27276 28960 27328
rect 29552 27276 29604 27328
rect 29920 27412 29972 27464
rect 30380 27412 30432 27464
rect 30012 27387 30064 27396
rect 30012 27353 30021 27387
rect 30021 27353 30055 27387
rect 30055 27353 30064 27387
rect 30012 27344 30064 27353
rect 34520 27412 34572 27464
rect 34796 27412 34848 27464
rect 34888 27455 34940 27464
rect 34888 27421 34897 27455
rect 34897 27421 34931 27455
rect 34931 27421 34940 27455
rect 34888 27412 34940 27421
rect 36452 27455 36504 27464
rect 36452 27421 36461 27455
rect 36461 27421 36495 27455
rect 36495 27421 36504 27455
rect 36452 27412 36504 27421
rect 37096 27480 37148 27532
rect 36820 27412 36872 27464
rect 34428 27344 34480 27396
rect 30932 27276 30984 27328
rect 34336 27276 34388 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 2780 27072 2832 27124
rect 5632 27115 5684 27124
rect 5632 27081 5641 27115
rect 5641 27081 5675 27115
rect 5675 27081 5684 27115
rect 5632 27072 5684 27081
rect 2136 26979 2188 26988
rect 2136 26945 2145 26979
rect 2145 26945 2179 26979
rect 2179 26945 2188 26979
rect 2136 26936 2188 26945
rect 3976 26979 4028 26988
rect 3976 26945 3985 26979
rect 3985 26945 4019 26979
rect 4019 26945 4028 26979
rect 3976 26936 4028 26945
rect 3424 26868 3476 26920
rect 4804 26936 4856 26988
rect 5908 26979 5960 26988
rect 5908 26945 5917 26979
rect 5917 26945 5951 26979
rect 5951 26945 5960 26979
rect 5908 26936 5960 26945
rect 6092 26979 6144 26988
rect 6092 26945 6101 26979
rect 6101 26945 6135 26979
rect 6135 26945 6144 26979
rect 6092 26936 6144 26945
rect 6184 26979 6236 26988
rect 6184 26945 6193 26979
rect 6193 26945 6227 26979
rect 6227 26945 6236 26979
rect 6184 26936 6236 26945
rect 6920 27004 6972 27056
rect 7564 27004 7616 27056
rect 7288 26936 7340 26988
rect 5540 26868 5592 26920
rect 6644 26911 6696 26920
rect 6644 26877 6653 26911
rect 6653 26877 6687 26911
rect 6687 26877 6696 26911
rect 6644 26868 6696 26877
rect 6920 26868 6972 26920
rect 7196 26868 7248 26920
rect 7656 26979 7708 26988
rect 7656 26945 7665 26979
rect 7665 26945 7699 26979
rect 7699 26945 7708 26979
rect 7656 26936 7708 26945
rect 8208 27115 8260 27124
rect 8208 27081 8217 27115
rect 8217 27081 8251 27115
rect 8251 27081 8260 27115
rect 8208 27072 8260 27081
rect 12440 27072 12492 27124
rect 15752 27072 15804 27124
rect 17500 27115 17552 27124
rect 9864 27004 9916 27056
rect 12992 27047 13044 27056
rect 12992 27013 13001 27047
rect 13001 27013 13035 27047
rect 13035 27013 13044 27047
rect 12992 27004 13044 27013
rect 13636 27004 13688 27056
rect 14096 27004 14148 27056
rect 8668 26979 8720 26988
rect 8668 26945 8677 26979
rect 8677 26945 8711 26979
rect 8711 26945 8720 26979
rect 8668 26936 8720 26945
rect 15384 26979 15436 26988
rect 15384 26945 15393 26979
rect 15393 26945 15427 26979
rect 15427 26945 15436 26979
rect 15384 26936 15436 26945
rect 16396 26979 16448 26988
rect 16396 26945 16405 26979
rect 16405 26945 16439 26979
rect 16439 26945 16448 26979
rect 16396 26936 16448 26945
rect 16948 26936 17000 26988
rect 17500 27081 17509 27115
rect 17509 27081 17543 27115
rect 17543 27081 17552 27115
rect 17500 27072 17552 27081
rect 18052 27072 18104 27124
rect 19248 27115 19300 27124
rect 19248 27081 19257 27115
rect 19257 27081 19291 27115
rect 19291 27081 19300 27115
rect 19248 27072 19300 27081
rect 19432 27072 19484 27124
rect 22560 27072 22612 27124
rect 25136 27072 25188 27124
rect 25228 27115 25280 27124
rect 25228 27081 25237 27115
rect 25237 27081 25271 27115
rect 25271 27081 25280 27115
rect 25228 27072 25280 27081
rect 25596 27072 25648 27124
rect 27068 27072 27120 27124
rect 27252 27072 27304 27124
rect 27436 27072 27488 27124
rect 28356 27115 28408 27124
rect 28356 27081 28365 27115
rect 28365 27081 28399 27115
rect 28399 27081 28408 27115
rect 28356 27072 28408 27081
rect 8024 26800 8076 26852
rect 12808 26868 12860 26920
rect 14188 26868 14240 26920
rect 18512 26868 18564 26920
rect 19432 26979 19484 26988
rect 19432 26945 19441 26979
rect 19441 26945 19475 26979
rect 19475 26945 19484 26979
rect 19432 26936 19484 26945
rect 19524 26979 19576 26988
rect 19524 26945 19533 26979
rect 19533 26945 19567 26979
rect 19567 26945 19576 26979
rect 19524 26936 19576 26945
rect 19616 26979 19668 26988
rect 19616 26945 19625 26979
rect 19625 26945 19659 26979
rect 19659 26945 19668 26979
rect 19616 26936 19668 26945
rect 19800 26979 19852 26988
rect 19800 26945 19809 26979
rect 19809 26945 19843 26979
rect 19843 26945 19852 26979
rect 19800 26936 19852 26945
rect 18788 26868 18840 26920
rect 20628 26936 20680 26988
rect 20720 26979 20772 26988
rect 20720 26945 20729 26979
rect 20729 26945 20763 26979
rect 20763 26945 20772 26979
rect 20720 26936 20772 26945
rect 22928 26979 22980 26988
rect 22928 26945 22937 26979
rect 22937 26945 22971 26979
rect 22971 26945 22980 26979
rect 22928 26936 22980 26945
rect 23020 26936 23072 26988
rect 20076 26868 20128 26920
rect 24584 26979 24636 26988
rect 24584 26945 24593 26979
rect 24593 26945 24627 26979
rect 24627 26945 24636 26979
rect 24584 26936 24636 26945
rect 24768 26936 24820 26988
rect 4068 26775 4120 26784
rect 4068 26741 4077 26775
rect 4077 26741 4111 26775
rect 4111 26741 4120 26775
rect 4068 26732 4120 26741
rect 4620 26732 4672 26784
rect 4804 26775 4856 26784
rect 4804 26741 4813 26775
rect 4813 26741 4847 26775
rect 4847 26741 4856 26775
rect 4804 26732 4856 26741
rect 5264 26775 5316 26784
rect 5264 26741 5273 26775
rect 5273 26741 5307 26775
rect 5307 26741 5316 26775
rect 5264 26732 5316 26741
rect 5908 26732 5960 26784
rect 6828 26775 6880 26784
rect 6828 26741 6837 26775
rect 6837 26741 6871 26775
rect 6871 26741 6880 26775
rect 6828 26732 6880 26741
rect 7288 26775 7340 26784
rect 7288 26741 7297 26775
rect 7297 26741 7331 26775
rect 7331 26741 7340 26775
rect 7288 26732 7340 26741
rect 7656 26732 7708 26784
rect 8208 26732 8260 26784
rect 9312 26732 9364 26784
rect 9404 26732 9456 26784
rect 14924 26775 14976 26784
rect 14924 26741 14933 26775
rect 14933 26741 14967 26775
rect 14967 26741 14976 26775
rect 14924 26732 14976 26741
rect 16304 26775 16356 26784
rect 16304 26741 16313 26775
rect 16313 26741 16347 26775
rect 16347 26741 16356 26775
rect 16304 26732 16356 26741
rect 17776 26732 17828 26784
rect 20996 26775 21048 26784
rect 20996 26741 21005 26775
rect 21005 26741 21039 26775
rect 21039 26741 21048 26775
rect 20996 26732 21048 26741
rect 23112 26800 23164 26852
rect 24124 26732 24176 26784
rect 25872 27004 25924 27056
rect 25136 26936 25188 26988
rect 25228 26979 25280 26988
rect 25228 26945 25237 26979
rect 25237 26945 25271 26979
rect 25271 26945 25280 26979
rect 25228 26936 25280 26945
rect 25964 26979 26016 26988
rect 25964 26945 25973 26979
rect 25973 26945 26007 26979
rect 26007 26945 26016 26979
rect 25964 26936 26016 26945
rect 26608 26979 26660 26988
rect 26608 26945 26617 26979
rect 26617 26945 26651 26979
rect 26651 26945 26660 26979
rect 26608 26936 26660 26945
rect 26792 26979 26844 26988
rect 26792 26945 26801 26979
rect 26801 26945 26835 26979
rect 26835 26945 26844 26979
rect 26792 26936 26844 26945
rect 25136 26800 25188 26852
rect 25228 26732 25280 26784
rect 27252 26936 27304 26988
rect 28724 27004 28776 27056
rect 27712 26979 27764 26988
rect 27712 26945 27721 26979
rect 27721 26945 27755 26979
rect 27755 26945 27764 26979
rect 27712 26936 27764 26945
rect 27896 26979 27948 26988
rect 27896 26945 27905 26979
rect 27905 26945 27939 26979
rect 27939 26945 27948 26979
rect 27896 26936 27948 26945
rect 27988 26979 28040 26988
rect 27988 26945 27997 26979
rect 27997 26945 28031 26979
rect 28031 26945 28040 26979
rect 27988 26936 28040 26945
rect 27160 26800 27212 26852
rect 27988 26800 28040 26852
rect 29184 26936 29236 26988
rect 30012 27004 30064 27056
rect 31300 27072 31352 27124
rect 32128 27072 32180 27124
rect 34888 27072 34940 27124
rect 30196 26979 30248 26988
rect 30196 26945 30205 26979
rect 30205 26945 30239 26979
rect 30239 26945 30248 26979
rect 30196 26936 30248 26945
rect 30472 26979 30524 26988
rect 30472 26945 30481 26979
rect 30481 26945 30515 26979
rect 30515 26945 30524 26979
rect 30472 26936 30524 26945
rect 25872 26732 25924 26784
rect 26148 26732 26200 26784
rect 27436 26732 27488 26784
rect 30288 26868 30340 26920
rect 30932 26936 30984 26988
rect 30748 26800 30800 26852
rect 31576 26979 31628 26988
rect 31576 26945 31585 26979
rect 31585 26945 31619 26979
rect 31619 26945 31628 26979
rect 31576 26936 31628 26945
rect 32404 26936 32456 26988
rect 33232 26979 33284 26988
rect 33232 26945 33241 26979
rect 33241 26945 33275 26979
rect 33275 26945 33284 26979
rect 33232 26936 33284 26945
rect 34428 27004 34480 27056
rect 33784 26979 33836 26988
rect 33784 26945 33794 26979
rect 33794 26945 33828 26979
rect 33828 26945 33836 26979
rect 33784 26936 33836 26945
rect 34060 26979 34112 26988
rect 34060 26945 34069 26979
rect 34069 26945 34103 26979
rect 34103 26945 34112 26979
rect 34060 26936 34112 26945
rect 36544 27072 36596 27124
rect 36176 27004 36228 27056
rect 36636 27004 36688 27056
rect 36728 27047 36780 27056
rect 36728 27013 36737 27047
rect 36737 27013 36771 27047
rect 36771 27013 36780 27047
rect 36728 27004 36780 27013
rect 34704 26979 34756 26988
rect 34704 26945 34713 26979
rect 34713 26945 34747 26979
rect 34747 26945 34756 26979
rect 34704 26936 34756 26945
rect 32772 26868 32824 26920
rect 32956 26911 33008 26920
rect 32956 26877 32965 26911
rect 32965 26877 32999 26911
rect 32999 26877 33008 26911
rect 32956 26868 33008 26877
rect 30380 26732 30432 26784
rect 30564 26732 30616 26784
rect 33140 26732 33192 26784
rect 33416 26732 33468 26784
rect 35348 26936 35400 26988
rect 35440 26979 35492 26988
rect 35440 26945 35449 26979
rect 35449 26945 35483 26979
rect 35483 26945 35492 26979
rect 35440 26936 35492 26945
rect 36820 26936 36872 26988
rect 35992 26868 36044 26920
rect 37004 26732 37056 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 2136 26528 2188 26580
rect 5540 26571 5592 26580
rect 5540 26537 5549 26571
rect 5549 26537 5583 26571
rect 5583 26537 5592 26571
rect 5540 26528 5592 26537
rect 6828 26528 6880 26580
rect 7288 26528 7340 26580
rect 8668 26528 8720 26580
rect 1400 26435 1452 26444
rect 1400 26401 1409 26435
rect 1409 26401 1443 26435
rect 1443 26401 1452 26435
rect 1400 26392 1452 26401
rect 3976 26460 4028 26512
rect 4804 26460 4856 26512
rect 4620 26392 4672 26444
rect 2780 26324 2832 26376
rect 4528 26299 4580 26308
rect 4528 26265 4537 26299
rect 4537 26265 4571 26299
rect 4571 26265 4580 26299
rect 9404 26460 9456 26512
rect 7012 26392 7064 26444
rect 8024 26392 8076 26444
rect 11244 26528 11296 26580
rect 13176 26528 13228 26580
rect 13268 26571 13320 26580
rect 13268 26537 13277 26571
rect 13277 26537 13311 26571
rect 13311 26537 13320 26571
rect 13268 26528 13320 26537
rect 15568 26528 15620 26580
rect 10416 26392 10468 26444
rect 12256 26392 12308 26444
rect 12440 26392 12492 26444
rect 7472 26324 7524 26376
rect 14096 26460 14148 26512
rect 19340 26528 19392 26580
rect 20628 26528 20680 26580
rect 20996 26528 21048 26580
rect 16856 26460 16908 26512
rect 16948 26460 17000 26512
rect 15200 26392 15252 26444
rect 16028 26392 16080 26444
rect 17316 26460 17368 26512
rect 18328 26435 18380 26444
rect 18328 26401 18337 26435
rect 18337 26401 18371 26435
rect 18371 26401 18380 26435
rect 18328 26392 18380 26401
rect 15016 26324 15068 26376
rect 16304 26324 16356 26376
rect 17040 26324 17092 26376
rect 4528 26256 4580 26265
rect 7932 26256 7984 26308
rect 5264 26188 5316 26240
rect 6828 26188 6880 26240
rect 9404 26231 9456 26240
rect 9404 26197 9413 26231
rect 9413 26197 9447 26231
rect 9447 26197 9456 26231
rect 9404 26188 9456 26197
rect 9864 26256 9916 26308
rect 12256 26256 12308 26308
rect 16488 26256 16540 26308
rect 17592 26367 17644 26376
rect 17592 26333 17601 26367
rect 17601 26333 17635 26367
rect 17635 26333 17644 26367
rect 17592 26324 17644 26333
rect 18052 26324 18104 26376
rect 18512 26324 18564 26376
rect 21364 26367 21416 26376
rect 21364 26333 21373 26367
rect 21373 26333 21407 26367
rect 21407 26333 21416 26367
rect 21364 26324 21416 26333
rect 17500 26188 17552 26240
rect 17868 26231 17920 26240
rect 17868 26197 17877 26231
rect 17877 26197 17911 26231
rect 17911 26197 17920 26231
rect 17868 26188 17920 26197
rect 18052 26188 18104 26240
rect 20720 26256 20772 26308
rect 22928 26528 22980 26580
rect 24400 26528 24452 26580
rect 25504 26528 25556 26580
rect 23296 26460 23348 26512
rect 23480 26392 23532 26444
rect 22376 26367 22428 26376
rect 22376 26333 22405 26367
rect 22405 26333 22428 26367
rect 23848 26460 23900 26512
rect 24768 26460 24820 26512
rect 22376 26324 22428 26333
rect 22192 26256 22244 26308
rect 23848 26367 23900 26376
rect 23848 26333 23857 26367
rect 23857 26333 23891 26367
rect 23891 26333 23900 26367
rect 23848 26324 23900 26333
rect 24216 26299 24268 26308
rect 24216 26265 24225 26299
rect 24225 26265 24259 26299
rect 24259 26265 24268 26299
rect 24216 26256 24268 26265
rect 25044 26324 25096 26376
rect 25412 26392 25464 26444
rect 25320 26367 25372 26376
rect 25320 26333 25329 26367
rect 25329 26333 25363 26367
rect 25363 26333 25372 26367
rect 25320 26324 25372 26333
rect 26332 26460 26384 26512
rect 26884 26460 26936 26512
rect 27712 26528 27764 26580
rect 27896 26528 27948 26580
rect 29184 26528 29236 26580
rect 29644 26528 29696 26580
rect 30288 26528 30340 26580
rect 32956 26571 33008 26580
rect 32956 26537 32965 26571
rect 32965 26537 32999 26571
rect 32999 26537 33008 26571
rect 32956 26528 33008 26537
rect 33416 26528 33468 26580
rect 34704 26528 34756 26580
rect 35440 26528 35492 26580
rect 36820 26571 36872 26580
rect 36820 26537 36829 26571
rect 36829 26537 36863 26571
rect 36863 26537 36872 26571
rect 36820 26528 36872 26537
rect 37004 26571 37056 26580
rect 37004 26537 37013 26571
rect 37013 26537 37047 26571
rect 37047 26537 37056 26571
rect 37004 26528 37056 26537
rect 26148 26367 26200 26376
rect 26148 26333 26157 26367
rect 26157 26333 26191 26367
rect 26191 26333 26200 26367
rect 26148 26324 26200 26333
rect 25688 26256 25740 26308
rect 26884 26324 26936 26376
rect 27160 26324 27212 26376
rect 27344 26367 27396 26376
rect 27344 26333 27353 26367
rect 27353 26333 27387 26367
rect 27387 26333 27396 26367
rect 27344 26324 27396 26333
rect 27436 26367 27488 26376
rect 27436 26333 27445 26367
rect 27445 26333 27479 26367
rect 27479 26333 27488 26367
rect 27436 26324 27488 26333
rect 28172 26324 28224 26376
rect 27896 26256 27948 26308
rect 28540 26392 28592 26444
rect 28724 26392 28776 26444
rect 28908 26369 28960 26376
rect 28908 26335 28917 26369
rect 28917 26335 28951 26369
rect 28951 26335 28960 26369
rect 31116 26392 31168 26444
rect 32496 26435 32548 26444
rect 32496 26401 32505 26435
rect 32505 26401 32539 26435
rect 32539 26401 32548 26435
rect 32496 26392 32548 26401
rect 28908 26324 28960 26335
rect 27252 26188 27304 26240
rect 28540 26231 28592 26240
rect 28540 26197 28549 26231
rect 28549 26197 28583 26231
rect 28583 26197 28592 26231
rect 28540 26188 28592 26197
rect 29368 26256 29420 26308
rect 29552 26299 29604 26308
rect 29552 26265 29561 26299
rect 29561 26265 29595 26299
rect 29595 26265 29604 26299
rect 29552 26256 29604 26265
rect 32220 26367 32272 26376
rect 32220 26333 32229 26367
rect 32229 26333 32263 26367
rect 32263 26333 32272 26367
rect 32220 26324 32272 26333
rect 32312 26256 32364 26308
rect 32956 26324 33008 26376
rect 33232 26392 33284 26444
rect 36728 26460 36780 26512
rect 33140 26324 33192 26376
rect 33416 26324 33468 26376
rect 34336 26324 34388 26376
rect 34244 26256 34296 26308
rect 36728 26324 36780 26376
rect 29184 26188 29236 26240
rect 31208 26188 31260 26240
rect 34336 26188 34388 26240
rect 37188 26188 37240 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 3424 26027 3476 26036
rect 3424 25993 3433 26027
rect 3433 25993 3467 26027
rect 3467 25993 3476 26027
rect 3424 25984 3476 25993
rect 1768 25959 1820 25968
rect 1768 25925 1777 25959
rect 1777 25925 1811 25959
rect 1811 25925 1820 25959
rect 1768 25916 1820 25925
rect 4528 25916 4580 25968
rect 5724 25984 5776 26036
rect 6920 25984 6972 26036
rect 9680 25984 9732 26036
rect 14648 25984 14700 26036
rect 7288 25916 7340 25968
rect 13360 25959 13412 25968
rect 13360 25925 13369 25959
rect 13369 25925 13403 25959
rect 13403 25925 13412 25959
rect 13360 25916 13412 25925
rect 940 25848 992 25900
rect 3332 25891 3384 25900
rect 3332 25857 3341 25891
rect 3341 25857 3375 25891
rect 3375 25857 3384 25891
rect 3332 25848 3384 25857
rect 4160 25848 4212 25900
rect 4620 25891 4672 25900
rect 4620 25857 4629 25891
rect 4629 25857 4663 25891
rect 4663 25857 4672 25891
rect 4620 25848 4672 25857
rect 5264 25848 5316 25900
rect 6368 25891 6420 25900
rect 6368 25857 6377 25891
rect 6377 25857 6411 25891
rect 6411 25857 6420 25891
rect 6368 25848 6420 25857
rect 7748 25848 7800 25900
rect 13176 25891 13228 25900
rect 13176 25857 13180 25891
rect 13180 25857 13214 25891
rect 13214 25857 13228 25891
rect 13176 25848 13228 25857
rect 13544 25891 13596 25900
rect 13544 25857 13553 25891
rect 13553 25857 13587 25891
rect 13587 25857 13596 25891
rect 13544 25848 13596 25857
rect 14188 25848 14240 25900
rect 14464 25848 14516 25900
rect 6644 25780 6696 25832
rect 4804 25712 4856 25764
rect 5448 25712 5500 25764
rect 14832 25959 14884 25968
rect 14832 25925 14841 25959
rect 14841 25925 14875 25959
rect 14875 25925 14884 25959
rect 14832 25916 14884 25925
rect 14740 25891 14792 25900
rect 14740 25857 14744 25891
rect 14744 25857 14778 25891
rect 14778 25857 14792 25891
rect 14740 25848 14792 25857
rect 15568 25848 15620 25900
rect 7288 25712 7340 25764
rect 15108 25712 15160 25764
rect 9680 25644 9732 25696
rect 14556 25687 14608 25696
rect 14556 25653 14565 25687
rect 14565 25653 14599 25687
rect 14599 25653 14608 25687
rect 14556 25644 14608 25653
rect 14740 25644 14792 25696
rect 15292 25644 15344 25696
rect 15660 25644 15712 25696
rect 15752 25687 15804 25696
rect 15752 25653 15761 25687
rect 15761 25653 15795 25687
rect 15795 25653 15804 25687
rect 15752 25644 15804 25653
rect 16212 25916 16264 25968
rect 16396 25916 16448 25968
rect 16580 25848 16632 25900
rect 17592 25848 17644 25900
rect 16488 25780 16540 25832
rect 19248 25891 19300 25900
rect 19248 25857 19257 25891
rect 19257 25857 19291 25891
rect 19291 25857 19300 25891
rect 19248 25848 19300 25857
rect 19340 25891 19392 25900
rect 19340 25857 19349 25891
rect 19349 25857 19383 25891
rect 19383 25857 19392 25891
rect 19340 25848 19392 25857
rect 19708 25916 19760 25968
rect 20628 25984 20680 26036
rect 23848 25984 23900 26036
rect 26332 25984 26384 26036
rect 28172 25984 28224 26036
rect 29092 25984 29144 26036
rect 30196 25984 30248 26036
rect 32220 25984 32272 26036
rect 32588 25984 32640 26036
rect 23204 25916 23256 25968
rect 20076 25848 20128 25900
rect 20168 25891 20220 25900
rect 20168 25857 20177 25891
rect 20177 25857 20211 25891
rect 20211 25857 20220 25891
rect 20168 25848 20220 25857
rect 22376 25848 22428 25900
rect 23480 25891 23532 25900
rect 23480 25857 23489 25891
rect 23489 25857 23523 25891
rect 23523 25857 23532 25891
rect 23480 25848 23532 25857
rect 17132 25712 17184 25764
rect 17316 25644 17368 25696
rect 17408 25644 17460 25696
rect 18788 25644 18840 25696
rect 18972 25687 19024 25696
rect 18972 25653 18981 25687
rect 18981 25653 19015 25687
rect 19015 25653 19024 25687
rect 18972 25644 19024 25653
rect 19708 25755 19760 25764
rect 19708 25721 19717 25755
rect 19717 25721 19751 25755
rect 19751 25721 19760 25755
rect 19708 25712 19760 25721
rect 26148 25891 26200 25900
rect 26148 25857 26157 25891
rect 26157 25857 26191 25891
rect 26191 25857 26200 25891
rect 26148 25848 26200 25857
rect 29184 25916 29236 25968
rect 30288 25916 30340 25968
rect 31024 25916 31076 25968
rect 32956 25984 33008 26036
rect 28540 25848 28592 25900
rect 30380 25848 30432 25900
rect 30840 25848 30892 25900
rect 31208 25891 31260 25900
rect 31208 25857 31217 25891
rect 31217 25857 31251 25891
rect 31251 25857 31260 25891
rect 31208 25848 31260 25857
rect 31392 25891 31444 25900
rect 31392 25857 31401 25891
rect 31401 25857 31435 25891
rect 31435 25857 31444 25891
rect 31392 25848 31444 25857
rect 31484 25891 31536 25900
rect 31484 25857 31493 25891
rect 31493 25857 31527 25891
rect 31527 25857 31536 25891
rect 31484 25848 31536 25857
rect 24860 25780 24912 25832
rect 29092 25780 29144 25832
rect 29552 25780 29604 25832
rect 30564 25780 30616 25832
rect 32220 25848 32272 25900
rect 32312 25891 32364 25900
rect 32312 25857 32321 25891
rect 32321 25857 32355 25891
rect 32355 25857 32364 25891
rect 32312 25848 32364 25857
rect 19984 25644 20036 25696
rect 31300 25712 31352 25764
rect 24124 25687 24176 25696
rect 24124 25653 24133 25687
rect 24133 25653 24167 25687
rect 24167 25653 24176 25687
rect 24124 25644 24176 25653
rect 27068 25644 27120 25696
rect 31944 25712 31996 25764
rect 32496 25823 32548 25832
rect 32496 25789 32505 25823
rect 32505 25789 32539 25823
rect 32539 25789 32548 25823
rect 32496 25780 32548 25789
rect 32864 25780 32916 25832
rect 33232 25780 33284 25832
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 7288 25440 7340 25492
rect 1400 25347 1452 25356
rect 1400 25313 1409 25347
rect 1409 25313 1443 25347
rect 1443 25313 1452 25347
rect 1400 25304 1452 25313
rect 4528 25304 4580 25356
rect 2780 25236 2832 25288
rect 4712 25236 4764 25288
rect 6828 25279 6880 25288
rect 6828 25245 6837 25279
rect 6837 25245 6871 25279
rect 6871 25245 6880 25279
rect 6828 25236 6880 25245
rect 6920 25236 6972 25288
rect 1676 25211 1728 25220
rect 1676 25177 1685 25211
rect 1685 25177 1719 25211
rect 1719 25177 1728 25211
rect 1676 25168 1728 25177
rect 5448 25168 5500 25220
rect 8300 25372 8352 25424
rect 9772 25372 9824 25424
rect 3792 25143 3844 25152
rect 3792 25109 3801 25143
rect 3801 25109 3835 25143
rect 3835 25109 3844 25143
rect 3792 25100 3844 25109
rect 5816 25100 5868 25152
rect 6460 25143 6512 25152
rect 6460 25109 6469 25143
rect 6469 25109 6503 25143
rect 6503 25109 6512 25143
rect 6460 25100 6512 25109
rect 10416 25347 10468 25356
rect 10416 25313 10425 25347
rect 10425 25313 10459 25347
rect 10459 25313 10468 25347
rect 10416 25304 10468 25313
rect 12900 25347 12952 25356
rect 12900 25313 12909 25347
rect 12909 25313 12943 25347
rect 12943 25313 12952 25347
rect 12900 25304 12952 25313
rect 8208 25236 8260 25288
rect 9496 25236 9548 25288
rect 12440 25236 12492 25288
rect 14740 25440 14792 25492
rect 14832 25440 14884 25492
rect 14924 25440 14976 25492
rect 17408 25440 17460 25492
rect 14280 25279 14332 25288
rect 14280 25245 14289 25279
rect 14289 25245 14323 25279
rect 14323 25245 14332 25279
rect 14280 25236 14332 25245
rect 16212 25372 16264 25424
rect 17316 25372 17368 25424
rect 17960 25483 18012 25492
rect 17960 25449 17969 25483
rect 17969 25449 18003 25483
rect 18003 25449 18012 25483
rect 17960 25440 18012 25449
rect 18052 25440 18104 25492
rect 18696 25483 18748 25492
rect 18696 25449 18705 25483
rect 18705 25449 18739 25483
rect 18739 25449 18748 25483
rect 18696 25440 18748 25449
rect 14740 25304 14792 25356
rect 15568 25304 15620 25356
rect 15016 25236 15068 25288
rect 15844 25279 15896 25288
rect 15844 25245 15848 25279
rect 15848 25245 15882 25279
rect 15882 25245 15896 25279
rect 15844 25236 15896 25245
rect 16028 25279 16080 25288
rect 16028 25245 16037 25279
rect 16037 25245 16071 25279
rect 16071 25245 16080 25279
rect 16028 25236 16080 25245
rect 19708 25440 19760 25492
rect 21364 25440 21416 25492
rect 26332 25440 26384 25492
rect 30288 25440 30340 25492
rect 31392 25440 31444 25492
rect 33048 25483 33100 25492
rect 33048 25449 33057 25483
rect 33057 25449 33091 25483
rect 33091 25449 33100 25483
rect 33048 25440 33100 25449
rect 36728 25483 36780 25492
rect 36728 25449 36737 25483
rect 36737 25449 36771 25483
rect 36771 25449 36780 25483
rect 36728 25440 36780 25449
rect 37188 25483 37240 25492
rect 37188 25449 37197 25483
rect 37197 25449 37231 25483
rect 37231 25449 37240 25483
rect 37188 25440 37240 25449
rect 19064 25372 19116 25424
rect 22192 25372 22244 25424
rect 16580 25236 16632 25288
rect 17040 25236 17092 25288
rect 17500 25236 17552 25288
rect 9864 25168 9916 25220
rect 9036 25100 9088 25152
rect 9588 25100 9640 25152
rect 11060 25143 11112 25152
rect 11060 25109 11069 25143
rect 11069 25109 11103 25143
rect 11103 25109 11112 25143
rect 11060 25100 11112 25109
rect 11428 25211 11480 25220
rect 11428 25177 11437 25211
rect 11437 25177 11471 25211
rect 11471 25177 11480 25211
rect 11428 25168 11480 25177
rect 13452 25168 13504 25220
rect 11612 25100 11664 25152
rect 14096 25143 14148 25152
rect 14096 25109 14105 25143
rect 14105 25109 14139 25143
rect 14139 25109 14148 25143
rect 14096 25100 14148 25109
rect 16488 25168 16540 25220
rect 18052 25279 18104 25288
rect 18052 25245 18061 25279
rect 18061 25245 18095 25279
rect 18095 25245 18104 25279
rect 18052 25236 18104 25245
rect 18144 25236 18196 25288
rect 19984 25347 20036 25356
rect 19984 25313 19993 25347
rect 19993 25313 20027 25347
rect 20027 25313 20036 25347
rect 19984 25304 20036 25313
rect 21916 25304 21968 25356
rect 32864 25372 32916 25424
rect 18512 25100 18564 25152
rect 19892 25279 19944 25288
rect 19892 25245 19901 25279
rect 19901 25245 19935 25279
rect 19935 25245 19944 25279
rect 19892 25236 19944 25245
rect 20536 25279 20588 25288
rect 20536 25245 20545 25279
rect 20545 25245 20579 25279
rect 20579 25245 20588 25279
rect 20536 25236 20588 25245
rect 23756 25236 23808 25288
rect 24676 25236 24728 25288
rect 25044 25279 25096 25288
rect 25044 25245 25053 25279
rect 25053 25245 25087 25279
rect 25087 25245 25096 25279
rect 25044 25236 25096 25245
rect 20812 25168 20864 25220
rect 23204 25168 23256 25220
rect 26700 25236 26752 25288
rect 27252 25279 27304 25288
rect 27252 25245 27261 25279
rect 27261 25245 27295 25279
rect 27295 25245 27304 25279
rect 27252 25236 27304 25245
rect 27344 25236 27396 25288
rect 30472 25279 30524 25288
rect 30472 25245 30481 25279
rect 30481 25245 30515 25279
rect 30515 25245 30524 25279
rect 30472 25236 30524 25245
rect 30748 25279 30800 25288
rect 30748 25245 30757 25279
rect 30757 25245 30791 25279
rect 30791 25245 30800 25279
rect 30748 25236 30800 25245
rect 30840 25279 30892 25288
rect 30840 25245 30849 25279
rect 30849 25245 30883 25279
rect 30883 25245 30892 25279
rect 30840 25236 30892 25245
rect 31116 25236 31168 25288
rect 32588 25236 32640 25288
rect 30380 25168 30432 25220
rect 32128 25168 32180 25220
rect 32956 25236 33008 25288
rect 33324 25279 33376 25288
rect 33324 25245 33333 25279
rect 33333 25245 33367 25279
rect 33367 25245 33376 25279
rect 33324 25236 33376 25245
rect 36452 25304 36504 25356
rect 33232 25168 33284 25220
rect 33692 25279 33744 25288
rect 33692 25245 33701 25279
rect 33701 25245 33735 25279
rect 33735 25245 33744 25279
rect 33692 25236 33744 25245
rect 37004 25279 37056 25288
rect 37004 25245 37013 25279
rect 37013 25245 37047 25279
rect 37047 25245 37056 25279
rect 37004 25236 37056 25245
rect 22008 25100 22060 25152
rect 22100 25100 22152 25152
rect 25320 25100 25372 25152
rect 27620 25100 27672 25152
rect 31484 25100 31536 25152
rect 32496 25100 32548 25152
rect 33508 25100 33560 25152
rect 33784 25100 33836 25152
rect 36636 25100 36688 25152
rect 36728 25100 36780 25152
rect 37188 25100 37240 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 1676 24896 1728 24948
rect 2780 24896 2832 24948
rect 3792 24896 3844 24948
rect 4804 24896 4856 24948
rect 8116 24896 8168 24948
rect 11060 24896 11112 24948
rect 11428 24896 11480 24948
rect 11612 24896 11664 24948
rect 14280 24896 14332 24948
rect 14924 24896 14976 24948
rect 15844 24896 15896 24948
rect 2964 24803 3016 24812
rect 2964 24769 2973 24803
rect 2973 24769 3007 24803
rect 3007 24769 3016 24803
rect 2964 24760 3016 24769
rect 4620 24760 4672 24812
rect 4804 24760 4856 24812
rect 6920 24760 6972 24812
rect 7656 24760 7708 24812
rect 10416 24828 10468 24880
rect 8024 24803 8076 24812
rect 8024 24769 8033 24803
rect 8033 24769 8067 24803
rect 8067 24769 8076 24803
rect 8024 24760 8076 24769
rect 14648 24828 14700 24880
rect 3700 24556 3752 24608
rect 5540 24735 5592 24744
rect 5540 24701 5549 24735
rect 5549 24701 5583 24735
rect 5583 24701 5592 24735
rect 5540 24692 5592 24701
rect 6552 24692 6604 24744
rect 6644 24735 6696 24744
rect 6644 24701 6653 24735
rect 6653 24701 6687 24735
rect 6687 24701 6696 24735
rect 6644 24692 6696 24701
rect 7104 24692 7156 24744
rect 7472 24735 7524 24744
rect 7472 24701 7481 24735
rect 7481 24701 7515 24735
rect 7515 24701 7524 24735
rect 7472 24692 7524 24701
rect 7564 24692 7616 24744
rect 5356 24624 5408 24676
rect 6828 24624 6880 24676
rect 8300 24735 8352 24744
rect 8300 24701 8309 24735
rect 8309 24701 8343 24735
rect 8343 24701 8352 24735
rect 8300 24692 8352 24701
rect 9036 24692 9088 24744
rect 10416 24692 10468 24744
rect 11888 24692 11940 24744
rect 13636 24692 13688 24744
rect 5264 24556 5316 24608
rect 5908 24556 5960 24608
rect 6184 24556 6236 24608
rect 7564 24556 7616 24608
rect 12164 24624 12216 24676
rect 14004 24803 14056 24812
rect 14004 24769 14013 24803
rect 14013 24769 14047 24803
rect 14047 24769 14056 24803
rect 14004 24760 14056 24769
rect 14188 24760 14240 24812
rect 14832 24803 14884 24812
rect 14832 24769 14841 24803
rect 14841 24769 14875 24803
rect 14875 24769 14884 24803
rect 14832 24760 14884 24769
rect 15200 24760 15252 24812
rect 15660 24828 15712 24880
rect 16212 24828 16264 24880
rect 17132 24828 17184 24880
rect 17316 24828 17368 24880
rect 17868 24828 17920 24880
rect 16856 24803 16908 24812
rect 16856 24769 16865 24803
rect 16865 24769 16899 24803
rect 16899 24769 16908 24803
rect 16856 24760 16908 24769
rect 17408 24760 17460 24812
rect 20536 24896 20588 24948
rect 22192 24939 22244 24948
rect 22192 24905 22201 24939
rect 22201 24905 22235 24939
rect 22235 24905 22244 24939
rect 22192 24896 22244 24905
rect 22836 24896 22888 24948
rect 28172 24896 28224 24948
rect 28540 24939 28592 24948
rect 28540 24905 28549 24939
rect 28549 24905 28583 24939
rect 28583 24905 28592 24939
rect 28540 24896 28592 24905
rect 29000 24896 29052 24948
rect 30288 24896 30340 24948
rect 18696 24828 18748 24880
rect 18144 24760 18196 24812
rect 18788 24760 18840 24812
rect 19340 24760 19392 24812
rect 20168 24760 20220 24812
rect 21180 24760 21232 24812
rect 22008 24760 22060 24812
rect 18052 24692 18104 24744
rect 18696 24735 18748 24744
rect 18696 24701 18705 24735
rect 18705 24701 18739 24735
rect 18739 24701 18748 24735
rect 18696 24692 18748 24701
rect 20812 24692 20864 24744
rect 21364 24624 21416 24676
rect 22928 24760 22980 24812
rect 23388 24828 23440 24880
rect 23848 24871 23900 24880
rect 23848 24837 23857 24871
rect 23857 24837 23891 24871
rect 23891 24837 23900 24871
rect 23848 24828 23900 24837
rect 23112 24803 23164 24812
rect 23112 24769 23121 24803
rect 23121 24769 23155 24803
rect 23155 24769 23164 24803
rect 23112 24760 23164 24769
rect 23388 24692 23440 24744
rect 23572 24760 23624 24812
rect 23756 24803 23808 24812
rect 23756 24769 23765 24803
rect 23765 24769 23799 24803
rect 23799 24769 23808 24803
rect 23756 24760 23808 24769
rect 24032 24803 24084 24812
rect 24032 24769 24041 24803
rect 24041 24769 24075 24803
rect 24075 24769 24084 24803
rect 24032 24760 24084 24769
rect 24124 24803 24176 24812
rect 24124 24769 24133 24803
rect 24133 24769 24167 24803
rect 24167 24769 24176 24803
rect 24124 24760 24176 24769
rect 26424 24828 26476 24880
rect 24400 24803 24452 24812
rect 24400 24769 24409 24803
rect 24409 24769 24443 24803
rect 24443 24769 24452 24803
rect 24400 24760 24452 24769
rect 24860 24760 24912 24812
rect 25872 24803 25924 24812
rect 25872 24769 25881 24803
rect 25881 24769 25915 24803
rect 25915 24769 25924 24803
rect 25872 24760 25924 24769
rect 24676 24735 24728 24744
rect 24676 24701 24702 24735
rect 24702 24701 24728 24735
rect 24676 24692 24728 24701
rect 26240 24692 26292 24744
rect 26424 24735 26476 24744
rect 26424 24701 26433 24735
rect 26433 24701 26467 24735
rect 26467 24701 26476 24735
rect 26424 24692 26476 24701
rect 26976 24803 27028 24812
rect 26976 24769 26985 24803
rect 26985 24769 27019 24803
rect 27019 24769 27028 24803
rect 26976 24760 27028 24769
rect 27160 24803 27212 24812
rect 27160 24769 27169 24803
rect 27169 24769 27203 24803
rect 27203 24769 27212 24803
rect 27160 24760 27212 24769
rect 27436 24803 27488 24812
rect 27436 24769 27445 24803
rect 27445 24769 27479 24803
rect 27479 24769 27488 24803
rect 27436 24760 27488 24769
rect 27528 24803 27580 24812
rect 27528 24769 27537 24803
rect 27537 24769 27571 24803
rect 27571 24769 27580 24803
rect 27528 24760 27580 24769
rect 28080 24828 28132 24880
rect 30564 24871 30616 24880
rect 30564 24837 30573 24871
rect 30573 24837 30607 24871
rect 30607 24837 30616 24871
rect 30564 24828 30616 24837
rect 31760 24896 31812 24948
rect 32220 24896 32272 24948
rect 33692 24896 33744 24948
rect 29276 24760 29328 24812
rect 28724 24735 28776 24744
rect 28724 24701 28733 24735
rect 28733 24701 28767 24735
rect 28767 24701 28776 24735
rect 28724 24692 28776 24701
rect 29184 24692 29236 24744
rect 32036 24760 32088 24812
rect 33968 24760 34020 24812
rect 34428 24803 34480 24812
rect 34428 24769 34437 24803
rect 34437 24769 34471 24803
rect 34471 24769 34480 24803
rect 34428 24760 34480 24769
rect 36176 24760 36228 24812
rect 13820 24556 13872 24608
rect 15016 24556 15068 24608
rect 17132 24556 17184 24608
rect 18512 24556 18564 24608
rect 19892 24556 19944 24608
rect 21640 24556 21692 24608
rect 22008 24556 22060 24608
rect 30748 24624 30800 24676
rect 31392 24624 31444 24676
rect 23112 24556 23164 24608
rect 23480 24599 23532 24608
rect 23480 24565 23489 24599
rect 23489 24565 23523 24599
rect 23523 24565 23532 24599
rect 23480 24556 23532 24565
rect 24400 24556 24452 24608
rect 25136 24556 25188 24608
rect 27068 24556 27120 24608
rect 29920 24556 29972 24608
rect 31024 24556 31076 24608
rect 31300 24556 31352 24608
rect 33048 24556 33100 24608
rect 33232 24599 33284 24608
rect 33232 24565 33241 24599
rect 33241 24565 33275 24599
rect 33275 24565 33284 24599
rect 33232 24556 33284 24565
rect 33416 24624 33468 24676
rect 36728 24692 36780 24744
rect 36912 24692 36964 24744
rect 33784 24556 33836 24608
rect 34244 24599 34296 24608
rect 34244 24565 34253 24599
rect 34253 24565 34287 24599
rect 34287 24565 34296 24599
rect 34244 24556 34296 24565
rect 36636 24556 36688 24608
rect 36820 24599 36872 24608
rect 36820 24565 36829 24599
rect 36829 24565 36863 24599
rect 36863 24565 36872 24599
rect 36820 24556 36872 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 4712 24352 4764 24404
rect 6736 24352 6788 24404
rect 6920 24352 6972 24404
rect 2964 24259 3016 24268
rect 2964 24225 2973 24259
rect 2973 24225 3007 24259
rect 3007 24225 3016 24259
rect 2964 24216 3016 24225
rect 3700 24216 3752 24268
rect 4620 24216 4672 24268
rect 2780 24148 2832 24200
rect 3792 24191 3844 24200
rect 3792 24157 3801 24191
rect 3801 24157 3835 24191
rect 3835 24157 3844 24191
rect 3792 24148 3844 24157
rect 3976 24148 4028 24200
rect 2320 24055 2372 24064
rect 2320 24021 2329 24055
rect 2329 24021 2363 24055
rect 2363 24021 2372 24055
rect 2320 24012 2372 24021
rect 4804 24012 4856 24064
rect 5632 24148 5684 24200
rect 6092 24148 6144 24200
rect 6644 24148 6696 24200
rect 6920 24191 6972 24200
rect 6920 24157 6929 24191
rect 6929 24157 6963 24191
rect 6963 24157 6972 24191
rect 6920 24148 6972 24157
rect 9772 24352 9824 24404
rect 11888 24395 11940 24404
rect 11888 24361 11897 24395
rect 11897 24361 11931 24395
rect 11931 24361 11940 24395
rect 11888 24352 11940 24361
rect 12164 24352 12216 24404
rect 12716 24352 12768 24404
rect 11980 24327 12032 24336
rect 11980 24293 11989 24327
rect 11989 24293 12023 24327
rect 12023 24293 12032 24327
rect 11980 24284 12032 24293
rect 12348 24284 12400 24336
rect 16212 24352 16264 24404
rect 19064 24352 19116 24404
rect 19708 24352 19760 24404
rect 17592 24284 17644 24336
rect 5540 24080 5592 24132
rect 6000 24080 6052 24132
rect 13728 24216 13780 24268
rect 9496 24191 9548 24200
rect 9496 24157 9505 24191
rect 9505 24157 9539 24191
rect 9539 24157 9548 24191
rect 9496 24148 9548 24157
rect 12348 24191 12400 24200
rect 12348 24157 12357 24191
rect 12357 24157 12391 24191
rect 12391 24157 12400 24191
rect 12348 24148 12400 24157
rect 5264 24012 5316 24064
rect 6644 24012 6696 24064
rect 7196 24012 7248 24064
rect 10232 24080 10284 24132
rect 13452 24191 13504 24200
rect 13452 24157 13461 24191
rect 13461 24157 13495 24191
rect 13495 24157 13504 24191
rect 13452 24148 13504 24157
rect 13544 24148 13596 24200
rect 14372 24216 14424 24268
rect 14740 24216 14792 24268
rect 15384 24191 15436 24200
rect 15384 24157 15392 24191
rect 15392 24157 15426 24191
rect 15426 24157 15436 24191
rect 15384 24148 15436 24157
rect 16856 24216 16908 24268
rect 20996 24216 21048 24268
rect 21824 24327 21876 24336
rect 21824 24293 21833 24327
rect 21833 24293 21867 24327
rect 21867 24293 21876 24327
rect 21824 24284 21876 24293
rect 22100 24284 22152 24336
rect 23020 24284 23072 24336
rect 23664 24327 23716 24336
rect 23664 24293 23673 24327
rect 23673 24293 23707 24327
rect 23707 24293 23716 24327
rect 23664 24284 23716 24293
rect 16028 24191 16080 24200
rect 9588 24012 9640 24064
rect 11520 24012 11572 24064
rect 11612 24012 11664 24064
rect 14648 24080 14700 24132
rect 16028 24157 16037 24191
rect 16037 24157 16071 24191
rect 16071 24157 16080 24191
rect 16028 24148 16080 24157
rect 16396 24191 16448 24200
rect 16396 24157 16405 24191
rect 16405 24157 16439 24191
rect 16439 24157 16448 24191
rect 16396 24148 16448 24157
rect 16764 24191 16816 24200
rect 16764 24157 16773 24191
rect 16773 24157 16807 24191
rect 16807 24157 16816 24191
rect 16764 24148 16816 24157
rect 18696 24148 18748 24200
rect 20168 24080 20220 24132
rect 20720 24148 20772 24200
rect 21364 24148 21416 24200
rect 22560 24259 22612 24268
rect 22560 24225 22585 24259
rect 22585 24225 22612 24259
rect 25872 24352 25924 24404
rect 26608 24352 26660 24404
rect 27436 24352 27488 24404
rect 27528 24352 27580 24404
rect 28632 24395 28684 24404
rect 28632 24361 28641 24395
rect 28641 24361 28675 24395
rect 28675 24361 28684 24395
rect 28632 24352 28684 24361
rect 29000 24352 29052 24404
rect 31576 24352 31628 24404
rect 33140 24395 33192 24404
rect 33140 24361 33149 24395
rect 33149 24361 33183 24395
rect 33183 24361 33192 24395
rect 33140 24352 33192 24361
rect 27620 24284 27672 24336
rect 22560 24216 22612 24225
rect 22284 24191 22336 24200
rect 22284 24157 22293 24191
rect 22293 24157 22327 24191
rect 22327 24157 22336 24191
rect 22284 24148 22336 24157
rect 22928 24148 22980 24200
rect 23204 24148 23256 24200
rect 24216 24148 24268 24200
rect 20628 24012 20680 24064
rect 22836 24123 22888 24132
rect 22836 24089 22845 24123
rect 22845 24089 22879 24123
rect 22879 24089 22888 24123
rect 22836 24080 22888 24089
rect 25044 24191 25096 24200
rect 25044 24157 25053 24191
rect 25053 24157 25087 24191
rect 25087 24157 25096 24191
rect 25044 24148 25096 24157
rect 25320 24191 25372 24200
rect 25320 24157 25329 24191
rect 25329 24157 25363 24191
rect 25363 24157 25372 24191
rect 25320 24148 25372 24157
rect 25596 24148 25648 24200
rect 26148 24191 26200 24200
rect 26148 24157 26157 24191
rect 26157 24157 26191 24191
rect 26191 24157 26200 24191
rect 26148 24148 26200 24157
rect 27896 24259 27948 24268
rect 27896 24225 27905 24259
rect 27905 24225 27939 24259
rect 27939 24225 27948 24259
rect 27896 24216 27948 24225
rect 21640 24012 21692 24064
rect 22468 24055 22520 24064
rect 22468 24021 22477 24055
rect 22477 24021 22511 24055
rect 22511 24021 22520 24055
rect 22468 24012 22520 24021
rect 24860 24012 24912 24064
rect 25780 24012 25832 24064
rect 27436 24012 27488 24064
rect 27804 24148 27856 24200
rect 27988 24191 28040 24200
rect 27988 24157 27997 24191
rect 27997 24157 28031 24191
rect 28031 24157 28040 24191
rect 27988 24148 28040 24157
rect 28172 24191 28224 24200
rect 28172 24157 28181 24191
rect 28181 24157 28215 24191
rect 28215 24157 28224 24191
rect 28172 24148 28224 24157
rect 29736 24284 29788 24336
rect 32220 24284 32272 24336
rect 28816 24216 28868 24268
rect 28724 24191 28776 24200
rect 28724 24157 28733 24191
rect 28733 24157 28767 24191
rect 28767 24157 28776 24191
rect 28724 24148 28776 24157
rect 28908 24191 28960 24200
rect 28908 24157 28917 24191
rect 28917 24157 28951 24191
rect 28951 24157 28960 24191
rect 28908 24148 28960 24157
rect 31392 24216 31444 24268
rect 30104 24148 30156 24200
rect 30472 24191 30524 24200
rect 30472 24157 30481 24191
rect 30481 24157 30515 24191
rect 30515 24157 30524 24191
rect 30472 24148 30524 24157
rect 30840 24191 30892 24200
rect 30840 24157 30849 24191
rect 30849 24157 30883 24191
rect 30883 24157 30892 24191
rect 30840 24148 30892 24157
rect 32036 24148 32088 24200
rect 32128 24148 32180 24200
rect 32864 24167 32873 24200
rect 32873 24167 32907 24200
rect 32907 24167 32916 24200
rect 32864 24148 32916 24167
rect 27620 24012 27672 24064
rect 29644 24080 29696 24132
rect 30564 24080 30616 24132
rect 30748 24123 30800 24132
rect 30748 24089 30757 24123
rect 30757 24089 30791 24123
rect 30791 24089 30800 24123
rect 30748 24080 30800 24089
rect 28908 24012 28960 24064
rect 29828 24012 29880 24064
rect 31944 24012 31996 24064
rect 32404 24055 32456 24064
rect 32404 24021 32413 24055
rect 32413 24021 32447 24055
rect 32447 24021 32456 24055
rect 32404 24012 32456 24021
rect 33048 24080 33100 24132
rect 33324 24080 33376 24132
rect 33784 24148 33836 24200
rect 34428 24148 34480 24200
rect 34612 24148 34664 24200
rect 34888 24191 34940 24200
rect 34888 24157 34897 24191
rect 34897 24157 34931 24191
rect 34931 24157 34940 24191
rect 34888 24148 34940 24157
rect 36268 24284 36320 24336
rect 35164 24191 35216 24200
rect 35164 24157 35203 24191
rect 35203 24157 35216 24191
rect 35164 24148 35216 24157
rect 36084 24148 36136 24200
rect 37004 24148 37056 24200
rect 37188 24191 37240 24200
rect 37188 24157 37197 24191
rect 37197 24157 37231 24191
rect 37231 24157 37240 24191
rect 37188 24148 37240 24157
rect 32772 24012 32824 24064
rect 36912 24080 36964 24132
rect 35256 24055 35308 24064
rect 35256 24021 35265 24055
rect 35265 24021 35299 24055
rect 35299 24021 35308 24055
rect 35256 24012 35308 24021
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 2320 23808 2372 23860
rect 3792 23808 3844 23860
rect 3884 23740 3936 23792
rect 4068 23740 4120 23792
rect 9496 23808 9548 23860
rect 9588 23808 9640 23860
rect 11428 23808 11480 23860
rect 11980 23808 12032 23860
rect 14004 23808 14056 23860
rect 16396 23808 16448 23860
rect 1768 23511 1820 23520
rect 1768 23477 1777 23511
rect 1777 23477 1811 23511
rect 1811 23477 1820 23511
rect 1768 23468 1820 23477
rect 3516 23647 3568 23656
rect 3516 23613 3525 23647
rect 3525 23613 3559 23647
rect 3559 23613 3568 23647
rect 3516 23604 3568 23613
rect 3976 23604 4028 23656
rect 5448 23715 5500 23724
rect 5448 23681 5457 23715
rect 5457 23681 5491 23715
rect 5491 23681 5500 23715
rect 5448 23672 5500 23681
rect 6828 23740 6880 23792
rect 7380 23740 7432 23792
rect 9404 23783 9456 23792
rect 9404 23749 9413 23783
rect 9413 23749 9447 23783
rect 9447 23749 9456 23783
rect 9404 23740 9456 23749
rect 11336 23740 11388 23792
rect 12348 23740 12400 23792
rect 13636 23740 13688 23792
rect 24032 23808 24084 23860
rect 21180 23740 21232 23792
rect 21364 23740 21416 23792
rect 23848 23783 23900 23792
rect 23848 23749 23857 23783
rect 23857 23749 23891 23783
rect 23891 23749 23900 23783
rect 23848 23740 23900 23749
rect 24216 23740 24268 23792
rect 27252 23808 27304 23860
rect 27344 23808 27396 23860
rect 29000 23808 29052 23860
rect 31944 23808 31996 23860
rect 32404 23808 32456 23860
rect 29276 23740 29328 23792
rect 29460 23740 29512 23792
rect 4620 23604 4672 23656
rect 4804 23604 4856 23656
rect 6920 23647 6972 23656
rect 6920 23613 6929 23647
rect 6929 23613 6963 23647
rect 6963 23613 6972 23647
rect 6920 23604 6972 23613
rect 9036 23604 9088 23656
rect 11520 23715 11572 23724
rect 11520 23681 11529 23715
rect 11529 23681 11563 23715
rect 11563 23681 11572 23715
rect 11520 23672 11572 23681
rect 11888 23647 11940 23656
rect 11888 23613 11897 23647
rect 11897 23613 11931 23647
rect 11931 23613 11940 23647
rect 11888 23604 11940 23613
rect 13268 23715 13320 23724
rect 13268 23681 13277 23715
rect 13277 23681 13311 23715
rect 13311 23681 13320 23715
rect 13268 23672 13320 23681
rect 14188 23672 14240 23724
rect 14648 23672 14700 23724
rect 17040 23715 17092 23724
rect 17040 23681 17049 23715
rect 17049 23681 17083 23715
rect 17083 23681 17092 23715
rect 17040 23672 17092 23681
rect 17592 23672 17644 23724
rect 2964 23468 3016 23520
rect 3792 23468 3844 23520
rect 4068 23468 4120 23520
rect 8392 23579 8444 23588
rect 8392 23545 8401 23579
rect 8401 23545 8435 23579
rect 8435 23545 8444 23579
rect 15936 23604 15988 23656
rect 17684 23604 17736 23656
rect 20628 23715 20680 23724
rect 20628 23681 20637 23715
rect 20637 23681 20671 23715
rect 20671 23681 20680 23715
rect 20628 23672 20680 23681
rect 20536 23604 20588 23656
rect 20996 23715 21048 23724
rect 20996 23681 21005 23715
rect 21005 23681 21039 23715
rect 21039 23681 21048 23715
rect 20996 23672 21048 23681
rect 23572 23672 23624 23724
rect 23756 23672 23808 23724
rect 21364 23604 21416 23656
rect 25596 23715 25648 23724
rect 25596 23681 25605 23715
rect 25605 23681 25639 23715
rect 25639 23681 25648 23715
rect 25596 23672 25648 23681
rect 28172 23672 28224 23724
rect 28816 23672 28868 23724
rect 30840 23672 30892 23724
rect 32772 23740 32824 23792
rect 33232 23808 33284 23860
rect 34888 23808 34940 23860
rect 25412 23647 25464 23656
rect 25412 23613 25421 23647
rect 25421 23613 25455 23647
rect 25455 23613 25464 23647
rect 25412 23604 25464 23613
rect 25964 23604 26016 23656
rect 27712 23604 27764 23656
rect 28080 23604 28132 23656
rect 29276 23604 29328 23656
rect 29644 23604 29696 23656
rect 30012 23604 30064 23656
rect 32128 23715 32180 23724
rect 32128 23681 32137 23715
rect 32137 23681 32171 23715
rect 32171 23681 32180 23715
rect 32128 23672 32180 23681
rect 32312 23715 32364 23724
rect 32312 23681 32319 23715
rect 32319 23681 32364 23715
rect 32312 23672 32364 23681
rect 32404 23715 32456 23724
rect 32404 23681 32413 23715
rect 32413 23681 32447 23715
rect 32447 23681 32456 23715
rect 32404 23672 32456 23681
rect 8392 23536 8444 23545
rect 20076 23536 20128 23588
rect 21640 23536 21692 23588
rect 5264 23468 5316 23520
rect 6644 23468 6696 23520
rect 11612 23468 11664 23520
rect 16672 23468 16724 23520
rect 17592 23468 17644 23520
rect 18328 23468 18380 23520
rect 24216 23511 24268 23520
rect 24216 23477 24225 23511
rect 24225 23477 24259 23511
rect 24259 23477 24268 23511
rect 24216 23468 24268 23477
rect 26148 23536 26200 23588
rect 29920 23536 29972 23588
rect 30472 23536 30524 23588
rect 32588 23715 32640 23724
rect 32588 23681 32602 23715
rect 32602 23681 32636 23715
rect 32636 23681 32640 23715
rect 32588 23672 32640 23681
rect 33140 23715 33192 23724
rect 33140 23681 33149 23715
rect 33149 23681 33183 23715
rect 33183 23681 33192 23715
rect 33140 23672 33192 23681
rect 34612 23740 34664 23792
rect 35992 23808 36044 23860
rect 36268 23851 36320 23860
rect 36268 23817 36277 23851
rect 36277 23817 36311 23851
rect 36311 23817 36320 23851
rect 36268 23808 36320 23817
rect 36636 23808 36688 23860
rect 36820 23808 36872 23860
rect 35256 23715 35308 23724
rect 35256 23681 35265 23715
rect 35265 23681 35299 23715
rect 35299 23681 35308 23715
rect 35256 23672 35308 23681
rect 35440 23672 35492 23724
rect 36912 23783 36964 23792
rect 36912 23749 36921 23783
rect 36921 23749 36955 23783
rect 36955 23749 36964 23783
rect 36912 23740 36964 23749
rect 34796 23604 34848 23656
rect 35348 23604 35400 23656
rect 36268 23647 36320 23656
rect 36268 23613 36277 23647
rect 36277 23613 36311 23647
rect 36311 23613 36320 23647
rect 36268 23604 36320 23613
rect 36728 23604 36780 23656
rect 26240 23468 26292 23520
rect 31208 23468 31260 23520
rect 34520 23468 34572 23520
rect 36084 23468 36136 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 2872 23264 2924 23316
rect 3516 23264 3568 23316
rect 3884 23307 3936 23316
rect 3884 23273 3893 23307
rect 3893 23273 3927 23307
rect 3927 23273 3936 23307
rect 3884 23264 3936 23273
rect 4620 23264 4672 23316
rect 6920 23264 6972 23316
rect 1768 23128 1820 23180
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 3700 23196 3752 23248
rect 7748 23196 7800 23248
rect 10232 23264 10284 23316
rect 15752 23264 15804 23316
rect 16672 23264 16724 23316
rect 16764 23307 16816 23316
rect 16764 23273 16773 23307
rect 16773 23273 16807 23307
rect 16807 23273 16816 23307
rect 16764 23264 16816 23273
rect 17040 23264 17092 23316
rect 8116 23128 8168 23180
rect 8392 23128 8444 23180
rect 10324 23196 10376 23248
rect 7288 23060 7340 23112
rect 13268 23196 13320 23248
rect 14372 23196 14424 23248
rect 18880 23264 18932 23316
rect 20168 23307 20220 23316
rect 20168 23273 20177 23307
rect 20177 23273 20211 23307
rect 20211 23273 20220 23307
rect 20168 23264 20220 23273
rect 20904 23264 20956 23316
rect 21364 23264 21416 23316
rect 22100 23264 22152 23316
rect 24584 23264 24636 23316
rect 27620 23307 27672 23316
rect 27620 23273 27629 23307
rect 27629 23273 27663 23307
rect 27663 23273 27672 23307
rect 27620 23264 27672 23273
rect 4712 22924 4764 22976
rect 11060 23103 11112 23112
rect 11060 23069 11069 23103
rect 11069 23069 11103 23103
rect 11103 23069 11112 23103
rect 11060 23060 11112 23069
rect 11612 23060 11664 23112
rect 8668 22992 8720 23044
rect 9772 22967 9824 22976
rect 9772 22933 9781 22967
rect 9781 22933 9815 22967
rect 9815 22933 9824 22967
rect 9772 22924 9824 22933
rect 10784 22992 10836 23044
rect 11520 23035 11572 23044
rect 11520 23001 11529 23035
rect 11529 23001 11563 23035
rect 11563 23001 11572 23035
rect 11520 22992 11572 23001
rect 12164 23060 12216 23112
rect 13544 23103 13596 23112
rect 13544 23069 13553 23103
rect 13553 23069 13587 23103
rect 13587 23069 13596 23103
rect 13544 23060 13596 23069
rect 13728 23103 13780 23112
rect 13728 23069 13737 23103
rect 13737 23069 13771 23103
rect 13771 23069 13780 23103
rect 13728 23060 13780 23069
rect 14464 23060 14516 23112
rect 14924 23103 14976 23112
rect 14924 23069 14933 23103
rect 14933 23069 14967 23103
rect 14967 23069 14976 23103
rect 14924 23060 14976 23069
rect 15108 23103 15160 23112
rect 15108 23069 15117 23103
rect 15117 23069 15151 23103
rect 15151 23069 15160 23103
rect 15108 23060 15160 23069
rect 15200 23060 15252 23112
rect 15660 23103 15712 23112
rect 15660 23069 15669 23103
rect 15669 23069 15703 23103
rect 15703 23069 15712 23103
rect 15660 23060 15712 23069
rect 15844 23103 15896 23112
rect 15844 23069 15853 23103
rect 15853 23069 15887 23103
rect 15887 23069 15896 23103
rect 15844 23060 15896 23069
rect 18328 23171 18380 23180
rect 18328 23137 18337 23171
rect 18337 23137 18371 23171
rect 18371 23137 18380 23171
rect 18328 23128 18380 23137
rect 17040 23060 17092 23112
rect 17316 23103 17368 23112
rect 17316 23069 17325 23103
rect 17325 23069 17359 23103
rect 17359 23069 17368 23103
rect 17316 23060 17368 23069
rect 17408 23103 17460 23112
rect 17408 23069 17417 23103
rect 17417 23069 17451 23103
rect 17451 23069 17460 23103
rect 17408 23060 17460 23069
rect 10232 22924 10284 22976
rect 10508 22924 10560 22976
rect 11612 22924 11664 22976
rect 12440 22967 12492 22976
rect 12440 22933 12449 22967
rect 12449 22933 12483 22967
rect 12483 22933 12492 22967
rect 12440 22924 12492 22933
rect 16028 22967 16080 22976
rect 16028 22933 16037 22967
rect 16037 22933 16071 22967
rect 16071 22933 16080 22967
rect 16028 22924 16080 22933
rect 16856 23035 16908 23044
rect 16856 23001 16865 23035
rect 16865 23001 16899 23035
rect 16899 23001 16908 23035
rect 16856 22992 16908 23001
rect 16948 22992 17000 23044
rect 18420 23060 18472 23112
rect 18604 23060 18656 23112
rect 18696 23103 18748 23112
rect 18696 23069 18705 23103
rect 18705 23069 18739 23103
rect 18739 23069 18748 23103
rect 18696 23060 18748 23069
rect 19708 23171 19760 23180
rect 19708 23137 19717 23171
rect 19717 23137 19751 23171
rect 19751 23137 19760 23171
rect 19708 23128 19760 23137
rect 20812 23128 20864 23180
rect 24860 23239 24912 23248
rect 24860 23205 24869 23239
rect 24869 23205 24903 23239
rect 24903 23205 24912 23239
rect 24860 23196 24912 23205
rect 28816 23264 28868 23316
rect 31300 23264 31352 23316
rect 32680 23264 32732 23316
rect 36268 23264 36320 23316
rect 23388 23128 23440 23180
rect 30748 23196 30800 23248
rect 32128 23196 32180 23248
rect 21364 23103 21416 23112
rect 21364 23069 21373 23103
rect 21373 23069 21407 23103
rect 21407 23069 21416 23103
rect 21364 23060 21416 23069
rect 23296 23060 23348 23112
rect 23848 23060 23900 23112
rect 25412 23060 25464 23112
rect 25780 23060 25832 23112
rect 26516 23103 26568 23112
rect 26516 23069 26525 23103
rect 26525 23069 26559 23103
rect 26559 23069 26568 23103
rect 26516 23060 26568 23069
rect 18236 22924 18288 22976
rect 18328 22924 18380 22976
rect 19616 22967 19668 22976
rect 19616 22933 19625 22967
rect 19625 22933 19659 22967
rect 19659 22933 19668 22967
rect 19616 22924 19668 22933
rect 21272 22992 21324 23044
rect 24400 22992 24452 23044
rect 26240 22992 26292 23044
rect 27436 23060 27488 23112
rect 27620 23060 27672 23112
rect 27804 23103 27856 23112
rect 27804 23069 27813 23103
rect 27813 23069 27847 23103
rect 27847 23069 27856 23103
rect 27804 23060 27856 23069
rect 28724 23128 28776 23180
rect 28816 23103 28868 23112
rect 28816 23069 28825 23103
rect 28825 23069 28859 23103
rect 28859 23069 28868 23103
rect 28816 23060 28868 23069
rect 29184 23171 29236 23180
rect 29184 23137 29193 23171
rect 29193 23137 29227 23171
rect 29227 23137 29236 23171
rect 29184 23128 29236 23137
rect 30472 23128 30524 23180
rect 31668 23171 31720 23180
rect 31668 23137 31677 23171
rect 31677 23137 31711 23171
rect 31711 23137 31720 23171
rect 31668 23128 31720 23137
rect 33876 23128 33928 23180
rect 34520 23128 34572 23180
rect 30104 23103 30156 23112
rect 30104 23069 30113 23103
rect 30113 23069 30147 23103
rect 30147 23069 30156 23103
rect 30104 23060 30156 23069
rect 30288 23103 30340 23112
rect 30288 23069 30297 23103
rect 30297 23069 30331 23103
rect 30331 23069 30340 23103
rect 30288 23060 30340 23069
rect 36820 23060 36872 23112
rect 22744 22967 22796 22976
rect 22744 22933 22753 22967
rect 22753 22933 22787 22967
rect 22787 22933 22796 22967
rect 22744 22924 22796 22933
rect 24860 22924 24912 22976
rect 25596 22924 25648 22976
rect 26332 22924 26384 22976
rect 27252 22924 27304 22976
rect 29184 22992 29236 23044
rect 29276 22992 29328 23044
rect 29644 23035 29696 23044
rect 29644 23001 29653 23035
rect 29653 23001 29687 23035
rect 29687 23001 29696 23035
rect 29644 22992 29696 23001
rect 31484 22992 31536 23044
rect 32220 22992 32272 23044
rect 32680 22992 32732 23044
rect 29736 22924 29788 22976
rect 30472 22967 30524 22976
rect 30472 22933 30481 22967
rect 30481 22933 30515 22967
rect 30515 22933 30524 22967
rect 30472 22924 30524 22933
rect 31024 22924 31076 22976
rect 33876 22924 33928 22976
rect 36728 22924 36780 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 5540 22720 5592 22772
rect 7104 22720 7156 22772
rect 9404 22720 9456 22772
rect 9772 22720 9824 22772
rect 10600 22720 10652 22772
rect 5356 22516 5408 22568
rect 7748 22652 7800 22704
rect 9312 22627 9364 22636
rect 9312 22593 9321 22627
rect 9321 22593 9355 22627
rect 9355 22593 9364 22627
rect 9312 22584 9364 22593
rect 9404 22627 9456 22636
rect 9404 22593 9413 22627
rect 9413 22593 9447 22627
rect 9447 22593 9456 22627
rect 9404 22584 9456 22593
rect 9680 22584 9732 22636
rect 9864 22584 9916 22636
rect 13544 22720 13596 22772
rect 13728 22720 13780 22772
rect 12440 22652 12492 22704
rect 7196 22516 7248 22568
rect 11612 22627 11664 22636
rect 11612 22593 11621 22627
rect 11621 22593 11655 22627
rect 11655 22593 11664 22627
rect 11612 22584 11664 22593
rect 11888 22516 11940 22568
rect 5540 22448 5592 22500
rect 5908 22448 5960 22500
rect 8300 22448 8352 22500
rect 6460 22423 6512 22432
rect 6460 22389 6469 22423
rect 6469 22389 6503 22423
rect 6503 22389 6512 22423
rect 6460 22380 6512 22389
rect 9772 22423 9824 22432
rect 9772 22389 9781 22423
rect 9781 22389 9815 22423
rect 9815 22389 9824 22423
rect 9772 22380 9824 22389
rect 12164 22448 12216 22500
rect 12900 22584 12952 22636
rect 15660 22720 15712 22772
rect 15936 22763 15988 22772
rect 15936 22729 15945 22763
rect 15945 22729 15979 22763
rect 15979 22729 15988 22763
rect 15936 22720 15988 22729
rect 16948 22720 17000 22772
rect 17224 22720 17276 22772
rect 17408 22720 17460 22772
rect 17592 22763 17644 22772
rect 17592 22729 17601 22763
rect 17601 22729 17635 22763
rect 17635 22729 17644 22763
rect 17592 22720 17644 22729
rect 19432 22720 19484 22772
rect 20168 22720 20220 22772
rect 15752 22695 15804 22704
rect 15752 22661 15761 22695
rect 15761 22661 15795 22695
rect 15795 22661 15804 22695
rect 15752 22652 15804 22661
rect 14372 22584 14424 22636
rect 14556 22584 14608 22636
rect 14924 22584 14976 22636
rect 16028 22584 16080 22636
rect 17040 22652 17092 22704
rect 16764 22516 16816 22568
rect 17316 22584 17368 22636
rect 18420 22627 18472 22636
rect 14188 22448 14240 22500
rect 14740 22448 14792 22500
rect 14924 22448 14976 22500
rect 15108 22448 15160 22500
rect 17040 22448 17092 22500
rect 17224 22448 17276 22500
rect 17592 22448 17644 22500
rect 17776 22516 17828 22568
rect 18420 22593 18429 22627
rect 18429 22593 18463 22627
rect 18463 22593 18472 22627
rect 18420 22584 18472 22593
rect 18328 22559 18380 22568
rect 18328 22525 18337 22559
rect 18337 22525 18371 22559
rect 18371 22525 18380 22559
rect 18328 22516 18380 22525
rect 11060 22380 11112 22432
rect 11704 22380 11756 22432
rect 12256 22380 12308 22432
rect 15844 22380 15896 22432
rect 18696 22448 18748 22500
rect 22100 22652 22152 22704
rect 20812 22584 20864 22636
rect 22008 22627 22060 22636
rect 22008 22593 22017 22627
rect 22017 22593 22051 22627
rect 22051 22593 22060 22627
rect 22008 22584 22060 22593
rect 21088 22559 21140 22568
rect 21088 22525 21097 22559
rect 21097 22525 21131 22559
rect 21131 22525 21140 22559
rect 21088 22516 21140 22525
rect 22284 22627 22336 22636
rect 22284 22593 22293 22627
rect 22293 22593 22327 22627
rect 22327 22593 22336 22627
rect 22284 22584 22336 22593
rect 22744 22695 22796 22704
rect 22744 22661 22753 22695
rect 22753 22661 22787 22695
rect 22787 22661 22796 22695
rect 22744 22652 22796 22661
rect 23848 22763 23900 22772
rect 23848 22729 23857 22763
rect 23857 22729 23891 22763
rect 23891 22729 23900 22763
rect 23848 22720 23900 22729
rect 24584 22720 24636 22772
rect 23020 22627 23072 22636
rect 23020 22593 23029 22627
rect 23029 22593 23063 22627
rect 23063 22593 23072 22627
rect 23020 22584 23072 22593
rect 23296 22584 23348 22636
rect 23388 22627 23440 22636
rect 23388 22593 23397 22627
rect 23397 22593 23431 22627
rect 23431 22593 23440 22627
rect 23388 22584 23440 22593
rect 23572 22584 23624 22636
rect 24124 22627 24176 22636
rect 24124 22593 24133 22627
rect 24133 22593 24167 22627
rect 24167 22593 24176 22627
rect 24124 22584 24176 22593
rect 24860 22627 24912 22636
rect 24860 22593 24869 22627
rect 24869 22593 24903 22627
rect 24903 22593 24912 22627
rect 24860 22584 24912 22593
rect 26056 22720 26108 22772
rect 26332 22720 26384 22772
rect 26516 22720 26568 22772
rect 25596 22652 25648 22704
rect 29184 22720 29236 22772
rect 25780 22627 25832 22636
rect 25780 22593 25789 22627
rect 25789 22593 25823 22627
rect 25823 22593 25832 22627
rect 25780 22584 25832 22593
rect 27344 22695 27396 22704
rect 27344 22661 27353 22695
rect 27353 22661 27387 22695
rect 27387 22661 27396 22695
rect 27344 22652 27396 22661
rect 27620 22652 27672 22704
rect 24768 22516 24820 22568
rect 22284 22448 22336 22500
rect 22376 22448 22428 22500
rect 25412 22516 25464 22568
rect 27804 22584 27856 22636
rect 27988 22584 28040 22636
rect 28264 22627 28316 22636
rect 28264 22593 28273 22627
rect 28273 22593 28307 22627
rect 28307 22593 28316 22627
rect 28264 22584 28316 22593
rect 29828 22652 29880 22704
rect 30012 22695 30064 22704
rect 30012 22661 30029 22695
rect 30029 22661 30064 22695
rect 30012 22652 30064 22661
rect 30288 22720 30340 22772
rect 30472 22720 30524 22772
rect 30748 22720 30800 22772
rect 31208 22720 31260 22772
rect 31300 22763 31352 22772
rect 31300 22729 31309 22763
rect 31309 22729 31343 22763
rect 31343 22729 31352 22763
rect 31300 22720 31352 22729
rect 31944 22720 31996 22772
rect 32588 22720 32640 22772
rect 33968 22720 34020 22772
rect 30196 22695 30248 22704
rect 30196 22661 30205 22695
rect 30205 22661 30239 22695
rect 30239 22661 30248 22695
rect 30196 22652 30248 22661
rect 17776 22380 17828 22432
rect 20260 22380 20312 22432
rect 23204 22380 23256 22432
rect 25780 22380 25832 22432
rect 29736 22584 29788 22636
rect 32312 22652 32364 22704
rect 31024 22584 31076 22636
rect 31208 22584 31260 22636
rect 31484 22627 31536 22636
rect 31484 22593 31493 22627
rect 31493 22593 31527 22627
rect 31527 22593 31536 22627
rect 31484 22584 31536 22593
rect 32036 22584 32088 22636
rect 32128 22627 32180 22636
rect 32128 22593 32137 22627
rect 32137 22593 32171 22627
rect 32171 22593 32180 22627
rect 32128 22584 32180 22593
rect 32220 22627 32272 22636
rect 32220 22593 32230 22627
rect 32230 22593 32264 22627
rect 32264 22593 32272 22627
rect 32220 22584 32272 22593
rect 32404 22627 32456 22636
rect 32404 22593 32413 22627
rect 32413 22593 32447 22627
rect 32447 22593 32456 22627
rect 32404 22584 32456 22593
rect 32496 22627 32548 22636
rect 32496 22593 32505 22627
rect 32505 22593 32539 22627
rect 32539 22593 32548 22627
rect 32496 22584 32548 22593
rect 32772 22584 32824 22636
rect 31944 22559 31996 22568
rect 31944 22525 31953 22559
rect 31953 22525 31987 22559
rect 31987 22525 31996 22559
rect 31944 22516 31996 22525
rect 30564 22448 30616 22500
rect 30656 22448 30708 22500
rect 28724 22380 28776 22432
rect 29736 22380 29788 22432
rect 33876 22627 33928 22636
rect 33876 22593 33885 22627
rect 33885 22593 33919 22627
rect 33919 22593 33928 22627
rect 33876 22584 33928 22593
rect 34336 22627 34388 22636
rect 34336 22593 34345 22627
rect 34345 22593 34379 22627
rect 34379 22593 34388 22627
rect 34336 22584 34388 22593
rect 34612 22720 34664 22772
rect 35348 22720 35400 22772
rect 35900 22720 35952 22772
rect 35992 22720 36044 22772
rect 34060 22516 34112 22568
rect 34428 22559 34480 22568
rect 34428 22525 34437 22559
rect 34437 22525 34471 22559
rect 34471 22525 34480 22559
rect 34428 22516 34480 22525
rect 34796 22584 34848 22636
rect 35532 22627 35584 22636
rect 35532 22593 35541 22627
rect 35541 22593 35575 22627
rect 35575 22593 35584 22627
rect 35532 22584 35584 22593
rect 35624 22627 35676 22636
rect 35624 22593 35633 22627
rect 35633 22593 35667 22627
rect 35667 22593 35676 22627
rect 35624 22584 35676 22593
rect 35716 22584 35768 22636
rect 36728 22695 36780 22704
rect 36728 22661 36737 22695
rect 36737 22661 36771 22695
rect 36771 22661 36780 22695
rect 36728 22652 36780 22661
rect 36268 22584 36320 22636
rect 36820 22627 36872 22636
rect 36820 22593 36829 22627
rect 36829 22593 36863 22627
rect 36863 22593 36872 22627
rect 36820 22584 36872 22593
rect 34888 22559 34940 22568
rect 34888 22525 34897 22559
rect 34897 22525 34931 22559
rect 34931 22525 34940 22559
rect 34888 22516 34940 22525
rect 33600 22448 33652 22500
rect 34704 22448 34756 22500
rect 36268 22448 36320 22500
rect 32956 22380 33008 22432
rect 35992 22380 36044 22432
rect 37280 22380 37332 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3792 22176 3844 22228
rect 7104 22176 7156 22228
rect 10968 22176 11020 22228
rect 13728 22176 13780 22228
rect 16764 22176 16816 22228
rect 16856 22176 16908 22228
rect 17776 22176 17828 22228
rect 17868 22176 17920 22228
rect 18144 22219 18196 22228
rect 18144 22185 18153 22219
rect 18153 22185 18187 22219
rect 18187 22185 18196 22219
rect 18144 22176 18196 22185
rect 18420 22176 18472 22228
rect 20628 22176 20680 22228
rect 23020 22176 23072 22228
rect 25044 22176 25096 22228
rect 3332 22040 3384 22092
rect 5356 22108 5408 22160
rect 9496 22151 9548 22160
rect 9496 22117 9505 22151
rect 9505 22117 9539 22151
rect 9539 22117 9548 22151
rect 9496 22108 9548 22117
rect 9864 22108 9916 22160
rect 11888 22108 11940 22160
rect 14924 22108 14976 22160
rect 5172 22040 5224 22092
rect 3148 21904 3200 21956
rect 2504 21879 2556 21888
rect 2504 21845 2513 21879
rect 2513 21845 2547 21879
rect 2547 21845 2556 21879
rect 2504 21836 2556 21845
rect 3056 21836 3108 21888
rect 5264 21972 5316 22024
rect 5448 21972 5500 22024
rect 4528 21836 4580 21888
rect 4620 21836 4672 21888
rect 7104 21972 7156 22024
rect 9312 22040 9364 22092
rect 6000 21947 6052 21956
rect 6000 21913 6009 21947
rect 6009 21913 6043 21947
rect 6043 21913 6052 21947
rect 6000 21904 6052 21913
rect 7748 21947 7800 21956
rect 7748 21913 7757 21947
rect 7757 21913 7791 21947
rect 7791 21913 7800 21947
rect 9036 21972 9088 22024
rect 7748 21904 7800 21913
rect 8852 21904 8904 21956
rect 6184 21836 6236 21888
rect 9220 21836 9272 21888
rect 9312 21879 9364 21888
rect 9312 21845 9321 21879
rect 9321 21845 9355 21879
rect 9355 21845 9364 21879
rect 9312 21836 9364 21845
rect 9772 21972 9824 22024
rect 10508 22040 10560 22092
rect 10876 22040 10928 22092
rect 15752 22108 15804 22160
rect 16212 22108 16264 22160
rect 16028 22040 16080 22092
rect 17040 22040 17092 22092
rect 17316 22040 17368 22092
rect 9864 21904 9916 21956
rect 10968 21904 11020 21956
rect 11980 21947 12032 21956
rect 11980 21913 11989 21947
rect 11989 21913 12023 21947
rect 12023 21913 12032 21947
rect 11980 21904 12032 21913
rect 12256 21904 12308 21956
rect 12440 21947 12492 21956
rect 12440 21913 12449 21947
rect 12449 21913 12483 21947
rect 12483 21913 12492 21947
rect 12440 21904 12492 21913
rect 9772 21836 9824 21888
rect 10048 21836 10100 21888
rect 12900 21879 12952 21888
rect 12900 21845 12909 21879
rect 12909 21845 12943 21879
rect 12943 21845 12952 21879
rect 12900 21836 12952 21845
rect 13544 21836 13596 21888
rect 14372 21904 14424 21956
rect 17500 21972 17552 22024
rect 17868 22015 17920 22024
rect 17868 21981 17877 22015
rect 17877 21981 17911 22015
rect 17911 21981 17920 22015
rect 17868 21972 17920 21981
rect 18052 21972 18104 22024
rect 19708 22108 19760 22160
rect 20076 22108 20128 22160
rect 22192 22108 22244 22160
rect 23296 22108 23348 22160
rect 20996 22040 21048 22092
rect 22008 22040 22060 22092
rect 20904 21972 20956 22024
rect 22100 22015 22152 22024
rect 22100 21981 22109 22015
rect 22109 21981 22143 22015
rect 22143 21981 22152 22015
rect 22100 21972 22152 21981
rect 22192 21972 22244 22024
rect 23388 22083 23440 22092
rect 23388 22049 23397 22083
rect 23397 22049 23431 22083
rect 23431 22049 23440 22083
rect 23388 22040 23440 22049
rect 28448 22176 28500 22228
rect 28540 22176 28592 22228
rect 26792 22108 26844 22160
rect 29000 22108 29052 22160
rect 29736 22108 29788 22160
rect 30104 22151 30156 22160
rect 30104 22117 30113 22151
rect 30113 22117 30147 22151
rect 30147 22117 30156 22151
rect 30104 22108 30156 22117
rect 32128 22176 32180 22228
rect 32680 22176 32732 22228
rect 33508 22219 33560 22228
rect 33508 22185 33517 22219
rect 33517 22185 33551 22219
rect 33551 22185 33560 22219
rect 33508 22176 33560 22185
rect 35256 22176 35308 22228
rect 35532 22176 35584 22228
rect 35900 22219 35952 22228
rect 35900 22185 35909 22219
rect 35909 22185 35943 22219
rect 35943 22185 35952 22219
rect 35900 22176 35952 22185
rect 15384 21904 15436 21956
rect 17040 21904 17092 21956
rect 17684 21904 17736 21956
rect 22376 21904 22428 21956
rect 23572 21904 23624 21956
rect 24124 21972 24176 22024
rect 24584 22015 24636 22024
rect 24584 21981 24593 22015
rect 24593 21981 24627 22015
rect 24627 21981 24636 22015
rect 24584 21972 24636 21981
rect 25780 22015 25832 22024
rect 25780 21981 25789 22015
rect 25789 21981 25823 22015
rect 25823 21981 25832 22015
rect 25780 21972 25832 21981
rect 26240 21972 26292 22024
rect 28540 22040 28592 22092
rect 28908 22040 28960 22092
rect 27252 21972 27304 22024
rect 28264 22015 28316 22024
rect 28264 21981 28273 22015
rect 28273 21981 28307 22015
rect 28307 21981 28316 22015
rect 28264 21972 28316 21981
rect 29276 21972 29328 22024
rect 29920 22015 29972 22024
rect 29920 21981 29929 22015
rect 29929 21981 29963 22015
rect 29963 21981 29972 22015
rect 29920 21972 29972 21981
rect 14832 21836 14884 21888
rect 15108 21836 15160 21888
rect 17776 21836 17828 21888
rect 20352 21836 20404 21888
rect 21088 21879 21140 21888
rect 21088 21845 21097 21879
rect 21097 21845 21131 21879
rect 21131 21845 21140 21879
rect 21088 21836 21140 21845
rect 25780 21836 25832 21888
rect 27528 21836 27580 21888
rect 27712 21836 27764 21888
rect 29828 21947 29880 21956
rect 29828 21913 29837 21947
rect 29837 21913 29871 21947
rect 29871 21913 29880 21947
rect 29828 21904 29880 21913
rect 31668 22040 31720 22092
rect 32036 22015 32088 22024
rect 32036 21981 32045 22015
rect 32045 21981 32079 22015
rect 32079 21981 32088 22015
rect 32036 21972 32088 21981
rect 31300 21904 31352 21956
rect 32404 21904 32456 21956
rect 32956 21972 33008 22024
rect 33508 21972 33560 22024
rect 33692 22015 33744 22024
rect 33692 21981 33701 22015
rect 33701 21981 33735 22015
rect 33735 21981 33744 22015
rect 33692 21972 33744 21981
rect 34060 21972 34112 22024
rect 34428 21972 34480 22024
rect 35716 22108 35768 22160
rect 34612 22040 34664 22092
rect 35164 22015 35216 22024
rect 35164 21981 35173 22015
rect 35173 21981 35207 22015
rect 35207 21981 35216 22015
rect 35164 21972 35216 21981
rect 30104 21836 30156 21888
rect 32496 21836 32548 21888
rect 34704 21836 34756 21888
rect 34796 21836 34848 21888
rect 35164 21836 35216 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 2504 21632 2556 21684
rect 5264 21632 5316 21684
rect 6000 21632 6052 21684
rect 9312 21632 9364 21684
rect 10692 21632 10744 21684
rect 1768 21539 1820 21548
rect 1768 21505 1777 21539
rect 1777 21505 1811 21539
rect 1811 21505 1820 21539
rect 1768 21496 1820 21505
rect 3056 21607 3108 21616
rect 3056 21573 3065 21607
rect 3065 21573 3099 21607
rect 3099 21573 3108 21607
rect 3056 21564 3108 21573
rect 3792 21564 3844 21616
rect 4528 21564 4580 21616
rect 2780 21539 2832 21548
rect 2780 21505 2789 21539
rect 2789 21505 2823 21539
rect 2823 21505 2832 21539
rect 2780 21496 2832 21505
rect 5540 21539 5592 21548
rect 5540 21505 5549 21539
rect 5549 21505 5583 21539
rect 5583 21505 5592 21539
rect 5540 21496 5592 21505
rect 6092 21496 6144 21548
rect 6552 21539 6604 21548
rect 6552 21505 6561 21539
rect 6561 21505 6595 21539
rect 6595 21505 6604 21539
rect 6552 21496 6604 21505
rect 9220 21564 9272 21616
rect 11520 21632 11572 21684
rect 8116 21428 8168 21480
rect 8208 21360 8260 21412
rect 8484 21360 8536 21412
rect 8576 21360 8628 21412
rect 9496 21496 9548 21548
rect 10968 21607 11020 21616
rect 10968 21573 10977 21607
rect 10977 21573 11011 21607
rect 11011 21573 11020 21607
rect 10968 21564 11020 21573
rect 10692 21539 10744 21548
rect 10692 21505 10701 21539
rect 10701 21505 10735 21539
rect 10735 21505 10744 21539
rect 10692 21496 10744 21505
rect 11704 21564 11756 21616
rect 13452 21607 13504 21616
rect 13452 21573 13461 21607
rect 13461 21573 13495 21607
rect 13495 21573 13504 21607
rect 13452 21564 13504 21573
rect 13728 21564 13780 21616
rect 14832 21632 14884 21684
rect 16028 21632 16080 21684
rect 17316 21675 17368 21684
rect 17316 21641 17325 21675
rect 17325 21641 17359 21675
rect 17359 21641 17368 21675
rect 17316 21632 17368 21641
rect 17500 21632 17552 21684
rect 18236 21675 18288 21684
rect 18236 21641 18245 21675
rect 18245 21641 18279 21675
rect 18279 21641 18288 21675
rect 18236 21632 18288 21641
rect 17868 21607 17920 21616
rect 9036 21360 9088 21412
rect 9772 21471 9824 21480
rect 9772 21437 9781 21471
rect 9781 21437 9815 21471
rect 9815 21437 9824 21471
rect 9772 21428 9824 21437
rect 9956 21471 10008 21480
rect 9956 21437 9965 21471
rect 9965 21437 9999 21471
rect 9999 21437 10008 21471
rect 9956 21428 10008 21437
rect 10324 21428 10376 21480
rect 10692 21360 10744 21412
rect 11612 21539 11664 21548
rect 11612 21505 11621 21539
rect 11621 21505 11655 21539
rect 11655 21505 11664 21539
rect 11612 21496 11664 21505
rect 11980 21539 12032 21548
rect 11980 21505 11989 21539
rect 11989 21505 12023 21539
rect 12023 21505 12032 21539
rect 11980 21496 12032 21505
rect 12256 21496 12308 21548
rect 13636 21539 13688 21548
rect 13636 21505 13645 21539
rect 13645 21505 13679 21539
rect 13679 21505 13688 21539
rect 13636 21496 13688 21505
rect 13820 21539 13872 21548
rect 13820 21505 13829 21539
rect 13829 21505 13863 21539
rect 13863 21505 13872 21539
rect 13820 21496 13872 21505
rect 11980 21360 12032 21412
rect 13820 21360 13872 21412
rect 14188 21496 14240 21548
rect 14924 21496 14976 21548
rect 15292 21496 15344 21548
rect 17868 21573 17877 21607
rect 17877 21573 17911 21607
rect 17911 21573 17920 21607
rect 17868 21564 17920 21573
rect 17500 21496 17552 21548
rect 20812 21632 20864 21684
rect 21180 21632 21232 21684
rect 23204 21632 23256 21684
rect 23388 21632 23440 21684
rect 24584 21632 24636 21684
rect 25780 21675 25832 21684
rect 25780 21641 25805 21675
rect 25805 21641 25832 21675
rect 25780 21632 25832 21641
rect 26516 21632 26568 21684
rect 26608 21675 26660 21684
rect 26608 21641 26617 21675
rect 26617 21641 26651 21675
rect 26651 21641 26660 21675
rect 26608 21632 26660 21641
rect 27160 21632 27212 21684
rect 27620 21675 27672 21684
rect 27620 21641 27629 21675
rect 27629 21641 27663 21675
rect 27663 21641 27672 21675
rect 27620 21632 27672 21641
rect 28264 21632 28316 21684
rect 29644 21632 29696 21684
rect 29920 21632 29972 21684
rect 34888 21632 34940 21684
rect 21916 21564 21968 21616
rect 15108 21360 15160 21412
rect 17316 21428 17368 21480
rect 16028 21360 16080 21412
rect 16120 21403 16172 21412
rect 16120 21369 16129 21403
rect 16129 21369 16163 21403
rect 16163 21369 16172 21403
rect 16120 21360 16172 21369
rect 19432 21539 19484 21548
rect 19432 21505 19441 21539
rect 19441 21505 19475 21539
rect 19475 21505 19484 21539
rect 19432 21496 19484 21505
rect 19708 21496 19760 21548
rect 20352 21496 20404 21548
rect 20628 21539 20680 21548
rect 20628 21505 20637 21539
rect 20637 21505 20671 21539
rect 20671 21505 20680 21539
rect 20628 21496 20680 21505
rect 20812 21539 20864 21548
rect 20812 21505 20821 21539
rect 20821 21505 20855 21539
rect 20855 21505 20864 21539
rect 20812 21496 20864 21505
rect 22744 21496 22796 21548
rect 23296 21539 23348 21548
rect 23296 21505 23305 21539
rect 23305 21505 23339 21539
rect 23339 21505 23348 21539
rect 23296 21496 23348 21505
rect 25136 21564 25188 21616
rect 25596 21607 25648 21616
rect 25596 21573 25605 21607
rect 25605 21573 25639 21607
rect 25639 21573 25648 21607
rect 25596 21564 25648 21573
rect 24860 21496 24912 21548
rect 25872 21496 25924 21548
rect 27252 21539 27304 21548
rect 27252 21505 27261 21539
rect 27261 21505 27295 21539
rect 27295 21505 27304 21539
rect 27252 21496 27304 21505
rect 27988 21539 28040 21548
rect 27988 21505 27997 21539
rect 27997 21505 28031 21539
rect 28031 21505 28040 21539
rect 27988 21496 28040 21505
rect 24124 21471 24176 21480
rect 940 21292 992 21344
rect 1860 21292 1912 21344
rect 7748 21292 7800 21344
rect 9956 21292 10008 21344
rect 10140 21335 10192 21344
rect 10140 21301 10149 21335
rect 10149 21301 10183 21335
rect 10183 21301 10192 21335
rect 10140 21292 10192 21301
rect 10600 21335 10652 21344
rect 10600 21301 10609 21335
rect 10609 21301 10643 21335
rect 10643 21301 10652 21335
rect 10600 21292 10652 21301
rect 11152 21335 11204 21344
rect 11152 21301 11161 21335
rect 11161 21301 11195 21335
rect 11195 21301 11204 21335
rect 11152 21292 11204 21301
rect 13636 21292 13688 21344
rect 14004 21292 14056 21344
rect 14648 21292 14700 21344
rect 16672 21335 16724 21344
rect 16672 21301 16681 21335
rect 16681 21301 16715 21335
rect 16715 21301 16724 21335
rect 16672 21292 16724 21301
rect 17500 21292 17552 21344
rect 18052 21292 18104 21344
rect 19800 21292 19852 21344
rect 21088 21360 21140 21412
rect 24124 21437 24133 21471
rect 24133 21437 24167 21471
rect 24167 21437 24176 21471
rect 24124 21428 24176 21437
rect 26240 21471 26292 21480
rect 26240 21437 26249 21471
rect 26249 21437 26283 21471
rect 26283 21437 26292 21471
rect 26240 21428 26292 21437
rect 26332 21471 26384 21480
rect 26332 21437 26341 21471
rect 26341 21437 26375 21471
rect 26375 21437 26384 21471
rect 26332 21428 26384 21437
rect 26516 21428 26568 21480
rect 28724 21539 28776 21548
rect 28724 21505 28733 21539
rect 28733 21505 28767 21539
rect 28767 21505 28776 21539
rect 28724 21496 28776 21505
rect 29000 21496 29052 21548
rect 29644 21539 29696 21548
rect 29644 21505 29653 21539
rect 29653 21505 29687 21539
rect 29687 21505 29696 21539
rect 29644 21496 29696 21505
rect 30840 21564 30892 21616
rect 35164 21632 35216 21684
rect 36820 21632 36872 21684
rect 31484 21496 31536 21548
rect 34520 21496 34572 21548
rect 36912 21539 36964 21548
rect 36912 21505 36921 21539
rect 36921 21505 36955 21539
rect 36955 21505 36964 21539
rect 36912 21496 36964 21505
rect 37096 21539 37148 21548
rect 37096 21505 37105 21539
rect 37105 21505 37139 21539
rect 37139 21505 37148 21539
rect 37096 21496 37148 21505
rect 37648 21539 37700 21548
rect 37648 21505 37657 21539
rect 37657 21505 37691 21539
rect 37691 21505 37700 21539
rect 37648 21496 37700 21505
rect 28632 21428 28684 21480
rect 28816 21428 28868 21480
rect 25596 21292 25648 21344
rect 27620 21360 27672 21412
rect 30104 21360 30156 21412
rect 27344 21292 27396 21344
rect 28448 21292 28500 21344
rect 31576 21292 31628 21344
rect 34152 21292 34204 21344
rect 37832 21335 37884 21344
rect 37832 21301 37841 21335
rect 37841 21301 37875 21335
rect 37875 21301 37884 21335
rect 37832 21292 37884 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1860 21088 1912 21140
rect 6092 21131 6144 21140
rect 6092 21097 6101 21131
rect 6101 21097 6135 21131
rect 6135 21097 6144 21131
rect 6092 21088 6144 21097
rect 8208 21088 8260 21140
rect 10692 21088 10744 21140
rect 11152 21088 11204 21140
rect 12900 21088 12952 21140
rect 13820 21088 13872 21140
rect 2780 21020 2832 21072
rect 10140 21020 10192 21072
rect 1400 20995 1452 21004
rect 1400 20961 1409 20995
rect 1409 20961 1443 20995
rect 1443 20961 1452 20995
rect 1400 20952 1452 20961
rect 4068 20952 4120 21004
rect 4620 20859 4672 20868
rect 4620 20825 4629 20859
rect 4629 20825 4663 20859
rect 4663 20825 4672 20859
rect 4620 20816 4672 20825
rect 8024 20927 8076 20936
rect 8024 20893 8033 20927
rect 8033 20893 8067 20927
rect 8067 20893 8076 20927
rect 8024 20884 8076 20893
rect 3148 20791 3200 20800
rect 3148 20757 3157 20791
rect 3157 20757 3191 20791
rect 3191 20757 3200 20791
rect 3148 20748 3200 20757
rect 3792 20748 3844 20800
rect 9036 20816 9088 20868
rect 10600 20884 10652 20936
rect 10876 20884 10928 20936
rect 11704 20952 11756 21004
rect 13544 20952 13596 21004
rect 14004 21020 14056 21072
rect 11612 20927 11664 20936
rect 11612 20893 11621 20927
rect 11621 20893 11655 20927
rect 11655 20893 11664 20927
rect 11612 20884 11664 20893
rect 10324 20816 10376 20868
rect 14372 20927 14424 20936
rect 14372 20893 14381 20927
rect 14381 20893 14415 20927
rect 14415 20893 14424 20927
rect 14372 20884 14424 20893
rect 14648 20927 14700 20936
rect 14648 20893 14656 20927
rect 14656 20893 14690 20927
rect 14690 20893 14700 20927
rect 14648 20884 14700 20893
rect 16672 21088 16724 21140
rect 20628 21088 20680 21140
rect 15292 20884 15344 20936
rect 21272 21088 21324 21140
rect 22560 21088 22612 21140
rect 25412 21131 25464 21140
rect 25412 21097 25421 21131
rect 25421 21097 25455 21131
rect 25455 21097 25464 21131
rect 25412 21088 25464 21097
rect 12348 20859 12400 20868
rect 12348 20825 12357 20859
rect 12357 20825 12391 20859
rect 12391 20825 12400 20859
rect 12348 20816 12400 20825
rect 14832 20816 14884 20868
rect 15476 20816 15528 20868
rect 20904 21020 20956 21072
rect 28724 21088 28776 21140
rect 30656 21088 30708 21140
rect 25596 21020 25648 21072
rect 27344 21020 27396 21072
rect 27620 21020 27672 21072
rect 28816 21020 28868 21072
rect 19340 20884 19392 20936
rect 6184 20748 6236 20800
rect 10416 20748 10468 20800
rect 11152 20748 11204 20800
rect 12256 20748 12308 20800
rect 19708 20884 19760 20936
rect 25136 20952 25188 21004
rect 25228 20995 25280 21004
rect 25228 20961 25237 20995
rect 25237 20961 25271 20995
rect 25271 20961 25280 20995
rect 25228 20952 25280 20961
rect 21088 20884 21140 20936
rect 21640 20884 21692 20936
rect 24032 20884 24084 20936
rect 24768 20816 24820 20868
rect 25780 20816 25832 20868
rect 30288 21020 30340 21072
rect 31852 21088 31904 21140
rect 32404 21088 32456 21140
rect 33692 21088 33744 21140
rect 29828 20952 29880 21004
rect 30196 20952 30248 21004
rect 27712 20884 27764 20936
rect 29644 20884 29696 20936
rect 31576 21020 31628 21072
rect 31760 21020 31812 21072
rect 15568 20748 15620 20800
rect 16304 20748 16356 20800
rect 17316 20748 17368 20800
rect 19432 20748 19484 20800
rect 20720 20748 20772 20800
rect 21456 20748 21508 20800
rect 22560 20748 22612 20800
rect 23480 20748 23532 20800
rect 24216 20748 24268 20800
rect 25504 20748 25556 20800
rect 26792 20748 26844 20800
rect 31024 20884 31076 20936
rect 31116 20927 31168 20936
rect 31116 20893 31125 20927
rect 31125 20893 31159 20927
rect 31159 20893 31168 20927
rect 31116 20884 31168 20893
rect 31300 20884 31352 20936
rect 33324 20995 33376 21004
rect 33324 20961 33333 20995
rect 33333 20961 33367 20995
rect 33367 20961 33376 20995
rect 33324 20952 33376 20961
rect 33876 20952 33928 21004
rect 34244 21020 34296 21072
rect 34428 21063 34480 21072
rect 34428 21029 34437 21063
rect 34437 21029 34471 21063
rect 34471 21029 34480 21063
rect 34428 21020 34480 21029
rect 34704 21131 34756 21140
rect 34704 21097 34713 21131
rect 34713 21097 34747 21131
rect 34747 21097 34756 21131
rect 34704 21088 34756 21097
rect 37188 21088 37240 21140
rect 32864 20884 32916 20936
rect 33232 20884 33284 20936
rect 33416 20927 33468 20936
rect 33416 20893 33425 20927
rect 33425 20893 33459 20927
rect 33459 20893 33468 20927
rect 33416 20884 33468 20893
rect 30564 20816 30616 20868
rect 31484 20859 31536 20868
rect 31484 20825 31493 20859
rect 31493 20825 31527 20859
rect 31527 20825 31536 20859
rect 31484 20816 31536 20825
rect 31576 20816 31628 20868
rect 34520 20952 34572 21004
rect 36912 21063 36964 21072
rect 36912 21029 36921 21063
rect 36921 21029 36955 21063
rect 36955 21029 36964 21063
rect 36912 21020 36964 21029
rect 36820 20995 36872 21004
rect 36820 20961 36829 20995
rect 36829 20961 36863 20995
rect 36863 20961 36872 20995
rect 36820 20952 36872 20961
rect 34152 20884 34204 20936
rect 34428 20884 34480 20936
rect 34612 20816 34664 20868
rect 35992 20884 36044 20936
rect 36912 20884 36964 20936
rect 37188 20927 37240 20936
rect 37188 20893 37197 20927
rect 37197 20893 37231 20927
rect 37231 20893 37240 20927
rect 37188 20884 37240 20893
rect 30380 20748 30432 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 9680 20544 9732 20596
rect 9772 20587 9824 20596
rect 9772 20553 9781 20587
rect 9781 20553 9815 20587
rect 9815 20553 9824 20587
rect 9772 20544 9824 20553
rect 10232 20544 10284 20596
rect 11612 20544 11664 20596
rect 17224 20544 17276 20596
rect 19524 20544 19576 20596
rect 20536 20544 20588 20596
rect 21272 20544 21324 20596
rect 21456 20544 21508 20596
rect 23940 20587 23992 20596
rect 23940 20553 23949 20587
rect 23949 20553 23983 20587
rect 23983 20553 23992 20587
rect 23940 20544 23992 20553
rect 24032 20587 24084 20596
rect 24032 20553 24041 20587
rect 24041 20553 24075 20587
rect 24075 20553 24084 20587
rect 24032 20544 24084 20553
rect 24400 20587 24452 20596
rect 24400 20553 24409 20587
rect 24409 20553 24443 20587
rect 24443 20553 24452 20587
rect 24400 20544 24452 20553
rect 24768 20544 24820 20596
rect 27804 20544 27856 20596
rect 28632 20544 28684 20596
rect 6828 20476 6880 20528
rect 7932 20476 7984 20528
rect 8300 20476 8352 20528
rect 8484 20519 8536 20528
rect 8484 20485 8493 20519
rect 8493 20485 8527 20519
rect 8527 20485 8536 20519
rect 8484 20476 8536 20485
rect 8208 20408 8260 20460
rect 9128 20340 9180 20392
rect 9404 20408 9456 20460
rect 10416 20408 10468 20460
rect 10876 20408 10928 20460
rect 10968 20408 11020 20460
rect 15200 20476 15252 20528
rect 12532 20408 12584 20460
rect 13084 20451 13136 20460
rect 13084 20417 13093 20451
rect 13093 20417 13127 20451
rect 13127 20417 13136 20451
rect 13084 20408 13136 20417
rect 8116 20272 8168 20324
rect 10784 20383 10836 20392
rect 10784 20349 10793 20383
rect 10793 20349 10827 20383
rect 10827 20349 10836 20383
rect 10784 20340 10836 20349
rect 13176 20340 13228 20392
rect 13912 20451 13964 20460
rect 13912 20417 13921 20451
rect 13921 20417 13955 20451
rect 13955 20417 13964 20451
rect 13912 20408 13964 20417
rect 15660 20451 15712 20460
rect 15660 20417 15669 20451
rect 15669 20417 15703 20451
rect 15703 20417 15712 20451
rect 15660 20408 15712 20417
rect 16120 20408 16172 20460
rect 19340 20476 19392 20528
rect 17132 20451 17184 20460
rect 17132 20417 17141 20451
rect 17141 20417 17175 20451
rect 17175 20417 17184 20451
rect 17132 20408 17184 20417
rect 17776 20451 17828 20460
rect 17776 20417 17785 20451
rect 17785 20417 17819 20451
rect 17819 20417 17828 20451
rect 17776 20408 17828 20417
rect 18144 20408 18196 20460
rect 6460 20247 6512 20256
rect 6460 20213 6469 20247
rect 6469 20213 6503 20247
rect 6503 20213 6512 20247
rect 6460 20204 6512 20213
rect 8024 20204 8076 20256
rect 8576 20204 8628 20256
rect 9128 20247 9180 20256
rect 9128 20213 9137 20247
rect 9137 20213 9171 20247
rect 9171 20213 9180 20247
rect 9128 20204 9180 20213
rect 12164 20272 12216 20324
rect 12440 20272 12492 20324
rect 12532 20272 12584 20324
rect 18604 20340 18656 20392
rect 19432 20451 19484 20460
rect 19432 20417 19441 20451
rect 19441 20417 19475 20451
rect 19475 20417 19484 20451
rect 19432 20408 19484 20417
rect 19616 20408 19668 20460
rect 19800 20408 19852 20460
rect 22560 20451 22612 20460
rect 22560 20417 22569 20451
rect 22569 20417 22603 20451
rect 22603 20417 22612 20451
rect 22560 20408 22612 20417
rect 20720 20383 20772 20392
rect 20720 20349 20729 20383
rect 20729 20349 20763 20383
rect 20763 20349 20772 20383
rect 20720 20340 20772 20349
rect 20904 20383 20956 20392
rect 20904 20349 20913 20383
rect 20913 20349 20947 20383
rect 20947 20349 20956 20383
rect 20904 20340 20956 20349
rect 25780 20476 25832 20528
rect 26056 20519 26108 20528
rect 26056 20485 26065 20519
rect 26065 20485 26099 20519
rect 26099 20485 26108 20519
rect 26056 20476 26108 20485
rect 24676 20408 24728 20460
rect 24860 20408 24912 20460
rect 26976 20408 27028 20460
rect 30012 20544 30064 20596
rect 30196 20587 30248 20596
rect 30196 20553 30205 20587
rect 30205 20553 30239 20587
rect 30239 20553 30248 20587
rect 30196 20544 30248 20553
rect 31576 20544 31628 20596
rect 31392 20476 31444 20528
rect 33508 20544 33560 20596
rect 33784 20544 33836 20596
rect 34060 20587 34112 20596
rect 34060 20553 34069 20587
rect 34069 20553 34103 20587
rect 34103 20553 34112 20587
rect 34060 20544 34112 20553
rect 37096 20587 37148 20596
rect 37096 20553 37105 20587
rect 37105 20553 37139 20587
rect 37139 20553 37148 20587
rect 37096 20544 37148 20553
rect 33324 20476 33376 20528
rect 33416 20476 33468 20528
rect 36820 20476 36872 20528
rect 36912 20519 36964 20528
rect 36912 20485 36937 20519
rect 36937 20485 36964 20519
rect 36912 20476 36964 20485
rect 24216 20340 24268 20392
rect 29460 20408 29512 20460
rect 29644 20408 29696 20460
rect 30012 20408 30064 20460
rect 30104 20451 30156 20460
rect 30104 20417 30113 20451
rect 30113 20417 30147 20451
rect 30147 20417 30156 20451
rect 30104 20408 30156 20417
rect 30288 20408 30340 20460
rect 30472 20451 30524 20460
rect 30472 20417 30481 20451
rect 30481 20417 30515 20451
rect 30515 20417 30524 20451
rect 30472 20408 30524 20417
rect 30656 20408 30708 20460
rect 31208 20408 31260 20460
rect 30932 20340 30984 20392
rect 31300 20340 31352 20392
rect 33968 20451 34020 20460
rect 33968 20417 33977 20451
rect 33977 20417 34011 20451
rect 34011 20417 34020 20451
rect 33968 20408 34020 20417
rect 11060 20247 11112 20256
rect 11060 20213 11069 20247
rect 11069 20213 11103 20247
rect 11103 20213 11112 20247
rect 11060 20204 11112 20213
rect 15844 20247 15896 20256
rect 15844 20213 15853 20247
rect 15853 20213 15887 20247
rect 15887 20213 15896 20247
rect 15844 20204 15896 20213
rect 17500 20247 17552 20256
rect 17500 20213 17509 20247
rect 17509 20213 17543 20247
rect 17543 20213 17552 20247
rect 17500 20204 17552 20213
rect 17592 20204 17644 20256
rect 19432 20204 19484 20256
rect 19984 20204 20036 20256
rect 21548 20204 21600 20256
rect 22192 20247 22244 20256
rect 22192 20213 22201 20247
rect 22201 20213 22235 20247
rect 22235 20213 22244 20247
rect 22192 20204 22244 20213
rect 22284 20204 22336 20256
rect 27068 20204 27120 20256
rect 30656 20204 30708 20256
rect 30932 20204 30984 20256
rect 31208 20272 31260 20324
rect 31852 20340 31904 20392
rect 33232 20340 33284 20392
rect 33784 20340 33836 20392
rect 33876 20340 33928 20392
rect 33140 20204 33192 20256
rect 33232 20204 33284 20256
rect 36544 20204 36596 20256
rect 37188 20204 37240 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 7932 20043 7984 20052
rect 7932 20009 7941 20043
rect 7941 20009 7975 20043
rect 7975 20009 7984 20043
rect 7932 20000 7984 20009
rect 9772 20000 9824 20052
rect 13912 20000 13964 20052
rect 14280 20000 14332 20052
rect 5448 19932 5500 19984
rect 3332 19864 3384 19916
rect 4068 19864 4120 19916
rect 6184 19907 6236 19916
rect 6184 19873 6193 19907
rect 6193 19873 6227 19907
rect 6227 19873 6236 19907
rect 6184 19864 6236 19873
rect 6460 19907 6512 19916
rect 6460 19873 6469 19907
rect 6469 19873 6503 19907
rect 6503 19873 6512 19907
rect 6460 19864 6512 19873
rect 9680 19796 9732 19848
rect 9772 19839 9824 19848
rect 9772 19805 9781 19839
rect 9781 19805 9815 19839
rect 9815 19805 9824 19839
rect 9772 19796 9824 19805
rect 9864 19839 9916 19848
rect 9864 19805 9873 19839
rect 9873 19805 9907 19839
rect 9907 19805 9916 19839
rect 9864 19796 9916 19805
rect 11060 19796 11112 19848
rect 11612 19796 11664 19848
rect 11888 19796 11940 19848
rect 13452 19932 13504 19984
rect 19800 20000 19852 20052
rect 20904 20000 20956 20052
rect 24216 20000 24268 20052
rect 24400 20000 24452 20052
rect 3332 19728 3384 19780
rect 4068 19771 4120 19780
rect 4068 19737 4077 19771
rect 4077 19737 4111 19771
rect 4111 19737 4120 19771
rect 4068 19728 4120 19737
rect 1952 19703 2004 19712
rect 1952 19669 1961 19703
rect 1961 19669 1995 19703
rect 1995 19669 2004 19703
rect 1952 19660 2004 19669
rect 3148 19660 3200 19712
rect 6000 19728 6052 19780
rect 4804 19660 4856 19712
rect 8300 19728 8352 19780
rect 9312 19728 9364 19780
rect 12532 19839 12584 19848
rect 12532 19805 12541 19839
rect 12541 19805 12575 19839
rect 12575 19805 12584 19839
rect 12532 19796 12584 19805
rect 13084 19839 13136 19848
rect 13084 19805 13093 19839
rect 13093 19805 13127 19839
rect 13127 19805 13136 19839
rect 13084 19796 13136 19805
rect 13176 19839 13228 19848
rect 13176 19805 13185 19839
rect 13185 19805 13219 19839
rect 13219 19805 13228 19839
rect 13176 19796 13228 19805
rect 17500 19932 17552 19984
rect 17868 19932 17920 19984
rect 19156 19932 19208 19984
rect 16948 19907 17000 19916
rect 10324 19703 10376 19712
rect 10324 19669 10333 19703
rect 10333 19669 10367 19703
rect 10367 19669 10376 19703
rect 10324 19660 10376 19669
rect 10416 19703 10468 19712
rect 10416 19669 10425 19703
rect 10425 19669 10459 19703
rect 10459 19669 10468 19703
rect 10416 19660 10468 19669
rect 16948 19873 16957 19907
rect 16957 19873 16991 19907
rect 16991 19873 17000 19907
rect 16948 19864 17000 19873
rect 19984 19907 20036 19916
rect 14372 19796 14424 19848
rect 15108 19839 15160 19848
rect 15108 19805 15117 19839
rect 15117 19805 15151 19839
rect 15151 19805 15160 19839
rect 15108 19796 15160 19805
rect 15660 19839 15712 19848
rect 14648 19660 14700 19712
rect 14832 19660 14884 19712
rect 15660 19805 15669 19839
rect 15669 19805 15703 19839
rect 15703 19805 15712 19839
rect 15660 19796 15712 19805
rect 16120 19839 16172 19848
rect 16120 19805 16129 19839
rect 16129 19805 16163 19839
rect 16163 19805 16172 19839
rect 16120 19796 16172 19805
rect 16488 19796 16540 19848
rect 19984 19873 19993 19907
rect 19993 19873 20027 19907
rect 20027 19873 20036 19907
rect 19984 19864 20036 19873
rect 20720 19932 20772 19984
rect 20996 19932 21048 19984
rect 17868 19839 17920 19848
rect 17868 19805 17877 19839
rect 17877 19805 17911 19839
rect 17911 19805 17920 19839
rect 17868 19796 17920 19805
rect 19064 19839 19116 19848
rect 19064 19805 19073 19839
rect 19073 19805 19107 19839
rect 19107 19805 19116 19839
rect 19064 19796 19116 19805
rect 19340 19796 19392 19848
rect 20628 19796 20680 19848
rect 17776 19728 17828 19780
rect 15476 19703 15528 19712
rect 15476 19669 15485 19703
rect 15485 19669 15519 19703
rect 15519 19669 15528 19703
rect 15476 19660 15528 19669
rect 15752 19660 15804 19712
rect 17224 19703 17276 19712
rect 17224 19669 17233 19703
rect 17233 19669 17267 19703
rect 17267 19669 17276 19703
rect 17224 19660 17276 19669
rect 17408 19660 17460 19712
rect 18328 19728 18380 19780
rect 19248 19728 19300 19780
rect 19616 19728 19668 19780
rect 19800 19728 19852 19780
rect 21180 19771 21232 19780
rect 21180 19737 21189 19771
rect 21189 19737 21223 19771
rect 21223 19737 21232 19771
rect 21180 19728 21232 19737
rect 19340 19660 19392 19712
rect 21824 19839 21876 19848
rect 21824 19805 21833 19839
rect 21833 19805 21867 19839
rect 21867 19805 21876 19839
rect 21824 19796 21876 19805
rect 24584 19907 24636 19916
rect 24584 19873 24593 19907
rect 24593 19873 24627 19907
rect 24627 19873 24636 19907
rect 24584 19864 24636 19873
rect 24860 19796 24912 19848
rect 27252 20000 27304 20052
rect 29184 20000 29236 20052
rect 30288 20000 30340 20052
rect 30380 20043 30432 20052
rect 30380 20009 30389 20043
rect 30389 20009 30423 20043
rect 30423 20009 30432 20043
rect 30380 20000 30432 20009
rect 30564 20043 30616 20052
rect 30564 20009 30573 20043
rect 30573 20009 30607 20043
rect 30607 20009 30616 20043
rect 30564 20000 30616 20009
rect 31116 20000 31168 20052
rect 26516 19932 26568 19984
rect 26240 19864 26292 19916
rect 25228 19839 25280 19848
rect 25228 19805 25237 19839
rect 25237 19805 25271 19839
rect 25271 19805 25280 19839
rect 25228 19796 25280 19805
rect 27252 19839 27304 19848
rect 27252 19805 27261 19839
rect 27261 19805 27295 19839
rect 27295 19805 27304 19839
rect 27252 19796 27304 19805
rect 27344 19796 27396 19848
rect 27804 19796 27856 19848
rect 29092 19932 29144 19984
rect 30748 19932 30800 19984
rect 28172 19864 28224 19916
rect 24032 19728 24084 19780
rect 24952 19728 25004 19780
rect 25044 19728 25096 19780
rect 28632 19839 28684 19848
rect 28632 19805 28641 19839
rect 28641 19805 28675 19839
rect 28675 19805 28684 19839
rect 28632 19796 28684 19805
rect 29460 19796 29512 19848
rect 30196 19864 30248 19916
rect 30104 19796 30156 19848
rect 31760 19932 31812 19984
rect 30932 19864 30984 19916
rect 23664 19660 23716 19712
rect 25136 19703 25188 19712
rect 25136 19669 25145 19703
rect 25145 19669 25179 19703
rect 25179 19669 25188 19703
rect 25136 19660 25188 19669
rect 26332 19660 26384 19712
rect 27252 19660 27304 19712
rect 30012 19728 30064 19780
rect 30288 19728 30340 19780
rect 31208 19907 31260 19916
rect 31208 19873 31217 19907
rect 31217 19873 31251 19907
rect 31251 19873 31260 19907
rect 31208 19864 31260 19873
rect 31300 19839 31352 19848
rect 31300 19805 31309 19839
rect 31309 19805 31343 19839
rect 31343 19805 31352 19839
rect 31300 19796 31352 19805
rect 33232 19975 33284 19984
rect 33232 19941 33241 19975
rect 33241 19941 33275 19975
rect 33275 19941 33284 19975
rect 33232 19932 33284 19941
rect 33968 20000 34020 20052
rect 34796 20043 34848 20052
rect 34796 20009 34805 20043
rect 34805 20009 34839 20043
rect 34839 20009 34848 20043
rect 34796 20000 34848 20009
rect 35348 20000 35400 20052
rect 35164 19932 35216 19984
rect 33876 19864 33928 19916
rect 34520 19864 34572 19916
rect 35256 19907 35308 19916
rect 35256 19873 35265 19907
rect 35265 19873 35299 19907
rect 35299 19873 35308 19907
rect 35256 19864 35308 19873
rect 31668 19728 31720 19780
rect 35072 19796 35124 19848
rect 36084 20043 36136 20052
rect 36084 20009 36093 20043
rect 36093 20009 36127 20043
rect 36127 20009 36136 20043
rect 36084 20000 36136 20009
rect 36544 20043 36596 20052
rect 36544 20009 36553 20043
rect 36553 20009 36587 20043
rect 36587 20009 36596 20043
rect 36544 20000 36596 20009
rect 36636 20000 36688 20052
rect 35992 19796 36044 19848
rect 30656 19660 30708 19712
rect 33416 19660 33468 19712
rect 35440 19660 35492 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 4068 19499 4120 19508
rect 4068 19465 4077 19499
rect 4077 19465 4111 19499
rect 4111 19465 4120 19499
rect 4068 19456 4120 19465
rect 1952 19388 2004 19440
rect 3148 19388 3200 19440
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 4804 19499 4856 19508
rect 4804 19465 4813 19499
rect 4813 19465 4847 19499
rect 4847 19465 4856 19499
rect 4804 19456 4856 19465
rect 5816 19456 5868 19508
rect 6828 19456 6880 19508
rect 11888 19456 11940 19508
rect 4712 19431 4764 19440
rect 4712 19397 4721 19431
rect 4721 19397 4755 19431
rect 4755 19397 4764 19431
rect 4712 19388 4764 19397
rect 9496 19388 9548 19440
rect 10692 19388 10744 19440
rect 11612 19388 11664 19440
rect 14556 19456 14608 19508
rect 15108 19456 15160 19508
rect 8024 19320 8076 19372
rect 9680 19363 9732 19372
rect 9680 19329 9689 19363
rect 9689 19329 9723 19363
rect 9723 19329 9732 19363
rect 9680 19320 9732 19329
rect 9772 19320 9824 19372
rect 3240 19252 3292 19304
rect 5356 19252 5408 19304
rect 9864 19252 9916 19304
rect 10140 19252 10192 19304
rect 11888 19320 11940 19372
rect 11980 19320 12032 19372
rect 12900 19363 12952 19372
rect 10508 19252 10560 19304
rect 10600 19252 10652 19304
rect 11060 19184 11112 19236
rect 3332 19116 3384 19168
rect 6368 19159 6420 19168
rect 6368 19125 6377 19159
rect 6377 19125 6411 19159
rect 6411 19125 6420 19159
rect 6368 19116 6420 19125
rect 7748 19116 7800 19168
rect 8484 19116 8536 19168
rect 11980 19159 12032 19168
rect 11980 19125 11989 19159
rect 11989 19125 12023 19159
rect 12023 19125 12032 19159
rect 11980 19116 12032 19125
rect 12900 19329 12909 19363
rect 12909 19329 12943 19363
rect 12943 19329 12952 19363
rect 12900 19320 12952 19329
rect 13176 19320 13228 19372
rect 13728 19388 13780 19440
rect 13452 19320 13504 19372
rect 15292 19363 15344 19372
rect 15292 19329 15301 19363
rect 15301 19329 15335 19363
rect 15335 19329 15344 19363
rect 15292 19320 15344 19329
rect 17224 19456 17276 19508
rect 15660 19388 15712 19440
rect 17592 19388 17644 19440
rect 18328 19388 18380 19440
rect 21824 19456 21876 19508
rect 22192 19456 22244 19508
rect 25044 19499 25096 19508
rect 25044 19465 25053 19499
rect 25053 19465 25087 19499
rect 25087 19465 25096 19499
rect 25044 19456 25096 19465
rect 25228 19456 25280 19508
rect 19064 19388 19116 19440
rect 26976 19499 27028 19508
rect 26976 19465 26985 19499
rect 26985 19465 27019 19499
rect 27019 19465 27028 19499
rect 26976 19456 27028 19465
rect 30380 19456 30432 19508
rect 30656 19456 30708 19508
rect 31208 19456 31260 19508
rect 35072 19499 35124 19508
rect 35072 19465 35081 19499
rect 35081 19465 35115 19499
rect 35115 19465 35124 19499
rect 35072 19456 35124 19465
rect 35164 19456 35216 19508
rect 35256 19456 35308 19508
rect 27160 19431 27212 19440
rect 18788 19320 18840 19372
rect 19524 19320 19576 19372
rect 22100 19320 22152 19372
rect 23664 19320 23716 19372
rect 25136 19320 25188 19372
rect 26148 19363 26200 19372
rect 26148 19329 26157 19363
rect 26157 19329 26191 19363
rect 26191 19329 26200 19363
rect 26148 19320 26200 19329
rect 27160 19397 27187 19431
rect 27187 19397 27212 19431
rect 27160 19388 27212 19397
rect 27804 19388 27856 19440
rect 30196 19388 30248 19440
rect 27436 19320 27488 19372
rect 28632 19320 28684 19372
rect 30748 19320 30800 19372
rect 31300 19320 31352 19372
rect 31668 19363 31720 19372
rect 31668 19329 31677 19363
rect 31677 19329 31711 19363
rect 31711 19329 31720 19363
rect 31668 19320 31720 19329
rect 33416 19320 33468 19372
rect 33876 19320 33928 19372
rect 34428 19363 34480 19372
rect 34428 19329 34437 19363
rect 34437 19329 34471 19363
rect 34471 19329 34480 19363
rect 34428 19320 34480 19329
rect 34612 19363 34664 19372
rect 34612 19329 34621 19363
rect 34621 19329 34655 19363
rect 34655 19329 34664 19363
rect 34612 19320 34664 19329
rect 35440 19363 35492 19372
rect 14556 19252 14608 19304
rect 17408 19252 17460 19304
rect 24584 19252 24636 19304
rect 15016 19184 15068 19236
rect 16672 19184 16724 19236
rect 18420 19184 18472 19236
rect 22284 19184 22336 19236
rect 26332 19252 26384 19304
rect 26424 19295 26476 19304
rect 26424 19261 26433 19295
rect 26433 19261 26467 19295
rect 26467 19261 26476 19295
rect 26424 19252 26476 19261
rect 26700 19252 26752 19304
rect 35440 19329 35449 19363
rect 35449 19329 35483 19363
rect 35483 19329 35492 19363
rect 35440 19320 35492 19329
rect 38292 19320 38344 19372
rect 35992 19252 36044 19304
rect 12348 19116 12400 19168
rect 12532 19116 12584 19168
rect 13912 19159 13964 19168
rect 13912 19125 13921 19159
rect 13921 19125 13955 19159
rect 13955 19125 13964 19159
rect 13912 19116 13964 19125
rect 14372 19116 14424 19168
rect 14740 19116 14792 19168
rect 18972 19116 19024 19168
rect 19248 19116 19300 19168
rect 20904 19116 20956 19168
rect 24584 19116 24636 19168
rect 25320 19116 25372 19168
rect 25688 19116 25740 19168
rect 26056 19116 26108 19168
rect 26240 19116 26292 19168
rect 37740 19159 37792 19168
rect 37740 19125 37749 19159
rect 37749 19125 37783 19159
rect 37783 19125 37792 19159
rect 37740 19116 37792 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 5908 18912 5960 18964
rect 8392 18912 8444 18964
rect 9680 18912 9732 18964
rect 9772 18912 9824 18964
rect 11152 18912 11204 18964
rect 11612 18912 11664 18964
rect 11980 18912 12032 18964
rect 3608 18776 3660 18828
rect 8208 18887 8260 18896
rect 8208 18853 8217 18887
rect 8217 18853 8251 18887
rect 8251 18853 8260 18887
rect 8208 18844 8260 18853
rect 5356 18776 5408 18828
rect 940 18708 992 18760
rect 2044 18572 2096 18624
rect 5448 18708 5500 18760
rect 6368 18708 6420 18760
rect 9496 18751 9548 18760
rect 9496 18717 9505 18751
rect 9505 18717 9539 18751
rect 9539 18717 9548 18751
rect 9496 18708 9548 18717
rect 9588 18708 9640 18760
rect 7748 18640 7800 18692
rect 10876 18844 10928 18896
rect 11060 18844 11112 18896
rect 13544 18844 13596 18896
rect 13728 18955 13780 18964
rect 13728 18921 13737 18955
rect 13737 18921 13771 18955
rect 13771 18921 13780 18955
rect 13728 18912 13780 18921
rect 13912 18912 13964 18964
rect 20720 18912 20772 18964
rect 22100 18912 22152 18964
rect 15384 18844 15436 18896
rect 16212 18844 16264 18896
rect 18420 18844 18472 18896
rect 5632 18615 5684 18624
rect 5632 18581 5641 18615
rect 5641 18581 5675 18615
rect 5675 18581 5684 18615
rect 5632 18572 5684 18581
rect 10048 18572 10100 18624
rect 10416 18708 10468 18760
rect 10324 18572 10376 18624
rect 10508 18615 10560 18624
rect 10508 18581 10517 18615
rect 10517 18581 10551 18615
rect 10551 18581 10560 18615
rect 10508 18572 10560 18581
rect 11888 18708 11940 18760
rect 12348 18776 12400 18828
rect 12900 18819 12952 18828
rect 12900 18785 12909 18819
rect 12909 18785 12943 18819
rect 12943 18785 12952 18819
rect 12900 18776 12952 18785
rect 12624 18708 12676 18760
rect 12808 18751 12860 18760
rect 12808 18717 12817 18751
rect 12817 18717 12851 18751
rect 12851 18717 12860 18751
rect 12808 18708 12860 18717
rect 13176 18751 13228 18760
rect 13176 18717 13185 18751
rect 13185 18717 13219 18751
rect 13219 18717 13228 18751
rect 13176 18708 13228 18717
rect 13636 18708 13688 18760
rect 13360 18615 13412 18624
rect 13360 18581 13369 18615
rect 13369 18581 13403 18615
rect 13403 18581 13412 18615
rect 13360 18572 13412 18581
rect 14372 18751 14424 18760
rect 14372 18717 14381 18751
rect 14381 18717 14415 18751
rect 14415 18717 14424 18751
rect 14372 18708 14424 18717
rect 14188 18640 14240 18692
rect 13912 18615 13964 18624
rect 13912 18581 13921 18615
rect 13921 18581 13955 18615
rect 13955 18581 13964 18615
rect 13912 18572 13964 18581
rect 14556 18572 14608 18624
rect 15292 18751 15344 18760
rect 15292 18717 15301 18751
rect 15301 18717 15335 18751
rect 15335 18717 15344 18751
rect 15292 18708 15344 18717
rect 16672 18776 16724 18828
rect 15844 18708 15896 18760
rect 18604 18751 18656 18760
rect 18604 18717 18613 18751
rect 18613 18717 18647 18751
rect 18647 18717 18656 18751
rect 18604 18708 18656 18717
rect 21088 18844 21140 18896
rect 24492 18912 24544 18964
rect 24676 18912 24728 18964
rect 29736 18912 29788 18964
rect 33416 18912 33468 18964
rect 34336 18912 34388 18964
rect 35348 18912 35400 18964
rect 37648 18912 37700 18964
rect 19340 18776 19392 18828
rect 20536 18776 20588 18828
rect 21548 18751 21600 18760
rect 21548 18717 21557 18751
rect 21557 18717 21591 18751
rect 21591 18717 21600 18751
rect 21548 18708 21600 18717
rect 22100 18751 22152 18760
rect 22100 18717 22109 18751
rect 22109 18717 22143 18751
rect 22143 18717 22152 18751
rect 22100 18708 22152 18717
rect 22284 18708 22336 18760
rect 22376 18751 22428 18760
rect 22376 18717 22385 18751
rect 22385 18717 22419 18751
rect 22419 18717 22428 18751
rect 22376 18708 22428 18717
rect 22468 18751 22520 18760
rect 22468 18717 22477 18751
rect 22477 18717 22511 18751
rect 22511 18717 22520 18751
rect 22468 18708 22520 18717
rect 22652 18776 22704 18828
rect 30656 18844 30708 18896
rect 23848 18708 23900 18760
rect 24676 18751 24728 18760
rect 24676 18717 24685 18751
rect 24685 18717 24719 18751
rect 24719 18717 24728 18751
rect 24676 18708 24728 18717
rect 25136 18776 25188 18828
rect 30104 18776 30156 18828
rect 33508 18844 33560 18896
rect 33784 18887 33836 18896
rect 33784 18853 33793 18887
rect 33793 18853 33827 18887
rect 33827 18853 33836 18887
rect 33784 18844 33836 18853
rect 34060 18844 34112 18896
rect 34612 18844 34664 18896
rect 17592 18640 17644 18692
rect 19984 18683 20036 18692
rect 19984 18649 19993 18683
rect 19993 18649 20027 18683
rect 20027 18649 20036 18683
rect 19984 18640 20036 18649
rect 16120 18572 16172 18624
rect 18328 18572 18380 18624
rect 19064 18615 19116 18624
rect 19064 18581 19073 18615
rect 19073 18581 19107 18615
rect 19107 18581 19116 18615
rect 19064 18572 19116 18581
rect 21272 18572 21324 18624
rect 23020 18572 23072 18624
rect 25044 18751 25096 18760
rect 25044 18717 25053 18751
rect 25053 18717 25087 18751
rect 25087 18717 25096 18751
rect 25044 18708 25096 18717
rect 25320 18708 25372 18760
rect 28816 18708 28868 18760
rect 29920 18708 29972 18760
rect 32404 18751 32456 18760
rect 32404 18717 32413 18751
rect 32413 18717 32447 18751
rect 32447 18717 32456 18751
rect 32404 18708 32456 18717
rect 33692 18776 33744 18828
rect 33416 18751 33468 18760
rect 33416 18717 33425 18751
rect 33425 18717 33459 18751
rect 33459 18717 33468 18751
rect 33416 18708 33468 18717
rect 33508 18751 33560 18760
rect 33508 18717 33517 18751
rect 33517 18717 33551 18751
rect 33551 18717 33560 18751
rect 34060 18751 34112 18760
rect 33508 18708 33560 18717
rect 34060 18717 34069 18751
rect 34069 18717 34103 18751
rect 34103 18717 34112 18751
rect 34060 18708 34112 18717
rect 33232 18640 33284 18692
rect 37372 18751 37424 18760
rect 37372 18717 37381 18751
rect 37381 18717 37415 18751
rect 37415 18717 37424 18751
rect 37372 18708 37424 18717
rect 27436 18572 27488 18624
rect 28724 18572 28776 18624
rect 28908 18615 28960 18624
rect 28908 18581 28917 18615
rect 28917 18581 28951 18615
rect 28951 18581 28960 18615
rect 28908 18572 28960 18581
rect 29276 18615 29328 18624
rect 29276 18581 29285 18615
rect 29285 18581 29319 18615
rect 29319 18581 29328 18615
rect 29276 18572 29328 18581
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 2044 18368 2096 18420
rect 3608 18368 3660 18420
rect 4712 18368 4764 18420
rect 5540 18368 5592 18420
rect 1400 18232 1452 18284
rect 3240 18232 3292 18284
rect 8852 18300 8904 18352
rect 5356 18164 5408 18216
rect 7748 18232 7800 18284
rect 8300 18232 8352 18284
rect 10324 18232 10376 18284
rect 10508 18368 10560 18420
rect 13176 18368 13228 18420
rect 13912 18368 13964 18420
rect 17776 18368 17828 18420
rect 19064 18368 19116 18420
rect 19984 18368 20036 18420
rect 22468 18368 22520 18420
rect 24676 18368 24728 18420
rect 11520 18300 11572 18352
rect 4804 18096 4856 18148
rect 3700 18071 3752 18080
rect 3700 18037 3709 18071
rect 3709 18037 3743 18071
rect 3743 18037 3752 18071
rect 3700 18028 3752 18037
rect 4896 18028 4948 18080
rect 11704 18164 11756 18216
rect 14280 18275 14332 18284
rect 14280 18241 14289 18275
rect 14289 18241 14323 18275
rect 14323 18241 14332 18275
rect 14280 18232 14332 18241
rect 14464 18275 14516 18284
rect 14464 18241 14473 18275
rect 14473 18241 14507 18275
rect 14507 18241 14516 18275
rect 14464 18232 14516 18241
rect 15568 18232 15620 18284
rect 15660 18164 15712 18216
rect 16304 18275 16356 18284
rect 16304 18241 16313 18275
rect 16313 18241 16347 18275
rect 16347 18241 16356 18275
rect 16304 18232 16356 18241
rect 16580 18232 16632 18284
rect 6460 18096 6512 18148
rect 14740 18096 14792 18148
rect 17040 18164 17092 18216
rect 7840 18028 7892 18080
rect 10232 18071 10284 18080
rect 10232 18037 10241 18071
rect 10241 18037 10275 18071
rect 10275 18037 10284 18071
rect 10232 18028 10284 18037
rect 11704 18028 11756 18080
rect 14648 18028 14700 18080
rect 15292 18028 15344 18080
rect 16488 18071 16540 18080
rect 16488 18037 16497 18071
rect 16497 18037 16531 18071
rect 16531 18037 16540 18071
rect 16488 18028 16540 18037
rect 16856 18028 16908 18080
rect 18420 18232 18472 18284
rect 19340 18343 19392 18352
rect 19340 18309 19349 18343
rect 19349 18309 19383 18343
rect 19383 18309 19392 18343
rect 19340 18300 19392 18309
rect 26056 18411 26108 18420
rect 26056 18377 26065 18411
rect 26065 18377 26099 18411
rect 26099 18377 26108 18411
rect 26056 18368 26108 18377
rect 28908 18368 28960 18420
rect 33232 18368 33284 18420
rect 33876 18368 33928 18420
rect 26608 18300 26660 18352
rect 17868 18207 17920 18216
rect 17868 18173 17877 18207
rect 17877 18173 17911 18207
rect 17911 18173 17920 18207
rect 17868 18164 17920 18173
rect 20444 18232 20496 18284
rect 21364 18232 21416 18284
rect 21824 18275 21876 18284
rect 21824 18241 21833 18275
rect 21833 18241 21867 18275
rect 21867 18241 21876 18275
rect 21824 18232 21876 18241
rect 20904 18164 20956 18216
rect 23848 18232 23900 18284
rect 25136 18232 25188 18284
rect 25228 18232 25280 18284
rect 26976 18275 27028 18284
rect 26976 18241 26985 18275
rect 26985 18241 27019 18275
rect 27019 18241 27028 18275
rect 26976 18232 27028 18241
rect 18512 18028 18564 18080
rect 18880 18071 18932 18080
rect 18880 18037 18889 18071
rect 18889 18037 18923 18071
rect 18923 18037 18932 18071
rect 18880 18028 18932 18037
rect 22928 18164 22980 18216
rect 23480 18164 23532 18216
rect 21088 18028 21140 18080
rect 21272 18028 21324 18080
rect 22192 18028 22244 18080
rect 23756 18028 23808 18080
rect 24676 18096 24728 18148
rect 29000 18207 29052 18216
rect 29000 18173 29009 18207
rect 29009 18173 29043 18207
rect 29043 18173 29052 18207
rect 29000 18164 29052 18173
rect 30380 18232 30432 18284
rect 31024 18207 31076 18216
rect 28632 18096 28684 18148
rect 26056 18028 26108 18080
rect 27160 18071 27212 18080
rect 27160 18037 27169 18071
rect 27169 18037 27203 18071
rect 27203 18037 27212 18071
rect 27160 18028 27212 18037
rect 27252 18028 27304 18080
rect 31024 18173 31033 18207
rect 31033 18173 31067 18207
rect 31067 18173 31076 18207
rect 31024 18164 31076 18173
rect 32220 18275 32272 18284
rect 32220 18241 32229 18275
rect 32229 18241 32263 18275
rect 32263 18241 32272 18275
rect 32220 18232 32272 18241
rect 32312 18275 32364 18284
rect 32312 18241 32321 18275
rect 32321 18241 32355 18275
rect 32355 18241 32364 18275
rect 32312 18232 32364 18241
rect 33508 18232 33560 18284
rect 33692 18207 33744 18216
rect 33692 18173 33701 18207
rect 33701 18173 33735 18207
rect 33735 18173 33744 18207
rect 33692 18164 33744 18173
rect 34336 18164 34388 18216
rect 37280 18164 37332 18216
rect 33140 18096 33192 18148
rect 33416 18139 33468 18148
rect 33416 18105 33425 18139
rect 33425 18105 33459 18139
rect 33459 18105 33468 18139
rect 33416 18096 33468 18105
rect 30472 18071 30524 18080
rect 30472 18037 30481 18071
rect 30481 18037 30515 18071
rect 30515 18037 30524 18071
rect 30472 18028 30524 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 4804 17824 4856 17876
rect 7748 17824 7800 17876
rect 7840 17824 7892 17876
rect 9496 17824 9548 17876
rect 10048 17824 10100 17876
rect 10692 17824 10744 17876
rect 13728 17824 13780 17876
rect 14096 17824 14148 17876
rect 17500 17824 17552 17876
rect 17776 17824 17828 17876
rect 18696 17824 18748 17876
rect 1400 17688 1452 17740
rect 1860 17688 1912 17740
rect 3976 17688 4028 17740
rect 4896 17620 4948 17672
rect 5632 17552 5684 17604
rect 4620 17527 4672 17536
rect 4620 17493 4629 17527
rect 4629 17493 4663 17527
rect 4663 17493 4672 17527
rect 4620 17484 4672 17493
rect 6184 17484 6236 17536
rect 7288 17620 7340 17672
rect 8116 17620 8168 17672
rect 9680 17620 9732 17672
rect 10048 17620 10100 17672
rect 8024 17595 8076 17604
rect 8024 17561 8033 17595
rect 8033 17561 8067 17595
rect 8067 17561 8076 17595
rect 8024 17552 8076 17561
rect 8392 17552 8444 17604
rect 10140 17552 10192 17604
rect 12164 17663 12216 17672
rect 12164 17629 12173 17663
rect 12173 17629 12207 17663
rect 12207 17629 12216 17663
rect 12164 17620 12216 17629
rect 12256 17663 12308 17672
rect 12256 17629 12265 17663
rect 12265 17629 12299 17663
rect 12299 17629 12308 17663
rect 12256 17620 12308 17629
rect 12532 17688 12584 17740
rect 13728 17620 13780 17672
rect 14740 17663 14792 17672
rect 10784 17552 10836 17604
rect 13452 17552 13504 17604
rect 7748 17484 7800 17536
rect 11612 17484 11664 17536
rect 11980 17484 12032 17536
rect 12256 17484 12308 17536
rect 12348 17484 12400 17536
rect 14740 17629 14749 17663
rect 14749 17629 14783 17663
rect 14783 17629 14792 17663
rect 14740 17620 14792 17629
rect 14832 17620 14884 17672
rect 15384 17663 15436 17672
rect 15384 17629 15393 17663
rect 15393 17629 15427 17663
rect 15427 17629 15436 17663
rect 15384 17620 15436 17629
rect 15660 17620 15712 17672
rect 17040 17688 17092 17740
rect 16212 17552 16264 17604
rect 16580 17620 16632 17672
rect 16856 17620 16908 17672
rect 17224 17663 17276 17672
rect 17224 17629 17233 17663
rect 17233 17629 17267 17663
rect 17267 17629 17276 17663
rect 17224 17620 17276 17629
rect 17776 17620 17828 17672
rect 18052 17663 18104 17672
rect 18052 17629 18061 17663
rect 18061 17629 18095 17663
rect 18095 17629 18104 17663
rect 18052 17620 18104 17629
rect 18236 17663 18288 17672
rect 18236 17629 18245 17663
rect 18245 17629 18279 17663
rect 18279 17629 18288 17663
rect 18236 17620 18288 17629
rect 18512 17620 18564 17672
rect 19156 17824 19208 17876
rect 20720 17824 20772 17876
rect 18972 17756 19024 17808
rect 24860 17824 24912 17876
rect 25228 17824 25280 17876
rect 16488 17552 16540 17604
rect 17040 17552 17092 17604
rect 18144 17552 18196 17604
rect 18972 17552 19024 17604
rect 19340 17620 19392 17672
rect 20352 17731 20404 17740
rect 20352 17697 20361 17731
rect 20361 17697 20395 17731
rect 20395 17697 20404 17731
rect 20352 17688 20404 17697
rect 20812 17663 20864 17672
rect 20812 17629 20821 17663
rect 20821 17629 20855 17663
rect 20855 17629 20864 17663
rect 20812 17620 20864 17629
rect 21088 17663 21140 17672
rect 21088 17629 21097 17663
rect 21097 17629 21131 17663
rect 21131 17629 21140 17663
rect 21088 17620 21140 17629
rect 21180 17620 21232 17672
rect 22284 17620 22336 17672
rect 20444 17484 20496 17536
rect 21180 17484 21232 17536
rect 23020 17620 23072 17672
rect 23848 17756 23900 17808
rect 23940 17688 23992 17740
rect 25136 17731 25188 17740
rect 25136 17697 25145 17731
rect 25145 17697 25179 17731
rect 25179 17697 25188 17731
rect 25136 17688 25188 17697
rect 25504 17756 25556 17808
rect 23480 17663 23532 17672
rect 23480 17629 23489 17663
rect 23489 17629 23523 17663
rect 23523 17629 23532 17663
rect 23480 17620 23532 17629
rect 22744 17552 22796 17604
rect 22928 17595 22980 17604
rect 22928 17561 22937 17595
rect 22937 17561 22971 17595
rect 22971 17561 22980 17595
rect 22928 17552 22980 17561
rect 25504 17620 25556 17672
rect 27160 17688 27212 17740
rect 24124 17552 24176 17604
rect 24952 17552 25004 17604
rect 25228 17552 25280 17604
rect 22468 17484 22520 17536
rect 22560 17484 22612 17536
rect 23848 17484 23900 17536
rect 24584 17484 24636 17536
rect 25964 17527 26016 17536
rect 25964 17493 25973 17527
rect 25973 17493 26007 17527
rect 26007 17493 26016 17527
rect 25964 17484 26016 17493
rect 26332 17484 26384 17536
rect 27528 17552 27580 17604
rect 29000 17824 29052 17876
rect 29276 17824 29328 17876
rect 37372 17824 37424 17876
rect 28816 17620 28868 17672
rect 30472 17688 30524 17740
rect 30840 17688 30892 17740
rect 30564 17663 30616 17672
rect 30564 17629 30573 17663
rect 30573 17629 30607 17663
rect 30607 17629 30616 17663
rect 30564 17620 30616 17629
rect 31208 17620 31260 17672
rect 31300 17552 31352 17604
rect 27436 17484 27488 17536
rect 28540 17527 28592 17536
rect 28540 17493 28549 17527
rect 28549 17493 28583 17527
rect 28583 17493 28592 17527
rect 28540 17484 28592 17493
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 3700 17280 3752 17332
rect 4620 17280 4672 17332
rect 8852 17280 8904 17332
rect 10692 17280 10744 17332
rect 6184 17212 6236 17264
rect 7840 17212 7892 17264
rect 3976 17144 4028 17196
rect 7932 17187 7984 17196
rect 7932 17153 7941 17187
rect 7941 17153 7975 17187
rect 7975 17153 7984 17187
rect 7932 17144 7984 17153
rect 2504 16940 2556 16992
rect 8208 16940 8260 16992
rect 9220 17187 9272 17196
rect 9220 17153 9229 17187
rect 9229 17153 9263 17187
rect 9263 17153 9272 17187
rect 9220 17144 9272 17153
rect 11060 17212 11112 17264
rect 11888 17323 11940 17332
rect 11888 17289 11897 17323
rect 11897 17289 11931 17323
rect 11931 17289 11940 17323
rect 11888 17280 11940 17289
rect 12164 17280 12216 17332
rect 12808 17280 12860 17332
rect 12256 17255 12308 17264
rect 12256 17221 12265 17255
rect 12265 17221 12299 17255
rect 12299 17221 12308 17255
rect 12256 17212 12308 17221
rect 12440 17255 12492 17264
rect 12440 17221 12449 17255
rect 12449 17221 12483 17255
rect 12483 17221 12492 17255
rect 12440 17212 12492 17221
rect 13084 17212 13136 17264
rect 9680 17187 9732 17196
rect 9680 17153 9689 17187
rect 9689 17153 9723 17187
rect 9723 17153 9732 17187
rect 9680 17144 9732 17153
rect 10232 17187 10284 17196
rect 10232 17153 10241 17187
rect 10241 17153 10275 17187
rect 10275 17153 10284 17187
rect 10232 17144 10284 17153
rect 10876 17144 10928 17196
rect 9772 17076 9824 17128
rect 10508 17076 10560 17128
rect 10692 17119 10744 17128
rect 10692 17085 10701 17119
rect 10701 17085 10735 17119
rect 10735 17085 10744 17119
rect 10692 17076 10744 17085
rect 11704 17144 11756 17196
rect 14648 17280 14700 17332
rect 14740 17280 14792 17332
rect 14004 17255 14056 17264
rect 14004 17221 14013 17255
rect 14013 17221 14047 17255
rect 14047 17221 14056 17255
rect 14004 17212 14056 17221
rect 14924 17212 14976 17264
rect 18696 17280 18748 17332
rect 11612 17076 11664 17128
rect 12624 17076 12676 17128
rect 14096 17187 14148 17196
rect 14096 17153 14110 17187
rect 14110 17153 14144 17187
rect 14144 17153 14148 17187
rect 14096 17144 14148 17153
rect 14464 17144 14516 17196
rect 14832 17144 14884 17196
rect 15660 17144 15712 17196
rect 16488 17212 16540 17264
rect 16856 17144 16908 17196
rect 17040 17187 17092 17196
rect 17040 17153 17049 17187
rect 17049 17153 17083 17187
rect 17083 17153 17092 17187
rect 17040 17144 17092 17153
rect 17224 17212 17276 17264
rect 20812 17323 20864 17332
rect 20812 17289 20821 17323
rect 20821 17289 20855 17323
rect 20855 17289 20864 17323
rect 20812 17280 20864 17289
rect 21180 17323 21232 17332
rect 21180 17289 21189 17323
rect 21189 17289 21223 17323
rect 21223 17289 21232 17323
rect 21180 17280 21232 17289
rect 22284 17212 22336 17264
rect 18972 17187 19024 17196
rect 18972 17153 18981 17187
rect 18981 17153 19015 17187
rect 19015 17153 19024 17187
rect 18972 17144 19024 17153
rect 20352 17144 20404 17196
rect 11704 17051 11756 17060
rect 11704 17017 11713 17051
rect 11713 17017 11747 17051
rect 11747 17017 11756 17051
rect 11704 17008 11756 17017
rect 11888 17008 11940 17060
rect 13544 17008 13596 17060
rect 19156 17076 19208 17128
rect 21548 17144 21600 17196
rect 22560 17144 22612 17196
rect 18880 17008 18932 17060
rect 22192 17076 22244 17128
rect 23020 17212 23072 17264
rect 24584 17280 24636 17332
rect 24676 17323 24728 17332
rect 24676 17289 24685 17323
rect 24685 17289 24719 17323
rect 24719 17289 24728 17323
rect 24676 17280 24728 17289
rect 25136 17280 25188 17332
rect 25872 17280 25924 17332
rect 25964 17280 26016 17332
rect 26976 17323 27028 17332
rect 26976 17289 26985 17323
rect 26985 17289 27019 17323
rect 27019 17289 27028 17323
rect 26976 17280 27028 17289
rect 9772 16940 9824 16992
rect 10784 16983 10836 16992
rect 10784 16949 10793 16983
rect 10793 16949 10827 16983
rect 10827 16949 10836 16983
rect 10784 16940 10836 16949
rect 10876 16940 10928 16992
rect 12440 16940 12492 16992
rect 14280 16983 14332 16992
rect 14280 16949 14289 16983
rect 14289 16949 14323 16983
rect 14323 16949 14332 16983
rect 14280 16940 14332 16949
rect 15384 16940 15436 16992
rect 15660 16940 15712 16992
rect 16948 16940 17000 16992
rect 17500 16940 17552 16992
rect 18604 16940 18656 16992
rect 20444 16983 20496 16992
rect 20444 16949 20453 16983
rect 20453 16949 20487 16983
rect 20487 16949 20496 16983
rect 20444 16940 20496 16949
rect 23204 17076 23256 17128
rect 23572 17076 23624 17128
rect 22836 17008 22888 17060
rect 23940 17076 23992 17128
rect 24400 17144 24452 17196
rect 25412 17187 25464 17196
rect 25412 17153 25421 17187
rect 25421 17153 25455 17187
rect 25455 17153 25464 17187
rect 25412 17144 25464 17153
rect 26332 17212 26384 17264
rect 28172 17280 28224 17332
rect 28540 17280 28592 17332
rect 24124 17008 24176 17060
rect 23204 16940 23256 16992
rect 23848 16940 23900 16992
rect 24768 16940 24820 16992
rect 30472 17212 30524 17264
rect 27988 17144 28040 17196
rect 37740 17212 37792 17264
rect 27528 17119 27580 17128
rect 27528 17085 27537 17119
rect 27537 17085 27571 17119
rect 27571 17085 27580 17119
rect 27528 17076 27580 17085
rect 33140 17144 33192 17196
rect 33232 17144 33284 17196
rect 26148 17008 26200 17060
rect 32220 17076 32272 17128
rect 33968 17119 34020 17128
rect 33968 17085 33977 17119
rect 33977 17085 34011 17119
rect 34011 17085 34020 17119
rect 33968 17076 34020 17085
rect 30932 16940 30984 16992
rect 33048 16940 33100 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 10600 16736 10652 16788
rect 1860 16643 1912 16652
rect 1860 16609 1869 16643
rect 1869 16609 1903 16643
rect 1903 16609 1912 16643
rect 1860 16600 1912 16609
rect 2504 16600 2556 16652
rect 4804 16600 4856 16652
rect 5540 16600 5592 16652
rect 3240 16532 3292 16584
rect 7104 16600 7156 16652
rect 7288 16643 7340 16652
rect 7288 16609 7297 16643
rect 7297 16609 7331 16643
rect 7331 16609 7340 16643
rect 7288 16600 7340 16609
rect 7748 16600 7800 16652
rect 8208 16643 8260 16652
rect 8208 16609 8217 16643
rect 8217 16609 8251 16643
rect 8251 16609 8260 16643
rect 8208 16600 8260 16609
rect 7840 16575 7892 16584
rect 7840 16541 7849 16575
rect 7849 16541 7883 16575
rect 7883 16541 7892 16575
rect 7840 16532 7892 16541
rect 8116 16532 8168 16584
rect 6184 16464 6236 16516
rect 9588 16668 9640 16720
rect 9220 16600 9272 16652
rect 10784 16600 10836 16652
rect 9128 16575 9180 16584
rect 9128 16541 9137 16575
rect 9137 16541 9171 16575
rect 9171 16541 9180 16575
rect 9128 16532 9180 16541
rect 9404 16532 9456 16584
rect 9496 16575 9548 16584
rect 9496 16541 9505 16575
rect 9505 16541 9539 16575
rect 9539 16541 9548 16575
rect 9496 16532 9548 16541
rect 9680 16575 9732 16584
rect 9680 16541 9687 16575
rect 9687 16541 9732 16575
rect 9680 16532 9732 16541
rect 9864 16575 9916 16584
rect 9864 16541 9873 16575
rect 9873 16541 9907 16575
rect 9907 16541 9916 16575
rect 9864 16532 9916 16541
rect 10416 16532 10468 16584
rect 10600 16575 10652 16584
rect 10600 16541 10604 16575
rect 10604 16541 10638 16575
rect 10638 16541 10652 16575
rect 10600 16532 10652 16541
rect 12348 16779 12400 16788
rect 12348 16745 12357 16779
rect 12357 16745 12391 16779
rect 12391 16745 12400 16779
rect 12348 16736 12400 16745
rect 15568 16736 15620 16788
rect 17500 16736 17552 16788
rect 18512 16736 18564 16788
rect 18880 16736 18932 16788
rect 23480 16736 23532 16788
rect 24768 16736 24820 16788
rect 24952 16736 25004 16788
rect 11612 16668 11664 16720
rect 6368 16439 6420 16448
rect 6368 16405 6377 16439
rect 6377 16405 6411 16439
rect 6411 16405 6420 16439
rect 6368 16396 6420 16405
rect 6736 16439 6788 16448
rect 6736 16405 6745 16439
rect 6745 16405 6779 16439
rect 6779 16405 6788 16439
rect 6736 16396 6788 16405
rect 7656 16396 7708 16448
rect 11060 16575 11112 16584
rect 11060 16541 11069 16575
rect 11069 16541 11103 16575
rect 11103 16541 11112 16575
rect 11060 16532 11112 16541
rect 11704 16532 11756 16584
rect 12256 16575 12308 16584
rect 12256 16541 12265 16575
rect 12265 16541 12299 16575
rect 12299 16541 12308 16575
rect 12256 16532 12308 16541
rect 12348 16532 12400 16584
rect 17960 16668 18012 16720
rect 18696 16668 18748 16720
rect 15384 16600 15436 16652
rect 13452 16532 13504 16584
rect 13544 16575 13596 16584
rect 13544 16541 13553 16575
rect 13553 16541 13587 16575
rect 13587 16541 13596 16575
rect 13544 16532 13596 16541
rect 14372 16575 14424 16584
rect 14372 16541 14381 16575
rect 14381 16541 14415 16575
rect 14415 16541 14424 16575
rect 14372 16532 14424 16541
rect 14464 16532 14516 16584
rect 15844 16532 15896 16584
rect 17408 16575 17460 16584
rect 17408 16541 17417 16575
rect 17417 16541 17451 16575
rect 17451 16541 17460 16575
rect 17408 16532 17460 16541
rect 19984 16600 20036 16652
rect 20812 16668 20864 16720
rect 9404 16396 9456 16448
rect 10140 16439 10192 16448
rect 10140 16405 10149 16439
rect 10149 16405 10183 16439
rect 10183 16405 10192 16439
rect 10140 16396 10192 16405
rect 10232 16396 10284 16448
rect 14648 16464 14700 16516
rect 11980 16396 12032 16448
rect 13912 16439 13964 16448
rect 13912 16405 13921 16439
rect 13921 16405 13955 16439
rect 13955 16405 13964 16439
rect 13912 16396 13964 16405
rect 16948 16507 17000 16516
rect 16948 16473 16957 16507
rect 16957 16473 16991 16507
rect 16991 16473 17000 16507
rect 16948 16464 17000 16473
rect 17224 16464 17276 16516
rect 18144 16464 18196 16516
rect 14924 16439 14976 16448
rect 14924 16405 14933 16439
rect 14933 16405 14967 16439
rect 14967 16405 14976 16439
rect 14924 16396 14976 16405
rect 17500 16396 17552 16448
rect 17684 16396 17736 16448
rect 19432 16532 19484 16584
rect 22100 16575 22152 16584
rect 22100 16541 22108 16575
rect 22108 16541 22142 16575
rect 22142 16541 22152 16575
rect 22100 16532 22152 16541
rect 22652 16600 22704 16652
rect 24124 16600 24176 16652
rect 22284 16575 22336 16584
rect 22284 16541 22293 16575
rect 22293 16541 22327 16575
rect 22327 16541 22336 16575
rect 22284 16532 22336 16541
rect 19616 16464 19668 16516
rect 20904 16464 20956 16516
rect 22560 16532 22612 16584
rect 22836 16575 22888 16584
rect 22836 16541 22844 16575
rect 22844 16541 22878 16575
rect 22878 16541 22888 16575
rect 22836 16532 22888 16541
rect 23020 16575 23072 16584
rect 23020 16541 23029 16575
rect 23029 16541 23063 16575
rect 23063 16541 23072 16575
rect 23020 16532 23072 16541
rect 23204 16575 23256 16584
rect 23204 16541 23213 16575
rect 23213 16541 23247 16575
rect 23247 16541 23256 16575
rect 23204 16532 23256 16541
rect 27068 16736 27120 16788
rect 29552 16736 29604 16788
rect 30748 16736 30800 16788
rect 30932 16779 30984 16788
rect 30932 16745 30962 16779
rect 30962 16745 30984 16779
rect 30932 16736 30984 16745
rect 32220 16736 32272 16788
rect 27620 16600 27672 16652
rect 26332 16575 26384 16584
rect 26332 16541 26341 16575
rect 26341 16541 26375 16575
rect 26375 16541 26384 16575
rect 26332 16532 26384 16541
rect 27160 16532 27212 16584
rect 33048 16600 33100 16652
rect 22652 16396 22704 16448
rect 22744 16396 22796 16448
rect 24124 16464 24176 16516
rect 25688 16464 25740 16516
rect 26424 16464 26476 16516
rect 25504 16396 25556 16448
rect 25872 16396 25924 16448
rect 26332 16396 26384 16448
rect 26792 16507 26844 16516
rect 26792 16473 26801 16507
rect 26801 16473 26835 16507
rect 26835 16473 26844 16507
rect 26792 16464 26844 16473
rect 29184 16464 29236 16516
rect 30104 16464 30156 16516
rect 32680 16575 32732 16584
rect 32680 16541 32689 16575
rect 32689 16541 32723 16575
rect 32723 16541 32732 16575
rect 32680 16532 32732 16541
rect 33968 16464 34020 16516
rect 27896 16396 27948 16448
rect 30196 16396 30248 16448
rect 31116 16396 31168 16448
rect 34428 16439 34480 16448
rect 34428 16405 34437 16439
rect 34437 16405 34471 16439
rect 34471 16405 34480 16439
rect 34428 16396 34480 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 940 16124 992 16176
rect 3976 16192 4028 16244
rect 6368 16192 6420 16244
rect 7288 16192 7340 16244
rect 7932 16192 7984 16244
rect 9220 16192 9272 16244
rect 9956 16192 10008 16244
rect 11612 16192 11664 16244
rect 11980 16192 12032 16244
rect 12348 16192 12400 16244
rect 9772 16167 9824 16176
rect 9772 16133 9781 16167
rect 9781 16133 9815 16167
rect 9815 16133 9824 16167
rect 9772 16124 9824 16133
rect 7656 16099 7708 16108
rect 7656 16065 7665 16099
rect 7665 16065 7699 16099
rect 7699 16065 7708 16099
rect 7656 16056 7708 16065
rect 7748 16056 7800 16108
rect 8116 16056 8168 16108
rect 8392 16099 8444 16108
rect 8392 16065 8401 16099
rect 8401 16065 8435 16099
rect 8435 16065 8444 16099
rect 8392 16056 8444 16065
rect 9404 16056 9456 16108
rect 9864 16099 9916 16108
rect 10692 16124 10744 16176
rect 9864 16065 9909 16099
rect 9909 16065 9916 16099
rect 9864 16056 9916 16065
rect 9680 15988 9732 16040
rect 10416 16099 10468 16108
rect 10416 16065 10425 16099
rect 10425 16065 10459 16099
rect 10459 16065 10468 16099
rect 10416 16056 10468 16065
rect 10600 16099 10652 16108
rect 10600 16065 10609 16099
rect 10609 16065 10643 16099
rect 10643 16065 10652 16099
rect 10600 16056 10652 16065
rect 11060 16056 11112 16108
rect 14004 16192 14056 16244
rect 14280 16192 14332 16244
rect 14464 16192 14516 16244
rect 15384 16192 15436 16244
rect 17592 16192 17644 16244
rect 19616 16192 19668 16244
rect 19708 16235 19760 16244
rect 19708 16201 19717 16235
rect 19717 16201 19751 16235
rect 19751 16201 19760 16235
rect 19708 16192 19760 16201
rect 12624 16124 12676 16176
rect 15660 16124 15712 16176
rect 12992 16056 13044 16108
rect 13268 16056 13320 16108
rect 13360 16099 13412 16108
rect 13360 16065 13369 16099
rect 13369 16065 13403 16099
rect 13403 16065 13412 16099
rect 13360 16056 13412 16065
rect 13912 16056 13964 16108
rect 14280 16056 14332 16108
rect 14096 15988 14148 16040
rect 14188 16031 14240 16040
rect 14188 15997 14197 16031
rect 14197 15997 14231 16031
rect 14231 15997 14240 16031
rect 14188 15988 14240 15997
rect 9864 15920 9916 15972
rect 12440 15963 12492 15972
rect 12440 15929 12449 15963
rect 12449 15929 12483 15963
rect 12483 15929 12492 15963
rect 12440 15920 12492 15929
rect 15936 16056 15988 16108
rect 14832 15988 14884 16040
rect 19340 16124 19392 16176
rect 16212 16056 16264 16108
rect 17224 16099 17276 16108
rect 17224 16065 17233 16099
rect 17233 16065 17267 16099
rect 17267 16065 17276 16099
rect 17224 16056 17276 16065
rect 17500 16099 17552 16108
rect 17500 16065 17509 16099
rect 17509 16065 17543 16099
rect 17543 16065 17552 16099
rect 17500 16056 17552 16065
rect 17316 15988 17368 16040
rect 18604 16056 18656 16108
rect 18328 15988 18380 16040
rect 15568 15920 15620 15972
rect 15844 15963 15896 15972
rect 15844 15929 15853 15963
rect 15853 15929 15887 15963
rect 15887 15929 15896 15963
rect 15844 15920 15896 15929
rect 19524 16056 19576 16108
rect 19616 16099 19668 16108
rect 19616 16065 19655 16099
rect 19655 16065 19668 16099
rect 19616 16056 19668 16065
rect 19340 15988 19392 16040
rect 19892 15988 19944 16040
rect 20536 16099 20588 16108
rect 20536 16065 20545 16099
rect 20545 16065 20579 16099
rect 20579 16065 20588 16099
rect 20536 16056 20588 16065
rect 20628 16099 20680 16108
rect 20628 16065 20637 16099
rect 20637 16065 20671 16099
rect 20671 16065 20680 16099
rect 20628 16056 20680 16065
rect 20904 16099 20956 16108
rect 20904 16065 20913 16099
rect 20913 16065 20947 16099
rect 20947 16065 20956 16099
rect 20904 16056 20956 16065
rect 21364 16056 21416 16108
rect 4068 15895 4120 15904
rect 4068 15861 4077 15895
rect 4077 15861 4111 15895
rect 4111 15861 4120 15895
rect 4068 15852 4120 15861
rect 5080 15852 5132 15904
rect 7748 15852 7800 15904
rect 9772 15852 9824 15904
rect 9956 15852 10008 15904
rect 10876 15852 10928 15904
rect 12900 15852 12952 15904
rect 13636 15852 13688 15904
rect 14556 15852 14608 15904
rect 15660 15852 15712 15904
rect 20076 15963 20128 15972
rect 20076 15929 20085 15963
rect 20085 15929 20119 15963
rect 20119 15929 20128 15963
rect 20076 15920 20128 15929
rect 22376 16192 22428 16244
rect 24124 16192 24176 16244
rect 21640 16124 21692 16176
rect 22100 16099 22152 16108
rect 22100 16065 22109 16099
rect 22109 16065 22143 16099
rect 22143 16065 22152 16099
rect 22100 16056 22152 16065
rect 22192 16099 22244 16108
rect 22192 16065 22201 16099
rect 22201 16065 22235 16099
rect 22235 16065 22244 16099
rect 22192 16056 22244 16065
rect 23756 16056 23808 16108
rect 24400 16192 24452 16244
rect 25044 16192 25096 16244
rect 26792 16192 26844 16244
rect 27436 16192 27488 16244
rect 29828 16192 29880 16244
rect 24676 16124 24728 16176
rect 24124 15920 24176 15972
rect 24308 15920 24360 15972
rect 24492 16099 24544 16108
rect 24492 16065 24506 16099
rect 24506 16065 24540 16099
rect 24540 16065 24544 16099
rect 24492 16056 24544 16065
rect 25044 16099 25096 16108
rect 25044 16065 25053 16099
rect 25053 16065 25087 16099
rect 25087 16065 25096 16099
rect 25044 16056 25096 16065
rect 25136 16056 25188 16108
rect 25780 16099 25832 16108
rect 25780 16065 25789 16099
rect 25789 16065 25823 16099
rect 25823 16065 25832 16099
rect 25780 16056 25832 16065
rect 25964 16099 26016 16108
rect 25964 16065 25971 16099
rect 25971 16065 26016 16099
rect 25964 16056 26016 16065
rect 26332 16124 26384 16176
rect 28540 16124 28592 16176
rect 24952 15988 25004 16040
rect 19616 15852 19668 15904
rect 19800 15852 19852 15904
rect 20904 15852 20956 15904
rect 21456 15852 21508 15904
rect 25872 15920 25924 15972
rect 26332 15920 26384 15972
rect 28632 16099 28684 16108
rect 28632 16065 28641 16099
rect 28641 16065 28675 16099
rect 28675 16065 28684 16099
rect 28632 16056 28684 16065
rect 29092 16099 29144 16108
rect 29092 16065 29101 16099
rect 29101 16065 29135 16099
rect 29135 16065 29144 16099
rect 29092 16056 29144 16065
rect 30104 16167 30156 16176
rect 30104 16133 30113 16167
rect 30113 16133 30147 16167
rect 30147 16133 30156 16167
rect 30104 16124 30156 16133
rect 30196 16167 30248 16176
rect 30196 16133 30205 16167
rect 30205 16133 30239 16167
rect 30239 16133 30248 16167
rect 30196 16124 30248 16133
rect 32680 16192 32732 16244
rect 33232 16235 33284 16244
rect 33232 16201 33241 16235
rect 33241 16201 33275 16235
rect 33275 16201 33284 16235
rect 33232 16192 33284 16201
rect 33324 16192 33376 16244
rect 33784 16192 33836 16244
rect 34428 16192 34480 16244
rect 29828 16099 29880 16108
rect 26608 15988 26660 16040
rect 27988 16031 28040 16040
rect 27988 15997 27997 16031
rect 27997 15997 28031 16031
rect 28031 15997 28040 16031
rect 27988 15988 28040 15997
rect 28080 15988 28132 16040
rect 29828 16065 29837 16099
rect 29837 16065 29871 16099
rect 29871 16065 29880 16099
rect 29828 16056 29880 16065
rect 30380 16056 30432 16108
rect 28356 15920 28408 15972
rect 25044 15852 25096 15904
rect 25320 15852 25372 15904
rect 27252 15852 27304 15904
rect 28264 15895 28316 15904
rect 28264 15861 28273 15895
rect 28273 15861 28307 15895
rect 28307 15861 28316 15895
rect 28264 15852 28316 15861
rect 28632 15852 28684 15904
rect 29276 15852 29328 15904
rect 29552 15963 29604 15972
rect 29552 15929 29561 15963
rect 29561 15929 29595 15963
rect 29595 15929 29604 15963
rect 29552 15920 29604 15929
rect 30564 16031 30616 16040
rect 30564 15997 30573 16031
rect 30573 15997 30607 16031
rect 30607 15997 30616 16031
rect 30564 15988 30616 15997
rect 30656 15988 30708 16040
rect 32036 16056 32088 16108
rect 33140 16056 33192 16108
rect 33876 16031 33928 16040
rect 33876 15997 33885 16031
rect 33885 15997 33919 16031
rect 33919 15997 33928 16031
rect 33876 15988 33928 15997
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 6736 15648 6788 15700
rect 9772 15691 9824 15700
rect 9772 15657 9781 15691
rect 9781 15657 9815 15691
rect 9815 15657 9824 15691
rect 9772 15648 9824 15657
rect 9864 15648 9916 15700
rect 12072 15648 12124 15700
rect 12440 15648 12492 15700
rect 12900 15691 12952 15700
rect 12900 15657 12909 15691
rect 12909 15657 12943 15691
rect 12943 15657 12952 15691
rect 12900 15648 12952 15657
rect 5080 15512 5132 15564
rect 3976 15444 4028 15496
rect 6184 15512 6236 15564
rect 8944 15512 8996 15564
rect 9312 15512 9364 15564
rect 9864 15555 9916 15564
rect 9864 15521 9873 15555
rect 9873 15521 9907 15555
rect 9907 15521 9916 15555
rect 9864 15512 9916 15521
rect 6828 15444 6880 15496
rect 9128 15444 9180 15496
rect 9956 15444 10008 15496
rect 11244 15512 11296 15564
rect 13360 15580 13412 15632
rect 13636 15580 13688 15632
rect 14096 15580 14148 15632
rect 14556 15580 14608 15632
rect 14924 15580 14976 15632
rect 10140 15444 10192 15496
rect 10232 15444 10284 15496
rect 12992 15512 13044 15564
rect 14188 15555 14240 15564
rect 14188 15521 14197 15555
rect 14197 15521 14231 15555
rect 14231 15521 14240 15555
rect 14188 15512 14240 15521
rect 7196 15308 7248 15360
rect 7748 15351 7800 15360
rect 7748 15317 7757 15351
rect 7757 15317 7791 15351
rect 7791 15317 7800 15351
rect 7748 15308 7800 15317
rect 10232 15351 10284 15360
rect 10232 15317 10241 15351
rect 10241 15317 10275 15351
rect 10275 15317 10284 15351
rect 10232 15308 10284 15317
rect 11612 15444 11664 15496
rect 11888 15487 11940 15496
rect 11888 15453 11897 15487
rect 11897 15453 11931 15487
rect 11931 15453 11940 15487
rect 11888 15444 11940 15453
rect 11980 15487 12032 15496
rect 11980 15453 11989 15487
rect 11989 15453 12023 15487
rect 12023 15453 12032 15487
rect 11980 15444 12032 15453
rect 12072 15487 12124 15496
rect 12072 15453 12081 15487
rect 12081 15453 12115 15487
rect 12115 15453 12124 15487
rect 12072 15444 12124 15453
rect 12624 15444 12676 15496
rect 14280 15487 14332 15496
rect 14280 15453 14289 15487
rect 14289 15453 14323 15487
rect 14323 15453 14332 15487
rect 14280 15444 14332 15453
rect 15384 15487 15436 15496
rect 15384 15453 15393 15487
rect 15393 15453 15427 15487
rect 15427 15453 15436 15487
rect 15384 15444 15436 15453
rect 15844 15444 15896 15496
rect 16028 15487 16080 15496
rect 16028 15453 16037 15487
rect 16037 15453 16071 15487
rect 16071 15453 16080 15487
rect 16028 15444 16080 15453
rect 18420 15580 18472 15632
rect 17224 15555 17276 15564
rect 17224 15521 17233 15555
rect 17233 15521 17267 15555
rect 17267 15521 17276 15555
rect 17224 15512 17276 15521
rect 19340 15648 19392 15700
rect 19064 15580 19116 15632
rect 19432 15580 19484 15632
rect 21456 15648 21508 15700
rect 21824 15648 21876 15700
rect 22192 15648 22244 15700
rect 22376 15648 22428 15700
rect 25320 15648 25372 15700
rect 26056 15648 26108 15700
rect 26424 15648 26476 15700
rect 26884 15691 26936 15700
rect 26884 15657 26893 15691
rect 26893 15657 26927 15691
rect 26927 15657 26936 15691
rect 26884 15648 26936 15657
rect 17408 15444 17460 15496
rect 17500 15487 17552 15496
rect 17500 15453 17509 15487
rect 17509 15453 17543 15487
rect 17543 15453 17552 15487
rect 17500 15444 17552 15453
rect 17960 15444 18012 15496
rect 15108 15419 15160 15428
rect 15108 15385 15117 15419
rect 15117 15385 15151 15419
rect 15151 15385 15160 15419
rect 15108 15376 15160 15385
rect 15568 15376 15620 15428
rect 16948 15419 17000 15428
rect 16948 15385 16957 15419
rect 16957 15385 16991 15419
rect 16991 15385 17000 15419
rect 16948 15376 17000 15385
rect 17132 15376 17184 15428
rect 11520 15308 11572 15360
rect 11704 15308 11756 15360
rect 18420 15444 18472 15496
rect 18604 15444 18656 15496
rect 20076 15580 20128 15632
rect 19616 15487 19668 15496
rect 19616 15453 19625 15487
rect 19625 15453 19659 15487
rect 19659 15453 19668 15487
rect 19616 15444 19668 15453
rect 19892 15487 19944 15496
rect 19892 15453 19901 15487
rect 19901 15453 19935 15487
rect 19935 15453 19944 15487
rect 19892 15444 19944 15453
rect 20260 15487 20312 15496
rect 20260 15453 20269 15487
rect 20269 15453 20303 15487
rect 20303 15453 20312 15487
rect 20260 15444 20312 15453
rect 21364 15580 21416 15632
rect 20536 15512 20588 15564
rect 22560 15555 22612 15564
rect 22560 15521 22569 15555
rect 22569 15521 22603 15555
rect 22603 15521 22612 15555
rect 22560 15512 22612 15521
rect 23388 15512 23440 15564
rect 25136 15512 25188 15564
rect 25320 15512 25372 15564
rect 25964 15580 26016 15632
rect 28356 15648 28408 15700
rect 28540 15648 28592 15700
rect 28264 15580 28316 15632
rect 20076 15419 20128 15428
rect 20076 15385 20085 15419
rect 20085 15385 20119 15419
rect 20119 15385 20128 15419
rect 20076 15376 20128 15385
rect 20536 15376 20588 15428
rect 20720 15419 20772 15428
rect 20720 15385 20729 15419
rect 20729 15385 20763 15419
rect 20763 15385 20772 15419
rect 20720 15376 20772 15385
rect 21272 15487 21324 15496
rect 21272 15453 21281 15487
rect 21281 15453 21315 15487
rect 21315 15453 21324 15487
rect 21272 15444 21324 15453
rect 22284 15444 22336 15496
rect 25596 15487 25648 15496
rect 25596 15453 25606 15487
rect 25606 15453 25640 15487
rect 25640 15453 25648 15487
rect 25596 15444 25648 15453
rect 26056 15444 26108 15496
rect 26792 15512 26844 15564
rect 29092 15691 29144 15700
rect 29092 15657 29101 15691
rect 29101 15657 29135 15691
rect 29135 15657 29144 15691
rect 29092 15648 29144 15657
rect 29276 15648 29328 15700
rect 30564 15648 30616 15700
rect 30380 15580 30432 15632
rect 26332 15444 26384 15496
rect 26424 15487 26476 15496
rect 26424 15453 26433 15487
rect 26433 15453 26467 15487
rect 26467 15453 26476 15487
rect 26424 15444 26476 15453
rect 19616 15308 19668 15360
rect 19800 15308 19852 15360
rect 20904 15308 20956 15360
rect 22836 15376 22888 15428
rect 23296 15376 23348 15428
rect 24032 15376 24084 15428
rect 25044 15419 25096 15428
rect 25044 15385 25053 15419
rect 25053 15385 25087 15419
rect 25087 15385 25096 15419
rect 25044 15376 25096 15385
rect 25780 15419 25832 15428
rect 25780 15385 25789 15419
rect 25789 15385 25823 15419
rect 25823 15385 25832 15419
rect 26608 15487 26660 15496
rect 26608 15453 26617 15487
rect 26617 15453 26651 15487
rect 26651 15453 26660 15487
rect 26608 15444 26660 15453
rect 26700 15444 26752 15496
rect 27068 15444 27120 15496
rect 25780 15376 25832 15385
rect 23848 15308 23900 15360
rect 24768 15308 24820 15360
rect 25136 15351 25188 15360
rect 25136 15317 25145 15351
rect 25145 15317 25179 15351
rect 25179 15317 25188 15351
rect 25136 15308 25188 15317
rect 25504 15308 25556 15360
rect 25964 15308 26016 15360
rect 27252 15308 27304 15360
rect 27528 15308 27580 15360
rect 27896 15487 27948 15496
rect 27896 15453 27906 15487
rect 27906 15453 27940 15487
rect 27940 15453 27948 15487
rect 27896 15444 27948 15453
rect 28172 15487 28224 15496
rect 28172 15453 28181 15487
rect 28181 15453 28215 15487
rect 28215 15453 28224 15487
rect 28172 15444 28224 15453
rect 28264 15487 28316 15496
rect 28264 15453 28278 15487
rect 28278 15453 28312 15487
rect 28312 15453 28316 15487
rect 28264 15444 28316 15453
rect 28724 15487 28776 15496
rect 28724 15453 28733 15487
rect 28733 15453 28767 15487
rect 28767 15453 28776 15487
rect 28724 15444 28776 15453
rect 28816 15444 28868 15496
rect 28908 15487 28960 15496
rect 28908 15453 28917 15487
rect 28917 15453 28951 15487
rect 28951 15453 28960 15487
rect 28908 15444 28960 15453
rect 33508 15512 33560 15564
rect 28080 15419 28132 15428
rect 28080 15385 28089 15419
rect 28089 15385 28123 15419
rect 28123 15385 28132 15419
rect 28080 15376 28132 15385
rect 28448 15376 28500 15428
rect 29092 15376 29144 15428
rect 30196 15444 30248 15496
rect 30564 15487 30616 15496
rect 30564 15453 30573 15487
rect 30573 15453 30607 15487
rect 30607 15453 30616 15487
rect 30564 15444 30616 15453
rect 30840 15487 30892 15496
rect 30840 15453 30849 15487
rect 30849 15453 30883 15487
rect 30883 15453 30892 15487
rect 30840 15444 30892 15453
rect 32404 15444 32456 15496
rect 33968 15376 34020 15428
rect 32588 15351 32640 15360
rect 32588 15317 32597 15351
rect 32597 15317 32631 15351
rect 32631 15317 32640 15351
rect 32588 15308 32640 15317
rect 33324 15308 33376 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 1768 15147 1820 15156
rect 1768 15113 1777 15147
rect 1777 15113 1811 15147
rect 1811 15113 1820 15147
rect 1768 15104 1820 15113
rect 9128 15147 9180 15156
rect 9128 15113 9137 15147
rect 9137 15113 9171 15147
rect 9171 15113 9180 15147
rect 9128 15104 9180 15113
rect 7748 15036 7800 15088
rect 9036 15036 9088 15088
rect 1952 15011 2004 15020
rect 1952 14977 1961 15011
rect 1961 14977 1995 15011
rect 1995 14977 2004 15011
rect 1952 14968 2004 14977
rect 11152 15104 11204 15156
rect 11888 15104 11940 15156
rect 16856 15104 16908 15156
rect 17684 15104 17736 15156
rect 17960 15104 18012 15156
rect 7196 14943 7248 14952
rect 7196 14909 7205 14943
rect 7205 14909 7239 14943
rect 7239 14909 7248 14943
rect 7196 14900 7248 14909
rect 8024 14900 8076 14952
rect 11704 15036 11756 15088
rect 10232 15011 10284 15020
rect 10232 14977 10241 15011
rect 10241 14977 10275 15011
rect 10275 14977 10284 15011
rect 10232 14968 10284 14977
rect 12256 15011 12308 15020
rect 12256 14977 12265 15011
rect 12265 14977 12299 15011
rect 12299 14977 12308 15011
rect 12256 14968 12308 14977
rect 12440 15011 12492 15020
rect 12440 14977 12449 15011
rect 12449 14977 12483 15011
rect 12483 14977 12492 15011
rect 12440 14968 12492 14977
rect 12808 14968 12860 15020
rect 11060 14832 11112 14884
rect 14556 14968 14608 15020
rect 14924 15011 14976 15020
rect 14924 14977 14933 15011
rect 14933 14977 14967 15011
rect 14967 14977 14976 15011
rect 14924 14968 14976 14977
rect 12900 14900 12952 14952
rect 15660 14968 15712 15020
rect 17132 15011 17184 15020
rect 17132 14977 17141 15011
rect 17141 14977 17175 15011
rect 17175 14977 17184 15011
rect 17132 14968 17184 14977
rect 15568 14900 15620 14952
rect 16396 14900 16448 14952
rect 17224 14832 17276 14884
rect 9588 14764 9640 14816
rect 12164 14764 12216 14816
rect 17776 14968 17828 15020
rect 17960 15011 18012 15020
rect 17960 14977 17969 15011
rect 17969 14977 18003 15011
rect 18003 14977 18012 15011
rect 17960 14968 18012 14977
rect 18236 14968 18288 15020
rect 18328 14968 18380 15020
rect 18420 15011 18472 15020
rect 18420 14977 18429 15011
rect 18429 14977 18463 15011
rect 18463 14977 18472 15011
rect 18420 14968 18472 14977
rect 19708 15104 19760 15156
rect 20352 15104 20404 15156
rect 20628 15104 20680 15156
rect 18696 15079 18748 15088
rect 18696 15045 18705 15079
rect 18705 15045 18739 15079
rect 18739 15045 18748 15079
rect 18696 15036 18748 15045
rect 19524 15036 19576 15088
rect 20812 15079 20864 15088
rect 20812 15045 20821 15079
rect 20821 15045 20855 15079
rect 20855 15045 20864 15079
rect 20812 15036 20864 15045
rect 20996 15104 21048 15156
rect 24400 15104 24452 15156
rect 24768 15104 24820 15156
rect 25228 15104 25280 15156
rect 19432 14968 19484 15020
rect 19616 15011 19668 15020
rect 19616 14977 19625 15011
rect 19625 14977 19659 15011
rect 19659 14977 19668 15011
rect 19616 14968 19668 14977
rect 19800 15011 19852 15020
rect 19800 14977 19817 15011
rect 19817 14977 19852 15011
rect 19800 14968 19852 14977
rect 20168 14968 20220 15020
rect 20536 15011 20588 15020
rect 20536 14977 20545 15011
rect 20545 14977 20579 15011
rect 20579 14977 20588 15011
rect 20536 14968 20588 14977
rect 20628 15011 20680 15020
rect 20628 14977 20637 15011
rect 20637 14977 20671 15011
rect 20671 14977 20680 15011
rect 20628 14968 20680 14977
rect 21732 14968 21784 15020
rect 21916 14968 21968 15020
rect 22284 14968 22336 15020
rect 23388 15011 23440 15020
rect 23388 14977 23397 15011
rect 23397 14977 23431 15011
rect 23431 14977 23440 15011
rect 23388 14968 23440 14977
rect 19708 14832 19760 14884
rect 21180 14900 21232 14952
rect 21272 14900 21324 14952
rect 20720 14832 20772 14884
rect 23572 14900 23624 14952
rect 24400 15011 24452 15020
rect 24400 14977 24409 15011
rect 24409 14977 24443 15011
rect 24443 14977 24452 15011
rect 24400 14968 24452 14977
rect 24584 15011 24636 15020
rect 24584 14977 24593 15011
rect 24593 14977 24627 15011
rect 24627 14977 24636 15011
rect 24584 14968 24636 14977
rect 25688 15104 25740 15156
rect 26148 15104 26200 15156
rect 26424 15104 26476 15156
rect 28540 15104 28592 15156
rect 28724 15104 28776 15156
rect 30564 15104 30616 15156
rect 30840 15104 30892 15156
rect 33968 15104 34020 15156
rect 25504 14968 25556 15020
rect 18512 14764 18564 14816
rect 19432 14764 19484 14816
rect 24952 14832 25004 14884
rect 25596 14832 25648 14884
rect 28356 15011 28408 15020
rect 28356 14977 28365 15011
rect 28365 14977 28399 15011
rect 28399 14977 28408 15011
rect 28356 14968 28408 14977
rect 26424 14900 26476 14952
rect 28172 14900 28224 14952
rect 28540 14968 28592 15020
rect 28816 14968 28868 15020
rect 30104 14943 30156 14952
rect 30104 14909 30113 14943
rect 30113 14909 30147 14943
rect 30147 14909 30156 14943
rect 30104 14900 30156 14909
rect 30472 14968 30524 15020
rect 31116 15011 31168 15020
rect 31116 14977 31125 15011
rect 31125 14977 31159 15011
rect 31159 14977 31168 15011
rect 31116 14968 31168 14977
rect 31668 14968 31720 15020
rect 32404 14968 32456 15020
rect 33048 15011 33100 15020
rect 33048 14977 33057 15011
rect 33057 14977 33091 15011
rect 33091 14977 33100 15011
rect 33048 14968 33100 14977
rect 32588 14900 32640 14952
rect 33324 14943 33376 14952
rect 33324 14909 33333 14943
rect 33333 14909 33367 14943
rect 33367 14909 33376 14943
rect 33324 14900 33376 14909
rect 28908 14832 28960 14884
rect 22192 14807 22244 14816
rect 22192 14773 22201 14807
rect 22201 14773 22235 14807
rect 22235 14773 22244 14807
rect 22192 14764 22244 14773
rect 22468 14764 22520 14816
rect 23204 14807 23256 14816
rect 23204 14773 23213 14807
rect 23213 14773 23247 14807
rect 23247 14773 23256 14807
rect 23204 14764 23256 14773
rect 29828 14764 29880 14816
rect 31116 14764 31168 14816
rect 33600 14764 33652 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 1952 14560 2004 14612
rect 5356 14424 5408 14476
rect 12256 14560 12308 14612
rect 12440 14560 12492 14612
rect 13912 14560 13964 14612
rect 17040 14560 17092 14612
rect 7196 14467 7248 14476
rect 7196 14433 7205 14467
rect 7205 14433 7239 14467
rect 7239 14433 7248 14467
rect 7196 14424 7248 14433
rect 8024 14467 8076 14476
rect 8024 14433 8033 14467
rect 8033 14433 8067 14467
rect 8067 14433 8076 14467
rect 8024 14424 8076 14433
rect 8208 14467 8260 14476
rect 8208 14433 8217 14467
rect 8217 14433 8251 14467
rect 8251 14433 8260 14467
rect 8208 14424 8260 14433
rect 9864 14492 9916 14544
rect 11704 14492 11756 14544
rect 17960 14560 18012 14612
rect 18420 14560 18472 14612
rect 19892 14560 19944 14612
rect 20996 14560 21048 14612
rect 21732 14603 21784 14612
rect 21732 14569 21741 14603
rect 21741 14569 21775 14603
rect 21775 14569 21784 14603
rect 21732 14560 21784 14569
rect 24308 14560 24360 14612
rect 25964 14560 26016 14612
rect 26516 14560 26568 14612
rect 28816 14560 28868 14612
rect 32496 14560 32548 14612
rect 33048 14560 33100 14612
rect 11060 14424 11112 14476
rect 4528 14399 4580 14408
rect 4528 14365 4537 14399
rect 4537 14365 4571 14399
rect 4571 14365 4580 14399
rect 4528 14356 4580 14365
rect 4620 14399 4672 14408
rect 4620 14365 4629 14399
rect 4629 14365 4663 14399
rect 4663 14365 4672 14399
rect 4620 14356 4672 14365
rect 7104 14356 7156 14408
rect 10048 14356 10100 14408
rect 10140 14356 10192 14408
rect 11612 14356 11664 14408
rect 12164 14424 12216 14476
rect 17224 14492 17276 14544
rect 20536 14492 20588 14544
rect 14648 14424 14700 14476
rect 19892 14424 19944 14476
rect 20168 14467 20220 14476
rect 20168 14433 20177 14467
rect 20177 14433 20211 14467
rect 20211 14433 20220 14467
rect 20168 14424 20220 14433
rect 6184 14288 6236 14340
rect 5264 14220 5316 14272
rect 6552 14263 6604 14272
rect 6552 14229 6561 14263
rect 6561 14229 6595 14263
rect 6595 14229 6604 14263
rect 6552 14220 6604 14229
rect 7564 14263 7616 14272
rect 7564 14229 7573 14263
rect 7573 14229 7607 14263
rect 7607 14229 7616 14263
rect 7564 14220 7616 14229
rect 8484 14288 8536 14340
rect 12624 14356 12676 14408
rect 15016 14399 15068 14408
rect 15016 14365 15025 14399
rect 15025 14365 15059 14399
rect 15059 14365 15068 14399
rect 15016 14356 15068 14365
rect 17316 14356 17368 14408
rect 17868 14399 17920 14408
rect 17868 14365 17877 14399
rect 17877 14365 17911 14399
rect 17911 14365 17920 14399
rect 17868 14356 17920 14365
rect 17960 14399 18012 14408
rect 17960 14365 17969 14399
rect 17969 14365 18003 14399
rect 18003 14365 18012 14399
rect 17960 14356 18012 14365
rect 18144 14356 18196 14408
rect 19248 14356 19300 14408
rect 19340 14356 19392 14408
rect 19984 14356 20036 14408
rect 20720 14356 20772 14408
rect 12532 14288 12584 14340
rect 16488 14288 16540 14340
rect 18604 14288 18656 14340
rect 9036 14220 9088 14272
rect 14280 14220 14332 14272
rect 14924 14263 14976 14272
rect 14924 14229 14933 14263
rect 14933 14229 14967 14263
rect 14967 14229 14976 14263
rect 14924 14220 14976 14229
rect 17684 14220 17736 14272
rect 17868 14220 17920 14272
rect 20444 14331 20496 14340
rect 20444 14297 20453 14331
rect 20453 14297 20487 14331
rect 20487 14297 20496 14331
rect 20444 14288 20496 14297
rect 20536 14288 20588 14340
rect 21916 14399 21968 14408
rect 21916 14365 21925 14399
rect 21925 14365 21959 14399
rect 21959 14365 21968 14399
rect 21916 14356 21968 14365
rect 22192 14356 22244 14408
rect 21180 14331 21232 14340
rect 21180 14297 21189 14331
rect 21189 14297 21223 14331
rect 21223 14297 21232 14331
rect 21180 14288 21232 14297
rect 21272 14331 21324 14340
rect 21272 14297 21281 14331
rect 21281 14297 21315 14331
rect 21315 14297 21324 14331
rect 21272 14288 21324 14297
rect 20904 14220 20956 14272
rect 21364 14220 21416 14272
rect 22100 14288 22152 14340
rect 23940 14492 23992 14544
rect 26424 14492 26476 14544
rect 29276 14492 29328 14544
rect 30196 14492 30248 14544
rect 23204 14424 23256 14476
rect 24676 14424 24728 14476
rect 25688 14424 25740 14476
rect 27528 14424 27580 14476
rect 29644 14424 29696 14476
rect 22468 14399 22520 14408
rect 22468 14365 22477 14399
rect 22477 14365 22511 14399
rect 22511 14365 22520 14399
rect 22468 14356 22520 14365
rect 27712 14399 27764 14408
rect 27712 14365 27721 14399
rect 27721 14365 27755 14399
rect 27755 14365 27764 14399
rect 27712 14356 27764 14365
rect 28264 14399 28316 14408
rect 28264 14365 28273 14399
rect 28273 14365 28307 14399
rect 28307 14365 28316 14399
rect 28264 14356 28316 14365
rect 29368 14356 29420 14408
rect 30288 14356 30340 14408
rect 23204 14288 23256 14340
rect 24768 14288 24820 14340
rect 27988 14288 28040 14340
rect 38292 14492 38344 14544
rect 33140 14424 33192 14476
rect 33324 14424 33376 14476
rect 33968 14424 34020 14476
rect 37648 14399 37700 14408
rect 37648 14365 37657 14399
rect 37657 14365 37691 14399
rect 37691 14365 37700 14399
rect 37648 14356 37700 14365
rect 31392 14331 31444 14340
rect 31392 14297 31401 14331
rect 31401 14297 31435 14331
rect 31435 14297 31444 14331
rect 31392 14288 31444 14297
rect 33508 14288 33560 14340
rect 24860 14220 24912 14272
rect 29092 14220 29144 14272
rect 30656 14220 30708 14272
rect 33784 14220 33836 14272
rect 35440 14263 35492 14272
rect 35440 14229 35449 14263
rect 35449 14229 35483 14263
rect 35483 14229 35492 14263
rect 35440 14220 35492 14229
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 4620 14016 4672 14068
rect 5264 14016 5316 14068
rect 6552 14016 6604 14068
rect 7564 14016 7616 14068
rect 6460 13948 6512 14000
rect 1492 13855 1544 13864
rect 1492 13821 1501 13855
rect 1501 13821 1535 13855
rect 1535 13821 1544 13855
rect 1492 13812 1544 13821
rect 9588 13948 9640 14000
rect 9772 13880 9824 13932
rect 9956 13880 10008 13932
rect 10140 13923 10192 13932
rect 10140 13889 10149 13923
rect 10149 13889 10183 13923
rect 10183 13889 10192 13923
rect 10140 13880 10192 13889
rect 10324 13923 10376 13932
rect 10324 13889 10333 13923
rect 10333 13889 10367 13923
rect 10367 13889 10376 13923
rect 10324 13880 10376 13889
rect 10508 13880 10560 13932
rect 4804 13744 4856 13796
rect 4528 13676 4580 13728
rect 5264 13676 5316 13728
rect 9128 13744 9180 13796
rect 10232 13812 10284 13864
rect 10600 13787 10652 13796
rect 10600 13753 10609 13787
rect 10609 13753 10643 13787
rect 10643 13753 10652 13787
rect 10600 13744 10652 13753
rect 11796 14016 11848 14068
rect 11612 13880 11664 13932
rect 11980 13880 12032 13932
rect 12348 13923 12400 13932
rect 12348 13889 12357 13923
rect 12357 13889 12391 13923
rect 12391 13889 12400 13923
rect 12348 13880 12400 13889
rect 14740 14016 14792 14068
rect 14924 14016 14976 14068
rect 15292 14016 15344 14068
rect 16396 14016 16448 14068
rect 14556 13880 14608 13932
rect 14648 13880 14700 13932
rect 17500 13991 17552 14000
rect 17500 13957 17509 13991
rect 17509 13957 17543 13991
rect 17543 13957 17552 13991
rect 17500 13948 17552 13957
rect 16120 13880 16172 13932
rect 7104 13676 7156 13728
rect 9680 13676 9732 13728
rect 9956 13676 10008 13728
rect 10048 13719 10100 13728
rect 10048 13685 10057 13719
rect 10057 13685 10091 13719
rect 10091 13685 10100 13719
rect 10048 13676 10100 13685
rect 13360 13676 13412 13728
rect 17776 13744 17828 13796
rect 18144 13923 18196 13932
rect 18144 13889 18153 13923
rect 18153 13889 18187 13923
rect 18187 13889 18196 13923
rect 18144 13880 18196 13889
rect 18236 13880 18288 13932
rect 18696 14016 18748 14068
rect 18604 13948 18656 14000
rect 21732 14016 21784 14068
rect 21916 14016 21968 14068
rect 22468 14016 22520 14068
rect 23388 14059 23440 14068
rect 23388 14025 23397 14059
rect 23397 14025 23431 14059
rect 23431 14025 23440 14059
rect 23388 14016 23440 14025
rect 23480 14016 23532 14068
rect 24308 14016 24360 14068
rect 25504 14016 25556 14068
rect 29184 14016 29236 14068
rect 31392 14059 31444 14068
rect 31392 14025 31401 14059
rect 31401 14025 31435 14059
rect 31435 14025 31444 14059
rect 31392 14016 31444 14025
rect 20168 13948 20220 14000
rect 20444 13948 20496 14000
rect 18512 13880 18564 13932
rect 19064 13923 19116 13932
rect 19064 13889 19073 13923
rect 19073 13889 19107 13923
rect 19107 13889 19116 13923
rect 19064 13880 19116 13889
rect 20904 13880 20956 13932
rect 20536 13812 20588 13864
rect 18604 13744 18656 13796
rect 18880 13744 18932 13796
rect 24124 13948 24176 14000
rect 26332 13948 26384 14000
rect 26700 13948 26752 14000
rect 21088 13923 21140 13932
rect 21088 13889 21097 13923
rect 21097 13889 21131 13923
rect 21131 13889 21140 13923
rect 21088 13880 21140 13889
rect 21364 13880 21416 13932
rect 21916 13880 21968 13932
rect 22284 13880 22336 13932
rect 22468 13880 22520 13932
rect 22652 13880 22704 13932
rect 27988 13948 28040 14000
rect 23480 13744 23532 13796
rect 24308 13744 24360 13796
rect 28816 13880 28868 13932
rect 28264 13812 28316 13864
rect 24952 13744 25004 13796
rect 14832 13676 14884 13728
rect 15200 13676 15252 13728
rect 16488 13719 16540 13728
rect 16488 13685 16497 13719
rect 16497 13685 16531 13719
rect 16531 13685 16540 13719
rect 16488 13676 16540 13685
rect 17040 13676 17092 13728
rect 24676 13676 24728 13728
rect 26792 13676 26844 13728
rect 27252 13676 27304 13728
rect 28356 13744 28408 13796
rect 29184 13880 29236 13932
rect 29276 13880 29328 13932
rect 29828 13923 29880 13932
rect 29828 13889 29837 13923
rect 29837 13889 29871 13923
rect 29871 13889 29880 13923
rect 29828 13880 29880 13889
rect 32496 14059 32548 14068
rect 32496 14025 32505 14059
rect 32505 14025 32539 14059
rect 32539 14025 32548 14059
rect 32496 14016 32548 14025
rect 33784 14016 33836 14068
rect 35440 14016 35492 14068
rect 33968 13880 34020 13932
rect 27804 13676 27856 13728
rect 29552 13719 29604 13728
rect 29552 13685 29561 13719
rect 29561 13685 29595 13719
rect 29595 13685 29604 13719
rect 29552 13676 29604 13685
rect 30380 13744 30432 13796
rect 31300 13744 31352 13796
rect 33600 13855 33652 13864
rect 33600 13821 33609 13855
rect 33609 13821 33643 13855
rect 33643 13821 33652 13855
rect 33600 13812 33652 13821
rect 32680 13676 32732 13728
rect 34060 13676 34112 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 8484 13515 8536 13524
rect 8484 13481 8493 13515
rect 8493 13481 8527 13515
rect 8527 13481 8536 13515
rect 8484 13472 8536 13481
rect 10048 13404 10100 13456
rect 10508 13447 10560 13456
rect 10508 13413 10517 13447
rect 10517 13413 10551 13447
rect 10551 13413 10560 13447
rect 10508 13404 10560 13413
rect 10600 13404 10652 13456
rect 5540 13336 5592 13388
rect 7104 13336 7156 13388
rect 9496 13336 9548 13388
rect 3976 13311 4028 13320
rect 3976 13277 3985 13311
rect 3985 13277 4019 13311
rect 4019 13277 4028 13311
rect 3976 13268 4028 13277
rect 5264 13311 5316 13320
rect 5264 13277 5273 13311
rect 5273 13277 5307 13311
rect 5307 13277 5316 13311
rect 5264 13268 5316 13277
rect 6460 13311 6512 13320
rect 6460 13277 6469 13311
rect 6469 13277 6503 13311
rect 6503 13277 6512 13311
rect 6460 13268 6512 13277
rect 9036 13268 9088 13320
rect 6920 13200 6972 13252
rect 10324 13268 10376 13320
rect 12348 13472 12400 13524
rect 13084 13472 13136 13524
rect 13268 13472 13320 13524
rect 15200 13515 15252 13524
rect 15200 13481 15209 13515
rect 15209 13481 15243 13515
rect 15243 13481 15252 13515
rect 15200 13472 15252 13481
rect 14556 13404 14608 13456
rect 14740 13404 14792 13456
rect 11888 13311 11940 13320
rect 11888 13277 11897 13311
rect 11897 13277 11931 13311
rect 11931 13277 11940 13311
rect 11888 13268 11940 13277
rect 3884 13175 3936 13184
rect 3884 13141 3893 13175
rect 3893 13141 3927 13175
rect 3927 13141 3936 13175
rect 3884 13132 3936 13141
rect 4712 13132 4764 13184
rect 9588 13132 9640 13184
rect 9772 13132 9824 13184
rect 12808 13336 12860 13388
rect 13268 13311 13320 13320
rect 13268 13277 13277 13311
rect 13277 13277 13311 13311
rect 13311 13277 13320 13311
rect 13268 13268 13320 13277
rect 13452 13268 13504 13320
rect 15752 13336 15804 13388
rect 13544 13243 13596 13252
rect 13544 13209 13553 13243
rect 13553 13209 13587 13243
rect 13587 13209 13596 13243
rect 13544 13200 13596 13209
rect 18144 13472 18196 13524
rect 18328 13472 18380 13524
rect 20720 13472 20772 13524
rect 22928 13472 22980 13524
rect 16028 13404 16080 13456
rect 16948 13404 17000 13456
rect 16120 13379 16172 13388
rect 16120 13345 16129 13379
rect 16129 13345 16163 13379
rect 16163 13345 16172 13379
rect 16120 13336 16172 13345
rect 16764 13336 16816 13388
rect 17592 13336 17644 13388
rect 16488 13268 16540 13320
rect 17132 13268 17184 13320
rect 17316 13311 17368 13320
rect 17316 13277 17326 13311
rect 17326 13277 17360 13311
rect 17360 13277 17368 13311
rect 17316 13268 17368 13277
rect 16948 13200 17000 13252
rect 17868 13200 17920 13252
rect 18236 13404 18288 13456
rect 25412 13404 25464 13456
rect 25596 13404 25648 13456
rect 25688 13404 25740 13456
rect 25964 13404 26016 13456
rect 20168 13379 20220 13388
rect 20168 13345 20177 13379
rect 20177 13345 20211 13379
rect 20211 13345 20220 13379
rect 20168 13336 20220 13345
rect 18420 13311 18472 13320
rect 18420 13277 18429 13311
rect 18429 13277 18463 13311
rect 18463 13277 18472 13311
rect 18420 13268 18472 13277
rect 24492 13336 24544 13388
rect 18972 13200 19024 13252
rect 12900 13132 12952 13184
rect 12992 13132 13044 13184
rect 17316 13132 17368 13184
rect 18236 13132 18288 13184
rect 18328 13175 18380 13184
rect 18328 13141 18337 13175
rect 18337 13141 18371 13175
rect 18371 13141 18380 13175
rect 22652 13268 22704 13320
rect 21364 13200 21416 13252
rect 24860 13243 24912 13252
rect 18328 13132 18380 13141
rect 19432 13132 19484 13184
rect 19708 13132 19760 13184
rect 20812 13132 20864 13184
rect 24860 13209 24869 13243
rect 24869 13209 24903 13243
rect 24903 13209 24912 13243
rect 24860 13200 24912 13209
rect 25228 13268 25280 13320
rect 25688 13311 25740 13320
rect 25688 13277 25698 13311
rect 25698 13277 25732 13311
rect 25732 13277 25740 13311
rect 25688 13268 25740 13277
rect 25504 13200 25556 13252
rect 25872 13243 25924 13252
rect 25872 13209 25881 13243
rect 25881 13209 25915 13243
rect 25915 13209 25924 13243
rect 25872 13200 25924 13209
rect 25780 13132 25832 13184
rect 26148 13200 26200 13252
rect 26608 13243 26660 13252
rect 26608 13209 26617 13243
rect 26617 13209 26651 13243
rect 26651 13209 26660 13243
rect 26608 13200 26660 13209
rect 26424 13132 26476 13184
rect 27344 13472 27396 13524
rect 28816 13472 28868 13524
rect 27344 13336 27396 13388
rect 27804 13311 27856 13320
rect 27804 13277 27813 13311
rect 27813 13277 27847 13311
rect 27847 13277 27856 13311
rect 27804 13268 27856 13277
rect 27896 13311 27948 13320
rect 27896 13277 27905 13311
rect 27905 13277 27939 13311
rect 27939 13277 27948 13311
rect 27896 13268 27948 13277
rect 29552 13404 29604 13456
rect 28448 13268 28500 13320
rect 28724 13243 28776 13252
rect 28724 13209 28733 13243
rect 28733 13209 28767 13243
rect 28767 13209 28776 13243
rect 28724 13200 28776 13209
rect 28908 13311 28960 13320
rect 28908 13277 28917 13311
rect 28917 13277 28951 13311
rect 28951 13277 28960 13311
rect 28908 13268 28960 13277
rect 29368 13268 29420 13320
rect 29000 13200 29052 13252
rect 29644 13200 29696 13252
rect 30288 13447 30340 13456
rect 30288 13413 30297 13447
rect 30297 13413 30331 13447
rect 30331 13413 30340 13447
rect 30288 13404 30340 13413
rect 30104 13268 30156 13320
rect 30288 13311 30340 13320
rect 30288 13277 30297 13311
rect 30297 13277 30331 13311
rect 30331 13277 30340 13311
rect 30288 13268 30340 13277
rect 34060 13472 34112 13524
rect 30656 13404 30708 13456
rect 30472 13336 30524 13388
rect 30564 13268 30616 13320
rect 30748 13200 30800 13252
rect 31484 13311 31536 13320
rect 31484 13277 31493 13311
rect 31493 13277 31527 13311
rect 31527 13277 31536 13311
rect 31484 13268 31536 13277
rect 27160 13132 27212 13184
rect 31116 13132 31168 13184
rect 31944 13268 31996 13320
rect 33600 13336 33652 13388
rect 33876 13379 33928 13388
rect 33876 13345 33885 13379
rect 33885 13345 33919 13379
rect 33919 13345 33928 13379
rect 33876 13336 33928 13345
rect 33232 13200 33284 13252
rect 32036 13132 32088 13184
rect 32312 13175 32364 13184
rect 32312 13141 32321 13175
rect 32321 13141 32355 13175
rect 32355 13141 32364 13175
rect 32312 13132 32364 13141
rect 33692 13175 33744 13184
rect 33692 13141 33701 13175
rect 33701 13141 33735 13175
rect 33735 13141 33744 13175
rect 33692 13132 33744 13141
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 3884 12928 3936 12980
rect 5264 12860 5316 12912
rect 6184 12860 6236 12912
rect 9680 12928 9732 12980
rect 9772 12971 9824 12980
rect 9772 12937 9781 12971
rect 9781 12937 9815 12971
rect 9815 12937 9824 12971
rect 9772 12928 9824 12937
rect 9588 12860 9640 12912
rect 12532 12928 12584 12980
rect 13084 12928 13136 12980
rect 4436 12724 4488 12776
rect 9128 12724 9180 12776
rect 9496 12835 9548 12844
rect 9496 12801 9505 12835
rect 9505 12801 9539 12835
rect 9539 12801 9548 12835
rect 9496 12792 9548 12801
rect 9864 12835 9916 12844
rect 9864 12801 9873 12835
rect 9873 12801 9907 12835
rect 9907 12801 9916 12835
rect 9864 12792 9916 12801
rect 10048 12792 10100 12844
rect 10232 12792 10284 12844
rect 13544 12928 13596 12980
rect 14648 12928 14700 12980
rect 10600 12792 10652 12844
rect 11980 12792 12032 12844
rect 9036 12656 9088 12708
rect 10968 12767 11020 12776
rect 10968 12733 10977 12767
rect 10977 12733 11011 12767
rect 11011 12733 11020 12767
rect 10968 12724 11020 12733
rect 12624 12792 12676 12844
rect 12808 12792 12860 12844
rect 13360 12860 13412 12912
rect 16212 12860 16264 12912
rect 14280 12792 14332 12844
rect 18328 12928 18380 12980
rect 19432 12928 19484 12980
rect 21364 12971 21416 12980
rect 21364 12937 21373 12971
rect 21373 12937 21407 12971
rect 21407 12937 21416 12971
rect 21364 12928 21416 12937
rect 24308 12928 24360 12980
rect 23204 12860 23256 12912
rect 22284 12835 22336 12844
rect 22284 12801 22293 12835
rect 22293 12801 22327 12835
rect 22327 12801 22336 12835
rect 22284 12792 22336 12801
rect 9772 12656 9824 12708
rect 18236 12724 18288 12776
rect 18788 12724 18840 12776
rect 19616 12767 19668 12776
rect 19616 12733 19625 12767
rect 19625 12733 19659 12767
rect 19659 12733 19668 12767
rect 19616 12724 19668 12733
rect 24308 12724 24360 12776
rect 9128 12588 9180 12640
rect 14372 12588 14424 12640
rect 15108 12588 15160 12640
rect 19524 12656 19576 12708
rect 24676 12835 24728 12844
rect 24676 12801 24686 12835
rect 24686 12801 24720 12835
rect 24720 12801 24728 12835
rect 24676 12792 24728 12801
rect 25044 12835 25096 12844
rect 25044 12801 25058 12835
rect 25058 12801 25092 12835
rect 25092 12801 25096 12835
rect 25044 12792 25096 12801
rect 25320 12928 25372 12980
rect 25412 12928 25464 12980
rect 26516 12903 26568 12912
rect 26516 12869 26525 12903
rect 26525 12869 26559 12903
rect 26559 12869 26568 12903
rect 26516 12860 26568 12869
rect 26976 12928 27028 12980
rect 27896 12971 27948 12980
rect 27896 12937 27905 12971
rect 27905 12937 27939 12971
rect 27939 12937 27948 12971
rect 27896 12928 27948 12937
rect 28724 12928 28776 12980
rect 28908 12928 28960 12980
rect 25044 12656 25096 12708
rect 16856 12588 16908 12640
rect 22192 12588 22244 12640
rect 23388 12588 23440 12640
rect 25780 12767 25832 12776
rect 25780 12733 25789 12767
rect 25789 12733 25823 12767
rect 25823 12733 25832 12767
rect 25780 12724 25832 12733
rect 26056 12792 26108 12844
rect 26792 12835 26844 12844
rect 26792 12801 26801 12835
rect 26801 12801 26835 12835
rect 26835 12801 26844 12835
rect 26792 12792 26844 12801
rect 26976 12792 27028 12844
rect 27252 12835 27304 12844
rect 27252 12801 27261 12835
rect 27261 12801 27295 12835
rect 27295 12801 27304 12835
rect 27252 12792 27304 12801
rect 26240 12656 26292 12708
rect 26608 12656 26660 12708
rect 26792 12656 26844 12708
rect 26884 12656 26936 12708
rect 27344 12656 27396 12708
rect 27804 12792 27856 12844
rect 28540 12860 28592 12912
rect 29000 12860 29052 12912
rect 29368 12835 29420 12844
rect 29368 12801 29377 12835
rect 29377 12801 29411 12835
rect 29411 12801 29420 12835
rect 29368 12792 29420 12801
rect 30288 12928 30340 12980
rect 31944 12971 31996 12980
rect 31944 12937 31953 12971
rect 31953 12937 31987 12971
rect 31987 12937 31996 12971
rect 31944 12928 31996 12937
rect 32036 12928 32088 12980
rect 32312 12928 32364 12980
rect 31484 12860 31536 12912
rect 30104 12792 30156 12844
rect 25596 12588 25648 12640
rect 25688 12588 25740 12640
rect 29000 12656 29052 12708
rect 31300 12767 31352 12776
rect 31300 12733 31309 12767
rect 31309 12733 31343 12767
rect 31343 12733 31352 12767
rect 31300 12724 31352 12733
rect 27896 12588 27948 12640
rect 28540 12588 28592 12640
rect 30288 12588 30340 12640
rect 31392 12588 31444 12640
rect 33968 12792 34020 12844
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 4620 12384 4672 12436
rect 9128 12384 9180 12436
rect 4804 12248 4856 12300
rect 4712 12180 4764 12232
rect 9128 12248 9180 12300
rect 10048 12316 10100 12368
rect 10692 12316 10744 12368
rect 10968 12316 11020 12368
rect 6460 12180 6512 12232
rect 9956 12180 10008 12232
rect 10784 12223 10836 12232
rect 10784 12189 10793 12223
rect 10793 12189 10827 12223
rect 10827 12189 10836 12223
rect 10784 12180 10836 12189
rect 5448 12155 5500 12164
rect 5448 12121 5457 12155
rect 5457 12121 5491 12155
rect 5491 12121 5500 12155
rect 5448 12112 5500 12121
rect 6184 12112 6236 12164
rect 6828 12112 6880 12164
rect 9680 12112 9732 12164
rect 10968 12180 11020 12232
rect 15384 12384 15436 12436
rect 15660 12384 15712 12436
rect 15844 12384 15896 12436
rect 15936 12384 15988 12436
rect 16304 12384 16356 12436
rect 16396 12384 16448 12436
rect 16856 12427 16908 12436
rect 16856 12393 16865 12427
rect 16865 12393 16899 12427
rect 16899 12393 16908 12427
rect 16856 12384 16908 12393
rect 11980 12180 12032 12232
rect 12992 12112 13044 12164
rect 15108 12112 15160 12164
rect 15660 12180 15712 12232
rect 16120 12248 16172 12300
rect 21180 12384 21232 12436
rect 17592 12316 17644 12368
rect 18052 12359 18104 12368
rect 18052 12325 18061 12359
rect 18061 12325 18095 12359
rect 18095 12325 18104 12359
rect 18052 12316 18104 12325
rect 19524 12316 19576 12368
rect 16488 12180 16540 12232
rect 16948 12223 17000 12232
rect 16948 12189 16957 12223
rect 16957 12189 16991 12223
rect 16991 12189 17000 12223
rect 16948 12180 17000 12189
rect 17316 12248 17368 12300
rect 17224 12180 17276 12232
rect 18604 12248 18656 12300
rect 19708 12248 19760 12300
rect 20812 12248 20864 12300
rect 22928 12316 22980 12368
rect 23940 12316 23992 12368
rect 24676 12316 24728 12368
rect 24308 12248 24360 12300
rect 25044 12359 25096 12368
rect 25044 12325 25053 12359
rect 25053 12325 25087 12359
rect 25087 12325 25096 12359
rect 25044 12316 25096 12325
rect 25688 12316 25740 12368
rect 15844 12112 15896 12164
rect 18696 12223 18748 12232
rect 18696 12189 18705 12223
rect 18705 12189 18739 12223
rect 18739 12189 18748 12223
rect 18696 12180 18748 12189
rect 18788 12180 18840 12232
rect 21272 12180 21324 12232
rect 22376 12223 22428 12232
rect 22376 12189 22385 12223
rect 22385 12189 22419 12223
rect 22419 12189 22428 12223
rect 22376 12180 22428 12189
rect 22560 12223 22612 12232
rect 22560 12189 22569 12223
rect 22569 12189 22603 12223
rect 22603 12189 22612 12223
rect 22560 12180 22612 12189
rect 12440 12087 12492 12096
rect 12440 12053 12449 12087
rect 12449 12053 12483 12087
rect 12483 12053 12492 12087
rect 12440 12044 12492 12053
rect 13360 12044 13412 12096
rect 15016 12044 15068 12096
rect 15568 12044 15620 12096
rect 16488 12044 16540 12096
rect 20720 12112 20772 12164
rect 20904 12112 20956 12164
rect 21180 12112 21232 12164
rect 22192 12112 22244 12164
rect 24124 12180 24176 12232
rect 24492 12180 24544 12232
rect 23940 12112 23992 12164
rect 24584 12155 24636 12164
rect 24584 12121 24593 12155
rect 24593 12121 24627 12155
rect 24627 12121 24636 12155
rect 24584 12112 24636 12121
rect 24860 12180 24912 12232
rect 25412 12155 25464 12164
rect 25412 12121 25421 12155
rect 25421 12121 25455 12155
rect 25455 12121 25464 12155
rect 25412 12112 25464 12121
rect 25872 12384 25924 12436
rect 26700 12384 26752 12436
rect 27252 12384 27304 12436
rect 29644 12384 29696 12436
rect 31300 12384 31352 12436
rect 26608 12316 26660 12368
rect 27988 12316 28040 12368
rect 31392 12316 31444 12368
rect 29276 12248 29328 12300
rect 29644 12248 29696 12300
rect 27344 12223 27396 12232
rect 27344 12189 27353 12223
rect 27353 12189 27387 12223
rect 27387 12189 27396 12223
rect 27344 12180 27396 12189
rect 30840 12248 30892 12300
rect 33416 12291 33468 12300
rect 33416 12257 33425 12291
rect 33425 12257 33459 12291
rect 33459 12257 33468 12291
rect 33416 12248 33468 12257
rect 33692 12316 33744 12368
rect 26884 12112 26936 12164
rect 27068 12112 27120 12164
rect 27896 12112 27948 12164
rect 30288 12155 30340 12164
rect 30288 12121 30297 12155
rect 30297 12121 30331 12155
rect 30331 12121 30340 12155
rect 30288 12112 30340 12121
rect 31024 12112 31076 12164
rect 31668 12112 31720 12164
rect 33600 12155 33652 12164
rect 33600 12121 33609 12155
rect 33609 12121 33643 12155
rect 33643 12121 33652 12155
rect 33600 12112 33652 12121
rect 17408 12044 17460 12096
rect 18512 12044 18564 12096
rect 23296 12044 23348 12096
rect 24676 12044 24728 12096
rect 24860 12044 24912 12096
rect 25044 12044 25096 12096
rect 25504 12044 25556 12096
rect 34152 12087 34204 12096
rect 34152 12053 34161 12087
rect 34161 12053 34195 12087
rect 34195 12053 34204 12087
rect 34152 12044 34204 12053
rect 34520 12087 34572 12096
rect 34520 12053 34529 12087
rect 34529 12053 34563 12087
rect 34563 12053 34572 12087
rect 34520 12044 34572 12053
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 5448 11840 5500 11892
rect 6828 11883 6880 11892
rect 6828 11849 6837 11883
rect 6837 11849 6871 11883
rect 6871 11849 6880 11883
rect 6828 11840 6880 11849
rect 8944 11840 8996 11892
rect 6920 11772 6972 11824
rect 10968 11772 11020 11824
rect 940 11704 992 11756
rect 2136 11747 2188 11756
rect 2136 11713 2145 11747
rect 2145 11713 2179 11747
rect 2179 11713 2188 11747
rect 2136 11704 2188 11713
rect 7380 11747 7432 11756
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7380 11704 7432 11713
rect 8024 11704 8076 11756
rect 9036 11747 9088 11756
rect 9036 11713 9045 11747
rect 9045 11713 9079 11747
rect 9079 11713 9088 11747
rect 9036 11704 9088 11713
rect 9496 11704 9548 11756
rect 6644 11636 6696 11688
rect 6920 11679 6972 11688
rect 6920 11645 6929 11679
rect 6929 11645 6963 11679
rect 6963 11645 6972 11679
rect 6920 11636 6972 11645
rect 7104 11500 7156 11552
rect 8944 11636 8996 11688
rect 9220 11636 9272 11688
rect 9956 11679 10008 11688
rect 9956 11645 9965 11679
rect 9965 11645 9999 11679
rect 9999 11645 10008 11679
rect 9956 11636 10008 11645
rect 10140 11747 10192 11756
rect 10140 11713 10149 11747
rect 10149 11713 10183 11747
rect 10183 11713 10192 11747
rect 10140 11704 10192 11713
rect 12440 11772 12492 11824
rect 12992 11772 13044 11824
rect 14004 11883 14056 11892
rect 14004 11849 14013 11883
rect 14013 11849 14047 11883
rect 14047 11849 14056 11883
rect 14004 11840 14056 11849
rect 14188 11772 14240 11824
rect 14464 11772 14516 11824
rect 15016 11772 15068 11824
rect 10508 11679 10560 11688
rect 10508 11645 10517 11679
rect 10517 11645 10551 11679
rect 10551 11645 10560 11679
rect 10508 11636 10560 11645
rect 10692 11636 10744 11688
rect 14280 11747 14332 11756
rect 14280 11713 14289 11747
rect 14289 11713 14323 11747
rect 14323 11713 14332 11747
rect 14280 11704 14332 11713
rect 14648 11704 14700 11756
rect 12624 11636 12676 11688
rect 12992 11636 13044 11688
rect 15476 11747 15528 11756
rect 15476 11713 15485 11747
rect 15485 11713 15519 11747
rect 15519 11713 15528 11747
rect 15476 11704 15528 11713
rect 18512 11840 18564 11892
rect 18696 11840 18748 11892
rect 22468 11883 22520 11892
rect 22468 11849 22477 11883
rect 22477 11849 22511 11883
rect 22511 11849 22520 11883
rect 22468 11840 22520 11849
rect 15936 11636 15988 11688
rect 16580 11636 16632 11688
rect 17316 11704 17368 11756
rect 17776 11772 17828 11824
rect 18236 11815 18288 11824
rect 18236 11781 18245 11815
rect 18245 11781 18279 11815
rect 18279 11781 18288 11815
rect 18236 11772 18288 11781
rect 18420 11772 18472 11824
rect 17500 11704 17552 11756
rect 17684 11704 17736 11756
rect 18052 11747 18104 11756
rect 18052 11713 18059 11747
rect 18059 11713 18104 11747
rect 18052 11704 18104 11713
rect 11520 11568 11572 11620
rect 10508 11500 10560 11552
rect 12256 11500 12308 11552
rect 13084 11500 13136 11552
rect 15200 11543 15252 11552
rect 15200 11509 15209 11543
rect 15209 11509 15243 11543
rect 15243 11509 15252 11543
rect 15200 11500 15252 11509
rect 16488 11568 16540 11620
rect 17408 11568 17460 11620
rect 18420 11636 18472 11688
rect 18972 11747 19024 11756
rect 18972 11713 18981 11747
rect 18981 11713 19015 11747
rect 19015 11713 19024 11747
rect 18972 11704 19024 11713
rect 20904 11772 20956 11824
rect 21548 11772 21600 11824
rect 22100 11772 22152 11824
rect 22192 11772 22244 11824
rect 22284 11772 22336 11824
rect 23480 11772 23532 11824
rect 24124 11772 24176 11824
rect 18880 11636 18932 11688
rect 23296 11704 23348 11756
rect 27068 11840 27120 11892
rect 28448 11840 28500 11892
rect 30012 11840 30064 11892
rect 30288 11840 30340 11892
rect 34152 11840 34204 11892
rect 25136 11772 25188 11824
rect 25320 11772 25372 11824
rect 29368 11772 29420 11824
rect 26792 11704 26844 11756
rect 27988 11704 28040 11756
rect 16856 11500 16908 11552
rect 17132 11500 17184 11552
rect 17316 11500 17368 11552
rect 18604 11568 18656 11620
rect 23480 11636 23532 11688
rect 24768 11636 24820 11688
rect 25504 11636 25556 11688
rect 27344 11636 27396 11688
rect 27620 11636 27672 11688
rect 28540 11636 28592 11688
rect 34060 11772 34112 11824
rect 34520 11772 34572 11824
rect 29828 11747 29880 11756
rect 29828 11713 29837 11747
rect 29837 11713 29871 11747
rect 29871 11713 29880 11747
rect 29828 11704 29880 11713
rect 29920 11747 29972 11756
rect 29920 11713 29929 11747
rect 29929 11713 29963 11747
rect 29963 11713 29972 11747
rect 29920 11704 29972 11713
rect 30288 11704 30340 11756
rect 31300 11747 31352 11756
rect 31300 11713 31309 11747
rect 31309 11713 31343 11747
rect 31343 11713 31352 11747
rect 31300 11704 31352 11713
rect 37648 11747 37700 11756
rect 37648 11713 37657 11747
rect 37657 11713 37691 11747
rect 37691 11713 37700 11747
rect 37648 11704 37700 11713
rect 30196 11636 30248 11688
rect 33600 11636 33652 11688
rect 18512 11543 18564 11552
rect 18512 11509 18521 11543
rect 18521 11509 18555 11543
rect 18555 11509 18564 11543
rect 18512 11500 18564 11509
rect 20812 11500 20864 11552
rect 22100 11500 22152 11552
rect 23112 11500 23164 11552
rect 23940 11500 23992 11552
rect 24308 11500 24360 11552
rect 24492 11500 24544 11552
rect 27068 11568 27120 11620
rect 30380 11568 30432 11620
rect 37832 11611 37884 11620
rect 37832 11577 37841 11611
rect 37841 11577 37875 11611
rect 37875 11577 37884 11611
rect 37832 11568 37884 11577
rect 27712 11500 27764 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 2136 11296 2188 11348
rect 10140 11296 10192 11348
rect 12624 11296 12676 11348
rect 12900 11296 12952 11348
rect 7104 11160 7156 11212
rect 5632 11092 5684 11144
rect 6460 11135 6512 11144
rect 6460 11101 6469 11135
rect 6469 11101 6503 11135
rect 6503 11101 6512 11135
rect 6460 11092 6512 11101
rect 10876 11203 10928 11212
rect 10876 11169 10885 11203
rect 10885 11169 10919 11203
rect 10919 11169 10928 11203
rect 10876 11160 10928 11169
rect 10692 11135 10744 11144
rect 10692 11101 10701 11135
rect 10701 11101 10735 11135
rect 10735 11101 10744 11135
rect 10692 11092 10744 11101
rect 11704 11092 11756 11144
rect 13084 11160 13136 11212
rect 5448 11024 5500 11076
rect 6920 11024 6972 11076
rect 7748 11024 7800 11076
rect 12164 11135 12216 11144
rect 12164 11101 12173 11135
rect 12173 11101 12207 11135
rect 12207 11101 12216 11135
rect 12164 11092 12216 11101
rect 13820 11160 13872 11212
rect 14096 11160 14148 11212
rect 15108 11296 15160 11348
rect 15660 11296 15712 11348
rect 13452 11092 13504 11144
rect 14004 11092 14056 11144
rect 14188 11135 14240 11144
rect 14188 11101 14197 11135
rect 14197 11101 14231 11135
rect 14231 11101 14240 11135
rect 14188 11092 14240 11101
rect 14280 11135 14332 11144
rect 14280 11101 14290 11135
rect 14290 11101 14324 11135
rect 14324 11101 14332 11135
rect 15200 11160 15252 11212
rect 14280 11092 14332 11101
rect 14924 11092 14976 11144
rect 13820 11024 13872 11076
rect 14096 11024 14148 11076
rect 14464 11067 14516 11076
rect 14464 11033 14473 11067
rect 14473 11033 14507 11067
rect 14507 11033 14516 11067
rect 14464 11024 14516 11033
rect 14556 11067 14608 11076
rect 14556 11033 14565 11067
rect 14565 11033 14599 11067
rect 14599 11033 14608 11067
rect 14556 11024 14608 11033
rect 15568 11135 15620 11144
rect 15568 11101 15577 11135
rect 15577 11101 15611 11135
rect 15611 11101 15620 11135
rect 15568 11092 15620 11101
rect 16028 11296 16080 11348
rect 16212 11296 16264 11348
rect 16764 11339 16816 11348
rect 16764 11305 16773 11339
rect 16773 11305 16807 11339
rect 16807 11305 16816 11339
rect 16764 11296 16816 11305
rect 18420 11296 18472 11348
rect 19156 11296 19208 11348
rect 20168 11296 20220 11348
rect 16212 11203 16264 11212
rect 16212 11169 16221 11203
rect 16221 11169 16255 11203
rect 16255 11169 16264 11203
rect 16212 11160 16264 11169
rect 8484 10999 8536 11008
rect 8484 10965 8493 10999
rect 8493 10965 8527 10999
rect 8527 10965 8536 10999
rect 8484 10956 8536 10965
rect 11612 10956 11664 11008
rect 11980 10956 12032 11008
rect 12532 10956 12584 11008
rect 14280 10956 14332 11008
rect 15108 10956 15160 11008
rect 15476 10956 15528 11008
rect 17040 11024 17092 11076
rect 16580 10956 16632 11008
rect 17316 11135 17368 11144
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 17408 11135 17460 11144
rect 17408 11101 17418 11135
rect 17418 11101 17452 11135
rect 17452 11101 17460 11135
rect 17408 11092 17460 11101
rect 17224 11024 17276 11076
rect 18328 11203 18380 11212
rect 18328 11169 18337 11203
rect 18337 11169 18371 11203
rect 18371 11169 18380 11203
rect 18328 11160 18380 11169
rect 18420 11203 18472 11212
rect 18420 11169 18429 11203
rect 18429 11169 18463 11203
rect 18463 11169 18472 11203
rect 18420 11160 18472 11169
rect 17776 11135 17828 11144
rect 17776 11101 17790 11135
rect 17790 11101 17824 11135
rect 17824 11101 17828 11135
rect 17776 11092 17828 11101
rect 18512 11092 18564 11144
rect 18604 11135 18656 11144
rect 18604 11101 18613 11135
rect 18613 11101 18647 11135
rect 18647 11101 18656 11135
rect 18604 11092 18656 11101
rect 18972 11160 19024 11212
rect 20076 11271 20128 11280
rect 20076 11237 20085 11271
rect 20085 11237 20119 11271
rect 20119 11237 20128 11271
rect 20076 11228 20128 11237
rect 19432 11135 19484 11144
rect 19432 11101 19441 11135
rect 19441 11101 19475 11135
rect 19475 11101 19484 11135
rect 19432 11092 19484 11101
rect 20720 11203 20772 11212
rect 20720 11169 20729 11203
rect 20729 11169 20763 11203
rect 20763 11169 20772 11203
rect 20720 11160 20772 11169
rect 21640 11228 21692 11280
rect 20904 11160 20956 11212
rect 21824 11228 21876 11280
rect 22928 11228 22980 11280
rect 24492 11296 24544 11348
rect 18236 11024 18288 11076
rect 19708 11024 19760 11076
rect 20904 11024 20956 11076
rect 21272 11092 21324 11144
rect 21824 11092 21876 11144
rect 22192 11135 22244 11144
rect 22192 11101 22201 11135
rect 22201 11101 22235 11135
rect 22235 11101 22244 11135
rect 22192 11092 22244 11101
rect 22560 11135 22612 11144
rect 22560 11101 22569 11135
rect 22569 11101 22603 11135
rect 22603 11101 22612 11135
rect 22560 11092 22612 11101
rect 23664 11228 23716 11280
rect 24216 11228 24268 11280
rect 27528 11296 27580 11348
rect 28356 11339 28408 11348
rect 28356 11305 28365 11339
rect 28365 11305 28399 11339
rect 28399 11305 28408 11339
rect 28356 11296 28408 11305
rect 28448 11296 28500 11348
rect 28540 11296 28592 11348
rect 27620 11228 27672 11280
rect 23296 11135 23348 11144
rect 23296 11101 23305 11135
rect 23305 11101 23339 11135
rect 23339 11101 23348 11135
rect 23296 11092 23348 11101
rect 17500 10956 17552 11008
rect 18880 10956 18932 11008
rect 19248 10999 19300 11008
rect 19248 10965 19257 10999
rect 19257 10965 19291 10999
rect 19291 10965 19300 10999
rect 19248 10956 19300 10965
rect 22836 11024 22888 11076
rect 23756 11092 23808 11144
rect 23940 11092 23992 11144
rect 23480 11024 23532 11076
rect 24032 11024 24084 11076
rect 24952 11135 25004 11144
rect 24952 11101 24961 11135
rect 24961 11101 24995 11135
rect 24995 11101 25004 11135
rect 24952 11092 25004 11101
rect 25136 11135 25188 11144
rect 25136 11101 25145 11135
rect 25145 11101 25179 11135
rect 25179 11101 25188 11135
rect 25136 11092 25188 11101
rect 25504 11135 25556 11144
rect 25504 11101 25513 11135
rect 25513 11101 25547 11135
rect 25547 11101 25556 11135
rect 25504 11092 25556 11101
rect 25780 11135 25832 11144
rect 25780 11101 25789 11135
rect 25789 11101 25823 11135
rect 25823 11101 25832 11135
rect 25780 11092 25832 11101
rect 25872 11135 25924 11144
rect 25872 11101 25881 11135
rect 25881 11101 25915 11135
rect 25915 11101 25924 11135
rect 25872 11092 25924 11101
rect 26424 11092 26476 11144
rect 26516 11135 26568 11144
rect 26516 11101 26525 11135
rect 26525 11101 26559 11135
rect 26559 11101 26568 11135
rect 26516 11092 26568 11101
rect 26608 11135 26660 11144
rect 26608 11101 26617 11135
rect 26617 11101 26651 11135
rect 26651 11101 26660 11135
rect 26608 11092 26660 11101
rect 27804 11135 27856 11144
rect 27804 11101 27813 11135
rect 27813 11101 27847 11135
rect 27847 11101 27856 11135
rect 27804 11092 27856 11101
rect 28264 11092 28316 11144
rect 29460 11296 29512 11348
rect 29736 11135 29788 11144
rect 29736 11101 29745 11135
rect 29745 11101 29779 11135
rect 29779 11101 29788 11135
rect 29736 11092 29788 11101
rect 29828 11135 29880 11144
rect 29828 11101 29837 11135
rect 29837 11101 29871 11135
rect 29871 11101 29880 11135
rect 29828 11092 29880 11101
rect 30564 11228 30616 11280
rect 30380 11203 30432 11212
rect 30380 11169 30389 11203
rect 30389 11169 30423 11203
rect 30423 11169 30432 11203
rect 30380 11160 30432 11169
rect 30748 11160 30800 11212
rect 24952 10956 25004 11008
rect 25688 10956 25740 11008
rect 26424 10956 26476 11008
rect 28172 10956 28224 11008
rect 30840 11092 30892 11144
rect 31116 11092 31168 11144
rect 32496 10956 32548 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 7380 10752 7432 10804
rect 8484 10752 8536 10804
rect 8576 10752 8628 10804
rect 11796 10752 11848 10804
rect 12164 10752 12216 10804
rect 6920 10684 6972 10736
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 8668 10616 8720 10668
rect 11152 10684 11204 10736
rect 11612 10684 11664 10736
rect 4712 10412 4764 10464
rect 5816 10480 5868 10532
rect 6644 10548 6696 10600
rect 11520 10659 11572 10668
rect 11520 10625 11529 10659
rect 11529 10625 11563 10659
rect 11563 10625 11572 10659
rect 11520 10616 11572 10625
rect 12348 10684 12400 10736
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 9496 10591 9548 10600
rect 9496 10557 9505 10591
rect 9505 10557 9539 10591
rect 9539 10557 9548 10591
rect 9496 10548 9548 10557
rect 9864 10591 9916 10600
rect 9864 10557 9873 10591
rect 9873 10557 9907 10591
rect 9907 10557 9916 10591
rect 9864 10548 9916 10557
rect 11244 10548 11296 10600
rect 11888 10659 11940 10668
rect 11888 10625 11897 10659
rect 11897 10625 11931 10659
rect 11931 10625 11940 10659
rect 11888 10616 11940 10625
rect 12808 10752 12860 10804
rect 14096 10752 14148 10804
rect 14188 10752 14240 10804
rect 12900 10684 12952 10736
rect 15476 10752 15528 10804
rect 17040 10752 17092 10804
rect 17132 10752 17184 10804
rect 17316 10752 17368 10804
rect 17408 10752 17460 10804
rect 16764 10684 16816 10736
rect 17224 10727 17276 10736
rect 17224 10693 17233 10727
rect 17233 10693 17267 10727
rect 17267 10693 17276 10727
rect 17224 10684 17276 10693
rect 18420 10752 18472 10804
rect 18604 10752 18656 10804
rect 18880 10752 18932 10804
rect 20536 10752 20588 10804
rect 20904 10795 20956 10804
rect 20904 10761 20913 10795
rect 20913 10761 20947 10795
rect 20947 10761 20956 10795
rect 20904 10752 20956 10761
rect 12624 10659 12676 10668
rect 12624 10625 12633 10659
rect 12633 10625 12667 10659
rect 12667 10625 12676 10659
rect 12624 10616 12676 10625
rect 6828 10480 6880 10532
rect 8208 10480 8260 10532
rect 13636 10548 13688 10600
rect 12348 10480 12400 10532
rect 13084 10480 13136 10532
rect 6368 10412 6420 10464
rect 11612 10412 11664 10464
rect 11796 10412 11848 10464
rect 14004 10616 14056 10668
rect 14372 10616 14424 10668
rect 14556 10616 14608 10668
rect 15200 10616 15252 10668
rect 15568 10616 15620 10668
rect 14096 10548 14148 10600
rect 14464 10548 14516 10600
rect 15936 10659 15988 10668
rect 15936 10625 15945 10659
rect 15945 10625 15979 10659
rect 15979 10625 15988 10659
rect 15936 10616 15988 10625
rect 16120 10659 16172 10668
rect 16120 10625 16129 10659
rect 16129 10625 16163 10659
rect 16163 10625 16172 10659
rect 16120 10616 16172 10625
rect 16212 10616 16264 10668
rect 17040 10659 17092 10668
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 17040 10616 17092 10625
rect 16856 10548 16908 10600
rect 17316 10659 17368 10668
rect 17316 10625 17325 10659
rect 17325 10625 17359 10659
rect 17359 10625 17368 10659
rect 17316 10616 17368 10625
rect 17408 10659 17460 10668
rect 17408 10625 17417 10659
rect 17417 10625 17451 10659
rect 17451 10625 17460 10659
rect 17408 10616 17460 10625
rect 17960 10659 18012 10668
rect 17960 10625 17969 10659
rect 17969 10625 18003 10659
rect 18003 10625 18012 10659
rect 17960 10616 18012 10625
rect 18144 10616 18196 10668
rect 18512 10659 18564 10668
rect 18512 10625 18521 10659
rect 18521 10625 18555 10659
rect 18555 10625 18564 10659
rect 18512 10616 18564 10625
rect 18604 10616 18656 10668
rect 20812 10684 20864 10736
rect 22744 10752 22796 10804
rect 22928 10752 22980 10804
rect 23296 10795 23348 10804
rect 23296 10761 23305 10795
rect 23305 10761 23339 10795
rect 23339 10761 23348 10795
rect 23296 10752 23348 10761
rect 24492 10752 24544 10804
rect 25412 10752 25464 10804
rect 19064 10659 19116 10668
rect 19064 10625 19073 10659
rect 19073 10625 19107 10659
rect 19107 10625 19116 10659
rect 19064 10616 19116 10625
rect 19248 10616 19300 10668
rect 20720 10616 20772 10668
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 21088 10616 21140 10625
rect 14188 10412 14240 10464
rect 17224 10480 17276 10532
rect 17592 10480 17644 10532
rect 17960 10480 18012 10532
rect 18880 10548 18932 10600
rect 19524 10548 19576 10600
rect 16580 10412 16632 10464
rect 17776 10412 17828 10464
rect 20536 10480 20588 10532
rect 21364 10659 21416 10668
rect 21364 10625 21373 10659
rect 21373 10625 21407 10659
rect 21407 10625 21416 10659
rect 21364 10616 21416 10625
rect 21548 10684 21600 10736
rect 22468 10684 22520 10736
rect 21732 10616 21784 10668
rect 22836 10659 22888 10668
rect 22836 10625 22845 10659
rect 22845 10625 22879 10659
rect 22879 10625 22888 10659
rect 22836 10616 22888 10625
rect 22928 10616 22980 10668
rect 26608 10752 26660 10804
rect 27804 10752 27856 10804
rect 29184 10752 29236 10804
rect 25228 10616 25280 10668
rect 25688 10659 25740 10668
rect 25688 10625 25698 10659
rect 25698 10625 25732 10659
rect 25732 10625 25740 10659
rect 25688 10616 25740 10625
rect 23480 10548 23532 10600
rect 24124 10548 24176 10600
rect 24768 10548 24820 10600
rect 25504 10548 25556 10600
rect 28172 10684 28224 10736
rect 28816 10727 28868 10736
rect 28816 10693 28825 10727
rect 28825 10693 28859 10727
rect 28859 10693 28868 10727
rect 28816 10684 28868 10693
rect 29828 10795 29880 10804
rect 29828 10761 29837 10795
rect 29837 10761 29871 10795
rect 29871 10761 29880 10795
rect 29828 10752 29880 10761
rect 31024 10752 31076 10804
rect 31576 10752 31628 10804
rect 25964 10659 26016 10668
rect 25964 10625 25973 10659
rect 25973 10625 26007 10659
rect 26007 10625 26016 10659
rect 25964 10616 26016 10625
rect 26148 10616 26200 10668
rect 27712 10616 27764 10668
rect 28356 10616 28408 10668
rect 28724 10616 28776 10668
rect 28080 10591 28132 10600
rect 28080 10557 28089 10591
rect 28089 10557 28123 10591
rect 28123 10557 28132 10591
rect 28080 10548 28132 10557
rect 28540 10548 28592 10600
rect 29000 10616 29052 10668
rect 24032 10480 24084 10532
rect 25412 10480 25464 10532
rect 22468 10412 22520 10464
rect 23204 10412 23256 10464
rect 25136 10412 25188 10464
rect 26884 10412 26936 10464
rect 27896 10412 27948 10464
rect 28172 10455 28224 10464
rect 28172 10421 28181 10455
rect 28181 10421 28215 10455
rect 28215 10421 28224 10455
rect 28172 10412 28224 10421
rect 28632 10412 28684 10464
rect 29552 10659 29604 10668
rect 29552 10625 29561 10659
rect 29561 10625 29595 10659
rect 29595 10625 29604 10659
rect 29552 10616 29604 10625
rect 29644 10659 29696 10668
rect 29644 10625 29653 10659
rect 29653 10625 29687 10659
rect 29687 10625 29696 10659
rect 29644 10616 29696 10625
rect 30012 10616 30064 10668
rect 32588 10684 32640 10736
rect 32496 10659 32548 10668
rect 32496 10625 32505 10659
rect 32505 10625 32539 10659
rect 32539 10625 32548 10659
rect 32496 10616 32548 10625
rect 32588 10591 32640 10600
rect 32588 10557 32597 10591
rect 32597 10557 32631 10591
rect 32631 10557 32640 10591
rect 32588 10548 32640 10557
rect 32680 10591 32732 10600
rect 32680 10557 32689 10591
rect 32689 10557 32723 10591
rect 32723 10557 32732 10591
rect 32680 10548 32732 10557
rect 33232 10591 33284 10600
rect 33232 10557 33241 10591
rect 33241 10557 33275 10591
rect 33275 10557 33284 10591
rect 33232 10548 33284 10557
rect 33324 10548 33376 10600
rect 29460 10480 29512 10532
rect 31300 10412 31352 10464
rect 34520 10412 34572 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 4712 10208 4764 10260
rect 3976 10072 4028 10124
rect 4620 10072 4672 10124
rect 6368 10115 6420 10124
rect 6368 10081 6377 10115
rect 6377 10081 6411 10115
rect 6411 10081 6420 10115
rect 6368 10072 6420 10081
rect 6736 10072 6788 10124
rect 8668 10208 8720 10260
rect 9404 10208 9456 10260
rect 12900 10208 12952 10260
rect 13084 10208 13136 10260
rect 15200 10208 15252 10260
rect 15384 10251 15436 10260
rect 15384 10217 15393 10251
rect 15393 10217 15427 10251
rect 15427 10217 15436 10251
rect 15384 10208 15436 10217
rect 15752 10208 15804 10260
rect 18144 10208 18196 10260
rect 19340 10208 19392 10260
rect 21088 10208 21140 10260
rect 22100 10251 22152 10260
rect 22100 10217 22109 10251
rect 22109 10217 22143 10251
rect 22143 10217 22152 10251
rect 22100 10208 22152 10217
rect 22836 10208 22888 10260
rect 23848 10208 23900 10260
rect 24124 10208 24176 10260
rect 25872 10208 25924 10260
rect 28080 10208 28132 10260
rect 28540 10208 28592 10260
rect 29736 10208 29788 10260
rect 32496 10208 32548 10260
rect 11612 10140 11664 10192
rect 11888 10140 11940 10192
rect 16948 10140 17000 10192
rect 17040 10140 17092 10192
rect 17960 10140 18012 10192
rect 8116 10072 8168 10124
rect 6184 9936 6236 9988
rect 6552 9911 6604 9920
rect 6552 9877 6561 9911
rect 6561 9877 6595 9911
rect 6595 9877 6604 9911
rect 6552 9868 6604 9877
rect 6828 9911 6880 9920
rect 6828 9877 6837 9911
rect 6837 9877 6871 9911
rect 6871 9877 6880 9911
rect 6828 9868 6880 9877
rect 8576 10004 8628 10056
rect 12624 10004 12676 10056
rect 15752 10072 15804 10124
rect 17316 10072 17368 10124
rect 13544 10004 13596 10056
rect 14556 10004 14608 10056
rect 14740 10004 14792 10056
rect 15200 10047 15252 10056
rect 15200 10013 15209 10047
rect 15209 10013 15243 10047
rect 15243 10013 15252 10047
rect 15200 10004 15252 10013
rect 8208 9868 8260 9920
rect 10968 9936 11020 9988
rect 11336 9936 11388 9988
rect 11612 9936 11664 9988
rect 16948 10004 17000 10056
rect 17408 10047 17460 10056
rect 17408 10013 17417 10047
rect 17417 10013 17451 10047
rect 17451 10013 17460 10047
rect 17408 10004 17460 10013
rect 17316 9936 17368 9988
rect 17868 10047 17920 10056
rect 17868 10013 17877 10047
rect 17877 10013 17911 10047
rect 17911 10013 17920 10047
rect 17868 10004 17920 10013
rect 18052 10047 18104 10056
rect 18052 10013 18061 10047
rect 18061 10013 18095 10047
rect 18095 10013 18104 10047
rect 18052 10004 18104 10013
rect 17960 9936 18012 9988
rect 21548 10140 21600 10192
rect 22928 10140 22980 10192
rect 26240 10140 26292 10192
rect 27252 10140 27304 10192
rect 28172 10140 28224 10192
rect 18880 10072 18932 10124
rect 23388 10072 23440 10124
rect 9496 9868 9548 9920
rect 10232 9868 10284 9920
rect 11520 9868 11572 9920
rect 11888 9868 11940 9920
rect 12164 9868 12216 9920
rect 15384 9868 15436 9920
rect 15568 9911 15620 9920
rect 15568 9877 15577 9911
rect 15577 9877 15611 9911
rect 15611 9877 15620 9911
rect 15568 9868 15620 9877
rect 15752 9868 15804 9920
rect 15936 9868 15988 9920
rect 19064 9868 19116 9920
rect 19156 9868 19208 9920
rect 19524 10004 19576 10056
rect 19616 10004 19668 10056
rect 19892 10004 19944 10056
rect 19524 9868 19576 9920
rect 20444 10047 20496 10056
rect 20444 10013 20458 10047
rect 20458 10013 20492 10047
rect 20492 10013 20496 10047
rect 20444 10004 20496 10013
rect 21640 10004 21692 10056
rect 22100 10004 22152 10056
rect 22560 10047 22612 10056
rect 22560 10013 22569 10047
rect 22569 10013 22603 10047
rect 22603 10013 22612 10047
rect 22560 10004 22612 10013
rect 23480 10004 23532 10056
rect 23848 10047 23900 10056
rect 23848 10013 23857 10047
rect 23857 10013 23891 10047
rect 23891 10013 23900 10047
rect 23848 10004 23900 10013
rect 23664 9936 23716 9988
rect 24032 10004 24084 10056
rect 24952 10047 25004 10056
rect 24952 10013 24961 10047
rect 24961 10013 24995 10047
rect 24995 10013 25004 10047
rect 24952 10004 25004 10013
rect 25688 10004 25740 10056
rect 27620 10072 27672 10124
rect 27804 10072 27856 10124
rect 27988 10004 28040 10056
rect 20444 9868 20496 9920
rect 22468 9911 22520 9920
rect 22468 9877 22477 9911
rect 22477 9877 22511 9911
rect 22511 9877 22520 9911
rect 22468 9868 22520 9877
rect 25964 9936 26016 9988
rect 25596 9868 25648 9920
rect 27620 9868 27672 9920
rect 28172 9979 28224 9988
rect 28172 9945 28181 9979
rect 28181 9945 28215 9979
rect 28215 9945 28224 9979
rect 29552 10140 29604 10192
rect 28448 10072 28500 10124
rect 28816 10004 28868 10056
rect 29000 10072 29052 10124
rect 29736 10072 29788 10124
rect 30380 10072 30432 10124
rect 30656 10072 30708 10124
rect 31300 10115 31352 10124
rect 31300 10081 31309 10115
rect 31309 10081 31343 10115
rect 31343 10081 31352 10115
rect 31300 10072 31352 10081
rect 31852 10072 31904 10124
rect 29184 10004 29236 10056
rect 33140 10004 33192 10056
rect 28172 9936 28224 9945
rect 31300 9936 31352 9988
rect 31576 9936 31628 9988
rect 28816 9911 28868 9920
rect 28816 9877 28841 9911
rect 28841 9877 28868 9911
rect 28816 9868 28868 9877
rect 29552 9868 29604 9920
rect 32772 9868 32824 9920
rect 35072 9868 35124 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 6552 9664 6604 9716
rect 6828 9664 6880 9716
rect 6920 9664 6972 9716
rect 8208 9664 8260 9716
rect 10784 9664 10836 9716
rect 7748 9528 7800 9580
rect 7932 9528 7984 9580
rect 9864 9596 9916 9648
rect 11612 9664 11664 9716
rect 11888 9664 11940 9716
rect 10968 9528 11020 9580
rect 6184 9460 6236 9512
rect 9864 9503 9916 9512
rect 9864 9469 9873 9503
rect 9873 9469 9907 9503
rect 9907 9469 9916 9503
rect 9864 9460 9916 9469
rect 10600 9460 10652 9512
rect 12164 9596 12216 9648
rect 13912 9639 13964 9648
rect 13912 9605 13921 9639
rect 13921 9605 13955 9639
rect 13955 9605 13964 9639
rect 13912 9596 13964 9605
rect 15568 9596 15620 9648
rect 16672 9664 16724 9716
rect 13360 9528 13412 9580
rect 15292 9528 15344 9580
rect 15660 9528 15712 9580
rect 15844 9571 15896 9580
rect 15844 9537 15853 9571
rect 15853 9537 15887 9571
rect 15887 9537 15896 9571
rect 15844 9528 15896 9537
rect 15936 9571 15988 9580
rect 15936 9537 15945 9571
rect 15945 9537 15979 9571
rect 15979 9537 15988 9571
rect 15936 9528 15988 9537
rect 16120 9571 16172 9580
rect 16120 9537 16129 9571
rect 16129 9537 16163 9571
rect 16163 9537 16172 9571
rect 16120 9528 16172 9537
rect 16948 9596 17000 9648
rect 10876 9392 10928 9444
rect 11520 9460 11572 9512
rect 12992 9460 13044 9512
rect 13268 9392 13320 9444
rect 14280 9392 14332 9444
rect 10416 9324 10468 9376
rect 11520 9324 11572 9376
rect 11796 9324 11848 9376
rect 12348 9324 12400 9376
rect 14464 9324 14516 9376
rect 16672 9528 16724 9580
rect 17500 9596 17552 9648
rect 17776 9707 17828 9716
rect 17776 9673 17785 9707
rect 17785 9673 17819 9707
rect 17819 9673 17828 9707
rect 17776 9664 17828 9673
rect 18512 9664 18564 9716
rect 20168 9664 20220 9716
rect 20904 9664 20956 9716
rect 21364 9664 21416 9716
rect 21548 9664 21600 9716
rect 19064 9596 19116 9648
rect 21272 9596 21324 9648
rect 22652 9664 22704 9716
rect 24216 9664 24268 9716
rect 23204 9596 23256 9648
rect 23940 9639 23992 9648
rect 23940 9605 23949 9639
rect 23949 9605 23983 9639
rect 23983 9605 23992 9639
rect 23940 9596 23992 9605
rect 24952 9664 25004 9716
rect 16764 9460 16816 9512
rect 16488 9392 16540 9444
rect 17040 9392 17092 9444
rect 16948 9324 17000 9376
rect 17408 9571 17460 9580
rect 17408 9537 17417 9571
rect 17417 9537 17451 9571
rect 17451 9537 17460 9571
rect 17408 9528 17460 9537
rect 18052 9528 18104 9580
rect 19340 9571 19392 9580
rect 19340 9537 19349 9571
rect 19349 9537 19383 9571
rect 19383 9537 19392 9571
rect 19340 9528 19392 9537
rect 20076 9528 20128 9580
rect 21824 9528 21876 9580
rect 22836 9528 22888 9580
rect 23572 9528 23624 9580
rect 23664 9571 23716 9580
rect 23664 9537 23673 9571
rect 23673 9537 23707 9571
rect 23707 9537 23716 9571
rect 23664 9528 23716 9537
rect 23756 9528 23808 9580
rect 24676 9639 24728 9648
rect 24676 9605 24685 9639
rect 24685 9605 24719 9639
rect 24719 9605 24728 9639
rect 24676 9596 24728 9605
rect 24860 9639 24912 9648
rect 24860 9605 24869 9639
rect 24869 9605 24903 9639
rect 24903 9605 24912 9639
rect 24860 9596 24912 9605
rect 26700 9596 26752 9648
rect 25872 9571 25924 9580
rect 25872 9537 25876 9571
rect 25876 9537 25910 9571
rect 25910 9537 25924 9571
rect 20260 9460 20312 9512
rect 20444 9460 20496 9512
rect 17500 9392 17552 9444
rect 22928 9435 22980 9444
rect 22928 9401 22937 9435
rect 22937 9401 22971 9435
rect 22971 9401 22980 9435
rect 22928 9392 22980 9401
rect 24676 9460 24728 9512
rect 25872 9528 25924 9537
rect 26148 9528 26200 9580
rect 26240 9571 26292 9580
rect 26240 9537 26248 9571
rect 26248 9537 26282 9571
rect 26282 9537 26292 9571
rect 26240 9528 26292 9537
rect 26608 9528 26660 9580
rect 26976 9528 27028 9580
rect 27160 9571 27212 9580
rect 27160 9537 27169 9571
rect 27169 9537 27203 9571
rect 27203 9537 27212 9571
rect 27160 9528 27212 9537
rect 28172 9664 28224 9716
rect 28080 9596 28132 9648
rect 28448 9664 28500 9716
rect 28816 9664 28868 9716
rect 33324 9707 33376 9716
rect 33324 9673 33333 9707
rect 33333 9673 33367 9707
rect 33367 9673 33376 9707
rect 33324 9664 33376 9673
rect 29368 9596 29420 9648
rect 30104 9596 30156 9648
rect 33508 9596 33560 9648
rect 34520 9596 34572 9648
rect 29460 9528 29512 9580
rect 28356 9460 28408 9512
rect 29920 9571 29972 9580
rect 29920 9537 29929 9571
rect 29929 9537 29963 9571
rect 29963 9537 29972 9571
rect 29920 9528 29972 9537
rect 30288 9528 30340 9580
rect 32772 9571 32824 9580
rect 32772 9537 32781 9571
rect 32781 9537 32815 9571
rect 32815 9537 32824 9571
rect 32772 9528 32824 9537
rect 31300 9460 31352 9512
rect 31944 9460 31996 9512
rect 24032 9392 24084 9444
rect 24584 9392 24636 9444
rect 25320 9392 25372 9444
rect 25780 9392 25832 9444
rect 26516 9392 26568 9444
rect 27252 9392 27304 9444
rect 29920 9392 29972 9444
rect 32588 9392 32640 9444
rect 17868 9324 17920 9376
rect 17960 9324 18012 9376
rect 19800 9324 19852 9376
rect 20628 9367 20680 9376
rect 20628 9333 20637 9367
rect 20637 9333 20671 9367
rect 20671 9333 20680 9367
rect 20628 9324 20680 9333
rect 20812 9324 20864 9376
rect 22284 9324 22336 9376
rect 22468 9367 22520 9376
rect 22468 9333 22477 9367
rect 22477 9333 22511 9367
rect 22511 9333 22520 9367
rect 22468 9324 22520 9333
rect 23480 9324 23532 9376
rect 30472 9324 30524 9376
rect 32404 9367 32456 9376
rect 32404 9333 32413 9367
rect 32413 9333 32447 9367
rect 32447 9333 32456 9367
rect 32404 9324 32456 9333
rect 32772 9324 32824 9376
rect 33324 9460 33376 9512
rect 33692 9528 33744 9580
rect 34428 9460 34480 9512
rect 35072 9503 35124 9512
rect 35072 9469 35081 9503
rect 35081 9469 35115 9503
rect 35115 9469 35124 9503
rect 35072 9460 35124 9469
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 9864 9120 9916 9172
rect 11152 9120 11204 9172
rect 12348 9120 12400 9172
rect 10968 9052 11020 9104
rect 12900 9052 12952 9104
rect 12992 9052 13044 9104
rect 15936 9120 15988 9172
rect 4620 8959 4672 8968
rect 4620 8925 4629 8959
rect 4629 8925 4663 8959
rect 4663 8925 4672 8959
rect 4620 8916 4672 8925
rect 4528 8823 4580 8832
rect 4528 8789 4537 8823
rect 4537 8789 4571 8823
rect 4571 8789 4580 8823
rect 4528 8780 4580 8789
rect 6920 8780 6972 8832
rect 10876 8916 10928 8968
rect 11336 8984 11388 9036
rect 12072 9027 12124 9036
rect 12072 8993 12081 9027
rect 12081 8993 12115 9027
rect 12115 8993 12124 9027
rect 12072 8984 12124 8993
rect 14924 9052 14976 9104
rect 15384 9052 15436 9104
rect 11152 8959 11204 8968
rect 11152 8925 11161 8959
rect 11161 8925 11195 8959
rect 11195 8925 11204 8959
rect 11152 8916 11204 8925
rect 11336 8848 11388 8900
rect 12992 8916 13044 8968
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 13636 8959 13688 8968
rect 13636 8925 13645 8959
rect 13645 8925 13679 8959
rect 13679 8925 13688 8959
rect 13636 8916 13688 8925
rect 13728 8959 13780 8968
rect 13728 8925 13737 8959
rect 13737 8925 13771 8959
rect 13771 8925 13780 8959
rect 13728 8916 13780 8925
rect 13912 8959 13964 8968
rect 13912 8925 13921 8959
rect 13921 8925 13955 8959
rect 13955 8925 13964 8959
rect 13912 8916 13964 8925
rect 14280 8916 14332 8968
rect 15200 8916 15252 8968
rect 17316 9052 17368 9104
rect 15660 8984 15712 9036
rect 15752 8959 15804 8968
rect 15752 8925 15761 8959
rect 15761 8925 15795 8959
rect 15795 8925 15804 8959
rect 15752 8916 15804 8925
rect 13820 8848 13872 8900
rect 17868 8959 17920 8968
rect 17868 8925 17877 8959
rect 17877 8925 17911 8959
rect 17911 8925 17920 8959
rect 17868 8916 17920 8925
rect 20444 9120 20496 9172
rect 18512 9095 18564 9104
rect 18512 9061 18521 9095
rect 18521 9061 18555 9095
rect 18555 9061 18564 9095
rect 18512 9052 18564 9061
rect 18696 9052 18748 9104
rect 19616 9095 19668 9104
rect 19616 9061 19625 9095
rect 19625 9061 19659 9095
rect 19659 9061 19668 9095
rect 19616 9052 19668 9061
rect 19800 9052 19852 9104
rect 18328 8916 18380 8968
rect 19616 8916 19668 8968
rect 20168 9052 20220 9104
rect 20536 9052 20588 9104
rect 20996 9163 21048 9172
rect 20996 9129 21005 9163
rect 21005 9129 21039 9163
rect 21039 9129 21048 9163
rect 20996 9120 21048 9129
rect 21640 9120 21692 9172
rect 23112 9120 23164 9172
rect 23664 9120 23716 9172
rect 25228 9120 25280 9172
rect 25320 9120 25372 9172
rect 28264 9120 28316 9172
rect 28816 9163 28868 9172
rect 28816 9129 28825 9163
rect 28825 9129 28859 9163
rect 28859 9129 28868 9163
rect 28816 9120 28868 9129
rect 29000 9163 29052 9172
rect 29000 9129 29009 9163
rect 29009 9129 29043 9163
rect 29043 9129 29052 9163
rect 29000 9120 29052 9129
rect 30104 9163 30156 9172
rect 30104 9129 30113 9163
rect 30113 9129 30147 9163
rect 30147 9129 30156 9163
rect 30104 9120 30156 9129
rect 19248 8848 19300 8900
rect 20536 8959 20588 8968
rect 20536 8925 20545 8959
rect 20545 8925 20579 8959
rect 20579 8925 20588 8959
rect 20536 8916 20588 8925
rect 21824 8984 21876 9036
rect 22836 9052 22888 9104
rect 28724 9052 28776 9104
rect 30840 9120 30892 9172
rect 31944 9163 31996 9172
rect 31944 9129 31953 9163
rect 31953 9129 31987 9163
rect 31987 9129 31996 9163
rect 31944 9120 31996 9129
rect 32404 9120 32456 9172
rect 34428 9163 34480 9172
rect 34428 9129 34437 9163
rect 34437 9129 34471 9163
rect 34471 9129 34480 9163
rect 34428 9120 34480 9129
rect 21180 8916 21232 8968
rect 21548 8959 21600 8968
rect 21548 8925 21557 8959
rect 21557 8925 21591 8959
rect 21591 8925 21600 8959
rect 21548 8916 21600 8925
rect 21916 8959 21968 8968
rect 21916 8925 21925 8959
rect 21925 8925 21959 8959
rect 21959 8925 21968 8959
rect 21916 8916 21968 8925
rect 24400 9027 24452 9036
rect 24400 8993 24409 9027
rect 24409 8993 24443 9027
rect 24443 8993 24452 9027
rect 24400 8984 24452 8993
rect 25044 8984 25096 9036
rect 20812 8848 20864 8900
rect 12348 8780 12400 8832
rect 12900 8780 12952 8832
rect 15384 8780 15436 8832
rect 18328 8780 18380 8832
rect 20444 8780 20496 8832
rect 21180 8780 21232 8832
rect 21824 8891 21876 8900
rect 21824 8857 21833 8891
rect 21833 8857 21867 8891
rect 21867 8857 21876 8891
rect 21824 8848 21876 8857
rect 22468 8891 22520 8900
rect 22468 8857 22477 8891
rect 22477 8857 22511 8891
rect 22511 8857 22520 8891
rect 22468 8848 22520 8857
rect 22560 8848 22612 8900
rect 22928 8916 22980 8968
rect 24584 8916 24636 8968
rect 26240 9027 26292 9036
rect 26240 8993 26249 9027
rect 26249 8993 26283 9027
rect 26283 8993 26292 9027
rect 26240 8984 26292 8993
rect 26424 8984 26476 9036
rect 28908 8984 28960 9036
rect 25780 8959 25832 8968
rect 25780 8925 25789 8959
rect 25789 8925 25823 8959
rect 25823 8925 25832 8959
rect 25780 8916 25832 8925
rect 25872 8916 25924 8968
rect 27436 8916 27488 8968
rect 28172 8916 28224 8968
rect 27896 8891 27948 8900
rect 27896 8857 27905 8891
rect 27905 8857 27939 8891
rect 27939 8857 27948 8891
rect 27896 8848 27948 8857
rect 29552 8959 29604 8968
rect 29552 8925 29561 8959
rect 29561 8925 29595 8959
rect 29595 8925 29604 8959
rect 29552 8916 29604 8925
rect 31576 9052 31628 9104
rect 30472 9027 30524 9036
rect 30472 8993 30481 9027
rect 30481 8993 30515 9027
rect 30515 8993 30524 9027
rect 30472 8984 30524 8993
rect 29920 8959 29972 8968
rect 29920 8925 29929 8959
rect 29929 8925 29963 8959
rect 29963 8925 29972 8959
rect 29920 8916 29972 8925
rect 30196 8959 30248 8968
rect 30196 8925 30205 8959
rect 30205 8925 30239 8959
rect 30239 8925 30248 8959
rect 30196 8916 30248 8925
rect 30564 8848 30616 8900
rect 33692 8984 33744 9036
rect 32680 8959 32732 8968
rect 32680 8925 32689 8959
rect 32689 8925 32723 8959
rect 32723 8925 32732 8959
rect 32680 8916 32732 8925
rect 22284 8780 22336 8832
rect 26148 8780 26200 8832
rect 33692 8848 33744 8900
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 4528 8576 4580 8628
rect 10416 8576 10468 8628
rect 12348 8576 12400 8628
rect 14096 8576 14148 8628
rect 6092 8508 6144 8560
rect 6184 8551 6236 8560
rect 6184 8517 6193 8551
rect 6193 8517 6227 8551
rect 6227 8517 6236 8551
rect 6184 8508 6236 8517
rect 11152 8508 11204 8560
rect 12072 8508 12124 8560
rect 14280 8508 14332 8560
rect 6920 8440 6972 8492
rect 14464 8440 14516 8492
rect 4896 8372 4948 8424
rect 10508 8372 10560 8424
rect 16120 8576 16172 8628
rect 17868 8576 17920 8628
rect 18420 8576 18472 8628
rect 19800 8576 19852 8628
rect 20812 8576 20864 8628
rect 21088 8576 21140 8628
rect 19156 8508 19208 8560
rect 20076 8551 20128 8560
rect 20076 8517 20085 8551
rect 20085 8517 20119 8551
rect 20119 8517 20128 8551
rect 20076 8508 20128 8517
rect 20352 8508 20404 8560
rect 15016 8483 15068 8492
rect 15016 8449 15025 8483
rect 15025 8449 15059 8483
rect 15059 8449 15068 8483
rect 15016 8440 15068 8449
rect 15108 8483 15160 8492
rect 15108 8449 15117 8483
rect 15117 8449 15151 8483
rect 15151 8449 15160 8483
rect 15108 8440 15160 8449
rect 16488 8440 16540 8492
rect 17040 8440 17092 8492
rect 17960 8440 18012 8492
rect 16212 8372 16264 8424
rect 17592 8372 17644 8424
rect 19616 8440 19668 8492
rect 20260 8483 20312 8492
rect 20260 8449 20274 8483
rect 20274 8449 20308 8483
rect 20308 8449 20312 8483
rect 20260 8440 20312 8449
rect 12164 8304 12216 8356
rect 13084 8304 13136 8356
rect 13452 8347 13504 8356
rect 13452 8313 13461 8347
rect 13461 8313 13495 8347
rect 13495 8313 13504 8347
rect 13452 8304 13504 8313
rect 13820 8304 13872 8356
rect 7196 8236 7248 8288
rect 11612 8236 11664 8288
rect 15016 8236 15068 8288
rect 15384 8279 15436 8288
rect 15384 8245 15393 8279
rect 15393 8245 15427 8279
rect 15427 8245 15436 8279
rect 15384 8236 15436 8245
rect 15660 8236 15712 8288
rect 16304 8236 16356 8288
rect 16856 8236 16908 8288
rect 19616 8236 19668 8288
rect 19892 8304 19944 8356
rect 20168 8304 20220 8356
rect 20904 8440 20956 8492
rect 21088 8483 21140 8492
rect 21088 8449 21097 8483
rect 21097 8449 21131 8483
rect 21131 8449 21140 8483
rect 21088 8440 21140 8449
rect 21456 8576 21508 8628
rect 21272 8551 21324 8560
rect 21272 8517 21281 8551
rect 21281 8517 21315 8551
rect 21315 8517 21324 8551
rect 21272 8508 21324 8517
rect 21916 8508 21968 8560
rect 22468 8576 22520 8628
rect 22652 8576 22704 8628
rect 22284 8508 22336 8560
rect 21456 8483 21508 8492
rect 21456 8449 21465 8483
rect 21465 8449 21499 8483
rect 21499 8449 21508 8483
rect 21456 8440 21508 8449
rect 21640 8440 21692 8492
rect 21916 8372 21968 8424
rect 22744 8483 22796 8492
rect 22744 8449 22753 8483
rect 22753 8449 22787 8483
rect 22787 8449 22796 8483
rect 22744 8440 22796 8449
rect 22836 8483 22888 8492
rect 22836 8449 22845 8483
rect 22845 8449 22879 8483
rect 22879 8449 22888 8483
rect 22836 8440 22888 8449
rect 23480 8551 23532 8560
rect 23480 8517 23489 8551
rect 23489 8517 23523 8551
rect 23523 8517 23532 8551
rect 23480 8508 23532 8517
rect 23112 8483 23164 8492
rect 23112 8449 23121 8483
rect 23121 8449 23155 8483
rect 23155 8449 23164 8483
rect 23112 8440 23164 8449
rect 23296 8440 23348 8492
rect 23572 8483 23624 8492
rect 23572 8449 23581 8483
rect 23581 8449 23615 8483
rect 23615 8449 23624 8483
rect 23572 8440 23624 8449
rect 23848 8483 23900 8492
rect 23848 8449 23857 8483
rect 23857 8449 23891 8483
rect 23891 8449 23900 8483
rect 23848 8440 23900 8449
rect 23940 8440 23992 8492
rect 24032 8440 24084 8492
rect 26056 8576 26108 8628
rect 26148 8576 26200 8628
rect 29920 8576 29972 8628
rect 30196 8576 30248 8628
rect 31668 8576 31720 8628
rect 32680 8576 32732 8628
rect 25780 8508 25832 8560
rect 22560 8304 22612 8356
rect 22652 8304 22704 8356
rect 25044 8372 25096 8424
rect 25964 8483 26016 8492
rect 25964 8449 25973 8483
rect 25973 8449 26007 8483
rect 26007 8449 26016 8483
rect 25964 8440 26016 8449
rect 26792 8551 26844 8560
rect 26792 8517 26801 8551
rect 26801 8517 26835 8551
rect 26835 8517 26844 8551
rect 26792 8508 26844 8517
rect 27896 8551 27948 8560
rect 27896 8517 27913 8551
rect 27913 8517 27948 8551
rect 27896 8508 27948 8517
rect 28724 8551 28776 8560
rect 28724 8517 28733 8551
rect 28733 8517 28767 8551
rect 28767 8517 28776 8551
rect 28724 8508 28776 8517
rect 28908 8551 28960 8560
rect 28908 8517 28917 8551
rect 28917 8517 28951 8551
rect 28951 8517 28960 8551
rect 28908 8508 28960 8517
rect 30932 8508 30984 8560
rect 26332 8440 26384 8492
rect 27436 8440 27488 8492
rect 27712 8483 27764 8492
rect 27712 8449 27721 8483
rect 27721 8449 27755 8483
rect 27755 8449 27764 8483
rect 27712 8440 27764 8449
rect 27988 8483 28040 8492
rect 27988 8449 27997 8483
rect 27997 8449 28031 8483
rect 28031 8449 28040 8483
rect 27988 8440 28040 8449
rect 28172 8483 28224 8492
rect 28172 8449 28181 8483
rect 28181 8449 28215 8483
rect 28215 8449 28224 8483
rect 28172 8440 28224 8449
rect 28264 8440 28316 8492
rect 28632 8483 28684 8492
rect 28632 8449 28641 8483
rect 28641 8449 28675 8483
rect 28675 8449 28684 8483
rect 28632 8440 28684 8449
rect 31852 8440 31904 8492
rect 28356 8304 28408 8356
rect 21180 8236 21232 8288
rect 23572 8236 23624 8288
rect 23756 8236 23808 8288
rect 31668 8236 31720 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 4896 8075 4948 8084
rect 4896 8041 4905 8075
rect 4905 8041 4939 8075
rect 4939 8041 4948 8075
rect 4896 8032 4948 8041
rect 6828 8032 6880 8084
rect 7932 8032 7984 8084
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 6184 7828 6236 7880
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 10968 8032 11020 8084
rect 11428 8032 11480 8084
rect 13912 8032 13964 8084
rect 14832 8032 14884 8084
rect 15108 8032 15160 8084
rect 16764 8075 16816 8084
rect 16764 8041 16773 8075
rect 16773 8041 16807 8075
rect 16807 8041 16816 8075
rect 16764 8032 16816 8041
rect 17316 8032 17368 8084
rect 9956 7964 10008 8016
rect 10232 7964 10284 8016
rect 8668 7896 8720 7948
rect 10324 7896 10376 7948
rect 15016 7964 15068 8016
rect 17040 7964 17092 8016
rect 7288 7803 7340 7812
rect 7288 7769 7297 7803
rect 7297 7769 7331 7803
rect 7331 7769 7340 7803
rect 7288 7760 7340 7769
rect 6552 7692 6604 7744
rect 8944 7692 8996 7744
rect 9312 7735 9364 7744
rect 9312 7701 9321 7735
rect 9321 7701 9355 7735
rect 9355 7701 9364 7735
rect 9312 7692 9364 7701
rect 9496 7735 9548 7744
rect 9496 7701 9505 7735
rect 9505 7701 9539 7735
rect 9539 7701 9548 7735
rect 9496 7692 9548 7701
rect 11612 7828 11664 7880
rect 11704 7871 11756 7880
rect 11704 7837 11713 7871
rect 11713 7837 11747 7871
rect 11747 7837 11756 7871
rect 11704 7828 11756 7837
rect 12900 7896 12952 7948
rect 11980 7871 12032 7880
rect 11980 7837 11989 7871
rect 11989 7837 12023 7871
rect 12023 7837 12032 7871
rect 11980 7828 12032 7837
rect 10140 7803 10192 7812
rect 10140 7769 10149 7803
rect 10149 7769 10183 7803
rect 10183 7769 10192 7803
rect 10140 7760 10192 7769
rect 12164 7871 12216 7880
rect 12164 7837 12173 7871
rect 12173 7837 12207 7871
rect 12207 7837 12216 7871
rect 12164 7828 12216 7837
rect 13544 7828 13596 7880
rect 12348 7760 12400 7812
rect 10876 7692 10928 7744
rect 11704 7692 11756 7744
rect 14832 7828 14884 7880
rect 15200 7828 15252 7880
rect 15476 7871 15528 7880
rect 15476 7837 15485 7871
rect 15485 7837 15519 7871
rect 15519 7837 15528 7871
rect 15476 7828 15528 7837
rect 16580 7896 16632 7948
rect 15844 7828 15896 7880
rect 16212 7828 16264 7880
rect 16304 7828 16356 7880
rect 16488 7871 16540 7880
rect 16488 7837 16497 7871
rect 16497 7837 16531 7871
rect 16531 7837 16540 7871
rect 16488 7828 16540 7837
rect 16856 7828 16908 7880
rect 17132 7828 17184 7880
rect 17960 8075 18012 8084
rect 17960 8041 17969 8075
rect 17969 8041 18003 8075
rect 18003 8041 18012 8075
rect 17960 8032 18012 8041
rect 18236 8032 18288 8084
rect 18696 8075 18748 8084
rect 18696 8041 18705 8075
rect 18705 8041 18739 8075
rect 18739 8041 18748 8075
rect 18696 8032 18748 8041
rect 17868 7828 17920 7880
rect 18236 7939 18288 7948
rect 18236 7905 18245 7939
rect 18245 7905 18279 7939
rect 18279 7905 18288 7939
rect 18236 7896 18288 7905
rect 15292 7803 15344 7812
rect 15292 7769 15301 7803
rect 15301 7769 15335 7803
rect 15335 7769 15344 7803
rect 15292 7760 15344 7769
rect 14096 7692 14148 7744
rect 15568 7760 15620 7812
rect 16304 7735 16356 7744
rect 16304 7701 16313 7735
rect 16313 7701 16347 7735
rect 16347 7701 16356 7735
rect 16304 7692 16356 7701
rect 17960 7760 18012 7812
rect 18512 7871 18564 7880
rect 18512 7837 18521 7871
rect 18521 7837 18555 7871
rect 18555 7837 18564 7871
rect 18512 7828 18564 7837
rect 20168 7964 20220 8016
rect 20536 8032 20588 8084
rect 21824 8032 21876 8084
rect 18696 7760 18748 7812
rect 20444 7828 20496 7880
rect 20536 7828 20588 7880
rect 22744 7964 22796 8016
rect 23848 8032 23900 8084
rect 24584 8032 24636 8084
rect 27988 8032 28040 8084
rect 28816 8032 28868 8084
rect 29736 8032 29788 8084
rect 30564 8075 30616 8084
rect 30564 8041 30573 8075
rect 30573 8041 30607 8075
rect 30607 8041 30616 8075
rect 30564 8032 30616 8041
rect 30932 8032 30984 8084
rect 23388 7964 23440 8016
rect 27252 7964 27304 8016
rect 21364 7896 21416 7948
rect 23112 7896 23164 7948
rect 21088 7828 21140 7880
rect 24952 7871 25004 7880
rect 24952 7837 24961 7871
rect 24961 7837 24995 7871
rect 24995 7837 25004 7871
rect 24952 7828 25004 7837
rect 25780 7896 25832 7948
rect 28908 7896 28960 7948
rect 25412 7828 25464 7880
rect 27804 7871 27856 7880
rect 27804 7837 27813 7871
rect 27813 7837 27847 7871
rect 27847 7837 27856 7871
rect 27804 7828 27856 7837
rect 20904 7760 20956 7812
rect 21916 7760 21968 7812
rect 22468 7760 22520 7812
rect 18420 7692 18472 7744
rect 19064 7692 19116 7744
rect 21272 7692 21324 7744
rect 29644 7828 29696 7880
rect 30012 7871 30064 7880
rect 30012 7837 30021 7871
rect 30021 7837 30055 7871
rect 30055 7837 30064 7871
rect 30012 7828 30064 7837
rect 30840 7896 30892 7948
rect 30472 7871 30524 7880
rect 30472 7837 30481 7871
rect 30481 7837 30515 7871
rect 30515 7837 30524 7871
rect 30472 7828 30524 7837
rect 31852 7828 31904 7880
rect 31668 7760 31720 7812
rect 33232 7760 33284 7812
rect 26148 7692 26200 7744
rect 27804 7692 27856 7744
rect 27896 7692 27948 7744
rect 29736 7692 29788 7744
rect 32312 7735 32364 7744
rect 32312 7701 32321 7735
rect 32321 7701 32355 7735
rect 32355 7701 32364 7735
rect 32312 7692 32364 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 7196 7488 7248 7540
rect 7288 7488 7340 7540
rect 8668 7488 8720 7540
rect 9312 7488 9364 7540
rect 9496 7488 9548 7540
rect 10324 7488 10376 7540
rect 6552 7420 6604 7472
rect 10968 7420 11020 7472
rect 6644 7216 6696 7268
rect 8300 7284 8352 7336
rect 11704 7488 11756 7540
rect 12164 7488 12216 7540
rect 12532 7488 12584 7540
rect 11796 7463 11848 7472
rect 11796 7429 11805 7463
rect 11805 7429 11839 7463
rect 11839 7429 11848 7463
rect 11796 7420 11848 7429
rect 12624 7420 12676 7472
rect 16488 7488 16540 7540
rect 16580 7488 16632 7540
rect 17316 7488 17368 7540
rect 16764 7420 16816 7472
rect 10140 7284 10192 7336
rect 10876 7327 10928 7336
rect 10876 7293 10885 7327
rect 10885 7293 10919 7327
rect 10919 7293 10928 7327
rect 15384 7395 15436 7404
rect 15384 7361 15393 7395
rect 15393 7361 15427 7395
rect 15427 7361 15436 7395
rect 15384 7352 15436 7361
rect 15476 7395 15528 7404
rect 15476 7361 15486 7395
rect 15486 7361 15520 7395
rect 15520 7361 15528 7395
rect 15476 7352 15528 7361
rect 15660 7395 15712 7404
rect 15660 7361 15669 7395
rect 15669 7361 15703 7395
rect 15703 7361 15712 7395
rect 15660 7352 15712 7361
rect 10876 7284 10928 7293
rect 5908 7191 5960 7200
rect 5908 7157 5917 7191
rect 5917 7157 5951 7191
rect 5951 7157 5960 7191
rect 5908 7148 5960 7157
rect 12808 7284 12860 7336
rect 14832 7284 14884 7336
rect 15200 7284 15252 7336
rect 16028 7352 16080 7404
rect 11980 7216 12032 7268
rect 12348 7216 12400 7268
rect 14740 7216 14792 7268
rect 15292 7216 15344 7268
rect 14096 7148 14148 7200
rect 16396 7352 16448 7404
rect 17040 7395 17092 7404
rect 17040 7361 17049 7395
rect 17049 7361 17083 7395
rect 17083 7361 17092 7395
rect 17040 7352 17092 7361
rect 17132 7352 17184 7404
rect 17224 7395 17276 7404
rect 17224 7361 17233 7395
rect 17233 7361 17267 7395
rect 17267 7361 17276 7395
rect 17224 7352 17276 7361
rect 18512 7488 18564 7540
rect 19800 7488 19852 7540
rect 19984 7488 20036 7540
rect 20536 7488 20588 7540
rect 21180 7488 21232 7540
rect 22376 7531 22428 7540
rect 22376 7497 22385 7531
rect 22385 7497 22419 7531
rect 22419 7497 22428 7531
rect 22376 7488 22428 7497
rect 22560 7488 22612 7540
rect 23020 7488 23072 7540
rect 23204 7488 23256 7540
rect 24952 7488 25004 7540
rect 25412 7488 25464 7540
rect 26332 7488 26384 7540
rect 28724 7488 28776 7540
rect 30012 7488 30064 7540
rect 30472 7488 30524 7540
rect 31392 7488 31444 7540
rect 31576 7531 31628 7540
rect 31576 7497 31585 7531
rect 31585 7497 31619 7531
rect 31619 7497 31628 7531
rect 31576 7488 31628 7497
rect 32312 7488 32364 7540
rect 17500 7352 17552 7404
rect 17684 7395 17736 7404
rect 17684 7361 17693 7395
rect 17693 7361 17727 7395
rect 17727 7361 17736 7395
rect 17684 7352 17736 7361
rect 17776 7395 17828 7404
rect 17776 7361 17786 7395
rect 17786 7361 17820 7395
rect 17820 7361 17828 7395
rect 17776 7352 17828 7361
rect 17868 7352 17920 7404
rect 18420 7395 18472 7404
rect 18420 7361 18449 7395
rect 18449 7361 18472 7395
rect 19156 7420 19208 7472
rect 20720 7420 20772 7472
rect 18420 7352 18472 7361
rect 16580 7216 16632 7268
rect 18972 7352 19024 7404
rect 19892 7352 19944 7404
rect 20536 7352 20588 7404
rect 19432 7284 19484 7336
rect 21272 7395 21324 7404
rect 21272 7361 21281 7395
rect 21281 7361 21315 7395
rect 21315 7361 21324 7395
rect 21272 7352 21324 7361
rect 21456 7352 21508 7404
rect 21824 7395 21876 7404
rect 21824 7361 21833 7395
rect 21833 7361 21867 7395
rect 21867 7361 21876 7395
rect 21824 7352 21876 7361
rect 21916 7352 21968 7404
rect 22192 7395 22244 7404
rect 22192 7361 22201 7395
rect 22201 7361 22235 7395
rect 22235 7361 22244 7395
rect 22192 7352 22244 7361
rect 22468 7352 22520 7404
rect 22284 7284 22336 7336
rect 23020 7395 23072 7404
rect 23020 7361 23029 7395
rect 23029 7361 23063 7395
rect 23063 7361 23072 7395
rect 23020 7352 23072 7361
rect 23112 7395 23164 7404
rect 23112 7361 23121 7395
rect 23121 7361 23155 7395
rect 23155 7361 23164 7395
rect 23112 7352 23164 7361
rect 24216 7352 24268 7404
rect 24676 7352 24728 7404
rect 25504 7395 25556 7404
rect 25504 7361 25508 7395
rect 25508 7361 25542 7395
rect 25542 7361 25556 7395
rect 25504 7352 25556 7361
rect 25596 7395 25648 7404
rect 25596 7361 25605 7395
rect 25605 7361 25639 7395
rect 25639 7361 25648 7395
rect 25596 7352 25648 7361
rect 25872 7395 25924 7404
rect 25872 7361 25880 7395
rect 25880 7361 25914 7395
rect 25914 7361 25924 7395
rect 25872 7352 25924 7361
rect 26056 7395 26108 7404
rect 26056 7361 26065 7395
rect 26065 7361 26099 7395
rect 26099 7361 26108 7395
rect 26056 7352 26108 7361
rect 29000 7463 29052 7472
rect 29000 7429 29009 7463
rect 29009 7429 29043 7463
rect 29043 7429 29052 7463
rect 29000 7420 29052 7429
rect 26516 7352 26568 7404
rect 26608 7352 26660 7404
rect 29920 7420 29972 7472
rect 19616 7216 19668 7268
rect 20076 7216 20128 7268
rect 18420 7148 18472 7200
rect 18972 7191 19024 7200
rect 18972 7157 18981 7191
rect 18981 7157 19015 7191
rect 19015 7157 19024 7191
rect 18972 7148 19024 7157
rect 19064 7148 19116 7200
rect 20260 7148 20312 7200
rect 20352 7148 20404 7200
rect 21088 7148 21140 7200
rect 22192 7148 22244 7200
rect 24308 7148 24360 7200
rect 24676 7191 24728 7200
rect 24676 7157 24685 7191
rect 24685 7157 24719 7191
rect 24719 7157 24728 7191
rect 24676 7148 24728 7157
rect 29552 7352 29604 7404
rect 29828 7395 29880 7404
rect 29828 7361 29838 7395
rect 29838 7361 29872 7395
rect 29872 7361 29880 7395
rect 32036 7420 32088 7472
rect 29828 7352 29880 7361
rect 30104 7395 30156 7404
rect 30104 7361 30113 7395
rect 30113 7361 30147 7395
rect 30147 7361 30156 7395
rect 30104 7352 30156 7361
rect 29644 7284 29696 7336
rect 31668 7352 31720 7404
rect 33692 7420 33744 7472
rect 25964 7216 26016 7268
rect 26148 7216 26200 7268
rect 28632 7216 28684 7268
rect 29092 7216 29144 7268
rect 29828 7216 29880 7268
rect 26240 7148 26292 7200
rect 27896 7148 27948 7200
rect 30104 7148 30156 7200
rect 31944 7191 31996 7200
rect 31944 7157 31953 7191
rect 31953 7157 31987 7191
rect 31987 7157 31996 7191
rect 31944 7148 31996 7157
rect 32404 7327 32456 7336
rect 32404 7293 32413 7327
rect 32413 7293 32447 7327
rect 32447 7293 32456 7327
rect 32404 7284 32456 7293
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 5908 6944 5960 6996
rect 7196 6987 7248 6996
rect 7196 6953 7205 6987
rect 7205 6953 7239 6987
rect 7239 6953 7248 6987
rect 7196 6944 7248 6953
rect 14740 6944 14792 6996
rect 14096 6851 14148 6860
rect 14096 6817 14105 6851
rect 14105 6817 14139 6851
rect 14139 6817 14148 6851
rect 16580 6876 16632 6928
rect 17776 6876 17828 6928
rect 18236 6944 18288 6996
rect 18696 6944 18748 6996
rect 20536 6944 20588 6996
rect 18420 6919 18472 6928
rect 18420 6885 18429 6919
rect 18429 6885 18463 6919
rect 18463 6885 18472 6919
rect 18420 6876 18472 6885
rect 21548 6876 21600 6928
rect 21640 6876 21692 6928
rect 22284 6944 22336 6996
rect 22836 6944 22888 6996
rect 14096 6808 14148 6817
rect 7748 6740 7800 6792
rect 7932 6740 7984 6792
rect 8944 6740 8996 6792
rect 6000 6672 6052 6724
rect 14188 6783 14240 6792
rect 14188 6749 14197 6783
rect 14197 6749 14231 6783
rect 14231 6749 14240 6783
rect 14188 6740 14240 6749
rect 14372 6783 14424 6792
rect 14372 6749 14381 6783
rect 14381 6749 14415 6783
rect 14415 6749 14424 6783
rect 14372 6740 14424 6749
rect 15476 6808 15528 6860
rect 15108 6783 15160 6792
rect 15108 6749 15122 6783
rect 15122 6749 15156 6783
rect 15156 6749 15160 6783
rect 15108 6740 15160 6749
rect 15660 6740 15712 6792
rect 18236 6808 18288 6860
rect 17592 6740 17644 6792
rect 18052 6740 18104 6792
rect 18328 6783 18380 6792
rect 18328 6749 18337 6783
rect 18337 6749 18371 6783
rect 18371 6749 18380 6783
rect 18328 6740 18380 6749
rect 18972 6808 19024 6860
rect 20260 6851 20312 6860
rect 20260 6817 20269 6851
rect 20269 6817 20303 6851
rect 20303 6817 20312 6851
rect 20260 6808 20312 6817
rect 21088 6808 21140 6860
rect 18696 6740 18748 6792
rect 20076 6783 20128 6792
rect 20076 6749 20085 6783
rect 20085 6749 20119 6783
rect 20119 6749 20128 6783
rect 20076 6740 20128 6749
rect 14832 6672 14884 6724
rect 17960 6672 18012 6724
rect 20628 6672 20680 6724
rect 20904 6672 20956 6724
rect 23296 6808 23348 6860
rect 22008 6740 22060 6792
rect 22192 6740 22244 6792
rect 22928 6740 22980 6792
rect 23020 6740 23072 6792
rect 26056 6944 26108 6996
rect 23572 6783 23624 6792
rect 23572 6749 23580 6783
rect 23580 6749 23614 6783
rect 23614 6749 23624 6783
rect 23572 6740 23624 6749
rect 23664 6783 23716 6792
rect 23664 6749 23673 6783
rect 23673 6749 23707 6783
rect 23707 6749 23716 6783
rect 23664 6740 23716 6749
rect 25688 6876 25740 6928
rect 26148 6876 26200 6928
rect 25228 6808 25280 6860
rect 22560 6715 22612 6724
rect 22560 6681 22569 6715
rect 22569 6681 22603 6715
rect 22603 6681 22612 6715
rect 22560 6672 22612 6681
rect 23296 6715 23348 6724
rect 23296 6681 23305 6715
rect 23305 6681 23339 6715
rect 23339 6681 23348 6715
rect 23296 6672 23348 6681
rect 24860 6672 24912 6724
rect 11796 6647 11848 6656
rect 11796 6613 11805 6647
rect 11805 6613 11839 6647
rect 11839 6613 11848 6647
rect 11796 6604 11848 6613
rect 12348 6604 12400 6656
rect 12532 6604 12584 6656
rect 14556 6604 14608 6656
rect 15752 6604 15804 6656
rect 16856 6604 16908 6656
rect 19800 6604 19852 6656
rect 21640 6604 21692 6656
rect 22192 6647 22244 6656
rect 22192 6613 22201 6647
rect 22201 6613 22235 6647
rect 22235 6613 22244 6647
rect 22192 6604 22244 6613
rect 22284 6604 22336 6656
rect 23020 6647 23072 6656
rect 23020 6613 23029 6647
rect 23029 6613 23063 6647
rect 23063 6613 23072 6647
rect 23020 6604 23072 6613
rect 23112 6604 23164 6656
rect 23940 6604 23992 6656
rect 25044 6647 25096 6656
rect 25044 6613 25053 6647
rect 25053 6613 25087 6647
rect 25087 6613 25096 6647
rect 25044 6604 25096 6613
rect 25780 6740 25832 6792
rect 26148 6783 26200 6792
rect 26148 6749 26157 6783
rect 26157 6749 26191 6783
rect 26191 6749 26200 6783
rect 26148 6740 26200 6749
rect 26240 6783 26292 6792
rect 26240 6749 26249 6783
rect 26249 6749 26283 6783
rect 26283 6749 26292 6783
rect 26240 6740 26292 6749
rect 26424 6783 26476 6792
rect 26424 6749 26432 6783
rect 26432 6749 26466 6783
rect 26466 6749 26476 6783
rect 26424 6740 26476 6749
rect 26516 6783 26568 6792
rect 26516 6749 26525 6783
rect 26525 6749 26559 6783
rect 26559 6749 26568 6783
rect 26516 6740 26568 6749
rect 27252 6783 27304 6792
rect 27252 6749 27261 6783
rect 27261 6749 27295 6783
rect 27295 6749 27304 6783
rect 27252 6740 27304 6749
rect 25412 6715 25464 6724
rect 25412 6681 25421 6715
rect 25421 6681 25455 6715
rect 25455 6681 25464 6715
rect 25412 6672 25464 6681
rect 25504 6715 25556 6724
rect 25504 6681 25513 6715
rect 25513 6681 25547 6715
rect 25547 6681 25556 6715
rect 25504 6672 25556 6681
rect 25596 6672 25648 6724
rect 26608 6672 26660 6724
rect 25320 6604 25372 6656
rect 26792 6604 26844 6656
rect 27160 6647 27212 6656
rect 27160 6613 27169 6647
rect 27169 6613 27203 6647
rect 27203 6613 27212 6647
rect 27160 6604 27212 6613
rect 28540 6944 28592 6996
rect 32404 6944 32456 6996
rect 28356 6876 28408 6928
rect 28724 6876 28776 6928
rect 29828 6876 29880 6928
rect 28080 6740 28132 6792
rect 28172 6740 28224 6792
rect 28724 6783 28776 6792
rect 28724 6749 28733 6783
rect 28733 6749 28767 6783
rect 28767 6749 28776 6783
rect 28724 6740 28776 6749
rect 29184 6740 29236 6792
rect 31944 6740 31996 6792
rect 27988 6604 28040 6656
rect 28080 6604 28132 6656
rect 30472 6672 30524 6724
rect 29552 6647 29604 6656
rect 29552 6613 29561 6647
rect 29561 6613 29595 6647
rect 29595 6613 29604 6647
rect 29552 6604 29604 6613
rect 29828 6604 29880 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 6000 6400 6052 6452
rect 11796 6400 11848 6452
rect 14096 6400 14148 6452
rect 14280 6400 14332 6452
rect 15568 6400 15620 6452
rect 16948 6400 17000 6452
rect 17408 6400 17460 6452
rect 17776 6400 17828 6452
rect 18328 6400 18380 6452
rect 20076 6400 20128 6452
rect 6736 6264 6788 6316
rect 8944 6307 8996 6316
rect 8944 6273 8953 6307
rect 8953 6273 8987 6307
rect 8987 6273 8996 6307
rect 8944 6264 8996 6273
rect 13636 6332 13688 6384
rect 13912 6375 13964 6384
rect 13912 6341 13921 6375
rect 13921 6341 13955 6375
rect 13955 6341 13964 6375
rect 13912 6332 13964 6341
rect 21456 6375 21508 6384
rect 21456 6341 21465 6375
rect 21465 6341 21499 6375
rect 21499 6341 21508 6375
rect 21456 6332 21508 6341
rect 22100 6400 22152 6452
rect 22192 6400 22244 6452
rect 22284 6400 22336 6452
rect 22376 6400 22428 6452
rect 13544 6264 13596 6316
rect 5448 6128 5500 6180
rect 11336 6128 11388 6180
rect 8668 6060 8720 6112
rect 10324 6060 10376 6112
rect 11888 6239 11940 6248
rect 11888 6205 11897 6239
rect 11897 6205 11931 6239
rect 11931 6205 11940 6239
rect 11888 6196 11940 6205
rect 14004 6239 14056 6248
rect 14004 6205 14013 6239
rect 14013 6205 14047 6239
rect 14047 6205 14056 6239
rect 14004 6196 14056 6205
rect 16672 6264 16724 6316
rect 17408 6264 17460 6316
rect 13820 6128 13872 6180
rect 17040 6196 17092 6248
rect 17592 6264 17644 6316
rect 17776 6307 17828 6316
rect 17776 6273 17785 6307
rect 17785 6273 17819 6307
rect 17819 6273 17828 6307
rect 17776 6264 17828 6273
rect 18052 6264 18104 6316
rect 18144 6196 18196 6248
rect 15476 6128 15528 6180
rect 16948 6128 17000 6180
rect 17960 6128 18012 6180
rect 21364 6307 21416 6316
rect 21364 6273 21373 6307
rect 21373 6273 21407 6307
rect 21407 6273 21416 6307
rect 21364 6264 21416 6273
rect 21916 6307 21968 6316
rect 21916 6273 21925 6307
rect 21925 6273 21959 6307
rect 21959 6273 21968 6307
rect 21916 6264 21968 6273
rect 22008 6264 22060 6316
rect 23020 6400 23072 6452
rect 23480 6443 23532 6452
rect 23480 6409 23489 6443
rect 23489 6409 23523 6443
rect 23523 6409 23532 6443
rect 23480 6400 23532 6409
rect 23848 6400 23900 6452
rect 24492 6443 24544 6452
rect 24492 6409 24501 6443
rect 24501 6409 24535 6443
rect 24535 6409 24544 6443
rect 24492 6400 24544 6409
rect 24860 6443 24912 6452
rect 24860 6409 24869 6443
rect 24869 6409 24903 6443
rect 24903 6409 24912 6443
rect 24860 6400 24912 6409
rect 25596 6400 25648 6452
rect 26424 6400 26476 6452
rect 27896 6400 27948 6452
rect 28724 6400 28776 6452
rect 29828 6400 29880 6452
rect 13452 6103 13504 6112
rect 13452 6069 13461 6103
rect 13461 6069 13495 6103
rect 13495 6069 13504 6103
rect 13452 6060 13504 6069
rect 14740 6060 14792 6112
rect 21548 6196 21600 6248
rect 23204 6307 23256 6316
rect 23204 6273 23213 6307
rect 23213 6273 23247 6307
rect 23247 6273 23256 6307
rect 23204 6264 23256 6273
rect 24308 6332 24360 6384
rect 26884 6332 26936 6384
rect 27160 6332 27212 6384
rect 24584 6307 24636 6316
rect 24584 6273 24593 6307
rect 24593 6273 24627 6307
rect 24627 6273 24636 6307
rect 24584 6264 24636 6273
rect 22836 6196 22888 6248
rect 25596 6307 25648 6316
rect 25596 6273 25605 6307
rect 25605 6273 25639 6307
rect 25639 6273 25648 6307
rect 25596 6264 25648 6273
rect 25872 6307 25924 6316
rect 25872 6273 25881 6307
rect 25881 6273 25915 6307
rect 25915 6273 25924 6307
rect 25872 6264 25924 6273
rect 25964 6307 26016 6316
rect 25964 6273 25973 6307
rect 25973 6273 26007 6307
rect 26007 6273 26016 6307
rect 25964 6264 26016 6273
rect 26148 6264 26200 6316
rect 26700 6196 26752 6248
rect 27252 6264 27304 6316
rect 27896 6307 27948 6316
rect 27896 6273 27905 6307
rect 27905 6273 27939 6307
rect 27939 6273 27948 6307
rect 27896 6264 27948 6273
rect 30196 6307 30248 6316
rect 30196 6273 30205 6307
rect 30205 6273 30239 6307
rect 30239 6273 30248 6307
rect 30196 6264 30248 6273
rect 28080 6196 28132 6248
rect 22284 6128 22336 6180
rect 26332 6128 26384 6180
rect 26792 6128 26844 6180
rect 27068 6128 27120 6180
rect 24952 6060 25004 6112
rect 25320 6060 25372 6112
rect 30012 6103 30064 6112
rect 30012 6069 30021 6103
rect 30021 6069 30055 6103
rect 30055 6069 30064 6103
rect 30012 6060 30064 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 10324 5856 10376 5908
rect 11888 5856 11940 5908
rect 14648 5856 14700 5908
rect 5724 5720 5776 5772
rect 8576 5720 8628 5772
rect 9128 5720 9180 5772
rect 5448 5652 5500 5704
rect 9772 5763 9824 5772
rect 9772 5729 9781 5763
rect 9781 5729 9815 5763
rect 9815 5729 9824 5763
rect 9772 5720 9824 5729
rect 9956 5763 10008 5772
rect 9956 5729 9965 5763
rect 9965 5729 9999 5763
rect 9999 5729 10008 5763
rect 9956 5720 10008 5729
rect 10600 5720 10652 5772
rect 11520 5720 11572 5772
rect 12256 5763 12308 5772
rect 12256 5729 12265 5763
rect 12265 5729 12299 5763
rect 12299 5729 12308 5763
rect 12256 5720 12308 5729
rect 6736 5584 6788 5636
rect 7012 5627 7064 5636
rect 7012 5593 7021 5627
rect 7021 5593 7055 5627
rect 7055 5593 7064 5627
rect 7012 5584 7064 5593
rect 7748 5584 7800 5636
rect 4160 5516 4212 5568
rect 8024 5516 8076 5568
rect 14832 5788 14884 5840
rect 13452 5720 13504 5772
rect 14924 5720 14976 5772
rect 23664 5856 23716 5908
rect 24952 5856 25004 5908
rect 31484 5856 31536 5908
rect 17408 5788 17460 5840
rect 17868 5788 17920 5840
rect 18512 5788 18564 5840
rect 23388 5788 23440 5840
rect 26424 5788 26476 5840
rect 15568 5763 15620 5772
rect 15568 5729 15577 5763
rect 15577 5729 15611 5763
rect 15611 5729 15620 5763
rect 15568 5720 15620 5729
rect 22560 5720 22612 5772
rect 25136 5720 25188 5772
rect 30012 5720 30064 5772
rect 12624 5652 12676 5704
rect 13912 5652 13964 5704
rect 10232 5584 10284 5636
rect 10600 5584 10652 5636
rect 15660 5652 15712 5704
rect 17408 5652 17460 5704
rect 17592 5695 17644 5704
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 19432 5695 19484 5704
rect 19432 5661 19441 5695
rect 19441 5661 19475 5695
rect 19475 5661 19484 5695
rect 19432 5652 19484 5661
rect 9036 5559 9088 5568
rect 9036 5525 9045 5559
rect 9045 5525 9079 5559
rect 9079 5525 9088 5559
rect 9036 5516 9088 5525
rect 12808 5516 12860 5568
rect 14096 5559 14148 5568
rect 14096 5525 14105 5559
rect 14105 5525 14139 5559
rect 14139 5525 14148 5559
rect 14096 5516 14148 5525
rect 14556 5559 14608 5568
rect 14556 5525 14565 5559
rect 14565 5525 14599 5559
rect 14599 5525 14608 5559
rect 14556 5516 14608 5525
rect 15200 5516 15252 5568
rect 16948 5584 17000 5636
rect 17040 5584 17092 5636
rect 21456 5652 21508 5704
rect 29644 5695 29696 5704
rect 29644 5661 29653 5695
rect 29653 5661 29687 5695
rect 29687 5661 29696 5695
rect 29644 5652 29696 5661
rect 31024 5652 31076 5704
rect 31484 5695 31536 5704
rect 31484 5661 31493 5695
rect 31493 5661 31527 5695
rect 31527 5661 31536 5695
rect 31484 5652 31536 5661
rect 22008 5584 22060 5636
rect 24584 5584 24636 5636
rect 31760 5627 31812 5636
rect 31760 5593 31769 5627
rect 31769 5593 31803 5627
rect 31803 5593 31812 5627
rect 31760 5584 31812 5593
rect 32036 5584 32088 5636
rect 17776 5559 17828 5568
rect 17776 5525 17785 5559
rect 17785 5525 17819 5559
rect 17819 5525 17828 5559
rect 17776 5516 17828 5525
rect 19248 5559 19300 5568
rect 19248 5525 19257 5559
rect 19257 5525 19291 5559
rect 19291 5525 19300 5559
rect 19248 5516 19300 5525
rect 19616 5559 19668 5568
rect 19616 5525 19625 5559
rect 19625 5525 19659 5559
rect 19659 5525 19668 5559
rect 19616 5516 19668 5525
rect 21364 5516 21416 5568
rect 24492 5516 24544 5568
rect 31392 5559 31444 5568
rect 31392 5525 31401 5559
rect 31401 5525 31435 5559
rect 31435 5525 31444 5559
rect 31392 5516 31444 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 18880 5312 18932 5364
rect 19616 5312 19668 5364
rect 22560 5312 22612 5364
rect 27344 5312 27396 5364
rect 28080 5312 28132 5364
rect 29644 5312 29696 5364
rect 30196 5312 30248 5364
rect 30472 5312 30524 5364
rect 31392 5312 31444 5364
rect 31484 5312 31536 5364
rect 32036 5312 32088 5364
rect 8576 5244 8628 5296
rect 9036 5244 9088 5296
rect 10232 5244 10284 5296
rect 11060 5244 11112 5296
rect 4160 5176 4212 5228
rect 6920 5108 6972 5160
rect 7012 5040 7064 5092
rect 8024 5108 8076 5160
rect 8300 5108 8352 5160
rect 8668 5151 8720 5160
rect 8668 5117 8677 5151
rect 8677 5117 8711 5151
rect 8711 5117 8720 5151
rect 8668 5108 8720 5117
rect 10600 5108 10652 5160
rect 11428 5108 11480 5160
rect 1768 5015 1820 5024
rect 1768 4981 1777 5015
rect 1777 4981 1811 5015
rect 1811 4981 1820 5015
rect 1768 4972 1820 4981
rect 12256 5244 12308 5296
rect 11888 5219 11940 5228
rect 11888 5185 11897 5219
rect 11897 5185 11931 5219
rect 11931 5185 11940 5219
rect 13176 5244 13228 5296
rect 13544 5244 13596 5296
rect 11888 5176 11940 5185
rect 12624 5108 12676 5160
rect 12808 5151 12860 5160
rect 12808 5117 12817 5151
rect 12817 5117 12851 5151
rect 12851 5117 12860 5151
rect 12808 5108 12860 5117
rect 13084 5151 13136 5160
rect 13084 5117 13093 5151
rect 13093 5117 13127 5151
rect 13127 5117 13136 5151
rect 13084 5108 13136 5117
rect 14556 5151 14608 5160
rect 14556 5117 14565 5151
rect 14565 5117 14599 5151
rect 14599 5117 14608 5151
rect 14556 5108 14608 5117
rect 14740 5151 14792 5160
rect 14740 5117 14749 5151
rect 14749 5117 14783 5151
rect 14783 5117 14792 5151
rect 14740 5108 14792 5117
rect 15016 5151 15068 5160
rect 15016 5117 15025 5151
rect 15025 5117 15059 5151
rect 15059 5117 15068 5151
rect 15016 5108 15068 5117
rect 15660 5108 15712 5160
rect 11060 4972 11112 5024
rect 14832 4972 14884 5024
rect 17684 5176 17736 5228
rect 22192 5244 22244 5296
rect 23296 5244 23348 5296
rect 23388 5244 23440 5296
rect 22284 5219 22336 5228
rect 22284 5185 22293 5219
rect 22293 5185 22327 5219
rect 22327 5185 22336 5219
rect 22284 5176 22336 5185
rect 22836 5176 22888 5228
rect 23940 5176 23992 5228
rect 19248 5151 19300 5160
rect 19248 5117 19257 5151
rect 19257 5117 19291 5151
rect 19291 5117 19300 5151
rect 19248 5108 19300 5117
rect 22560 5151 22612 5160
rect 22560 5117 22569 5151
rect 22569 5117 22603 5151
rect 22603 5117 22612 5151
rect 22560 5108 22612 5117
rect 23664 5151 23716 5160
rect 23664 5117 23673 5151
rect 23673 5117 23707 5151
rect 23707 5117 23716 5151
rect 23664 5108 23716 5117
rect 26976 5219 27028 5228
rect 26976 5185 26985 5219
rect 26985 5185 27019 5219
rect 27019 5185 27028 5219
rect 26976 5176 27028 5185
rect 27252 5219 27304 5228
rect 27252 5185 27261 5219
rect 27261 5185 27295 5219
rect 27295 5185 27304 5219
rect 27252 5176 27304 5185
rect 26516 5108 26568 5160
rect 27620 5108 27672 5160
rect 27896 5176 27948 5228
rect 28264 5176 28316 5228
rect 30288 5176 30340 5228
rect 19892 4972 19944 5024
rect 20720 5015 20772 5024
rect 20720 4981 20729 5015
rect 20729 4981 20763 5015
rect 20763 4981 20772 5015
rect 20720 4972 20772 4981
rect 21916 5015 21968 5024
rect 21916 4981 21925 5015
rect 21925 4981 21959 5015
rect 21959 4981 21968 5015
rect 21916 4972 21968 4981
rect 22744 4972 22796 5024
rect 24768 5040 24820 5092
rect 27896 5040 27948 5092
rect 24216 5015 24268 5024
rect 24216 4981 24225 5015
rect 24225 4981 24259 5015
rect 24259 4981 24268 5015
rect 24216 4972 24268 4981
rect 27160 5015 27212 5024
rect 27160 4981 27169 5015
rect 27169 4981 27203 5015
rect 27203 4981 27212 5015
rect 27160 4972 27212 4981
rect 27528 4972 27580 5024
rect 27804 4972 27856 5024
rect 31760 5040 31812 5092
rect 31576 4972 31628 5024
rect 32680 5151 32732 5160
rect 32680 5117 32689 5151
rect 32689 5117 32723 5151
rect 32723 5117 32732 5151
rect 32680 5108 32732 5117
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 6276 4768 6328 4820
rect 9772 4768 9824 4820
rect 19340 4768 19392 4820
rect 22836 4811 22888 4820
rect 22836 4777 22845 4811
rect 22845 4777 22879 4811
rect 22879 4777 22888 4811
rect 22836 4768 22888 4777
rect 12624 4700 12676 4752
rect 13084 4700 13136 4752
rect 14096 4700 14148 4752
rect 15016 4743 15068 4752
rect 15016 4709 15025 4743
rect 15025 4709 15059 4743
rect 15059 4709 15068 4743
rect 15016 4700 15068 4709
rect 15200 4700 15252 4752
rect 17040 4700 17092 4752
rect 940 4496 992 4548
rect 19892 4675 19944 4684
rect 19892 4641 19901 4675
rect 19901 4641 19935 4675
rect 19935 4641 19944 4675
rect 19892 4632 19944 4641
rect 23388 4632 23440 4684
rect 19432 4564 19484 4616
rect 20168 4564 20220 4616
rect 20720 4564 20772 4616
rect 9036 4428 9088 4480
rect 9128 4471 9180 4480
rect 9128 4437 9137 4471
rect 9137 4437 9171 4471
rect 9171 4437 9180 4471
rect 9128 4428 9180 4437
rect 9956 4428 10008 4480
rect 15844 4428 15896 4480
rect 16672 4428 16724 4480
rect 19708 4471 19760 4480
rect 19708 4437 19717 4471
rect 19717 4437 19751 4471
rect 19751 4437 19760 4471
rect 19708 4428 19760 4437
rect 23572 4564 23624 4616
rect 24216 4768 24268 4820
rect 24308 4768 24360 4820
rect 27252 4768 27304 4820
rect 27344 4768 27396 4820
rect 29092 4700 29144 4752
rect 32680 4700 32732 4752
rect 26516 4675 26568 4684
rect 26516 4641 26525 4675
rect 26525 4641 26559 4675
rect 26559 4641 26568 4675
rect 26516 4632 26568 4641
rect 21364 4539 21416 4548
rect 21364 4505 21373 4539
rect 21373 4505 21407 4539
rect 21407 4505 21416 4539
rect 21364 4496 21416 4505
rect 22652 4496 22704 4548
rect 22744 4428 22796 4480
rect 22928 4471 22980 4480
rect 22928 4437 22937 4471
rect 22937 4437 22971 4471
rect 22971 4437 22980 4471
rect 22928 4428 22980 4437
rect 23296 4428 23348 4480
rect 25780 4564 25832 4616
rect 27068 4564 27120 4616
rect 27436 4607 27488 4616
rect 27436 4573 27445 4607
rect 27445 4573 27479 4607
rect 27479 4573 27488 4607
rect 27436 4564 27488 4573
rect 27620 4496 27672 4548
rect 26792 4471 26844 4480
rect 26792 4437 26801 4471
rect 26801 4437 26835 4471
rect 26835 4437 26844 4471
rect 26792 4428 26844 4437
rect 27160 4428 27212 4480
rect 28540 4428 28592 4480
rect 29460 4428 29512 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 11796 4224 11848 4276
rect 12716 4224 12768 4276
rect 16212 4224 16264 4276
rect 21364 4224 21416 4276
rect 22192 4224 22244 4276
rect 22652 4224 22704 4276
rect 23388 4224 23440 4276
rect 25780 4224 25832 4276
rect 26792 4224 26844 4276
rect 26976 4267 27028 4276
rect 26976 4233 26985 4267
rect 26985 4233 27019 4267
rect 27019 4233 27028 4267
rect 26976 4224 27028 4233
rect 27068 4224 27120 4276
rect 29736 4224 29788 4276
rect 11428 4156 11480 4208
rect 13452 4156 13504 4208
rect 16120 4156 16172 4208
rect 20996 4156 21048 4208
rect 25320 4156 25372 4208
rect 12348 4088 12400 4140
rect 12808 4088 12860 4140
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 19340 4088 19392 4140
rect 21548 4088 21600 4140
rect 21916 4088 21968 4140
rect 24768 4088 24820 4140
rect 29460 4156 29512 4208
rect 31024 4156 31076 4208
rect 11060 3952 11112 4004
rect 11980 3952 12032 4004
rect 14556 3952 14608 4004
rect 16672 4063 16724 4072
rect 16672 4029 16681 4063
rect 16681 4029 16715 4063
rect 16715 4029 16724 4063
rect 16672 4020 16724 4029
rect 12164 3927 12216 3936
rect 12164 3893 12173 3927
rect 12173 3893 12207 3927
rect 12207 3893 12216 3927
rect 12164 3884 12216 3893
rect 12256 3884 12308 3936
rect 14648 3884 14700 3936
rect 17500 3884 17552 3936
rect 20352 3952 20404 4004
rect 19800 3884 19852 3936
rect 27804 4063 27856 4072
rect 27804 4029 27813 4063
rect 27813 4029 27847 4063
rect 27847 4029 27856 4063
rect 27804 4020 27856 4029
rect 28080 4063 28132 4072
rect 28080 4029 28089 4063
rect 28089 4029 28123 4063
rect 28123 4029 28132 4063
rect 28080 4020 28132 4029
rect 29092 3884 29144 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 9772 3680 9824 3732
rect 12164 3680 12216 3732
rect 14556 3680 14608 3732
rect 12256 3544 12308 3596
rect 14372 3544 14424 3596
rect 6920 3519 6972 3528
rect 6920 3485 6929 3519
rect 6929 3485 6963 3519
rect 6963 3485 6972 3519
rect 6920 3476 6972 3485
rect 9036 3519 9088 3528
rect 9036 3485 9045 3519
rect 9045 3485 9079 3519
rect 9079 3485 9088 3519
rect 9036 3476 9088 3485
rect 11428 3476 11480 3528
rect 11612 3519 11664 3528
rect 11612 3485 11621 3519
rect 11621 3485 11655 3519
rect 11655 3485 11664 3519
rect 11612 3476 11664 3485
rect 11704 3519 11756 3528
rect 11704 3485 11713 3519
rect 11713 3485 11747 3519
rect 11747 3485 11756 3519
rect 11704 3476 11756 3485
rect 13452 3476 13504 3528
rect 14280 3519 14332 3528
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14280 3476 14332 3485
rect 14648 3519 14700 3528
rect 14648 3485 14657 3519
rect 14657 3485 14691 3519
rect 14691 3485 14700 3519
rect 14648 3476 14700 3485
rect 15844 3587 15896 3596
rect 15844 3553 15853 3587
rect 15853 3553 15887 3587
rect 15887 3553 15896 3587
rect 15844 3544 15896 3553
rect 16304 3680 16356 3732
rect 17960 3655 18012 3664
rect 17960 3621 17969 3655
rect 17969 3621 18003 3655
rect 18003 3621 18012 3655
rect 17960 3612 18012 3621
rect 18788 3587 18840 3596
rect 18788 3553 18797 3587
rect 18797 3553 18831 3587
rect 18831 3553 18840 3587
rect 18788 3544 18840 3553
rect 19800 3587 19852 3596
rect 19800 3553 19809 3587
rect 19809 3553 19843 3587
rect 19843 3553 19852 3587
rect 19800 3544 19852 3553
rect 9496 3408 9548 3460
rect 9588 3451 9640 3460
rect 9588 3417 9597 3451
rect 9597 3417 9631 3451
rect 9631 3417 9640 3451
rect 9588 3408 9640 3417
rect 11244 3408 11296 3460
rect 13912 3451 13964 3460
rect 13912 3417 13921 3451
rect 13921 3417 13955 3451
rect 13955 3417 13964 3451
rect 13912 3408 13964 3417
rect 18604 3519 18656 3528
rect 18604 3485 18613 3519
rect 18613 3485 18647 3519
rect 18647 3485 18656 3519
rect 18604 3476 18656 3485
rect 18880 3476 18932 3528
rect 20628 3476 20680 3528
rect 22928 3476 22980 3528
rect 24584 3587 24636 3596
rect 24584 3553 24593 3587
rect 24593 3553 24627 3587
rect 24627 3553 24636 3587
rect 24584 3544 24636 3553
rect 24768 3587 24820 3596
rect 24768 3553 24777 3587
rect 24777 3553 24811 3587
rect 24811 3553 24820 3587
rect 24768 3544 24820 3553
rect 25228 3544 25280 3596
rect 25320 3587 25372 3596
rect 25320 3553 25329 3587
rect 25329 3553 25363 3587
rect 25363 3553 25372 3587
rect 25320 3544 25372 3553
rect 29368 3680 29420 3732
rect 26332 3612 26384 3664
rect 26792 3544 26844 3596
rect 24676 3408 24728 3460
rect 27712 3476 27764 3528
rect 28264 3476 28316 3528
rect 31208 3544 31260 3596
rect 37464 3519 37516 3528
rect 37464 3485 37473 3519
rect 37473 3485 37507 3519
rect 37507 3485 37516 3519
rect 37464 3476 37516 3485
rect 9220 3340 9272 3392
rect 12348 3340 12400 3392
rect 12440 3340 12492 3392
rect 14648 3340 14700 3392
rect 14740 3383 14792 3392
rect 14740 3349 14749 3383
rect 14749 3349 14783 3383
rect 14783 3349 14792 3383
rect 14740 3340 14792 3349
rect 14924 3383 14976 3392
rect 14924 3349 14933 3383
rect 14933 3349 14967 3383
rect 14967 3349 14976 3383
rect 14924 3340 14976 3349
rect 15568 3383 15620 3392
rect 15568 3349 15577 3383
rect 15577 3349 15611 3383
rect 15611 3349 15620 3383
rect 15568 3340 15620 3349
rect 16304 3340 16356 3392
rect 16948 3383 17000 3392
rect 16948 3349 16957 3383
rect 16957 3349 16991 3383
rect 16991 3349 17000 3383
rect 16948 3340 17000 3349
rect 17500 3383 17552 3392
rect 17500 3349 17509 3383
rect 17509 3349 17543 3383
rect 17543 3349 17552 3383
rect 17500 3340 17552 3349
rect 17592 3383 17644 3392
rect 17592 3349 17601 3383
rect 17601 3349 17635 3383
rect 17635 3349 17644 3383
rect 17592 3340 17644 3349
rect 19708 3340 19760 3392
rect 20352 3340 20404 3392
rect 20904 3383 20956 3392
rect 20904 3349 20913 3383
rect 20913 3349 20947 3383
rect 20947 3349 20956 3383
rect 20904 3340 20956 3349
rect 22008 3383 22060 3392
rect 22008 3349 22017 3383
rect 22017 3349 22051 3383
rect 22051 3349 22060 3383
rect 22008 3340 22060 3349
rect 22192 3383 22244 3392
rect 22192 3349 22201 3383
rect 22201 3349 22235 3383
rect 22235 3349 22244 3383
rect 22192 3340 22244 3349
rect 24032 3383 24084 3392
rect 24032 3349 24041 3383
rect 24041 3349 24075 3383
rect 24075 3349 24084 3383
rect 24032 3340 24084 3349
rect 24860 3383 24912 3392
rect 24860 3349 24869 3383
rect 24869 3349 24903 3383
rect 24903 3349 24912 3383
rect 24860 3340 24912 3349
rect 25228 3383 25280 3392
rect 25228 3349 25237 3383
rect 25237 3349 25271 3383
rect 25271 3349 25280 3383
rect 25228 3340 25280 3349
rect 25688 3383 25740 3392
rect 25688 3349 25697 3383
rect 25697 3349 25731 3383
rect 25731 3349 25740 3383
rect 25688 3340 25740 3349
rect 26516 3340 26568 3392
rect 26700 3383 26752 3392
rect 26700 3349 26709 3383
rect 26709 3349 26743 3383
rect 26743 3349 26752 3383
rect 26700 3340 26752 3349
rect 27160 3383 27212 3392
rect 27160 3349 27169 3383
rect 27169 3349 27203 3383
rect 27203 3349 27212 3383
rect 27160 3340 27212 3349
rect 36912 3340 36964 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 9220 3136 9272 3188
rect 9496 3136 9548 3188
rect 1768 3111 1820 3120
rect 1768 3077 1777 3111
rect 1777 3077 1811 3111
rect 1811 3077 1820 3111
rect 1768 3068 1820 3077
rect 9588 3068 9640 3120
rect 1492 2839 1544 2848
rect 1492 2805 1501 2839
rect 1501 2805 1535 2839
rect 1535 2805 1544 2839
rect 1492 2796 1544 2805
rect 1952 2839 2004 2848
rect 1952 2805 1961 2839
rect 1961 2805 1995 2839
rect 1995 2805 2004 2839
rect 1952 2796 2004 2805
rect 6920 2796 6972 2848
rect 12440 3068 12492 3120
rect 14648 3136 14700 3188
rect 14740 3136 14792 3188
rect 14464 3111 14516 3120
rect 14464 3077 14473 3111
rect 14473 3077 14507 3111
rect 14507 3077 14516 3111
rect 14464 3068 14516 3077
rect 14924 3136 14976 3188
rect 16948 3136 17000 3188
rect 10968 2975 11020 2984
rect 10968 2941 10977 2975
rect 10977 2941 11011 2975
rect 11011 2941 11020 2975
rect 10968 2932 11020 2941
rect 11244 2932 11296 2984
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 11612 3043 11664 3052
rect 11612 3009 11621 3043
rect 11621 3009 11655 3043
rect 11655 3009 11664 3043
rect 11612 3000 11664 3009
rect 11796 3043 11848 3052
rect 11796 3009 11805 3043
rect 11805 3009 11839 3043
rect 11839 3009 11848 3043
rect 11796 3000 11848 3009
rect 11888 3000 11940 3052
rect 11980 2975 12032 2984
rect 11980 2941 11989 2975
rect 11989 2941 12023 2975
rect 12023 2941 12032 2975
rect 11980 2932 12032 2941
rect 13912 3000 13964 3052
rect 16120 3068 16172 3120
rect 17960 3136 18012 3188
rect 18236 3136 18288 3188
rect 19524 3136 19576 3188
rect 17684 3068 17736 3120
rect 20904 3136 20956 3188
rect 22008 3136 22060 3188
rect 22192 3136 22244 3188
rect 23572 3179 23624 3188
rect 23572 3145 23581 3179
rect 23581 3145 23615 3179
rect 23615 3145 23624 3179
rect 23572 3136 23624 3145
rect 24032 3136 24084 3188
rect 24860 3136 24912 3188
rect 20352 3068 20404 3120
rect 15568 2932 15620 2984
rect 12808 2864 12860 2916
rect 13912 2864 13964 2916
rect 12532 2796 12584 2848
rect 18236 2932 18288 2984
rect 18604 2932 18656 2984
rect 19340 2975 19392 2984
rect 19340 2941 19349 2975
rect 19349 2941 19383 2975
rect 19383 2941 19392 2975
rect 19340 2932 19392 2941
rect 18696 2864 18748 2916
rect 16304 2839 16356 2848
rect 16304 2805 16313 2839
rect 16313 2805 16347 2839
rect 16347 2805 16356 2839
rect 20628 2932 20680 2984
rect 23388 3068 23440 3120
rect 27344 3136 27396 3188
rect 25136 2932 25188 2984
rect 25688 3000 25740 3052
rect 26700 3000 26752 3052
rect 27160 3068 27212 3120
rect 28540 3068 28592 3120
rect 31024 3043 31076 3052
rect 31024 3009 31033 3043
rect 31033 3009 31067 3043
rect 31067 3009 31076 3043
rect 31024 3000 31076 3009
rect 25780 2932 25832 2984
rect 16304 2796 16356 2805
rect 19708 2839 19760 2848
rect 19708 2805 19717 2839
rect 19717 2805 19751 2839
rect 19751 2805 19760 2839
rect 19708 2796 19760 2805
rect 19800 2796 19852 2848
rect 26332 2864 26384 2916
rect 26516 2864 26568 2916
rect 32128 3000 32180 3052
rect 36912 3043 36964 3052
rect 36912 3009 36921 3043
rect 36921 3009 36955 3043
rect 36955 3009 36964 3043
rect 36912 3000 36964 3009
rect 26424 2796 26476 2848
rect 37280 2796 37332 2848
rect 37832 2839 37884 2848
rect 37832 2805 37841 2839
rect 37841 2805 37875 2839
rect 37875 2805 37884 2839
rect 37832 2796 37884 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 1952 2388 2004 2440
rect 9128 2592 9180 2644
rect 11612 2592 11664 2644
rect 11520 2524 11572 2576
rect 19800 2592 19852 2644
rect 25136 2635 25188 2644
rect 25136 2601 25145 2635
rect 25145 2601 25179 2635
rect 25179 2601 25188 2635
rect 25136 2592 25188 2601
rect 8944 2456 8996 2508
rect 6920 2431 6972 2440
rect 6920 2397 6929 2431
rect 6929 2397 6963 2431
rect 6963 2397 6972 2431
rect 6920 2388 6972 2397
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 13360 2456 13412 2508
rect 14372 2499 14424 2508
rect 14372 2465 14381 2499
rect 14381 2465 14415 2499
rect 14415 2465 14424 2499
rect 14372 2456 14424 2465
rect 12440 2431 12492 2440
rect 12440 2397 12449 2431
rect 12449 2397 12483 2431
rect 12483 2397 12492 2431
rect 12440 2388 12492 2397
rect 12532 2431 12584 2440
rect 12532 2397 12541 2431
rect 12541 2397 12575 2431
rect 12575 2397 12584 2431
rect 12532 2388 12584 2397
rect 12992 2431 13044 2440
rect 12992 2397 13001 2431
rect 13001 2397 13035 2431
rect 13035 2397 13044 2431
rect 12992 2388 13044 2397
rect 20 2320 72 2372
rect 2044 2363 2096 2372
rect 2044 2329 2053 2363
rect 2053 2329 2087 2363
rect 2087 2329 2096 2363
rect 2044 2320 2096 2329
rect 3976 2363 4028 2372
rect 3976 2329 3985 2363
rect 3985 2329 4019 2363
rect 4019 2329 4028 2363
rect 3976 2320 4028 2329
rect 6552 2363 6604 2372
rect 6552 2329 6561 2363
rect 6561 2329 6595 2363
rect 6595 2329 6604 2363
rect 6552 2320 6604 2329
rect 31024 2524 31076 2576
rect 14372 2320 14424 2372
rect 16212 2456 16264 2508
rect 19708 2456 19760 2508
rect 25228 2456 25280 2508
rect 31116 2456 31168 2508
rect 24676 2431 24728 2440
rect 24676 2397 24685 2431
rect 24685 2397 24719 2431
rect 24719 2397 24728 2431
rect 24676 2388 24728 2397
rect 26700 2388 26752 2440
rect 31024 2431 31076 2440
rect 31024 2397 31033 2431
rect 31033 2397 31067 2431
rect 31067 2397 31076 2431
rect 31024 2388 31076 2397
rect 35532 2431 35584 2440
rect 35532 2397 35541 2431
rect 35541 2397 35575 2431
rect 35575 2397 35584 2431
rect 35532 2388 35584 2397
rect 37280 2388 37332 2440
rect 15568 2363 15620 2372
rect 15568 2329 15577 2363
rect 15577 2329 15611 2363
rect 15611 2329 15620 2363
rect 15568 2320 15620 2329
rect 11152 2252 11204 2304
rect 20260 2295 20312 2304
rect 20260 2261 20269 2295
rect 20269 2261 20303 2295
rect 20303 2261 20312 2295
rect 20260 2252 20312 2261
rect 24584 2252 24636 2304
rect 26424 2252 26476 2304
rect 35716 2295 35768 2304
rect 35716 2261 35725 2295
rect 35725 2261 35759 2295
rect 35759 2261 35768 2295
rect 35716 2252 35768 2261
rect 37740 2252 37792 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
<< metal2 >>
rect 662 40765 718 41565
rect 2594 40765 2650 41565
rect 5170 40765 5226 41565
rect 7102 40765 7158 41565
rect 9678 40882 9734 41565
rect 9678 40854 9812 40882
rect 9678 40765 9734 40854
rect 676 39098 704 40765
rect 1122 39536 1178 39545
rect 1122 39471 1178 39480
rect 664 39092 716 39098
rect 664 39034 716 39040
rect 1136 39030 1164 39471
rect 1124 39024 1176 39030
rect 1124 38966 1176 38972
rect 1768 38956 1820 38962
rect 1768 38898 1820 38904
rect 2044 38956 2096 38962
rect 2044 38898 2096 38904
rect 1780 37670 1808 38898
rect 2056 38554 2084 38898
rect 2044 38548 2096 38554
rect 2044 38490 2096 38496
rect 940 37664 992 37670
rect 940 37606 992 37612
rect 1768 37664 1820 37670
rect 1768 37606 1820 37612
rect 952 37505 980 37606
rect 938 37496 994 37505
rect 938 37431 994 37440
rect 2608 37330 2636 40765
rect 5184 39794 5212 40765
rect 5184 39766 5304 39794
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 4874 39131 5182 39140
rect 5276 39098 5304 39766
rect 9784 39098 9812 40854
rect 11610 40765 11666 41565
rect 14186 40765 14242 41565
rect 16118 40765 16174 41565
rect 18694 40765 18750 41565
rect 20626 40765 20682 41565
rect 23202 40765 23258 41565
rect 25134 40765 25190 41565
rect 27066 40882 27122 41565
rect 27066 40854 27384 40882
rect 27066 40765 27122 40854
rect 14200 39098 14228 40765
rect 20640 39114 20668 40765
rect 5264 39092 5316 39098
rect 5264 39034 5316 39040
rect 9772 39092 9824 39098
rect 9772 39034 9824 39040
rect 14188 39092 14240 39098
rect 14188 39034 14240 39040
rect 17592 39092 17644 39098
rect 20640 39086 20760 39114
rect 23216 39098 23244 40765
rect 25148 39098 25176 40765
rect 27356 39098 27384 40854
rect 29642 40765 29698 41565
rect 31574 40765 31630 41565
rect 34150 40765 34206 41565
rect 36082 40882 36138 41565
rect 36082 40854 36400 40882
rect 36082 40765 36138 40854
rect 31588 39114 31616 40765
rect 31588 39098 31892 39114
rect 34164 39098 34192 40765
rect 35594 39196 35902 39205
rect 35594 39194 35600 39196
rect 35656 39194 35680 39196
rect 35736 39194 35760 39196
rect 35816 39194 35840 39196
rect 35896 39194 35902 39196
rect 35656 39142 35658 39194
rect 35838 39142 35840 39194
rect 35594 39140 35600 39142
rect 35656 39140 35680 39142
rect 35736 39140 35760 39142
rect 35816 39140 35840 39142
rect 35896 39140 35902 39142
rect 35594 39131 35902 39140
rect 36372 39098 36400 40854
rect 38658 40765 38714 41565
rect 37186 40216 37242 40225
rect 37186 40151 37242 40160
rect 17592 39034 17644 39040
rect 9680 38956 9732 38962
rect 9680 38898 9732 38904
rect 10140 38956 10192 38962
rect 10140 38898 10192 38904
rect 14740 38956 14792 38962
rect 14740 38898 14792 38904
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 9692 38554 9720 38898
rect 9680 38548 9732 38554
rect 9680 38490 9732 38496
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 10152 38010 10180 38898
rect 13912 38820 13964 38826
rect 13912 38762 13964 38768
rect 11612 38344 11664 38350
rect 11612 38286 11664 38292
rect 10324 38208 10376 38214
rect 10324 38150 10376 38156
rect 10336 38010 10364 38150
rect 10140 38004 10192 38010
rect 10140 37946 10192 37952
rect 10324 38004 10376 38010
rect 10324 37946 10376 37952
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 11624 37466 11652 38286
rect 12072 37868 12124 37874
rect 12072 37810 12124 37816
rect 12992 37868 13044 37874
rect 13044 37828 13124 37856
rect 12992 37810 13044 37816
rect 12084 37466 12112 37810
rect 11612 37460 11664 37466
rect 11612 37402 11664 37408
rect 12072 37460 12124 37466
rect 12072 37402 12124 37408
rect 2596 37324 2648 37330
rect 2596 37266 2648 37272
rect 8484 37324 8536 37330
rect 8484 37266 8536 37272
rect 11980 37324 12032 37330
rect 12032 37284 12204 37312
rect 11980 37266 12032 37272
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 8300 36168 8352 36174
rect 8300 36110 8352 36116
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 8208 35692 8260 35698
rect 8312 35680 8340 36110
rect 8260 35652 8340 35680
rect 8208 35634 8260 35640
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 940 35012 992 35018
rect 940 34954 992 34960
rect 6000 35012 6052 35018
rect 6000 34954 6052 34960
rect 952 34785 980 34954
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 938 34776 994 34785
rect 4874 34779 5182 34788
rect 938 34711 994 34720
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4068 33992 4120 33998
rect 4068 33934 4120 33940
rect 4080 33454 4108 33934
rect 5724 33924 5776 33930
rect 5724 33866 5776 33872
rect 5356 33856 5408 33862
rect 5356 33798 5408 33804
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 5368 33590 5396 33798
rect 5736 33658 5764 33866
rect 5724 33652 5776 33658
rect 5724 33594 5776 33600
rect 4620 33584 4672 33590
rect 4620 33526 4672 33532
rect 5356 33584 5408 33590
rect 5356 33526 5408 33532
rect 4068 33448 4120 33454
rect 4068 33390 4120 33396
rect 4080 31890 4108 33390
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4632 33114 4660 33526
rect 4620 33108 4672 33114
rect 4620 33050 4672 33056
rect 5368 32994 5396 33526
rect 5816 33312 5868 33318
rect 5816 33254 5868 33260
rect 5368 32966 5488 32994
rect 5356 32904 5408 32910
rect 5356 32846 5408 32852
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4804 32020 4856 32026
rect 4804 31962 4856 31968
rect 4068 31884 4120 31890
rect 4068 31826 4120 31832
rect 3332 31816 3384 31822
rect 3332 31758 3384 31764
rect 4160 31816 4212 31822
rect 4160 31758 4212 31764
rect 3344 31346 3372 31758
rect 4172 31346 4200 31758
rect 3332 31340 3384 31346
rect 3332 31282 3384 31288
rect 4160 31340 4212 31346
rect 4160 31282 4212 31288
rect 3056 31272 3108 31278
rect 3056 31214 3108 31220
rect 3424 31272 3476 31278
rect 3424 31214 3476 31220
rect 4620 31272 4672 31278
rect 4620 31214 4672 31220
rect 3068 30938 3096 31214
rect 3056 30932 3108 30938
rect 3056 30874 3108 30880
rect 3332 30728 3384 30734
rect 3332 30670 3384 30676
rect 3344 30258 3372 30670
rect 3436 30258 3464 31214
rect 4068 31136 4120 31142
rect 4068 31078 4120 31084
rect 4080 30938 4108 31078
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4632 30938 4660 31214
rect 4068 30932 4120 30938
rect 4068 30874 4120 30880
rect 4620 30932 4672 30938
rect 4620 30874 4672 30880
rect 4528 30864 4580 30870
rect 4528 30806 4580 30812
rect 3976 30728 4028 30734
rect 3976 30670 4028 30676
rect 4344 30728 4396 30734
rect 4344 30670 4396 30676
rect 3332 30252 3384 30258
rect 3332 30194 3384 30200
rect 3424 30252 3476 30258
rect 3424 30194 3476 30200
rect 3516 30252 3568 30258
rect 3516 30194 3568 30200
rect 1768 29708 1820 29714
rect 1768 29650 1820 29656
rect 1676 29572 1728 29578
rect 1676 29514 1728 29520
rect 1688 29306 1716 29514
rect 1676 29300 1728 29306
rect 1676 29242 1728 29248
rect 1780 28626 1808 29650
rect 2688 29640 2740 29646
rect 2688 29582 2740 29588
rect 2780 29640 2832 29646
rect 2780 29582 2832 29588
rect 1768 28620 1820 28626
rect 1768 28562 1820 28568
rect 2136 28620 2188 28626
rect 2136 28562 2188 28568
rect 1768 27872 1820 27878
rect 1768 27814 1820 27820
rect 1400 26444 1452 26450
rect 1400 26386 1452 26392
rect 938 25936 994 25945
rect 938 25871 940 25880
rect 992 25871 994 25880
rect 940 25842 992 25848
rect 1412 25362 1440 26386
rect 1780 25974 1808 27814
rect 2148 26994 2176 28562
rect 2700 28082 2728 29582
rect 2792 28490 2820 29582
rect 3528 28762 3556 30194
rect 3608 30184 3660 30190
rect 3608 30126 3660 30132
rect 3620 29782 3648 30126
rect 3988 30054 4016 30670
rect 4068 30660 4120 30666
rect 4068 30602 4120 30608
rect 4080 30394 4108 30602
rect 4068 30388 4120 30394
rect 4068 30330 4120 30336
rect 4356 30054 4384 30670
rect 4436 30592 4488 30598
rect 4436 30534 4488 30540
rect 4448 30394 4476 30534
rect 4540 30394 4568 30806
rect 4816 30734 4844 31962
rect 5264 31748 5316 31754
rect 5264 31690 5316 31696
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 5276 31482 5304 31690
rect 5264 31476 5316 31482
rect 5264 31418 5316 31424
rect 4988 31340 5040 31346
rect 4988 31282 5040 31288
rect 4804 30728 4856 30734
rect 4804 30670 4856 30676
rect 4712 30660 4764 30666
rect 4712 30602 4764 30608
rect 4436 30388 4488 30394
rect 4436 30330 4488 30336
rect 4528 30388 4580 30394
rect 4528 30330 4580 30336
rect 4620 30252 4672 30258
rect 4620 30194 4672 30200
rect 3976 30048 4028 30054
rect 3976 29990 4028 29996
rect 4344 30048 4396 30054
rect 4344 29990 4396 29996
rect 3608 29776 3660 29782
rect 3608 29718 3660 29724
rect 3988 29306 4016 29990
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4528 29640 4580 29646
rect 4528 29582 4580 29588
rect 4344 29572 4396 29578
rect 4344 29514 4396 29520
rect 3976 29300 4028 29306
rect 3976 29242 4028 29248
rect 4356 29102 4384 29514
rect 4540 29306 4568 29582
rect 4528 29300 4580 29306
rect 4528 29242 4580 29248
rect 4632 29209 4660 30194
rect 4724 30122 4752 30602
rect 4816 30122 4844 30670
rect 5000 30666 5028 31282
rect 5080 31272 5132 31278
rect 5080 31214 5132 31220
rect 5092 30938 5120 31214
rect 5264 31136 5316 31142
rect 5264 31078 5316 31084
rect 5080 30932 5132 30938
rect 5080 30874 5132 30880
rect 4988 30660 5040 30666
rect 4988 30602 5040 30608
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 5276 30326 5304 31078
rect 5264 30320 5316 30326
rect 5264 30262 5316 30268
rect 4988 30184 5040 30190
rect 4988 30126 5040 30132
rect 4712 30116 4764 30122
rect 4712 30058 4764 30064
rect 4804 30116 4856 30122
rect 4804 30058 4856 30064
rect 4724 29578 4752 30058
rect 4816 29782 4844 30058
rect 5000 30054 5028 30126
rect 4988 30048 5040 30054
rect 4988 29990 5040 29996
rect 5000 29782 5028 29990
rect 4804 29776 4856 29782
rect 4804 29718 4856 29724
rect 4988 29776 5040 29782
rect 4988 29718 5040 29724
rect 4712 29572 4764 29578
rect 4712 29514 4764 29520
rect 4618 29200 4674 29209
rect 4618 29135 4674 29144
rect 4724 29152 4752 29514
rect 4816 29288 4844 29718
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 5080 29300 5132 29306
rect 4816 29260 5028 29288
rect 5000 29170 5028 29260
rect 5080 29242 5132 29248
rect 5092 29209 5120 29242
rect 5078 29200 5134 29209
rect 4804 29164 4856 29170
rect 4724 29124 4804 29152
rect 4804 29106 4856 29112
rect 4988 29164 5040 29170
rect 5078 29135 5134 29144
rect 5264 29164 5316 29170
rect 4988 29106 5040 29112
rect 5264 29106 5316 29112
rect 4344 29096 4396 29102
rect 4344 29038 4396 29044
rect 4620 29028 4672 29034
rect 4620 28970 4672 28976
rect 4988 29028 5040 29034
rect 4988 28970 5040 28976
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4632 28762 4660 28970
rect 4712 28960 4764 28966
rect 4712 28902 4764 28908
rect 3516 28756 3568 28762
rect 3516 28698 3568 28704
rect 4620 28756 4672 28762
rect 4620 28698 4672 28704
rect 2780 28484 2832 28490
rect 2780 28426 2832 28432
rect 2688 28076 2740 28082
rect 2688 28018 2740 28024
rect 2792 27130 2820 28426
rect 4724 28150 4752 28902
rect 5000 28558 5028 28970
rect 5276 28762 5304 29106
rect 5264 28756 5316 28762
rect 5264 28698 5316 28704
rect 4988 28552 5040 28558
rect 4988 28494 5040 28500
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4712 28144 4764 28150
rect 4712 28086 4764 28092
rect 5264 27872 5316 27878
rect 5264 27814 5316 27820
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4804 27668 4856 27674
rect 4804 27610 4856 27616
rect 4160 27600 4212 27606
rect 4160 27542 4212 27548
rect 2780 27124 2832 27130
rect 2780 27066 2832 27072
rect 2136 26988 2188 26994
rect 2136 26930 2188 26936
rect 2148 26586 2176 26930
rect 2136 26580 2188 26586
rect 2136 26522 2188 26528
rect 2792 26382 2820 27066
rect 3976 26988 4028 26994
rect 3976 26930 4028 26936
rect 3424 26920 3476 26926
rect 3424 26862 3476 26868
rect 2780 26376 2832 26382
rect 2780 26318 2832 26324
rect 1768 25968 1820 25974
rect 1768 25910 1820 25916
rect 1400 25356 1452 25362
rect 1400 25298 1452 25304
rect 2792 25294 2820 26318
rect 3436 26042 3464 26862
rect 3988 26518 4016 26930
rect 4172 26874 4200 27542
rect 4620 27328 4672 27334
rect 4620 27270 4672 27276
rect 4712 27328 4764 27334
rect 4712 27270 4764 27276
rect 4080 26846 4200 26874
rect 4080 26790 4108 26846
rect 4632 26790 4660 27270
rect 4068 26784 4120 26790
rect 4068 26726 4120 26732
rect 4620 26784 4672 26790
rect 4620 26726 4672 26732
rect 3976 26512 4028 26518
rect 3976 26454 4028 26460
rect 4080 26466 4108 26726
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4080 26438 4200 26466
rect 4632 26450 4660 26726
rect 3424 26036 3476 26042
rect 3424 25978 3476 25984
rect 4172 25906 4200 26438
rect 4620 26444 4672 26450
rect 4620 26386 4672 26392
rect 4528 26308 4580 26314
rect 4528 26250 4580 26256
rect 4540 25974 4568 26250
rect 4528 25968 4580 25974
rect 4528 25910 4580 25916
rect 3332 25900 3384 25906
rect 3332 25842 3384 25848
rect 4160 25900 4212 25906
rect 4160 25842 4212 25848
rect 4620 25900 4672 25906
rect 4620 25842 4672 25848
rect 2780 25288 2832 25294
rect 2832 25248 2912 25276
rect 2780 25230 2832 25236
rect 1676 25220 1728 25226
rect 1676 25162 1728 25168
rect 1688 24954 1716 25162
rect 1676 24948 1728 24954
rect 1676 24890 1728 24896
rect 2780 24948 2832 24954
rect 2780 24890 2832 24896
rect 2792 24206 2820 24890
rect 2780 24200 2832 24206
rect 2780 24142 2832 24148
rect 2320 24064 2372 24070
rect 2320 24006 2372 24012
rect 2332 23866 2360 24006
rect 2320 23860 2372 23866
rect 2320 23802 2372 23808
rect 1768 23520 1820 23526
rect 1768 23462 1820 23468
rect 2884 23474 2912 25248
rect 2964 24812 3016 24818
rect 2964 24754 3016 24760
rect 2976 24274 3004 24754
rect 2964 24268 3016 24274
rect 2964 24210 3016 24216
rect 2964 23520 3016 23526
rect 2884 23468 2964 23474
rect 2884 23462 3016 23468
rect 1780 23186 1808 23462
rect 2884 23446 3004 23462
rect 2884 23322 2912 23446
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 1768 23180 1820 23186
rect 1768 23122 1820 23128
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 940 21344 992 21350
rect 940 21286 992 21292
rect 952 21185 980 21286
rect 938 21176 994 21185
rect 938 21111 994 21120
rect 1412 21010 1440 23054
rect 3344 22098 3372 25842
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4528 25356 4580 25362
rect 4528 25298 4580 25304
rect 3792 25152 3844 25158
rect 3792 25094 3844 25100
rect 3804 24954 3832 25094
rect 3792 24948 3844 24954
rect 3792 24890 3844 24896
rect 4540 24698 4568 25298
rect 4632 24834 4660 25842
rect 4724 25294 4752 27270
rect 4816 26994 4844 27610
rect 5276 27334 5304 27814
rect 5264 27328 5316 27334
rect 5264 27270 5316 27276
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4804 26988 4856 26994
rect 4804 26930 4856 26936
rect 5276 26790 5304 27270
rect 4804 26784 4856 26790
rect 4804 26726 4856 26732
rect 5264 26784 5316 26790
rect 5264 26726 5316 26732
rect 4816 26518 4844 26726
rect 4804 26512 4856 26518
rect 4804 26454 4856 26460
rect 5276 26246 5304 26726
rect 5264 26240 5316 26246
rect 5264 26182 5316 26188
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 5276 25906 5304 26182
rect 5264 25900 5316 25906
rect 5264 25842 5316 25848
rect 4804 25764 4856 25770
rect 4804 25706 4856 25712
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 4816 24954 4844 25706
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4804 24948 4856 24954
rect 4804 24890 4856 24896
rect 4632 24818 4752 24834
rect 4620 24812 4752 24818
rect 4672 24806 4752 24812
rect 4620 24754 4672 24760
rect 4540 24670 4660 24698
rect 3700 24608 3752 24614
rect 3700 24550 3752 24556
rect 3712 24274 3740 24550
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4632 24274 4660 24670
rect 4724 24410 4752 24806
rect 4804 24812 4856 24818
rect 4804 24754 4856 24760
rect 4712 24404 4764 24410
rect 4712 24346 4764 24352
rect 4816 24290 4844 24754
rect 5368 24682 5396 32846
rect 5460 31686 5488 32966
rect 5828 32910 5856 33254
rect 5816 32904 5868 32910
rect 5816 32846 5868 32852
rect 5724 32768 5776 32774
rect 5724 32710 5776 32716
rect 5448 31680 5500 31686
rect 5448 31622 5500 31628
rect 5448 30252 5500 30258
rect 5448 30194 5500 30200
rect 5460 25770 5488 30194
rect 5540 28552 5592 28558
rect 5540 28494 5592 28500
rect 5552 27674 5580 28494
rect 5632 28416 5684 28422
rect 5632 28358 5684 28364
rect 5540 27668 5592 27674
rect 5540 27610 5592 27616
rect 5644 27130 5672 28358
rect 5632 27124 5684 27130
rect 5632 27066 5684 27072
rect 5540 26920 5592 26926
rect 5540 26862 5592 26868
rect 5552 26586 5580 26862
rect 5540 26580 5592 26586
rect 5540 26522 5592 26528
rect 5736 26042 5764 32710
rect 6012 28540 6040 34954
rect 6920 34128 6972 34134
rect 6920 34070 6972 34076
rect 6092 33516 6144 33522
rect 6092 33458 6144 33464
rect 6736 33516 6788 33522
rect 6736 33458 6788 33464
rect 6104 33114 6132 33458
rect 6748 33114 6776 33458
rect 6092 33108 6144 33114
rect 6092 33050 6144 33056
rect 6736 33108 6788 33114
rect 6736 33050 6788 33056
rect 6932 32910 6960 34070
rect 8300 33652 8352 33658
rect 8300 33594 8352 33600
rect 7012 33448 7064 33454
rect 7012 33390 7064 33396
rect 6920 32904 6972 32910
rect 6920 32846 6972 32852
rect 6736 32768 6788 32774
rect 6736 32710 6788 32716
rect 6644 31748 6696 31754
rect 6644 31690 6696 31696
rect 6656 31482 6684 31690
rect 6644 31476 6696 31482
rect 6644 31418 6696 31424
rect 6460 31408 6512 31414
rect 6460 31350 6512 31356
rect 6184 28960 6236 28966
rect 6184 28902 6236 28908
rect 6196 28558 6224 28902
rect 6092 28552 6144 28558
rect 6012 28512 6092 28540
rect 5816 28484 5868 28490
rect 5816 28426 5868 28432
rect 5828 28218 5856 28426
rect 5816 28212 5868 28218
rect 5816 28154 5868 28160
rect 5908 26988 5960 26994
rect 5908 26930 5960 26936
rect 5920 26790 5948 26930
rect 6012 26874 6040 28512
rect 6092 28494 6144 28500
rect 6184 28552 6236 28558
rect 6184 28494 6236 28500
rect 6368 28552 6420 28558
rect 6368 28494 6420 28500
rect 6092 27872 6144 27878
rect 6092 27814 6144 27820
rect 6104 26994 6132 27814
rect 6196 26994 6224 28494
rect 6092 26988 6144 26994
rect 6092 26930 6144 26936
rect 6184 26988 6236 26994
rect 6184 26930 6236 26936
rect 6012 26846 6132 26874
rect 5908 26784 5960 26790
rect 5908 26726 5960 26732
rect 5724 26036 5776 26042
rect 5644 25996 5724 26024
rect 5448 25764 5500 25770
rect 5448 25706 5500 25712
rect 5448 25220 5500 25226
rect 5448 25162 5500 25168
rect 5356 24676 5408 24682
rect 5356 24618 5408 24624
rect 5264 24608 5316 24614
rect 5264 24550 5316 24556
rect 3700 24268 3752 24274
rect 3700 24210 3752 24216
rect 4620 24268 4672 24274
rect 4620 24210 4672 24216
rect 4724 24262 4844 24290
rect 3516 23656 3568 23662
rect 3516 23598 3568 23604
rect 3528 23322 3556 23598
rect 3516 23316 3568 23322
rect 3516 23258 3568 23264
rect 3712 23254 3740 24210
rect 3792 24200 3844 24206
rect 3792 24142 3844 24148
rect 3976 24200 4028 24206
rect 3976 24142 4028 24148
rect 3804 23866 3832 24142
rect 3792 23860 3844 23866
rect 3792 23802 3844 23808
rect 3884 23792 3936 23798
rect 3884 23734 3936 23740
rect 3792 23520 3844 23526
rect 3792 23462 3844 23468
rect 3700 23248 3752 23254
rect 3700 23190 3752 23196
rect 3804 22234 3832 23462
rect 3896 23322 3924 23734
rect 3988 23662 4016 24142
rect 4068 23792 4120 23798
rect 4068 23734 4120 23740
rect 3976 23656 4028 23662
rect 3976 23598 4028 23604
rect 4080 23526 4108 23734
rect 4620 23656 4672 23662
rect 4620 23598 4672 23604
rect 4068 23520 4120 23526
rect 4068 23462 4120 23468
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23322 4660 23598
rect 3884 23316 3936 23322
rect 3884 23258 3936 23264
rect 4620 23316 4672 23322
rect 4620 23258 4672 23264
rect 4724 22982 4752 24262
rect 5276 24070 5304 24550
rect 4804 24064 4856 24070
rect 4804 24006 4856 24012
rect 5264 24064 5316 24070
rect 5264 24006 5316 24012
rect 4816 23662 4844 24006
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4804 23656 4856 23662
rect 4804 23598 4856 23604
rect 5276 23526 5304 24006
rect 5264 23520 5316 23526
rect 5264 23462 5316 23468
rect 4712 22976 4764 22982
rect 4712 22918 4764 22924
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 5368 22692 5396 24618
rect 5460 23848 5488 25162
rect 5540 24744 5592 24750
rect 5540 24686 5592 24692
rect 5552 24138 5580 24686
rect 5644 24206 5672 25996
rect 5724 25978 5776 25984
rect 5816 25152 5868 25158
rect 5816 25094 5868 25100
rect 5632 24200 5684 24206
rect 5632 24142 5684 24148
rect 5540 24132 5592 24138
rect 5540 24074 5592 24080
rect 5460 23820 5580 23848
rect 5448 23724 5500 23730
rect 5448 23666 5500 23672
rect 5184 22664 5396 22692
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 3792 22228 3844 22234
rect 3792 22170 3844 22176
rect 3332 22092 3384 22098
rect 3332 22034 3384 22040
rect 3148 21956 3200 21962
rect 3148 21898 3200 21904
rect 2504 21888 2556 21894
rect 2504 21830 2556 21836
rect 3056 21888 3108 21894
rect 3056 21830 3108 21836
rect 2516 21690 2544 21830
rect 2504 21684 2556 21690
rect 2504 21626 2556 21632
rect 3068 21622 3096 21830
rect 3056 21616 3108 21622
rect 3056 21558 3108 21564
rect 1768 21548 1820 21554
rect 1768 21490 1820 21496
rect 2780 21548 2832 21554
rect 2780 21490 2832 21496
rect 1400 21004 1452 21010
rect 1400 20946 1452 20952
rect 1412 19378 1440 20946
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 940 18760 992 18766
rect 940 18702 992 18708
rect 952 18465 980 18702
rect 938 18456 994 18465
rect 938 18391 994 18400
rect 1412 18290 1440 19314
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1412 17746 1440 18226
rect 1400 17740 1452 17746
rect 1400 17682 1452 17688
rect 938 16416 994 16425
rect 938 16351 994 16360
rect 952 16182 980 16351
rect 940 16176 992 16182
rect 940 16118 992 16124
rect 1780 15162 1808 21490
rect 1860 21344 1912 21350
rect 1860 21286 1912 21292
rect 1872 21146 1900 21286
rect 1860 21140 1912 21146
rect 1860 21082 1912 21088
rect 2792 21078 2820 21490
rect 2780 21072 2832 21078
rect 2780 21014 2832 21020
rect 3160 20913 3188 21898
rect 3146 20904 3202 20913
rect 3146 20839 3202 20848
rect 3160 20806 3188 20839
rect 3148 20800 3200 20806
rect 3148 20742 3200 20748
rect 3344 19922 3372 22034
rect 3804 21622 3832 22170
rect 5184 22098 5212 22664
rect 5356 22568 5408 22574
rect 5356 22510 5408 22516
rect 5368 22166 5396 22510
rect 5356 22160 5408 22166
rect 5356 22102 5408 22108
rect 5172 22092 5224 22098
rect 5172 22034 5224 22040
rect 5264 22024 5316 22030
rect 5264 21966 5316 21972
rect 4528 21888 4580 21894
rect 4528 21830 4580 21836
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 4540 21622 4568 21830
rect 3792 21616 3844 21622
rect 3792 21558 3844 21564
rect 4528 21616 4580 21622
rect 4528 21558 4580 21564
rect 3804 20806 3832 21558
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 3792 20800 3844 20806
rect 3792 20742 3844 20748
rect 4080 19922 4108 20946
rect 4632 20874 4660 21830
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5276 21690 5304 21966
rect 5264 21684 5316 21690
rect 5264 21626 5316 21632
rect 4620 20868 4672 20874
rect 4620 20810 4672 20816
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3332 19916 3384 19922
rect 3252 19876 3332 19904
rect 1952 19712 2004 19718
rect 1952 19654 2004 19660
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 1964 19446 1992 19654
rect 3160 19446 3188 19654
rect 1952 19440 2004 19446
rect 3148 19440 3200 19446
rect 1952 19382 2004 19388
rect 3146 19408 3148 19417
rect 3200 19408 3202 19417
rect 3146 19343 3202 19352
rect 3252 19310 3280 19876
rect 3332 19858 3384 19864
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 3332 19780 3384 19786
rect 3332 19722 3384 19728
rect 4068 19780 4120 19786
rect 4068 19722 4120 19728
rect 3240 19304 3292 19310
rect 3240 19246 3292 19252
rect 3344 19174 3372 19722
rect 4080 19514 4108 19722
rect 4804 19712 4856 19718
rect 4804 19654 4856 19660
rect 4816 19514 4844 19654
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 4712 19440 4764 19446
rect 4712 19382 4764 19388
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 2044 18624 2096 18630
rect 2044 18566 2096 18572
rect 2056 18426 2084 18566
rect 2044 18420 2096 18426
rect 2044 18362 2096 18368
rect 3240 18284 3292 18290
rect 3344 18272 3372 19110
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3608 18828 3660 18834
rect 3608 18770 3660 18776
rect 3620 18426 3648 18770
rect 4724 18426 4752 19382
rect 5368 19310 5396 22102
rect 5460 22030 5488 23666
rect 5552 22778 5580 23820
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 5540 22500 5592 22506
rect 5540 22442 5592 22448
rect 5448 22024 5500 22030
rect 5448 21966 5500 21972
rect 5552 21672 5580 22442
rect 5460 21644 5580 21672
rect 5460 19990 5488 21644
rect 5540 21548 5592 21554
rect 5644 21536 5672 24142
rect 5592 21508 5672 21536
rect 5540 21490 5592 21496
rect 5448 19984 5500 19990
rect 5448 19926 5500 19932
rect 5356 19304 5408 19310
rect 5356 19246 5408 19252
rect 5368 18834 5396 19246
rect 5356 18828 5408 18834
rect 5356 18770 5408 18776
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 4712 18420 4764 18426
rect 4712 18362 4764 18368
rect 3292 18244 3372 18272
rect 3240 18226 3292 18232
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 1872 16658 1900 17682
rect 2504 16992 2556 16998
rect 2504 16934 2556 16940
rect 2516 16658 2544 16934
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 2504 16652 2556 16658
rect 2504 16594 2556 16600
rect 3252 16590 3280 18226
rect 5368 18222 5396 18770
rect 5460 18766 5488 19926
rect 5448 18760 5500 18766
rect 5448 18702 5500 18708
rect 5552 18426 5580 21490
rect 5828 19514 5856 25094
rect 5908 24608 5960 24614
rect 5908 24550 5960 24556
rect 5920 22506 5948 24550
rect 6104 24206 6132 26846
rect 6196 24614 6224 26930
rect 6380 25906 6408 28494
rect 6472 28422 6500 31350
rect 6552 30660 6604 30666
rect 6552 30602 6604 30608
rect 6564 30190 6592 30602
rect 6552 30184 6604 30190
rect 6552 30126 6604 30132
rect 6748 28490 6776 32710
rect 7024 31890 7052 33390
rect 7472 32972 7524 32978
rect 7472 32914 7524 32920
rect 7104 32904 7156 32910
rect 7104 32846 7156 32852
rect 7012 31884 7064 31890
rect 7012 31826 7064 31832
rect 6920 31272 6972 31278
rect 6920 31214 6972 31220
rect 6828 29164 6880 29170
rect 6828 29106 6880 29112
rect 6840 28762 6868 29106
rect 6932 29102 6960 31214
rect 7024 30802 7052 31826
rect 7012 30796 7064 30802
rect 7012 30738 7064 30744
rect 6920 29096 6972 29102
rect 6920 29038 6972 29044
rect 6828 28756 6880 28762
rect 6828 28698 6880 28704
rect 6828 28620 6880 28626
rect 6828 28562 6880 28568
rect 6736 28484 6788 28490
rect 6736 28426 6788 28432
rect 6460 28416 6512 28422
rect 6460 28358 6512 28364
rect 6368 25900 6420 25906
rect 6368 25842 6420 25848
rect 6472 25158 6500 28358
rect 6644 26920 6696 26926
rect 6564 26868 6644 26874
rect 6564 26862 6696 26868
rect 6564 26846 6684 26862
rect 6460 25152 6512 25158
rect 6460 25094 6512 25100
rect 6564 24750 6592 26846
rect 6644 25832 6696 25838
rect 6644 25774 6696 25780
rect 6656 24857 6684 25774
rect 6642 24848 6698 24857
rect 6642 24783 6698 24792
rect 6656 24750 6684 24783
rect 6552 24744 6604 24750
rect 6552 24686 6604 24692
rect 6644 24744 6696 24750
rect 6644 24686 6696 24692
rect 6184 24608 6236 24614
rect 6184 24550 6236 24556
rect 6656 24392 6684 24686
rect 6748 24410 6776 28426
rect 6840 27878 6868 28562
rect 6828 27872 6880 27878
rect 6828 27814 6880 27820
rect 6932 27674 6960 29038
rect 6920 27668 6972 27674
rect 6920 27610 6972 27616
rect 7012 27668 7064 27674
rect 7012 27610 7064 27616
rect 6920 27464 6972 27470
rect 6840 27424 6920 27452
rect 6840 26790 6868 27424
rect 6920 27406 6972 27412
rect 6920 27056 6972 27062
rect 7024 27044 7052 27610
rect 7116 27606 7144 32846
rect 7484 31754 7512 32914
rect 8312 32910 8340 33594
rect 8300 32904 8352 32910
rect 8300 32846 8352 32852
rect 7932 32836 7984 32842
rect 7932 32778 7984 32784
rect 7944 32366 7972 32778
rect 8208 32768 8260 32774
rect 8208 32710 8260 32716
rect 8220 32570 8248 32710
rect 8208 32564 8260 32570
rect 8208 32506 8260 32512
rect 7656 32360 7708 32366
rect 7656 32302 7708 32308
rect 7932 32360 7984 32366
rect 7932 32302 7984 32308
rect 7668 31890 7696 32302
rect 8496 31890 8524 37266
rect 11612 37120 11664 37126
rect 11612 37062 11664 37068
rect 10692 36712 10744 36718
rect 10692 36654 10744 36660
rect 9864 36236 9916 36242
rect 9864 36178 9916 36184
rect 9220 36168 9272 36174
rect 9220 36110 9272 36116
rect 8944 35624 8996 35630
rect 8944 35566 8996 35572
rect 8956 35290 8984 35566
rect 8944 35284 8996 35290
rect 8944 35226 8996 35232
rect 8944 33516 8996 33522
rect 8944 33458 8996 33464
rect 8956 32502 8984 33458
rect 9232 33454 9260 36110
rect 9772 36100 9824 36106
rect 9772 36042 9824 36048
rect 9784 35834 9812 36042
rect 9772 35828 9824 35834
rect 9772 35770 9824 35776
rect 9876 35766 9904 36178
rect 9864 35760 9916 35766
rect 9864 35702 9916 35708
rect 9876 35034 9904 35702
rect 9956 35624 10008 35630
rect 9956 35566 10008 35572
rect 9968 35290 9996 35566
rect 10704 35494 10732 36654
rect 11624 36106 11652 37062
rect 11612 36100 11664 36106
rect 11612 36042 11664 36048
rect 11244 36032 11296 36038
rect 11244 35974 11296 35980
rect 11256 35834 11284 35974
rect 11244 35828 11296 35834
rect 11244 35770 11296 35776
rect 11256 35630 11284 35770
rect 11060 35624 11112 35630
rect 11060 35566 11112 35572
rect 11244 35624 11296 35630
rect 11244 35566 11296 35572
rect 10692 35488 10744 35494
rect 10692 35430 10744 35436
rect 9956 35284 10008 35290
rect 9956 35226 10008 35232
rect 10704 35154 10732 35430
rect 11072 35290 11100 35566
rect 11624 35329 11652 36042
rect 11796 35556 11848 35562
rect 11796 35498 11848 35504
rect 11610 35320 11666 35329
rect 11060 35284 11112 35290
rect 11808 35290 11836 35498
rect 11888 35488 11940 35494
rect 11888 35430 11940 35436
rect 11900 35290 11928 35430
rect 11610 35255 11666 35264
rect 11796 35284 11848 35290
rect 11060 35226 11112 35232
rect 11796 35226 11848 35232
rect 11888 35284 11940 35290
rect 11888 35226 11940 35232
rect 10692 35148 10744 35154
rect 10692 35090 10744 35096
rect 9876 35006 9996 35034
rect 9864 34944 9916 34950
rect 9864 34886 9916 34892
rect 9876 34746 9904 34886
rect 9864 34740 9916 34746
rect 9864 34682 9916 34688
rect 9968 33590 9996 35006
rect 9772 33584 9824 33590
rect 9772 33526 9824 33532
rect 9956 33584 10008 33590
rect 9956 33526 10008 33532
rect 9220 33448 9272 33454
rect 9220 33390 9272 33396
rect 8944 32496 8996 32502
rect 8680 32444 8944 32450
rect 8680 32438 8996 32444
rect 8680 32422 8984 32438
rect 7656 31884 7708 31890
rect 7656 31826 7708 31832
rect 8484 31884 8536 31890
rect 8484 31826 8536 31832
rect 7392 31726 7512 31754
rect 7392 31278 7420 31726
rect 7668 31482 7696 31826
rect 8680 31822 8708 32422
rect 8668 31816 8720 31822
rect 8668 31758 8720 31764
rect 8116 31680 8168 31686
rect 8116 31622 8168 31628
rect 7656 31476 7708 31482
rect 7656 31418 7708 31424
rect 7472 31408 7524 31414
rect 7472 31350 7524 31356
rect 7380 31272 7432 31278
rect 7380 31214 7432 31220
rect 7392 30802 7420 31214
rect 7380 30796 7432 30802
rect 7380 30738 7432 30744
rect 7288 30660 7340 30666
rect 7288 30602 7340 30608
rect 7300 30394 7328 30602
rect 7288 30388 7340 30394
rect 7288 30330 7340 30336
rect 7288 29572 7340 29578
rect 7288 29514 7340 29520
rect 7300 29306 7328 29514
rect 7288 29300 7340 29306
rect 7288 29242 7340 29248
rect 7288 29096 7340 29102
rect 7288 29038 7340 29044
rect 7300 27606 7328 29038
rect 7380 28552 7432 28558
rect 7380 28494 7432 28500
rect 7392 28082 7420 28494
rect 7380 28076 7432 28082
rect 7380 28018 7432 28024
rect 7104 27600 7156 27606
rect 7104 27542 7156 27548
rect 7288 27600 7340 27606
rect 7288 27542 7340 27548
rect 6972 27016 7052 27044
rect 6920 26998 6972 27004
rect 6920 26920 6972 26926
rect 6920 26862 6972 26868
rect 6828 26784 6880 26790
rect 6828 26726 6880 26732
rect 6840 26586 6868 26726
rect 6828 26580 6880 26586
rect 6828 26522 6880 26528
rect 6840 26246 6868 26522
rect 6828 26240 6880 26246
rect 6828 26182 6880 26188
rect 6840 25294 6868 26182
rect 6932 26042 6960 26862
rect 7024 26450 7052 27016
rect 7012 26444 7064 26450
rect 7012 26386 7064 26392
rect 6920 26036 6972 26042
rect 6920 25978 6972 25984
rect 6828 25288 6880 25294
rect 6828 25230 6880 25236
rect 6920 25288 6972 25294
rect 6920 25230 6972 25236
rect 6932 24818 6960 25230
rect 6920 24812 6972 24818
rect 6920 24754 6972 24760
rect 6828 24676 6880 24682
rect 6828 24618 6880 24624
rect 6288 24364 6684 24392
rect 6736 24404 6788 24410
rect 6092 24200 6144 24206
rect 6092 24142 6144 24148
rect 6000 24132 6052 24138
rect 6000 24074 6052 24080
rect 5908 22500 5960 22506
rect 5908 22442 5960 22448
rect 6012 22094 6040 24074
rect 5920 22066 6040 22094
rect 5816 19508 5868 19514
rect 5816 19450 5868 19456
rect 5920 18970 5948 22066
rect 6000 21956 6052 21962
rect 6000 21898 6052 21904
rect 6012 21690 6040 21898
rect 6184 21888 6236 21894
rect 6184 21830 6236 21836
rect 6000 21684 6052 21690
rect 6000 21626 6052 21632
rect 6090 21584 6146 21593
rect 6090 21519 6092 21528
rect 6144 21519 6146 21528
rect 6092 21490 6144 21496
rect 6104 21146 6132 21490
rect 6092 21140 6144 21146
rect 6092 21082 6144 21088
rect 6196 20806 6224 21830
rect 6184 20800 6236 20806
rect 6184 20742 6236 20748
rect 6196 19922 6224 20742
rect 6184 19916 6236 19922
rect 6184 19858 6236 19864
rect 6000 19780 6052 19786
rect 6000 19722 6052 19728
rect 6012 19334 6040 19722
rect 6012 19306 6224 19334
rect 5908 18964 5960 18970
rect 5908 18906 5960 18912
rect 5632 18624 5684 18630
rect 5632 18566 5684 18572
rect 5540 18420 5592 18426
rect 5540 18362 5592 18368
rect 5356 18216 5408 18222
rect 5356 18158 5408 18164
rect 4804 18148 4856 18154
rect 4804 18090 4856 18096
rect 3700 18080 3752 18086
rect 3700 18022 3752 18028
rect 3712 17338 3740 18022
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4816 17882 4844 18090
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 3700 17332 3752 17338
rect 3700 17274 3752 17280
rect 3988 17202 4016 17682
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 4632 17338 4660 17478
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 3988 16250 4016 17138
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4816 16658 4844 17818
rect 4908 17678 4936 18022
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 5644 17610 5672 18566
rect 5632 17604 5684 17610
rect 5632 17546 5684 17552
rect 6196 17542 6224 19306
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 6196 17270 6224 17478
rect 6184 17264 6236 17270
rect 6184 17206 6236 17212
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 5080 15904 5132 15910
rect 5080 15846 5132 15852
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 1768 15156 1820 15162
rect 1768 15098 1820 15104
rect 1952 15020 2004 15026
rect 1952 14962 2004 14968
rect 1964 14618 1992 14962
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 1504 13705 1532 13806
rect 1490 13696 1546 13705
rect 1490 13631 1546 13640
rect 3988 13326 4016 15438
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 3896 12986 3924 13126
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 940 11756 992 11762
rect 940 11698 992 11704
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 952 11665 980 11698
rect 938 11656 994 11665
rect 938 11591 994 11600
rect 2148 11354 2176 11698
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 3988 10130 4016 13262
rect 4080 11665 4108 15846
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 5092 15570 5120 15846
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 5368 14482 5488 14498
rect 5356 14476 5488 14482
rect 5408 14470 5488 14476
rect 5356 14418 5408 14424
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4540 13734 4568 14350
rect 4632 14074 4660 14350
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 5276 14074 5304 14214
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 4804 13796 4856 13802
rect 4804 13738 4856 13744
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4436 12776 4488 12782
rect 4488 12724 4660 12730
rect 4436 12718 4660 12724
rect 4448 12702 4660 12718
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12442 4660 12702
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 4724 12238 4752 13126
rect 4816 12306 4844 13738
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5276 13326 5304 13670
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 5276 12918 5304 13262
rect 5264 12912 5316 12918
rect 5264 12854 5316 12860
rect 5460 12434 5488 14470
rect 5552 13394 5580 16594
rect 6196 16522 6224 17206
rect 6184 16516 6236 16522
rect 6184 16458 6236 16464
rect 6196 15570 6224 16458
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6196 14346 6224 15506
rect 6184 14340 6236 14346
rect 6184 14282 6236 14288
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5368 12406 5488 12434
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 5368 11778 5396 12406
rect 5448 12164 5500 12170
rect 5448 12106 5500 12112
rect 5460 11898 5488 12106
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5368 11750 5488 11778
rect 4066 11656 4122 11665
rect 4066 11591 4122 11600
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 5460 11082 5488 11750
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4724 10266 4752 10406
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 3976 10124 4028 10130
rect 3976 10066 4028 10072
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 8974 4660 10066
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4540 8634 4568 8774
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4908 8090 4936 8366
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5460 6186 5488 11018
rect 5552 10520 5580 13330
rect 6196 12918 6224 14282
rect 6184 12912 6236 12918
rect 6184 12854 6236 12860
rect 6196 12170 6224 12854
rect 6184 12164 6236 12170
rect 6184 12106 6236 12112
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 5644 10674 5672 11086
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5816 10532 5868 10538
rect 5552 10492 5816 10520
rect 5816 10474 5868 10480
rect 6184 9988 6236 9994
rect 6184 9930 6236 9936
rect 6196 9518 6224 9930
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6196 8650 6224 9454
rect 6104 8622 6224 8650
rect 6104 8566 6132 8622
rect 6092 8560 6144 8566
rect 6092 8502 6144 8508
rect 6184 8560 6236 8566
rect 6184 8502 6236 8508
rect 6196 7886 6224 8502
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 5460 5710 5488 6122
rect 5736 5778 5764 7822
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 5920 7002 5948 7142
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 6000 6724 6052 6730
rect 6000 6666 6052 6672
rect 6012 6458 6040 6666
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4172 5234 4200 5510
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 940 4548 992 4554
rect 940 4490 992 4496
rect 952 4185 980 4490
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 1780 3126 1808 4966
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 6288 4826 6316 24364
rect 6736 24346 6788 24352
rect 6644 24200 6696 24206
rect 6644 24142 6696 24148
rect 6656 24070 6684 24142
rect 6644 24064 6696 24070
rect 6644 24006 6696 24012
rect 6656 23526 6684 24006
rect 6644 23520 6696 23526
rect 6644 23462 6696 23468
rect 6460 22432 6512 22438
rect 6460 22374 6512 22380
rect 6472 22094 6500 22374
rect 6748 22094 6776 24346
rect 6840 23798 6868 24618
rect 6932 24410 6960 24754
rect 6920 24404 6972 24410
rect 6920 24346 6972 24352
rect 6920 24200 6972 24206
rect 7024 24188 7052 26386
rect 7116 24750 7144 27542
rect 7288 27328 7340 27334
rect 7288 27270 7340 27276
rect 7300 26994 7328 27270
rect 7288 26988 7340 26994
rect 7288 26930 7340 26936
rect 7196 26920 7248 26926
rect 7196 26862 7248 26868
rect 7104 24744 7156 24750
rect 7104 24686 7156 24692
rect 6972 24160 7052 24188
rect 6920 24142 6972 24148
rect 6828 23792 6880 23798
rect 6932 23769 6960 24142
rect 6828 23734 6880 23740
rect 6918 23760 6974 23769
rect 6918 23695 6974 23704
rect 6920 23656 6972 23662
rect 6920 23598 6972 23604
rect 6932 23322 6960 23598
rect 6920 23316 6972 23322
rect 6920 23258 6972 23264
rect 7116 23066 7144 24686
rect 7208 24070 7236 26862
rect 7300 26790 7328 26930
rect 7288 26784 7340 26790
rect 7288 26726 7340 26732
rect 7300 26586 7328 26726
rect 7288 26580 7340 26586
rect 7288 26522 7340 26528
rect 7300 25974 7328 26522
rect 7392 26194 7420 28018
rect 7484 26382 7512 31350
rect 8128 31346 8156 31622
rect 8116 31340 8168 31346
rect 8116 31282 8168 31288
rect 8680 30734 8708 31758
rect 9232 31482 9260 33390
rect 9784 33114 9812 33526
rect 9968 33454 9996 33526
rect 9956 33448 10008 33454
rect 9956 33390 10008 33396
rect 9772 33108 9824 33114
rect 9772 33050 9824 33056
rect 10704 32978 10732 35090
rect 11980 35080 12032 35086
rect 11980 35022 12032 35028
rect 11704 35012 11756 35018
rect 11704 34954 11756 34960
rect 11612 34944 11664 34950
rect 11612 34886 11664 34892
rect 11624 34610 11652 34886
rect 11716 34746 11744 34954
rect 11992 34785 12020 35022
rect 11978 34776 12034 34785
rect 11704 34740 11756 34746
rect 11704 34682 11756 34688
rect 11808 34734 11978 34762
rect 11612 34604 11664 34610
rect 11612 34546 11664 34552
rect 11808 33658 11836 34734
rect 11978 34711 12034 34720
rect 11980 34468 12032 34474
rect 11980 34410 12032 34416
rect 11796 33652 11848 33658
rect 11796 33594 11848 33600
rect 11992 33590 12020 34410
rect 11980 33584 12032 33590
rect 12032 33544 12112 33572
rect 11980 33526 12032 33532
rect 11704 33516 11756 33522
rect 11704 33458 11756 33464
rect 11796 33516 11848 33522
rect 11796 33458 11848 33464
rect 11888 33516 11940 33522
rect 11888 33458 11940 33464
rect 11612 33448 11664 33454
rect 11612 33390 11664 33396
rect 10968 33312 11020 33318
rect 10968 33254 11020 33260
rect 11520 33312 11572 33318
rect 11520 33254 11572 33260
rect 10692 32972 10744 32978
rect 10692 32914 10744 32920
rect 10980 32774 11008 33254
rect 11532 32978 11560 33254
rect 11624 32978 11652 33390
rect 11716 33114 11744 33458
rect 11808 33114 11836 33458
rect 11704 33108 11756 33114
rect 11704 33050 11756 33056
rect 11796 33108 11848 33114
rect 11796 33050 11848 33056
rect 11520 32972 11572 32978
rect 11520 32914 11572 32920
rect 11612 32972 11664 32978
rect 11612 32914 11664 32920
rect 10784 32768 10836 32774
rect 10784 32710 10836 32716
rect 10968 32768 11020 32774
rect 10968 32710 11020 32716
rect 9588 31816 9640 31822
rect 9588 31758 9640 31764
rect 9220 31476 9272 31482
rect 9220 31418 9272 31424
rect 9232 31346 9260 31418
rect 9600 31396 9628 31758
rect 10796 31754 10824 32710
rect 11336 32428 11388 32434
rect 11336 32370 11388 32376
rect 10796 31726 10916 31754
rect 9864 31408 9916 31414
rect 9600 31368 9864 31396
rect 9864 31350 9916 31356
rect 9220 31340 9272 31346
rect 9220 31282 9272 31288
rect 9588 31272 9640 31278
rect 9588 31214 9640 31220
rect 9404 31136 9456 31142
rect 9404 31078 9456 31084
rect 9416 30802 9444 31078
rect 9600 30938 9628 31214
rect 9588 30932 9640 30938
rect 9588 30874 9640 30880
rect 10888 30802 10916 31726
rect 11152 31340 11204 31346
rect 11152 31282 11204 31288
rect 11060 31136 11112 31142
rect 11060 31078 11112 31084
rect 9404 30796 9456 30802
rect 9404 30738 9456 30744
rect 10876 30796 10928 30802
rect 10876 30738 10928 30744
rect 8668 30728 8720 30734
rect 8668 30670 8720 30676
rect 8944 30592 8996 30598
rect 8944 30534 8996 30540
rect 9312 30592 9364 30598
rect 9312 30534 9364 30540
rect 8956 30394 8984 30534
rect 8944 30388 8996 30394
rect 8944 30330 8996 30336
rect 8024 29708 8076 29714
rect 8024 29650 8076 29656
rect 8036 29102 8064 29650
rect 8300 29504 8352 29510
rect 8300 29446 8352 29452
rect 8760 29504 8812 29510
rect 8760 29446 8812 29452
rect 8024 29096 8076 29102
rect 8024 29038 8076 29044
rect 8036 28014 8064 29038
rect 8312 28150 8340 29446
rect 8772 29238 8800 29446
rect 8760 29232 8812 29238
rect 8760 29174 8812 29180
rect 9036 28212 9088 28218
rect 8772 28172 9036 28200
rect 8300 28144 8352 28150
rect 8300 28086 8352 28092
rect 8576 28144 8628 28150
rect 8576 28086 8628 28092
rect 8024 28008 8076 28014
rect 8024 27950 8076 27956
rect 8300 28008 8352 28014
rect 8300 27950 8352 27956
rect 7656 27464 7708 27470
rect 7656 27406 7708 27412
rect 7564 27328 7616 27334
rect 7564 27270 7616 27276
rect 7576 27062 7604 27270
rect 7564 27056 7616 27062
rect 7564 26998 7616 27004
rect 7668 26994 7696 27406
rect 7656 26988 7708 26994
rect 7656 26930 7708 26936
rect 7668 26790 7696 26930
rect 8036 26858 8064 27950
rect 8312 27674 8340 27950
rect 8588 27674 8616 28086
rect 8300 27668 8352 27674
rect 8300 27610 8352 27616
rect 8576 27668 8628 27674
rect 8576 27610 8628 27616
rect 8208 27396 8260 27402
rect 8208 27338 8260 27344
rect 8220 27130 8248 27338
rect 8208 27124 8260 27130
rect 8208 27066 8260 27072
rect 8668 26988 8720 26994
rect 8668 26930 8720 26936
rect 8024 26852 8076 26858
rect 8024 26794 8076 26800
rect 7656 26784 7708 26790
rect 7656 26726 7708 26732
rect 8036 26450 8064 26794
rect 8208 26784 8260 26790
rect 8208 26726 8260 26732
rect 8024 26444 8076 26450
rect 8024 26386 8076 26392
rect 7472 26376 7524 26382
rect 7472 26318 7524 26324
rect 7932 26308 7984 26314
rect 7932 26250 7984 26256
rect 7392 26166 7512 26194
rect 7288 25968 7340 25974
rect 7288 25910 7340 25916
rect 7288 25764 7340 25770
rect 7288 25706 7340 25712
rect 7300 25498 7328 25706
rect 7288 25492 7340 25498
rect 7288 25434 7340 25440
rect 7484 24750 7512 26166
rect 7748 25900 7800 25906
rect 7748 25842 7800 25848
rect 7656 24812 7708 24818
rect 7656 24754 7708 24760
rect 7472 24744 7524 24750
rect 7472 24686 7524 24692
rect 7564 24744 7616 24750
rect 7564 24686 7616 24692
rect 7484 24585 7512 24686
rect 7576 24614 7604 24686
rect 7564 24608 7616 24614
rect 7470 24576 7526 24585
rect 7564 24550 7616 24556
rect 7470 24511 7526 24520
rect 7668 24426 7696 24754
rect 7392 24398 7696 24426
rect 7196 24064 7248 24070
rect 7196 24006 7248 24012
rect 7392 23798 7420 24398
rect 7380 23792 7432 23798
rect 7380 23734 7432 23740
rect 7288 23112 7340 23118
rect 7116 23060 7288 23066
rect 7116 23054 7340 23060
rect 7116 23038 7328 23054
rect 7116 22778 7144 23038
rect 7104 22772 7156 22778
rect 7104 22714 7156 22720
rect 7196 22568 7248 22574
rect 7024 22516 7196 22522
rect 7024 22510 7248 22516
rect 7024 22494 7236 22510
rect 6472 22066 6592 22094
rect 6748 22066 6868 22094
rect 6564 21554 6592 22066
rect 6552 21548 6604 21554
rect 6552 21490 6604 21496
rect 6840 20534 6868 22066
rect 6828 20528 6880 20534
rect 6828 20470 6880 20476
rect 6460 20256 6512 20262
rect 6460 20198 6512 20204
rect 6472 19922 6500 20198
rect 6460 19916 6512 19922
rect 6460 19858 6512 19864
rect 6840 19514 6868 20470
rect 6828 19508 6880 19514
rect 6828 19450 6880 19456
rect 6368 19168 6420 19174
rect 6368 19110 6420 19116
rect 6380 18766 6408 19110
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 6460 18148 6512 18154
rect 6460 18090 6512 18096
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 6380 16250 6408 16390
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6472 14006 6500 18090
rect 6736 16448 6788 16454
rect 6736 16390 6788 16396
rect 6748 15706 6776 16390
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6564 14074 6592 14214
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6472 12238 6500 13262
rect 6840 12434 6868 15438
rect 7024 14906 7052 22494
rect 7392 22386 7420 23734
rect 7760 23254 7788 25842
rect 7748 23248 7800 23254
rect 7748 23190 7800 23196
rect 7748 22704 7800 22710
rect 7748 22646 7800 22652
rect 7116 22358 7420 22386
rect 7116 22234 7144 22358
rect 7104 22228 7156 22234
rect 7104 22170 7156 22176
rect 7116 22030 7144 22170
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 7760 21962 7788 22646
rect 7944 22094 7972 26250
rect 8036 24818 8064 26386
rect 8220 25294 8248 26726
rect 8680 26586 8708 26930
rect 8668 26580 8720 26586
rect 8668 26522 8720 26528
rect 8300 25424 8352 25430
rect 8300 25366 8352 25372
rect 8208 25288 8260 25294
rect 8208 25230 8260 25236
rect 8116 24948 8168 24954
rect 8116 24890 8168 24896
rect 8024 24812 8076 24818
rect 8024 24754 8076 24760
rect 8128 23186 8156 24890
rect 8312 24750 8340 25366
rect 8300 24744 8352 24750
rect 8300 24686 8352 24692
rect 8392 23588 8444 23594
rect 8392 23530 8444 23536
rect 8404 23186 8432 23530
rect 8116 23180 8168 23186
rect 8116 23122 8168 23128
rect 8392 23180 8444 23186
rect 8392 23122 8444 23128
rect 7944 22066 8064 22094
rect 7748 21956 7800 21962
rect 7748 21898 7800 21904
rect 7760 21350 7788 21898
rect 7748 21344 7800 21350
rect 7748 21286 7800 21292
rect 8036 20942 8064 22066
rect 8128 21486 8156 23122
rect 8668 23044 8720 23050
rect 8668 22986 8720 22992
rect 8300 22500 8352 22506
rect 8300 22442 8352 22448
rect 8116 21480 8168 21486
rect 8116 21422 8168 21428
rect 8024 20936 8076 20942
rect 8024 20878 8076 20884
rect 7932 20528 7984 20534
rect 7930 20496 7932 20505
rect 7984 20496 7986 20505
rect 7930 20431 7986 20440
rect 7944 20058 7972 20431
rect 8128 20330 8156 21422
rect 8208 21412 8260 21418
rect 8208 21354 8260 21360
rect 8220 21146 8248 21354
rect 8208 21140 8260 21146
rect 8208 21082 8260 21088
rect 8220 20466 8248 21082
rect 8312 20534 8340 22442
rect 8484 21412 8536 21418
rect 8484 21354 8536 21360
rect 8576 21412 8628 21418
rect 8576 21354 8628 21360
rect 8496 20534 8524 21354
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 8484 20528 8536 20534
rect 8484 20470 8536 20476
rect 8208 20460 8260 20466
rect 8208 20402 8260 20408
rect 8116 20324 8168 20330
rect 8116 20266 8168 20272
rect 8024 20256 8076 20262
rect 8024 20198 8076 20204
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 8036 19378 8064 20198
rect 8312 19938 8340 20470
rect 8312 19910 8432 19938
rect 8298 19816 8354 19825
rect 8298 19751 8300 19760
rect 8352 19751 8354 19760
rect 8300 19722 8352 19728
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7760 18698 7788 19110
rect 7748 18692 7800 18698
rect 7748 18634 7800 18640
rect 7760 18290 7788 18634
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 7760 17882 7788 18226
rect 7840 18080 7892 18086
rect 7840 18022 7892 18028
rect 7852 17882 7880 18022
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 7300 16658 7328 17614
rect 7760 17542 7788 17818
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 7760 16658 7788 17478
rect 7852 17270 7880 17818
rect 8036 17610 8064 19314
rect 8404 18970 8432 19910
rect 8496 19174 8524 20470
rect 8588 20262 8616 21354
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 8208 18896 8260 18902
rect 8208 18838 8260 18844
rect 8220 18442 8248 18838
rect 8128 18414 8340 18442
rect 8128 17678 8156 18414
rect 8312 18290 8340 18414
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 8116 17672 8168 17678
rect 8116 17614 8168 17620
rect 8024 17604 8076 17610
rect 8024 17546 8076 17552
rect 8392 17604 8444 17610
rect 8392 17546 8444 17552
rect 7840 17264 7892 17270
rect 7840 17206 7892 17212
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 7748 16652 7800 16658
rect 7748 16594 7800 16600
rect 6932 14878 7052 14906
rect 6932 13258 6960 14878
rect 7116 14414 7144 16594
rect 7300 16250 7328 16594
rect 7656 16448 7708 16454
rect 7656 16390 7708 16396
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 7668 16114 7696 16390
rect 7760 16114 7788 16594
rect 7852 16590 7880 17206
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 7840 16584 7892 16590
rect 7840 16526 7892 16532
rect 7944 16250 7972 17138
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 8220 16658 8248 16934
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 8128 16114 8156 16526
rect 8404 16114 8432 17546
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 7760 15910 7788 16050
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 7208 14958 7236 15302
rect 7760 15094 7788 15302
rect 7748 15088 7800 15094
rect 7748 15030 7800 15036
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 8036 14482 8064 14894
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 8024 14476 8076 14482
rect 8024 14418 8076 14424
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7116 13394 7144 13670
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 6748 12406 6868 12434
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6472 11150 6500 12174
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6656 10606 6684 11630
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6380 10130 6408 10406
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6564 9722 6592 9862
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6564 7478 6592 7686
rect 6552 7472 6604 7478
rect 6552 7414 6604 7420
rect 6656 7274 6684 10542
rect 6748 10130 6776 12406
rect 6828 12164 6880 12170
rect 6828 12106 6880 12112
rect 6840 11898 6868 12106
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 6932 11830 6960 13194
rect 6920 11824 6972 11830
rect 6920 11766 6972 11772
rect 6920 11688 6972 11694
rect 7208 11676 7236 14418
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7576 14074 7604 14214
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 8220 12481 8248 14418
rect 8484 14340 8536 14346
rect 8484 14282 8536 14288
rect 8496 13530 8524 14282
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8206 12472 8262 12481
rect 8128 12416 8206 12434
rect 8128 12407 8262 12416
rect 8128 12406 8248 12407
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 6972 11648 7236 11676
rect 6920 11630 6972 11636
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 7116 11218 7144 11494
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6932 10742 6960 11018
rect 7392 10810 7420 11698
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 6828 10532 6880 10538
rect 6828 10474 6880 10480
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 6748 7886 6776 10066
rect 6840 10010 6868 10474
rect 6840 9982 6960 10010
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6840 9722 6868 9862
rect 6932 9722 6960 9982
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6932 9602 6960 9658
rect 6840 9574 6960 9602
rect 7760 9586 7788 11018
rect 7748 9580 7800 9586
rect 6840 8090 6868 9574
rect 7748 9522 7800 9528
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 8498 6960 8774
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6644 7268 6696 7274
rect 6644 7210 6696 7216
rect 6748 6322 6776 7822
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6748 5642 6776 6258
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 6932 5166 6960 8434
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7208 7546 7236 8230
rect 7944 8090 7972 9522
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 7288 7812 7340 7818
rect 7288 7754 7340 7760
rect 7300 7546 7328 7754
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7208 7002 7236 7482
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7944 6798 7972 8026
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7760 5642 7788 6734
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 6932 3534 6960 5102
rect 7024 5098 7052 5578
rect 8036 5574 8064 11698
rect 8128 10130 8156 12406
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8496 10810 8524 10950
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 8128 9602 8156 10066
rect 8220 9926 8248 10474
rect 8588 10062 8616 10746
rect 8680 10674 8708 22986
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8680 10266 8708 10610
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8220 9722 8248 9862
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8128 9574 8340 9602
rect 8312 7342 8340 9574
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8680 7546 8708 7890
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 8036 5166 8064 5510
rect 8312 5166 8340 7278
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8588 5302 8616 5714
rect 8576 5296 8628 5302
rect 8576 5238 8628 5244
rect 8680 5166 8708 6054
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 7012 5092 7064 5098
rect 7012 5034 7064 5040
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 1768 3120 1820 3126
rect 1768 3062 1820 3068
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 1952 2848 2004 2854
rect 1952 2790 2004 2796
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 32 800 60 2314
rect 1504 2145 1532 2790
rect 1964 2446 1992 2790
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 6932 2446 6960 2790
rect 8772 2774 8800 28172
rect 9036 28154 9088 28160
rect 8944 28008 8996 28014
rect 8944 27950 8996 27956
rect 8850 21992 8906 22001
rect 8850 21927 8852 21936
rect 8904 21927 8906 21936
rect 8852 21898 8904 21904
rect 8852 18352 8904 18358
rect 8852 18294 8904 18300
rect 8864 17338 8892 18294
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8956 15688 8984 27950
rect 9324 26790 9352 30534
rect 10600 30048 10652 30054
rect 10600 29990 10652 29996
rect 9680 29504 9732 29510
rect 9680 29446 9732 29452
rect 9692 29238 9720 29446
rect 9680 29232 9732 29238
rect 9680 29174 9732 29180
rect 9864 29232 9916 29238
rect 9864 29174 9916 29180
rect 9588 27872 9640 27878
rect 9588 27814 9640 27820
rect 9772 27872 9824 27878
rect 9772 27814 9824 27820
rect 9600 27334 9628 27814
rect 9784 27606 9812 27814
rect 9876 27674 9904 29174
rect 9864 27668 9916 27674
rect 9864 27610 9916 27616
rect 9772 27600 9824 27606
rect 9772 27542 9824 27548
rect 9680 27532 9732 27538
rect 9680 27474 9732 27480
rect 9588 27328 9640 27334
rect 9588 27270 9640 27276
rect 9312 26784 9364 26790
rect 9312 26726 9364 26732
rect 9404 26784 9456 26790
rect 9404 26726 9456 26732
rect 9324 26330 9352 26726
rect 9416 26518 9444 26726
rect 9404 26512 9456 26518
rect 9404 26454 9456 26460
rect 9324 26302 9444 26330
rect 9416 26246 9444 26302
rect 9404 26240 9456 26246
rect 9404 26182 9456 26188
rect 9496 25288 9548 25294
rect 9496 25230 9548 25236
rect 9036 25152 9088 25158
rect 9036 25094 9088 25100
rect 9048 24750 9076 25094
rect 9036 24744 9088 24750
rect 9036 24686 9088 24692
rect 9508 24206 9536 25230
rect 9600 25158 9628 27270
rect 9692 26042 9720 27474
rect 9876 27062 9904 27610
rect 9864 27056 9916 27062
rect 9864 26998 9916 27004
rect 9876 26314 9904 26998
rect 10416 26444 10468 26450
rect 10416 26386 10468 26392
rect 9864 26308 9916 26314
rect 9864 26250 9916 26256
rect 9680 26036 9732 26042
rect 9680 25978 9732 25984
rect 9876 25922 9904 26250
rect 9876 25894 10272 25922
rect 9680 25696 9732 25702
rect 9680 25638 9732 25644
rect 9588 25152 9640 25158
rect 9588 25094 9640 25100
rect 9496 24200 9548 24206
rect 9496 24142 9548 24148
rect 9508 23866 9536 24142
rect 9588 24064 9640 24070
rect 9588 24006 9640 24012
rect 9600 23866 9628 24006
rect 9496 23860 9548 23866
rect 9496 23802 9548 23808
rect 9588 23860 9640 23866
rect 9588 23802 9640 23808
rect 9404 23792 9456 23798
rect 9404 23734 9456 23740
rect 9036 23656 9088 23662
rect 9036 23598 9088 23604
rect 9048 22030 9076 23598
rect 9416 22794 9444 23734
rect 9416 22778 9628 22794
rect 9404 22772 9628 22778
rect 9456 22766 9628 22772
rect 9404 22714 9456 22720
rect 9312 22636 9364 22642
rect 9312 22578 9364 22584
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9324 22098 9352 22578
rect 9312 22092 9364 22098
rect 9312 22034 9364 22040
rect 9036 22024 9088 22030
rect 9036 21966 9088 21972
rect 9048 21418 9076 21966
rect 9220 21888 9272 21894
rect 9220 21830 9272 21836
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9232 21622 9260 21830
rect 9324 21690 9352 21830
rect 9312 21684 9364 21690
rect 9312 21626 9364 21632
rect 9220 21616 9272 21622
rect 9220 21558 9272 21564
rect 9036 21412 9088 21418
rect 9036 21354 9088 21360
rect 9048 20874 9076 21354
rect 9036 20868 9088 20874
rect 9036 20810 9088 20816
rect 9416 20466 9444 22578
rect 9496 22160 9548 22166
rect 9496 22102 9548 22108
rect 9508 21554 9536 22102
rect 9496 21548 9548 21554
rect 9496 21490 9548 21496
rect 9404 20460 9456 20466
rect 9404 20402 9456 20408
rect 9128 20392 9180 20398
rect 9128 20334 9180 20340
rect 9140 20262 9168 20334
rect 9128 20256 9180 20262
rect 9128 20198 9180 20204
rect 9140 16590 9168 20198
rect 9312 19780 9364 19786
rect 9312 19722 9364 19728
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9232 16658 9260 17138
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9232 16250 9260 16594
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 8864 15660 8984 15688
rect 8864 11676 8892 15660
rect 9324 15570 9352 19722
rect 9496 19440 9548 19446
rect 9496 19382 9548 19388
rect 9508 18766 9536 19382
rect 9600 18766 9628 22766
rect 9692 22642 9720 25638
rect 9772 25424 9824 25430
rect 9772 25366 9824 25372
rect 9784 24410 9812 25366
rect 9864 25220 9916 25226
rect 9864 25162 9916 25168
rect 9772 24404 9824 24410
rect 9772 24346 9824 24352
rect 9772 22976 9824 22982
rect 9772 22918 9824 22924
rect 9784 22778 9812 22918
rect 9772 22772 9824 22778
rect 9772 22714 9824 22720
rect 9876 22642 9904 25162
rect 10244 24138 10272 25894
rect 10428 25362 10456 26386
rect 10416 25356 10468 25362
rect 10416 25298 10468 25304
rect 10428 24886 10456 25298
rect 10416 24880 10468 24886
rect 10416 24822 10468 24828
rect 10416 24744 10468 24750
rect 10416 24686 10468 24692
rect 10232 24132 10284 24138
rect 10232 24074 10284 24080
rect 10232 23316 10284 23322
rect 10232 23258 10284 23264
rect 10244 22982 10272 23258
rect 10324 23248 10376 23254
rect 10324 23190 10376 23196
rect 10232 22976 10284 22982
rect 10232 22918 10284 22924
rect 9680 22636 9732 22642
rect 9680 22578 9732 22584
rect 9864 22636 9916 22642
rect 9864 22578 9916 22584
rect 9876 22522 9904 22578
rect 9692 22494 9904 22522
rect 9692 20602 9720 22494
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9784 22250 9812 22374
rect 9784 22222 9996 22250
rect 9864 22160 9916 22166
rect 9864 22102 9916 22108
rect 9772 22024 9824 22030
rect 9772 21966 9824 21972
rect 9784 21894 9812 21966
rect 9876 21962 9904 22102
rect 9864 21956 9916 21962
rect 9864 21898 9916 21904
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9772 21480 9824 21486
rect 9772 21422 9824 21428
rect 9784 20602 9812 21422
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9772 20596 9824 20602
rect 9772 20538 9824 20544
rect 9692 19854 9720 20538
rect 9784 20058 9812 20538
rect 9772 20052 9824 20058
rect 9772 19994 9824 20000
rect 9876 19938 9904 21898
rect 9968 21486 9996 22222
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 9956 21480 10008 21486
rect 9956 21422 10008 21428
rect 9956 21344 10008 21350
rect 9956 21286 10008 21292
rect 9784 19910 9904 19938
rect 9784 19854 9812 19910
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9692 18970 9720 19314
rect 9784 18970 9812 19314
rect 9876 19310 9904 19790
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9588 18760 9640 18766
rect 9640 18708 9720 18714
rect 9588 18702 9720 18708
rect 9508 17882 9536 18702
rect 9600 18686 9720 18702
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9692 17678 9720 18686
rect 9968 18612 9996 21286
rect 10060 19334 10088 21830
rect 10336 21570 10364 23190
rect 10428 22001 10456 24686
rect 10508 22976 10560 22982
rect 10508 22918 10560 22924
rect 10520 22098 10548 22918
rect 10612 22778 10640 29990
rect 10888 29714 10916 30738
rect 11072 30734 11100 31078
rect 11164 30870 11192 31282
rect 11152 30864 11204 30870
rect 11152 30806 11204 30812
rect 11060 30728 11112 30734
rect 11060 30670 11112 30676
rect 10692 29708 10744 29714
rect 10692 29650 10744 29656
rect 10876 29708 10928 29714
rect 10876 29650 10928 29656
rect 10704 27538 10732 29650
rect 11164 29646 11192 30806
rect 11152 29640 11204 29646
rect 11152 29582 11204 29588
rect 10876 29572 10928 29578
rect 10876 29514 10928 29520
rect 10888 29306 10916 29514
rect 10876 29300 10928 29306
rect 10876 29242 10928 29248
rect 11164 29170 11192 29582
rect 11152 29164 11204 29170
rect 11152 29106 11204 29112
rect 10692 27532 10744 27538
rect 10692 27474 10744 27480
rect 11244 27328 11296 27334
rect 11244 27270 11296 27276
rect 11256 26586 11284 27270
rect 11244 26580 11296 26586
rect 11244 26522 11296 26528
rect 11348 26466 11376 32370
rect 11624 32366 11652 32914
rect 11704 32904 11756 32910
rect 11704 32846 11756 32852
rect 11612 32360 11664 32366
rect 11612 32302 11664 32308
rect 11520 31816 11572 31822
rect 11520 31758 11572 31764
rect 11532 31346 11560 31758
rect 11716 31754 11744 32846
rect 11796 31816 11848 31822
rect 11796 31758 11848 31764
rect 11704 31748 11756 31754
rect 11704 31690 11756 31696
rect 11520 31340 11572 31346
rect 11520 31282 11572 31288
rect 11520 31136 11572 31142
rect 11520 31078 11572 31084
rect 11532 30938 11560 31078
rect 11520 30932 11572 30938
rect 11520 30874 11572 30880
rect 11716 30666 11744 31690
rect 11808 30938 11836 31758
rect 11900 31414 11928 33458
rect 11980 32768 12032 32774
rect 11980 32710 12032 32716
rect 11992 31822 12020 32710
rect 11980 31816 12032 31822
rect 11980 31758 12032 31764
rect 11888 31408 11940 31414
rect 11888 31350 11940 31356
rect 11796 30932 11848 30938
rect 11796 30874 11848 30880
rect 11704 30660 11756 30666
rect 11704 30602 11756 30608
rect 11520 29504 11572 29510
rect 11520 29446 11572 29452
rect 11796 29504 11848 29510
rect 11796 29446 11848 29452
rect 11532 29306 11560 29446
rect 11808 29306 11836 29446
rect 11520 29300 11572 29306
rect 11520 29242 11572 29248
rect 11796 29300 11848 29306
rect 11796 29242 11848 29248
rect 11900 29238 11928 31350
rect 11992 30666 12020 31758
rect 12084 31346 12112 33544
rect 12176 31414 12204 37284
rect 12440 37256 12492 37262
rect 12440 37198 12492 37204
rect 12716 37256 12768 37262
rect 12716 37198 12768 37204
rect 12348 36780 12400 36786
rect 12348 36722 12400 36728
rect 12360 35494 12388 36722
rect 12452 35873 12480 37198
rect 12728 36922 12756 37198
rect 12900 37120 12952 37126
rect 12900 37062 12952 37068
rect 12912 36922 12940 37062
rect 12716 36916 12768 36922
rect 12716 36858 12768 36864
rect 12900 36916 12952 36922
rect 12900 36858 12952 36864
rect 12992 36848 13044 36854
rect 12992 36790 13044 36796
rect 12716 36712 12768 36718
rect 12716 36654 12768 36660
rect 12624 36032 12676 36038
rect 12624 35974 12676 35980
rect 12438 35864 12494 35873
rect 12636 35834 12664 35974
rect 12728 35834 12756 36654
rect 13004 36310 13032 36790
rect 12992 36304 13044 36310
rect 12992 36246 13044 36252
rect 12438 35799 12494 35808
rect 12624 35828 12676 35834
rect 12624 35770 12676 35776
rect 12716 35828 12768 35834
rect 12716 35770 12768 35776
rect 12440 35692 12492 35698
rect 12440 35634 12492 35640
rect 12348 35488 12400 35494
rect 12348 35430 12400 35436
rect 12360 35086 12388 35430
rect 12452 35290 12480 35634
rect 12532 35624 12584 35630
rect 12532 35566 12584 35572
rect 12440 35284 12492 35290
rect 12440 35226 12492 35232
rect 12544 35170 12572 35566
rect 12636 35290 12664 35770
rect 12992 35624 13044 35630
rect 12990 35592 12992 35601
rect 13044 35592 13046 35601
rect 12990 35527 13046 35536
rect 12624 35284 12676 35290
rect 12624 35226 12676 35232
rect 12452 35142 12572 35170
rect 12900 35148 12952 35154
rect 12452 35086 12480 35142
rect 12900 35090 12952 35096
rect 12348 35080 12400 35086
rect 12348 35022 12400 35028
rect 12440 35080 12492 35086
rect 12440 35022 12492 35028
rect 12348 34672 12400 34678
rect 12348 34614 12400 34620
rect 12256 34604 12308 34610
rect 12256 34546 12308 34552
rect 12268 33658 12296 34546
rect 12256 33652 12308 33658
rect 12256 33594 12308 33600
rect 12360 33318 12388 34614
rect 12452 34066 12480 35022
rect 12532 35012 12584 35018
rect 12532 34954 12584 34960
rect 12440 34060 12492 34066
rect 12440 34002 12492 34008
rect 12440 33448 12492 33454
rect 12440 33390 12492 33396
rect 12348 33312 12400 33318
rect 12348 33254 12400 33260
rect 12256 32836 12308 32842
rect 12256 32778 12308 32784
rect 12268 31822 12296 32778
rect 12360 32502 12388 33254
rect 12348 32496 12400 32502
rect 12348 32438 12400 32444
rect 12256 31816 12308 31822
rect 12256 31758 12308 31764
rect 12348 31816 12400 31822
rect 12348 31758 12400 31764
rect 12164 31408 12216 31414
rect 12164 31350 12216 31356
rect 12072 31340 12124 31346
rect 12072 31282 12124 31288
rect 11980 30660 12032 30666
rect 11980 30602 12032 30608
rect 12084 29782 12112 31282
rect 12072 29776 12124 29782
rect 12072 29718 12124 29724
rect 12176 29458 12204 31350
rect 12360 31210 12388 31758
rect 12452 31482 12480 33390
rect 12544 31822 12572 34954
rect 12716 34944 12768 34950
rect 12716 34886 12768 34892
rect 12728 34474 12756 34886
rect 12716 34468 12768 34474
rect 12716 34410 12768 34416
rect 12912 34406 12940 35090
rect 12992 35080 13044 35086
rect 12992 35022 13044 35028
rect 13004 34610 13032 35022
rect 12992 34604 13044 34610
rect 12992 34546 13044 34552
rect 12624 34400 12676 34406
rect 12624 34342 12676 34348
rect 12900 34400 12952 34406
rect 12900 34342 12952 34348
rect 12636 32842 12664 34342
rect 12992 34060 13044 34066
rect 12992 34002 13044 34008
rect 12900 33924 12952 33930
rect 12900 33866 12952 33872
rect 12912 33658 12940 33866
rect 12900 33652 12952 33658
rect 12900 33594 12952 33600
rect 13004 33538 13032 34002
rect 12716 33516 12768 33522
rect 12716 33458 12768 33464
rect 12912 33510 13032 33538
rect 12728 32910 12756 33458
rect 12716 32904 12768 32910
rect 12716 32846 12768 32852
rect 12624 32836 12676 32842
rect 12624 32778 12676 32784
rect 12808 32428 12860 32434
rect 12808 32370 12860 32376
rect 12624 32224 12676 32230
rect 12624 32166 12676 32172
rect 12532 31816 12584 31822
rect 12532 31758 12584 31764
rect 12636 31482 12664 32166
rect 12440 31476 12492 31482
rect 12440 31418 12492 31424
rect 12624 31476 12676 31482
rect 12624 31418 12676 31424
rect 12348 31204 12400 31210
rect 12348 31146 12400 31152
rect 12348 29776 12400 29782
rect 12348 29718 12400 29724
rect 11992 29430 12204 29458
rect 11888 29232 11940 29238
rect 11888 29174 11940 29180
rect 11796 29164 11848 29170
rect 11796 29106 11848 29112
rect 11704 28076 11756 28082
rect 11704 28018 11756 28024
rect 11716 27402 11744 28018
rect 11808 28014 11836 29106
rect 11796 28008 11848 28014
rect 11796 27950 11848 27956
rect 11992 27826 12020 29430
rect 12164 29300 12216 29306
rect 12164 29242 12216 29248
rect 12176 29073 12204 29242
rect 12360 29238 12388 29718
rect 12256 29232 12308 29238
rect 12256 29174 12308 29180
rect 12348 29232 12400 29238
rect 12348 29174 12400 29180
rect 12162 29064 12218 29073
rect 11808 27798 12020 27826
rect 12084 29022 12162 29050
rect 11704 27396 11756 27402
rect 11704 27338 11756 27344
rect 11256 26438 11376 26466
rect 11060 25152 11112 25158
rect 11060 25094 11112 25100
rect 11072 24954 11100 25094
rect 11060 24948 11112 24954
rect 11060 24890 11112 24896
rect 11060 23112 11112 23118
rect 11060 23054 11112 23060
rect 10784 23044 10836 23050
rect 10784 22986 10836 22992
rect 10600 22772 10652 22778
rect 10600 22714 10652 22720
rect 10508 22092 10560 22098
rect 10508 22034 10560 22040
rect 10414 21992 10470 22001
rect 10414 21927 10470 21936
rect 10244 21542 10364 21570
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 10152 21078 10180 21286
rect 10140 21072 10192 21078
rect 10140 21014 10192 21020
rect 10244 20602 10272 21542
rect 10324 21480 10376 21486
rect 10324 21422 10376 21428
rect 10428 21434 10456 21927
rect 10506 21448 10562 21457
rect 10336 20874 10364 21422
rect 10428 21406 10506 21434
rect 10506 21383 10562 21392
rect 10324 20868 10376 20874
rect 10324 20810 10376 20816
rect 10416 20800 10468 20806
rect 10416 20742 10468 20748
rect 10232 20596 10284 20602
rect 10232 20538 10284 20544
rect 10244 19802 10272 20538
rect 10428 20466 10456 20742
rect 10416 20460 10468 20466
rect 10416 20402 10468 20408
rect 10244 19774 10364 19802
rect 10336 19718 10364 19774
rect 10428 19718 10456 20402
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 10520 19394 10548 21383
rect 10612 21350 10640 22714
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 10704 21554 10732 21626
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10692 21412 10744 21418
rect 10692 21354 10744 21360
rect 10600 21344 10652 21350
rect 10600 21286 10652 21292
rect 10704 21146 10732 21354
rect 10692 21140 10744 21146
rect 10692 21082 10744 21088
rect 10600 20936 10652 20942
rect 10600 20878 10652 20884
rect 10428 19366 10548 19394
rect 10060 19310 10180 19334
rect 10060 19306 10192 19310
rect 10140 19304 10192 19306
rect 10140 19246 10192 19252
rect 10048 18624 10100 18630
rect 9968 18584 10048 18612
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9692 17202 9720 17614
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9772 17128 9824 17134
rect 9692 17076 9772 17082
rect 9692 17070 9824 17076
rect 9692 17054 9812 17070
rect 9588 16720 9640 16726
rect 9416 16668 9588 16674
rect 9416 16662 9640 16668
rect 9416 16646 9628 16662
rect 9416 16590 9444 16646
rect 9692 16590 9720 17054
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9404 16584 9456 16590
rect 9404 16526 9456 16532
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 9416 16114 9444 16390
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9508 16028 9536 16526
rect 9784 16182 9812 16934
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 9772 16176 9824 16182
rect 9772 16118 9824 16124
rect 9876 16114 9904 16526
rect 9968 16250 9996 18584
rect 10048 18566 10100 18572
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 10060 17678 10088 17818
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 10152 17610 10180 19246
rect 10428 18766 10456 19366
rect 10612 19310 10640 20878
rect 10704 19446 10732 21082
rect 10796 20398 10824 22986
rect 11072 22438 11100 23054
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 10968 22228 11020 22234
rect 10968 22170 11020 22176
rect 10876 22092 10928 22098
rect 10876 22034 10928 22040
rect 10888 20942 10916 22034
rect 10980 21962 11008 22170
rect 10968 21956 11020 21962
rect 10968 21898 11020 21904
rect 10980 21622 11008 21898
rect 10968 21616 11020 21622
rect 10968 21558 11020 21564
rect 11152 21344 11204 21350
rect 11152 21286 11204 21292
rect 11164 21146 11192 21286
rect 11152 21140 11204 21146
rect 11152 21082 11204 21088
rect 10876 20936 10928 20942
rect 10928 20896 11008 20924
rect 10876 20878 10928 20884
rect 10980 20466 11008 20896
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 10692 19440 10744 19446
rect 10692 19382 10744 19388
rect 10508 19304 10560 19310
rect 10508 19246 10560 19252
rect 10600 19304 10652 19310
rect 10600 19246 10652 19252
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10336 18290 10364 18566
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 10140 17604 10192 17610
rect 10140 17546 10192 17552
rect 10244 17202 10272 18022
rect 10428 17954 10456 18702
rect 10520 18630 10548 19246
rect 10508 18624 10560 18630
rect 10508 18566 10560 18572
rect 10520 18426 10548 18566
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10428 17926 10548 17954
rect 10414 17776 10470 17785
rect 10336 17734 10414 17762
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9680 16040 9732 16046
rect 9508 16000 9680 16028
rect 9680 15982 9732 15988
rect 9864 15972 9916 15978
rect 9864 15914 9916 15920
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 9784 15706 9812 15846
rect 9876 15706 9904 15914
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 8956 11898 8984 15506
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9140 15162 9168 15438
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 9036 15088 9088 15094
rect 9036 15030 9088 15036
rect 9048 14278 9076 15030
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 9048 13326 9076 14214
rect 9600 14006 9628 14758
rect 9588 14000 9640 14006
rect 9416 13960 9588 13988
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 9140 12782 9168 13738
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 9048 11762 9076 12650
rect 9140 12646 9168 12718
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9140 12442 9168 12582
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 8944 11688 8996 11694
rect 8864 11648 8944 11676
rect 8944 11630 8996 11636
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8956 6798 8984 7686
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 8956 6322 8984 6734
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 9140 5778 9168 12242
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 9416 11642 9444 13960
rect 9588 13942 9640 13948
rect 9784 13938 9812 15642
rect 9968 15586 9996 15846
rect 9876 15570 10088 15586
rect 9864 15564 10088 15570
rect 9916 15558 10088 15564
rect 9864 15506 9916 15512
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9864 14544 9916 14550
rect 9864 14486 9916 14492
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9508 12850 9536 13330
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9600 12918 9628 13126
rect 9692 12986 9720 13670
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9784 12986 9812 13126
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9508 12730 9536 12786
rect 9508 12702 9628 12730
rect 9600 12220 9628 12702
rect 9508 12192 9628 12220
rect 9508 11762 9536 12192
rect 9692 12170 9720 12922
rect 9876 12850 9904 14486
rect 9968 13938 9996 15438
rect 10060 14414 10088 15558
rect 10152 15502 10180 16390
rect 10244 15502 10272 16390
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10152 14414 10180 15438
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10244 15026 10272 15302
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 10048 14408 10100 14414
rect 10048 14350 10100 14356
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9968 13734 9996 13874
rect 10060 13818 10088 14350
rect 10152 13938 10180 14350
rect 10336 13938 10364 17734
rect 10414 17711 10470 17720
rect 10520 17377 10548 17926
rect 10506 17368 10562 17377
rect 10506 17303 10562 17312
rect 10520 17134 10548 17303
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10612 16794 10640 19246
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10704 17338 10732 17818
rect 10796 17610 10824 20334
rect 10888 19009 10916 20402
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 11072 19854 11100 20198
rect 11060 19848 11112 19854
rect 11060 19790 11112 19796
rect 10966 19272 11022 19281
rect 10966 19207 11022 19216
rect 11060 19236 11112 19242
rect 10874 19000 10930 19009
rect 10874 18935 10930 18944
rect 10888 18902 10916 18935
rect 10876 18896 10928 18902
rect 10876 18838 10928 18844
rect 10784 17604 10836 17610
rect 10784 17546 10836 17552
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10704 17134 10732 17274
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10428 16114 10456 16526
rect 10612 16114 10640 16526
rect 10704 16182 10732 17070
rect 10888 16998 10916 17138
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10796 16658 10824 16934
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10692 16176 10744 16182
rect 10692 16118 10744 16124
rect 10416 16108 10468 16114
rect 10416 16050 10468 16056
rect 10600 16108 10652 16114
rect 10600 16050 10652 16056
rect 10980 15994 11008 19207
rect 11060 19178 11112 19184
rect 11072 18902 11100 19178
rect 11164 18970 11192 20742
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 11060 18896 11112 18902
rect 11060 18838 11112 18844
rect 11150 18048 11206 18057
rect 11150 17983 11206 17992
rect 11060 17264 11112 17270
rect 11058 17232 11060 17241
rect 11112 17232 11114 17241
rect 11058 17167 11114 17176
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 11072 16114 11100 16526
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 10888 15966 11008 15994
rect 10888 15910 10916 15966
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 11164 15162 11192 17983
rect 11256 15570 11284 26438
rect 11428 25220 11480 25226
rect 11428 25162 11480 25168
rect 11440 24954 11468 25162
rect 11612 25152 11664 25158
rect 11612 25094 11664 25100
rect 11624 24954 11652 25094
rect 11428 24948 11480 24954
rect 11428 24890 11480 24896
rect 11612 24948 11664 24954
rect 11612 24890 11664 24896
rect 11520 24064 11572 24070
rect 11520 24006 11572 24012
rect 11612 24064 11664 24070
rect 11612 24006 11664 24012
rect 11428 23860 11480 23866
rect 11428 23802 11480 23808
rect 11336 23792 11388 23798
rect 11336 23734 11388 23740
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11152 15156 11204 15162
rect 11152 15098 11204 15104
rect 11058 15056 11114 15065
rect 11058 14991 11114 15000
rect 11072 14890 11100 14991
rect 11060 14884 11112 14890
rect 11060 14826 11112 14832
rect 11072 14482 11100 14826
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10232 13864 10284 13870
rect 10060 13812 10232 13818
rect 10060 13806 10284 13812
rect 10060 13790 10272 13806
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 10060 13462 10088 13670
rect 10048 13456 10100 13462
rect 10048 13398 10100 13404
rect 10336 13326 10364 13874
rect 10520 13462 10548 13874
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 10612 13462 10640 13738
rect 10874 13696 10930 13705
rect 10874 13631 10930 13640
rect 10508 13456 10560 13462
rect 10508 13398 10560 13404
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10232 12844 10284 12850
rect 10336 12832 10364 13262
rect 10612 12850 10640 13398
rect 10782 13288 10838 13297
rect 10782 13223 10838 13232
rect 10284 12804 10364 12832
rect 10232 12786 10284 12792
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 9048 5302 9076 5510
rect 9036 5296 9088 5302
rect 9036 5238 9088 5244
rect 9126 4584 9182 4593
rect 9126 4519 9182 4528
rect 9140 4486 9168 4519
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9048 3534 9076 4422
rect 9232 4298 9260 11630
rect 9416 11614 9536 11642
rect 9508 10606 9536 11614
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9416 10266 9444 10542
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9508 9926 9536 10542
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9324 7546 9352 7686
rect 9508 7546 9536 7686
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9784 5778 9812 12650
rect 9876 12220 9904 12786
rect 10060 12374 10088 12786
rect 10336 12434 10364 12804
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10336 12406 10548 12434
rect 10048 12368 10100 12374
rect 10048 12310 10100 12316
rect 9956 12232 10008 12238
rect 9876 12192 9956 12220
rect 9956 12174 10008 12180
rect 9968 11694 9996 12174
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 10152 11354 10180 11698
rect 10520 11694 10548 12406
rect 10692 12368 10744 12374
rect 10692 12310 10744 12316
rect 10704 11694 10732 12310
rect 10796 12238 10824 13223
rect 10888 12481 10916 13631
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10874 12472 10930 12481
rect 10874 12407 10930 12416
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10520 11558 10548 11630
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9876 9654 9904 10542
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 9876 9178 9904 9454
rect 9864 9172 9916 9178
rect 9864 9114 9916 9120
rect 10138 8256 10194 8265
rect 10138 8191 10194 8200
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 9968 5778 9996 7958
rect 10152 7818 10180 8191
rect 10244 8022 10272 9862
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10428 8634 10456 9318
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10520 8430 10548 11494
rect 10704 11150 10732 11630
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10796 9722 10824 12174
rect 10888 11218 10916 12407
rect 10980 12374 11008 12718
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10980 11830 11008 12174
rect 10968 11824 11020 11830
rect 10968 11766 11020 11772
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10232 8016 10284 8022
rect 10232 7958 10284 7964
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 10152 7342 10180 7754
rect 10336 7546 10364 7890
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10336 5914 10364 6054
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10612 5778 10640 9454
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9140 4270 9260 4298
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 8772 2746 8984 2774
rect 8956 2514 8984 2746
rect 9140 2650 9168 4270
rect 9784 3738 9812 4762
rect 9968 4486 9996 5714
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10244 5302 10272 5578
rect 10232 5296 10284 5302
rect 10232 5238 10284 5244
rect 10612 5166 10640 5578
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 10796 3482 10824 9658
rect 10980 9586 11008 9930
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10888 8974 10916 9386
rect 10980 9110 11008 9522
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10980 8090 11008 9046
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10888 7342 10916 7686
rect 10980 7478 11008 8026
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 11072 5302 11100 14418
rect 11152 10736 11204 10742
rect 11150 10704 11152 10713
rect 11204 10704 11206 10713
rect 11150 10639 11206 10648
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11256 9674 11284 10542
rect 11348 9994 11376 23734
rect 11336 9988 11388 9994
rect 11336 9930 11388 9936
rect 11256 9646 11376 9674
rect 11150 9616 11206 9625
rect 11150 9551 11206 9560
rect 11164 9178 11192 9551
rect 11242 9480 11298 9489
rect 11242 9415 11298 9424
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11164 8566 11192 8910
rect 11152 8560 11204 8566
rect 11152 8502 11204 8508
rect 11256 6168 11284 9415
rect 11348 9042 11376 9646
rect 11440 9489 11468 23802
rect 11532 23730 11560 24006
rect 11520 23724 11572 23730
rect 11520 23666 11572 23672
rect 11532 23202 11560 23666
rect 11624 23526 11652 24006
rect 11612 23520 11664 23526
rect 11612 23462 11664 23468
rect 11532 23174 11652 23202
rect 11624 23118 11652 23174
rect 11612 23112 11664 23118
rect 11612 23054 11664 23060
rect 11520 23044 11572 23050
rect 11520 22986 11572 22992
rect 11532 21690 11560 22986
rect 11612 22976 11664 22982
rect 11612 22918 11664 22924
rect 11624 22642 11652 22918
rect 11612 22636 11664 22642
rect 11612 22578 11664 22584
rect 11704 22432 11756 22438
rect 11704 22374 11756 22380
rect 11716 22094 11744 22374
rect 11624 22066 11744 22094
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 11532 18358 11560 21626
rect 11624 21554 11652 22066
rect 11704 21616 11756 21622
rect 11704 21558 11756 21564
rect 11612 21548 11664 21554
rect 11612 21490 11664 21496
rect 11716 21457 11744 21558
rect 11702 21448 11758 21457
rect 11702 21383 11758 21392
rect 11704 21004 11756 21010
rect 11704 20946 11756 20952
rect 11612 20936 11664 20942
rect 11612 20878 11664 20884
rect 11624 20602 11652 20878
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 11624 19854 11652 20538
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11610 19680 11666 19689
rect 11610 19615 11666 19624
rect 11624 19446 11652 19615
rect 11612 19440 11664 19446
rect 11612 19382 11664 19388
rect 11716 19145 11744 20946
rect 11702 19136 11758 19145
rect 11702 19071 11758 19080
rect 11612 18964 11664 18970
rect 11612 18906 11664 18912
rect 11520 18352 11572 18358
rect 11520 18294 11572 18300
rect 11624 17542 11652 18906
rect 11716 18222 11744 19071
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11612 17536 11664 17542
rect 11612 17478 11664 17484
rect 11624 17134 11652 17478
rect 11716 17202 11744 18022
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11612 17128 11664 17134
rect 11612 17070 11664 17076
rect 11704 17060 11756 17066
rect 11704 17002 11756 17008
rect 11612 16720 11664 16726
rect 11612 16662 11664 16668
rect 11624 16250 11652 16662
rect 11716 16590 11744 17002
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11520 15360 11572 15366
rect 11520 15302 11572 15308
rect 11532 14793 11560 15302
rect 11518 14784 11574 14793
rect 11518 14719 11574 14728
rect 11624 14414 11652 15438
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11716 15201 11744 15302
rect 11702 15192 11758 15201
rect 11702 15127 11758 15136
rect 11704 15088 11756 15094
rect 11704 15030 11756 15036
rect 11716 14550 11744 15030
rect 11704 14544 11756 14550
rect 11704 14486 11756 14492
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11624 13938 11652 14350
rect 11808 14074 11836 27798
rect 11888 24744 11940 24750
rect 11888 24686 11940 24692
rect 11900 24410 11928 24686
rect 11888 24404 11940 24410
rect 11888 24346 11940 24352
rect 11980 24336 12032 24342
rect 11980 24278 12032 24284
rect 11992 23866 12020 24278
rect 11980 23860 12032 23866
rect 11980 23802 12032 23808
rect 11888 23656 11940 23662
rect 11888 23598 11940 23604
rect 11900 22574 11928 23598
rect 12084 22794 12112 29022
rect 12268 29034 12296 29174
rect 12162 28999 12218 29008
rect 12256 29028 12308 29034
rect 12256 28970 12308 28976
rect 12360 27470 12388 29174
rect 12348 27464 12400 27470
rect 12348 27406 12400 27412
rect 12256 26444 12308 26450
rect 12256 26386 12308 26392
rect 12268 26314 12296 26386
rect 12256 26308 12308 26314
rect 12256 26250 12308 26256
rect 12164 24676 12216 24682
rect 12164 24618 12216 24624
rect 12176 24410 12204 24618
rect 12164 24404 12216 24410
rect 12164 24346 12216 24352
rect 12360 24342 12388 27406
rect 12452 27130 12480 31418
rect 12820 31346 12848 32370
rect 12532 31340 12584 31346
rect 12532 31282 12584 31288
rect 12808 31340 12860 31346
rect 12808 31282 12860 31288
rect 12544 30870 12572 31282
rect 12716 31204 12768 31210
rect 12716 31146 12768 31152
rect 12532 30864 12584 30870
rect 12532 30806 12584 30812
rect 12728 30734 12756 31146
rect 12820 30734 12848 31282
rect 12716 30728 12768 30734
rect 12716 30670 12768 30676
rect 12808 30728 12860 30734
rect 12808 30670 12860 30676
rect 12532 30660 12584 30666
rect 12532 30602 12584 30608
rect 12544 30433 12572 30602
rect 12716 30592 12768 30598
rect 12716 30534 12768 30540
rect 12530 30424 12586 30433
rect 12530 30359 12586 30368
rect 12624 30048 12676 30054
rect 12624 29990 12676 29996
rect 12636 28218 12664 29990
rect 12728 29782 12756 30534
rect 12808 29844 12860 29850
rect 12808 29786 12860 29792
rect 12716 29776 12768 29782
rect 12716 29718 12768 29724
rect 12716 29572 12768 29578
rect 12716 29514 12768 29520
rect 12728 28558 12756 29514
rect 12820 29306 12848 29786
rect 12912 29646 12940 33510
rect 12992 31884 13044 31890
rect 12992 31826 13044 31832
rect 12900 29640 12952 29646
rect 12900 29582 12952 29588
rect 12900 29504 12952 29510
rect 12900 29446 12952 29452
rect 12808 29300 12860 29306
rect 12808 29242 12860 29248
rect 12808 29028 12860 29034
rect 12808 28970 12860 28976
rect 12716 28552 12768 28558
rect 12716 28494 12768 28500
rect 12820 28404 12848 28970
rect 12912 28490 12940 29446
rect 12900 28484 12952 28490
rect 12900 28426 12952 28432
rect 12728 28376 12848 28404
rect 12624 28212 12676 28218
rect 12624 28154 12676 28160
rect 12532 27940 12584 27946
rect 12532 27882 12584 27888
rect 12544 27470 12572 27882
rect 12728 27606 12756 28376
rect 12716 27600 12768 27606
rect 12716 27542 12768 27548
rect 12720 27526 12756 27542
rect 12532 27464 12584 27470
rect 12720 27452 12748 27526
rect 12912 27452 12940 28426
rect 12720 27424 12756 27452
rect 12532 27406 12584 27412
rect 12440 27124 12492 27130
rect 12440 27066 12492 27072
rect 12440 26444 12492 26450
rect 12440 26386 12492 26392
rect 12452 25294 12480 26386
rect 12440 25288 12492 25294
rect 12440 25230 12492 25236
rect 12728 24410 12756 27424
rect 12820 27424 12940 27452
rect 12820 26926 12848 27424
rect 13004 27062 13032 31826
rect 13096 27606 13124 37828
rect 13544 37188 13596 37194
rect 13544 37130 13596 37136
rect 13556 36106 13584 37130
rect 13544 36100 13596 36106
rect 13544 36042 13596 36048
rect 13360 35828 13412 35834
rect 13360 35770 13412 35776
rect 13176 35488 13228 35494
rect 13228 35448 13308 35476
rect 13176 35430 13228 35436
rect 13280 35154 13308 35448
rect 13372 35290 13400 35770
rect 13452 35760 13504 35766
rect 13452 35702 13504 35708
rect 13360 35284 13412 35290
rect 13360 35226 13412 35232
rect 13268 35148 13320 35154
rect 13268 35090 13320 35096
rect 13464 35086 13492 35702
rect 13452 35080 13504 35086
rect 13452 35022 13504 35028
rect 13464 34746 13492 35022
rect 13452 34740 13504 34746
rect 13452 34682 13504 34688
rect 13556 33590 13584 36042
rect 13924 35714 13952 38762
rect 14648 38752 14700 38758
rect 14648 38694 14700 38700
rect 14188 38344 14240 38350
rect 14188 38286 14240 38292
rect 14004 37936 14056 37942
rect 14004 37878 14056 37884
rect 14016 37806 14044 37878
rect 14004 37800 14056 37806
rect 14004 37742 14056 37748
rect 14016 36156 14044 37742
rect 14096 36780 14148 36786
rect 14096 36722 14148 36728
rect 14108 36378 14136 36722
rect 14200 36582 14228 38286
rect 14464 37324 14516 37330
rect 14464 37266 14516 37272
rect 14188 36576 14240 36582
rect 14188 36518 14240 36524
rect 14096 36372 14148 36378
rect 14096 36314 14148 36320
rect 14096 36168 14148 36174
rect 14016 36128 14096 36156
rect 14096 36110 14148 36116
rect 13924 35686 14044 35714
rect 13636 35556 13688 35562
rect 13636 35498 13688 35504
rect 13648 35018 13676 35498
rect 13636 35012 13688 35018
rect 13636 34954 13688 34960
rect 13648 34678 13676 34954
rect 13636 34672 13688 34678
rect 13636 34614 13688 34620
rect 13544 33584 13596 33590
rect 13544 33526 13596 33532
rect 13176 33516 13228 33522
rect 13176 33458 13228 33464
rect 13188 30870 13216 33458
rect 13544 32904 13596 32910
rect 13544 32846 13596 32852
rect 13268 32836 13320 32842
rect 13268 32778 13320 32784
rect 13280 32366 13308 32778
rect 13556 32434 13584 32846
rect 13544 32428 13596 32434
rect 13544 32370 13596 32376
rect 13268 32360 13320 32366
rect 13268 32302 13320 32308
rect 14016 31754 14044 35686
rect 14108 33998 14136 36110
rect 14200 35630 14228 36518
rect 14476 36174 14504 37266
rect 14556 36576 14608 36582
rect 14556 36518 14608 36524
rect 14464 36168 14516 36174
rect 14384 36128 14464 36156
rect 14188 35624 14240 35630
rect 14188 35566 14240 35572
rect 14200 34066 14228 35566
rect 14384 34746 14412 36128
rect 14464 36110 14516 36116
rect 14464 35624 14516 35630
rect 14464 35566 14516 35572
rect 14476 35290 14504 35566
rect 14464 35284 14516 35290
rect 14464 35226 14516 35232
rect 14568 35018 14596 36518
rect 14556 35012 14608 35018
rect 14556 34954 14608 34960
rect 14372 34740 14424 34746
rect 14372 34682 14424 34688
rect 14188 34060 14240 34066
rect 14188 34002 14240 34008
rect 14096 33992 14148 33998
rect 14096 33934 14148 33940
rect 13924 31726 14044 31754
rect 14108 31754 14136 33934
rect 14200 33658 14228 34002
rect 14384 33998 14412 34682
rect 14372 33992 14424 33998
rect 14372 33934 14424 33940
rect 14188 33652 14240 33658
rect 14188 33594 14240 33600
rect 14372 32768 14424 32774
rect 14372 32710 14424 32716
rect 14464 32768 14516 32774
rect 14464 32710 14516 32716
rect 14556 32768 14608 32774
rect 14556 32710 14608 32716
rect 14384 32298 14412 32710
rect 14372 32292 14424 32298
rect 14372 32234 14424 32240
rect 14108 31726 14228 31754
rect 13820 31680 13872 31686
rect 13820 31622 13872 31628
rect 13726 31512 13782 31521
rect 13544 31476 13596 31482
rect 13544 31418 13596 31424
rect 13648 31470 13726 31498
rect 13176 30864 13228 30870
rect 13176 30806 13228 30812
rect 13188 29714 13216 30806
rect 13452 30592 13504 30598
rect 13452 30534 13504 30540
rect 13464 30394 13492 30534
rect 13452 30388 13504 30394
rect 13452 30330 13504 30336
rect 13556 30326 13584 31418
rect 13648 31346 13676 31470
rect 13726 31447 13782 31456
rect 13832 31346 13860 31622
rect 13636 31340 13688 31346
rect 13636 31282 13688 31288
rect 13728 31340 13780 31346
rect 13728 31282 13780 31288
rect 13820 31340 13872 31346
rect 13820 31282 13872 31288
rect 13740 30938 13768 31282
rect 13820 31204 13872 31210
rect 13820 31146 13872 31152
rect 13832 31113 13860 31146
rect 13818 31104 13874 31113
rect 13818 31039 13874 31048
rect 13728 30932 13780 30938
rect 13728 30874 13780 30880
rect 13544 30320 13596 30326
rect 13544 30262 13596 30268
rect 13268 30252 13320 30258
rect 13268 30194 13320 30200
rect 13176 29708 13228 29714
rect 13176 29650 13228 29656
rect 13280 29646 13308 30194
rect 13360 29708 13412 29714
rect 13360 29650 13412 29656
rect 13268 29640 13320 29646
rect 13268 29582 13320 29588
rect 13280 28608 13308 29582
rect 13372 29238 13400 29650
rect 13452 29504 13504 29510
rect 13452 29446 13504 29452
rect 13464 29306 13492 29446
rect 13452 29300 13504 29306
rect 13452 29242 13504 29248
rect 13360 29232 13412 29238
rect 13360 29174 13412 29180
rect 13360 29096 13412 29102
rect 13556 29084 13584 30262
rect 13820 30252 13872 30258
rect 13820 30194 13872 30200
rect 13728 30116 13780 30122
rect 13728 30058 13780 30064
rect 13636 30048 13688 30054
rect 13636 29990 13688 29996
rect 13412 29056 13584 29084
rect 13360 29038 13412 29044
rect 13280 28580 13400 28608
rect 13176 28416 13228 28422
rect 13176 28358 13228 28364
rect 13188 28218 13216 28358
rect 13176 28212 13228 28218
rect 13176 28154 13228 28160
rect 13084 27600 13136 27606
rect 13084 27542 13136 27548
rect 13268 27396 13320 27402
rect 13268 27338 13320 27344
rect 13176 27328 13228 27334
rect 13176 27270 13228 27276
rect 12992 27056 13044 27062
rect 12992 26998 13044 27004
rect 12808 26920 12860 26926
rect 12808 26862 12860 26868
rect 12716 24404 12768 24410
rect 12716 24346 12768 24352
rect 12348 24336 12400 24342
rect 12348 24278 12400 24284
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12360 23798 12388 24142
rect 12348 23792 12400 23798
rect 12348 23734 12400 23740
rect 12164 23112 12216 23118
rect 12164 23054 12216 23060
rect 11992 22766 12112 22794
rect 11888 22568 11940 22574
rect 11888 22510 11940 22516
rect 11900 22166 11928 22510
rect 11888 22160 11940 22166
rect 11888 22102 11940 22108
rect 11900 21842 11928 22102
rect 11992 22094 12020 22766
rect 12176 22506 12204 23054
rect 12440 22976 12492 22982
rect 12440 22918 12492 22924
rect 12452 22710 12480 22918
rect 12440 22704 12492 22710
rect 12440 22646 12492 22652
rect 12164 22500 12216 22506
rect 12164 22442 12216 22448
rect 12256 22432 12308 22438
rect 12256 22374 12308 22380
rect 11992 22066 12112 22094
rect 11978 21992 12034 22001
rect 11978 21927 11980 21936
rect 12032 21927 12034 21936
rect 11980 21898 12032 21904
rect 11900 21814 12020 21842
rect 11992 21554 12020 21814
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 11980 21412 12032 21418
rect 11980 21354 12032 21360
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 11900 19514 11928 19790
rect 11888 19508 11940 19514
rect 11888 19450 11940 19456
rect 11992 19378 12020 21354
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11980 19372 12032 19378
rect 11980 19314 12032 19320
rect 11900 18766 11928 19314
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 11992 18970 12020 19110
rect 11980 18964 12032 18970
rect 11980 18906 12032 18912
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11900 17338 11928 18702
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 11900 17066 11928 17274
rect 11888 17060 11940 17066
rect 11888 17002 11940 17008
rect 11992 16454 12020 17478
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 11992 16250 12020 16390
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 12084 15706 12112 22066
rect 12268 21962 12296 22374
rect 12256 21956 12308 21962
rect 12256 21898 12308 21904
rect 12440 21956 12492 21962
rect 12440 21898 12492 21904
rect 12268 21554 12296 21898
rect 12256 21548 12308 21554
rect 12256 21490 12308 21496
rect 12268 20806 12296 21490
rect 12348 20868 12400 20874
rect 12348 20810 12400 20816
rect 12256 20800 12308 20806
rect 12360 20777 12388 20810
rect 12256 20742 12308 20748
rect 12346 20768 12402 20777
rect 12346 20703 12402 20712
rect 12452 20330 12480 21898
rect 12532 20460 12584 20466
rect 12532 20402 12584 20408
rect 12544 20330 12572 20402
rect 12164 20324 12216 20330
rect 12164 20266 12216 20272
rect 12440 20324 12492 20330
rect 12440 20266 12492 20272
rect 12532 20324 12584 20330
rect 12532 20266 12584 20272
rect 12176 17762 12204 20266
rect 12544 20210 12572 20266
rect 12452 20182 12572 20210
rect 12452 19281 12480 20182
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12438 19272 12494 19281
rect 12438 19207 12494 19216
rect 12544 19174 12572 19790
rect 12820 19334 12848 26862
rect 13188 26586 13216 27270
rect 13280 26586 13308 27338
rect 13176 26580 13228 26586
rect 13176 26522 13228 26528
rect 13268 26580 13320 26586
rect 13268 26522 13320 26528
rect 13372 25974 13400 28580
rect 13648 28082 13676 29990
rect 13740 29714 13768 30058
rect 13728 29708 13780 29714
rect 13728 29650 13780 29656
rect 13832 29102 13860 30194
rect 13820 29096 13872 29102
rect 13820 29038 13872 29044
rect 13832 28082 13860 29038
rect 13636 28076 13688 28082
rect 13636 28018 13688 28024
rect 13820 28076 13872 28082
rect 13820 28018 13872 28024
rect 13648 27062 13676 28018
rect 13636 27056 13688 27062
rect 13636 26998 13688 27004
rect 13360 25968 13412 25974
rect 13360 25910 13412 25916
rect 13176 25900 13228 25906
rect 13176 25842 13228 25848
rect 13544 25900 13596 25906
rect 13544 25842 13596 25848
rect 13188 25809 13216 25842
rect 13174 25800 13230 25809
rect 13174 25735 13230 25744
rect 12898 25392 12954 25401
rect 12898 25327 12900 25336
rect 12952 25327 12954 25336
rect 12900 25298 12952 25304
rect 13452 25220 13504 25226
rect 13452 25162 13504 25168
rect 13464 24206 13492 25162
rect 13556 24206 13584 25842
rect 13636 24744 13688 24750
rect 13636 24686 13688 24692
rect 13452 24200 13504 24206
rect 13452 24142 13504 24148
rect 13544 24200 13596 24206
rect 13544 24142 13596 24148
rect 13648 23798 13676 24686
rect 13820 24608 13872 24614
rect 13924 24585 13952 31726
rect 14096 31680 14148 31686
rect 14096 31622 14148 31628
rect 14108 31414 14136 31622
rect 14096 31408 14148 31414
rect 14096 31350 14148 31356
rect 14200 31226 14228 31726
rect 14280 31476 14332 31482
rect 14280 31418 14332 31424
rect 14108 31198 14228 31226
rect 14108 30258 14136 31198
rect 14292 30938 14320 31418
rect 14476 31328 14504 32710
rect 14568 31958 14596 32710
rect 14556 31952 14608 31958
rect 14556 31894 14608 31900
rect 14556 31340 14608 31346
rect 14476 31300 14556 31328
rect 14556 31282 14608 31288
rect 14280 30932 14332 30938
rect 14280 30874 14332 30880
rect 14096 30252 14148 30258
rect 14096 30194 14148 30200
rect 14188 29572 14240 29578
rect 14188 29514 14240 29520
rect 14200 29306 14228 29514
rect 14188 29300 14240 29306
rect 14188 29242 14240 29248
rect 14464 28076 14516 28082
rect 14464 28018 14516 28024
rect 14372 27464 14424 27470
rect 14372 27406 14424 27412
rect 14096 27396 14148 27402
rect 14096 27338 14148 27344
rect 14108 27062 14136 27338
rect 14188 27328 14240 27334
rect 14188 27270 14240 27276
rect 14096 27056 14148 27062
rect 14096 26998 14148 27004
rect 14108 26518 14136 26998
rect 14200 26926 14228 27270
rect 14188 26920 14240 26926
rect 14188 26862 14240 26868
rect 14096 26512 14148 26518
rect 14096 26454 14148 26460
rect 14188 25900 14240 25906
rect 14188 25842 14240 25848
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 14004 24812 14056 24818
rect 14004 24754 14056 24760
rect 13820 24550 13872 24556
rect 13910 24576 13966 24585
rect 13728 24268 13780 24274
rect 13728 24210 13780 24216
rect 13636 23792 13688 23798
rect 13636 23734 13688 23740
rect 13268 23724 13320 23730
rect 13268 23666 13320 23672
rect 13280 23254 13308 23666
rect 13268 23248 13320 23254
rect 13268 23190 13320 23196
rect 13740 23118 13768 24210
rect 13544 23112 13596 23118
rect 13544 23054 13596 23060
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 13556 22778 13584 23054
rect 13740 22778 13768 23054
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 13728 22772 13780 22778
rect 13728 22714 13780 22720
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 12912 21894 12940 22578
rect 13740 22234 13768 22714
rect 13728 22228 13780 22234
rect 13728 22170 13780 22176
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 13544 21888 13596 21894
rect 13544 21830 13596 21836
rect 13740 21842 13768 22170
rect 13832 21944 13860 24550
rect 13910 24511 13966 24520
rect 14016 23866 14044 24754
rect 14004 23860 14056 23866
rect 14004 23802 14056 23808
rect 13832 21916 13952 21944
rect 12912 21146 12940 21830
rect 13452 21616 13504 21622
rect 13452 21558 13504 21564
rect 12900 21140 12952 21146
rect 12900 21082 12952 21088
rect 13084 20460 13136 20466
rect 13084 20402 13136 20408
rect 13096 19854 13124 20402
rect 13176 20392 13228 20398
rect 13176 20334 13228 20340
rect 13188 19854 13216 20334
rect 13464 19990 13492 21558
rect 13556 21010 13584 21830
rect 13740 21814 13860 21842
rect 13728 21616 13780 21622
rect 13728 21558 13780 21564
rect 13636 21548 13688 21554
rect 13636 21490 13688 21496
rect 13648 21350 13676 21490
rect 13636 21344 13688 21350
rect 13636 21286 13688 21292
rect 13544 21004 13596 21010
rect 13544 20946 13596 20952
rect 13452 19984 13504 19990
rect 13452 19926 13504 19932
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 13176 19848 13228 19854
rect 13228 19808 13308 19836
rect 13176 19790 13228 19796
rect 12728 19306 12848 19334
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 12348 19168 12400 19174
rect 12348 19110 12400 19116
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12360 18834 12388 19110
rect 12348 18828 12400 18834
rect 12348 18770 12400 18776
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 12636 17762 12664 18702
rect 12176 17734 12296 17762
rect 12544 17746 12664 17762
rect 12268 17678 12296 17734
rect 12532 17740 12664 17746
rect 12584 17734 12664 17740
rect 12532 17682 12584 17688
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 12176 17338 12204 17614
rect 12268 17542 12296 17614
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12256 17264 12308 17270
rect 12256 17206 12308 17212
rect 12268 16590 12296 17206
rect 12360 16794 12388 17478
rect 12440 17264 12492 17270
rect 12440 17206 12492 17212
rect 12452 16998 12480 17206
rect 12636 17134 12664 17734
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 12360 16250 12388 16526
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12636 16182 12664 17070
rect 12624 16176 12676 16182
rect 12624 16118 12676 16124
rect 12440 15972 12492 15978
rect 12440 15914 12492 15920
rect 12452 15706 12480 15914
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12636 15502 12664 16118
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11980 15496 12032 15502
rect 12072 15496 12124 15502
rect 11980 15438 12032 15444
rect 12070 15464 12072 15473
rect 12624 15496 12676 15502
rect 12124 15464 12126 15473
rect 11900 15162 11928 15438
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11992 13938 12020 15438
rect 12624 15438 12676 15444
rect 12070 15399 12126 15408
rect 12256 15020 12308 15026
rect 12256 14962 12308 14968
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 12176 14482 12204 14758
rect 12268 14618 12296 14962
rect 12452 14618 12480 14962
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12532 14340 12584 14346
rect 12532 14282 12584 14288
rect 11612 13932 11664 13938
rect 11980 13932 12032 13938
rect 11612 13874 11664 13880
rect 11808 13892 11980 13920
rect 11520 11620 11572 11626
rect 11624 11608 11652 13874
rect 11572 11580 11652 11608
rect 11520 11562 11572 11568
rect 11532 10674 11560 11562
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11624 10742 11652 10950
rect 11612 10736 11664 10742
rect 11612 10678 11664 10684
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11532 9926 11560 10610
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11624 10198 11652 10406
rect 11612 10192 11664 10198
rect 11612 10134 11664 10140
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11532 9518 11560 9862
rect 11624 9722 11652 9930
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11520 9512 11572 9518
rect 11426 9480 11482 9489
rect 11520 9454 11572 9460
rect 11426 9415 11482 9424
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11348 8906 11468 8922
rect 11336 8900 11468 8906
rect 11388 8894 11468 8900
rect 11336 8842 11388 8848
rect 11440 8090 11468 8894
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11532 7426 11560 9318
rect 11716 9160 11744 11086
rect 11808 10810 11836 13892
rect 11980 13874 12032 13880
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12360 13530 12388 13874
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 11886 13424 11942 13433
rect 11886 13359 11942 13368
rect 11900 13326 11928 13359
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 12544 12986 12572 14282
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 11978 12880 12034 12889
rect 11978 12815 11980 12824
rect 12032 12815 12034 12824
rect 11980 12786 12032 12792
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 11992 11014 12020 12174
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12452 11830 12480 12038
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 12268 11098 12296 11494
rect 12544 11234 12572 12922
rect 12636 12850 12664 14350
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12636 11354 12664 11630
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12544 11206 12664 11234
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 12176 10810 12204 11086
rect 12268 11070 12480 11098
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11794 10568 11850 10577
rect 11794 10503 11850 10512
rect 11808 10470 11836 10503
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11808 9382 11836 10406
rect 11900 10198 11928 10610
rect 12360 10538 12388 10678
rect 12348 10532 12400 10538
rect 12348 10474 12400 10480
rect 11888 10192 11940 10198
rect 12452 10146 12480 11070
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 11888 10134 11940 10140
rect 12360 10118 12480 10146
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 11900 9722 11928 9862
rect 11888 9716 11940 9722
rect 11888 9658 11940 9664
rect 12176 9654 12204 9862
rect 12360 9674 12388 10118
rect 12164 9648 12216 9654
rect 12360 9646 12480 9674
rect 12164 9590 12216 9596
rect 11978 9480 12034 9489
rect 11978 9415 12034 9424
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11716 9132 11836 9160
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11624 7886 11652 8230
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11704 7880 11756 7886
rect 11808 7868 11836 9132
rect 11992 8956 12020 9415
rect 12348 9376 12400 9382
rect 12452 9353 12480 9646
rect 12348 9318 12400 9324
rect 12438 9344 12494 9353
rect 12070 9208 12126 9217
rect 12360 9178 12388 9318
rect 12438 9279 12494 9288
rect 12070 9143 12126 9152
rect 12348 9172 12400 9178
rect 12084 9042 12112 9143
rect 12348 9114 12400 9120
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 11756 7840 11836 7868
rect 11900 8928 12020 8956
rect 11704 7822 11756 7828
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11716 7546 11744 7686
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11796 7472 11848 7478
rect 11532 7398 11744 7426
rect 11900 7460 11928 8928
rect 12084 8566 12112 8978
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12360 8634 12388 8774
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12072 8560 12124 8566
rect 12072 8502 12124 8508
rect 12164 8356 12216 8362
rect 12164 8298 12216 8304
rect 12176 7970 12204 8298
rect 12176 7942 12296 7970
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 11848 7432 11928 7460
rect 11796 7414 11848 7420
rect 11336 6180 11388 6186
rect 11256 6140 11336 6168
rect 11336 6122 11388 6128
rect 11060 5296 11112 5302
rect 11060 5238 11112 5244
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 11072 4010 11100 4966
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 10966 3496 11022 3505
rect 9496 3460 9548 3466
rect 9496 3402 9548 3408
rect 9588 3460 9640 3466
rect 10796 3454 10966 3482
rect 10966 3431 11022 3440
rect 11244 3460 11296 3466
rect 9588 3402 9640 3408
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 9232 3194 9260 3334
rect 9508 3194 9536 3402
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9600 3126 9628 3402
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 10980 2990 11008 3431
rect 11244 3402 11296 3408
rect 11256 2990 11284 3402
rect 11348 3040 11376 6122
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 11440 4214 11468 5102
rect 11428 4208 11480 4214
rect 11428 4150 11480 4156
rect 11440 3534 11468 4150
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 11532 3380 11560 5714
rect 11610 3904 11666 3913
rect 11610 3839 11666 3848
rect 11624 3534 11652 3839
rect 11716 3534 11744 7398
rect 11992 7274 12020 7822
rect 12176 7546 12204 7822
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 11980 7268 12032 7274
rect 11980 7210 12032 7216
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11808 6458 11836 6598
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11900 5914 11928 6190
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 12268 5778 12296 7942
rect 12348 7812 12400 7818
rect 12348 7754 12400 7760
rect 12360 7274 12388 7754
rect 12544 7546 12572 10950
rect 12636 10674 12664 11206
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12636 10305 12664 10610
rect 12622 10296 12678 10305
rect 12622 10231 12678 10240
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12348 7268 12400 7274
rect 12348 7210 12400 7216
rect 12544 6662 12572 7482
rect 12636 7478 12664 9998
rect 12624 7472 12676 7478
rect 12624 7414 12676 7420
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12256 5772 12308 5778
rect 12256 5714 12308 5720
rect 12268 5302 12296 5714
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 11532 3352 11652 3380
rect 11624 3058 11652 3352
rect 11808 3058 11836 4218
rect 11900 3058 11928 5170
rect 12360 4146 12388 6598
rect 12636 5710 12664 7414
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12636 4758 12664 5102
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12728 4282 12756 19306
rect 12912 18834 12940 19314
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12820 17377 12848 18702
rect 12806 17368 12862 17377
rect 12806 17303 12808 17312
rect 12860 17303 12862 17312
rect 12808 17274 12860 17280
rect 13096 17270 13124 19790
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 13188 18766 13216 19314
rect 13176 18760 13228 18766
rect 13176 18702 13228 18708
rect 13188 18426 13216 18702
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 13174 18320 13230 18329
rect 13174 18255 13230 18264
rect 13084 17264 13136 17270
rect 13084 17206 13136 17212
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12912 15706 12940 15846
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 13004 15570 13032 16050
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 12820 13394 12848 14962
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12912 13190 12940 14894
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12820 10810 12848 12786
rect 12912 11354 12940 13126
rect 13004 12170 13032 13126
rect 13096 12986 13124 13466
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 12992 11824 13044 11830
rect 12992 11766 13044 11772
rect 13004 11694 13032 11766
rect 12992 11688 13044 11694
rect 12992 11630 13044 11636
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12820 7342 12848 10746
rect 12900 10736 12952 10742
rect 12900 10678 12952 10684
rect 12912 10266 12940 10678
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 13004 9518 13032 11630
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 13096 11218 13124 11494
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 13096 10266 13124 10474
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 13082 10160 13138 10169
rect 13082 10095 13138 10104
rect 12992 9512 13044 9518
rect 12912 9472 12992 9500
rect 12912 9110 12940 9472
rect 12992 9454 13044 9460
rect 12900 9104 12952 9110
rect 12900 9046 12952 9052
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 13004 8974 13032 9046
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12912 7954 12940 8774
rect 13096 8362 13124 10095
rect 13084 8356 13136 8362
rect 13084 8298 13136 8304
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12820 5166 12848 5510
rect 13188 5302 13216 18255
rect 13280 16114 13308 19808
rect 13464 19378 13492 19926
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 13556 18902 13584 20946
rect 13740 19446 13768 21558
rect 13832 21554 13860 21814
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13820 21412 13872 21418
rect 13820 21354 13872 21360
rect 13832 21146 13860 21354
rect 13820 21140 13872 21146
rect 13820 21082 13872 21088
rect 13924 20584 13952 21916
rect 14004 21344 14056 21350
rect 14004 21286 14056 21292
rect 14016 21078 14044 21286
rect 14004 21072 14056 21078
rect 14004 21014 14056 21020
rect 13832 20556 13952 20584
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 13740 19122 13768 19382
rect 13648 19094 13768 19122
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 13648 18766 13676 19094
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 13636 18760 13688 18766
rect 13636 18702 13688 18708
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 13372 16114 13400 18566
rect 13452 17604 13504 17610
rect 13452 17546 13504 17552
rect 13464 16590 13492 17546
rect 13542 17096 13598 17105
rect 13542 17031 13544 17040
rect 13596 17031 13598 17040
rect 13544 17002 13596 17008
rect 13556 16590 13584 17002
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13372 15638 13400 16050
rect 13648 15910 13676 18702
rect 13740 17882 13768 18906
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13740 17678 13768 17818
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13360 15632 13412 15638
rect 13360 15574 13412 15580
rect 13636 15632 13688 15638
rect 13636 15574 13688 15580
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13280 13326 13308 13466
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13372 12918 13400 13670
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13372 10713 13400 12038
rect 13464 11150 13492 13262
rect 13544 13252 13596 13258
rect 13544 13194 13596 13200
rect 13556 12986 13584 13194
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13648 11801 13676 15574
rect 13832 12434 13860 20556
rect 13912 20460 13964 20466
rect 13912 20402 13964 20408
rect 13924 20058 13952 20402
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 13912 19168 13964 19174
rect 13912 19110 13964 19116
rect 13924 18970 13952 19110
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13924 18426 13952 18566
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 14108 18057 14136 25094
rect 14200 24818 14228 25842
rect 14280 25288 14332 25294
rect 14280 25230 14332 25236
rect 14292 24954 14320 25230
rect 14280 24948 14332 24954
rect 14280 24890 14332 24896
rect 14188 24812 14240 24818
rect 14188 24754 14240 24760
rect 14200 23730 14228 24754
rect 14384 24274 14412 27406
rect 14476 25922 14504 28018
rect 14660 26042 14688 38694
rect 14752 34202 14780 38898
rect 14832 38888 14884 38894
rect 14832 38830 14884 38836
rect 14844 36378 14872 38830
rect 17604 38282 17632 39034
rect 20732 39030 20760 39086
rect 23204 39092 23256 39098
rect 23204 39034 23256 39040
rect 25136 39092 25188 39098
rect 25136 39034 25188 39040
rect 27344 39092 27396 39098
rect 31588 39092 31904 39098
rect 31588 39086 31852 39092
rect 27344 39034 27396 39040
rect 31852 39034 31904 39040
rect 34152 39092 34204 39098
rect 34152 39034 34204 39040
rect 36360 39092 36412 39098
rect 36360 39034 36412 39040
rect 37200 39030 37228 40151
rect 20720 39024 20772 39030
rect 20720 38966 20772 38972
rect 23940 39024 23992 39030
rect 23940 38966 23992 38972
rect 37188 39024 37240 39030
rect 37188 38966 37240 38972
rect 17776 38956 17828 38962
rect 17776 38898 17828 38904
rect 23388 38956 23440 38962
rect 23388 38898 23440 38904
rect 15292 38276 15344 38282
rect 15292 38218 15344 38224
rect 15844 38276 15896 38282
rect 15844 38218 15896 38224
rect 17592 38276 17644 38282
rect 17592 38218 17644 38224
rect 15304 38010 15332 38218
rect 15292 38004 15344 38010
rect 15292 37946 15344 37952
rect 15856 36786 15884 38218
rect 16764 38208 16816 38214
rect 16764 38150 16816 38156
rect 16776 38010 16804 38150
rect 17788 38010 17816 38898
rect 19432 38548 19484 38554
rect 19432 38490 19484 38496
rect 21088 38548 21140 38554
rect 21088 38490 21140 38496
rect 17960 38412 18012 38418
rect 17960 38354 18012 38360
rect 16396 38004 16448 38010
rect 16396 37946 16448 37952
rect 16764 38004 16816 38010
rect 16764 37946 16816 37952
rect 17776 38004 17828 38010
rect 17776 37946 17828 37952
rect 16408 37874 16436 37946
rect 16120 37868 16172 37874
rect 16120 37810 16172 37816
rect 16212 37868 16264 37874
rect 16212 37810 16264 37816
rect 16304 37868 16356 37874
rect 16304 37810 16356 37816
rect 16396 37868 16448 37874
rect 16396 37810 16448 37816
rect 16132 37466 16160 37810
rect 16120 37460 16172 37466
rect 16120 37402 16172 37408
rect 16224 37346 16252 37810
rect 16316 37466 16344 37810
rect 16304 37460 16356 37466
rect 16304 37402 16356 37408
rect 16132 37330 16252 37346
rect 16120 37324 16252 37330
rect 16172 37318 16252 37324
rect 16120 37266 16172 37272
rect 16776 37262 16804 37946
rect 17684 37936 17736 37942
rect 17684 37878 17736 37884
rect 17132 37800 17184 37806
rect 17132 37742 17184 37748
rect 17316 37800 17368 37806
rect 17316 37742 17368 37748
rect 16304 37256 16356 37262
rect 16304 37198 16356 37204
rect 16764 37256 16816 37262
rect 16764 37198 16816 37204
rect 15844 36780 15896 36786
rect 15844 36722 15896 36728
rect 14832 36372 14884 36378
rect 14832 36314 14884 36320
rect 15384 36236 15436 36242
rect 15384 36178 15436 36184
rect 15200 36168 15252 36174
rect 15200 36110 15252 36116
rect 14924 36032 14976 36038
rect 14924 35974 14976 35980
rect 14936 35086 14964 35974
rect 14924 35080 14976 35086
rect 14924 35022 14976 35028
rect 15212 34406 15240 36110
rect 15396 35290 15424 36178
rect 15752 36168 15804 36174
rect 15752 36110 15804 36116
rect 15764 35494 15792 36110
rect 15856 35766 15884 36722
rect 16316 36174 16344 37198
rect 17144 36378 17172 37742
rect 17132 36372 17184 36378
rect 17132 36314 17184 36320
rect 17328 36310 17356 37742
rect 17316 36304 17368 36310
rect 17316 36246 17368 36252
rect 16580 36236 16632 36242
rect 16580 36178 16632 36184
rect 16304 36168 16356 36174
rect 16304 36110 16356 36116
rect 15844 35760 15896 35766
rect 16316 35748 16344 36110
rect 16592 35834 16620 36178
rect 16764 36168 16816 36174
rect 16764 36110 16816 36116
rect 16580 35828 16632 35834
rect 16580 35770 16632 35776
rect 16396 35760 16448 35766
rect 16316 35720 16396 35748
rect 15844 35702 15896 35708
rect 16396 35702 16448 35708
rect 15752 35488 15804 35494
rect 15752 35430 15804 35436
rect 15384 35284 15436 35290
rect 15384 35226 15436 35232
rect 15292 35012 15344 35018
rect 15292 34954 15344 34960
rect 15304 34610 15332 34954
rect 15292 34604 15344 34610
rect 15292 34546 15344 34552
rect 15200 34400 15252 34406
rect 15200 34342 15252 34348
rect 14740 34196 14792 34202
rect 14740 34138 14792 34144
rect 15108 33924 15160 33930
rect 15108 33866 15160 33872
rect 14832 33516 14884 33522
rect 14832 33458 14884 33464
rect 15016 33516 15068 33522
rect 15016 33458 15068 33464
rect 14844 33046 14872 33458
rect 15028 33046 15056 33458
rect 14832 33040 14884 33046
rect 14832 32982 14884 32988
rect 15016 33040 15068 33046
rect 15016 32982 15068 32988
rect 14832 31816 14884 31822
rect 14832 31758 14884 31764
rect 14844 31346 14872 31758
rect 14832 31340 14884 31346
rect 14832 31282 14884 31288
rect 15016 31340 15068 31346
rect 15016 31282 15068 31288
rect 14830 31240 14886 31249
rect 14830 31175 14832 31184
rect 14884 31175 14886 31184
rect 14832 31146 14884 31152
rect 15028 30802 15056 31282
rect 15016 30796 15068 30802
rect 15016 30738 15068 30744
rect 15120 29782 15148 33866
rect 15200 33312 15252 33318
rect 15200 33254 15252 33260
rect 15212 32910 15240 33254
rect 15200 32904 15252 32910
rect 15200 32846 15252 32852
rect 15304 31754 15332 34546
rect 15384 33992 15436 33998
rect 15384 33934 15436 33940
rect 15476 33992 15528 33998
rect 15476 33934 15528 33940
rect 15396 33658 15424 33934
rect 15384 33652 15436 33658
rect 15384 33594 15436 33600
rect 15384 33312 15436 33318
rect 15384 33254 15436 33260
rect 15396 32756 15424 33254
rect 15488 32910 15516 33934
rect 15660 33924 15712 33930
rect 15660 33866 15712 33872
rect 15672 33658 15700 33866
rect 15660 33652 15712 33658
rect 15660 33594 15712 33600
rect 15476 32904 15528 32910
rect 15476 32846 15528 32852
rect 15396 32728 15516 32756
rect 15304 31726 15424 31754
rect 15292 31680 15344 31686
rect 15292 31622 15344 31628
rect 15304 31210 15332 31622
rect 15292 31204 15344 31210
rect 15292 31146 15344 31152
rect 15200 31136 15252 31142
rect 15198 31104 15200 31113
rect 15252 31104 15254 31113
rect 15198 31039 15254 31048
rect 15396 30274 15424 31726
rect 15488 31686 15516 32728
rect 15476 31680 15528 31686
rect 15476 31622 15528 31628
rect 15304 30246 15424 30274
rect 15108 29776 15160 29782
rect 15160 29736 15240 29764
rect 15108 29718 15160 29724
rect 15108 29028 15160 29034
rect 15108 28970 15160 28976
rect 15120 28558 15148 28970
rect 15108 28552 15160 28558
rect 15108 28494 15160 28500
rect 15016 28008 15068 28014
rect 15016 27950 15068 27956
rect 15028 27674 15056 27950
rect 15016 27668 15068 27674
rect 15016 27610 15068 27616
rect 14832 27600 14884 27606
rect 14832 27542 14884 27548
rect 14844 27470 14872 27542
rect 14832 27464 14884 27470
rect 14832 27406 14884 27412
rect 14648 26036 14700 26042
rect 14648 25978 14700 25984
rect 14844 25974 14872 27406
rect 14924 26784 14976 26790
rect 14924 26726 14976 26732
rect 14936 26353 14964 26726
rect 15028 26382 15056 27610
rect 15212 26450 15240 29736
rect 15200 26444 15252 26450
rect 15200 26386 15252 26392
rect 15016 26376 15068 26382
rect 14922 26344 14978 26353
rect 15016 26318 15068 26324
rect 14922 26279 14978 26288
rect 14832 25968 14884 25974
rect 14554 25936 14610 25945
rect 14476 25906 14554 25922
rect 14464 25900 14554 25906
rect 14516 25894 14554 25900
rect 14832 25910 14884 25916
rect 14740 25900 14792 25906
rect 14554 25871 14610 25880
rect 14464 25842 14516 25848
rect 14660 25860 14740 25888
rect 14556 25696 14608 25702
rect 14556 25638 14608 25644
rect 14372 24268 14424 24274
rect 14372 24210 14424 24216
rect 14188 23724 14240 23730
rect 14188 23666 14240 23672
rect 14568 23497 14596 25638
rect 14660 24886 14688 25860
rect 14740 25842 14792 25848
rect 14740 25696 14792 25702
rect 14740 25638 14792 25644
rect 14752 25498 14780 25638
rect 14844 25498 14872 25910
rect 14740 25492 14792 25498
rect 14740 25434 14792 25440
rect 14832 25492 14884 25498
rect 14832 25434 14884 25440
rect 14924 25492 14976 25498
rect 14924 25434 14976 25440
rect 14740 25356 14792 25362
rect 14740 25298 14792 25304
rect 14648 24880 14700 24886
rect 14648 24822 14700 24828
rect 14752 24274 14780 25298
rect 14936 24954 14964 25434
rect 15028 25294 15056 26318
rect 15108 25764 15160 25770
rect 15108 25706 15160 25712
rect 15016 25288 15068 25294
rect 15016 25230 15068 25236
rect 14924 24948 14976 24954
rect 14924 24890 14976 24896
rect 14832 24812 14884 24818
rect 14936 24800 14964 24890
rect 14884 24772 14964 24800
rect 14832 24754 14884 24760
rect 15120 24721 15148 25706
rect 15304 25702 15332 30246
rect 15384 28416 15436 28422
rect 15384 28358 15436 28364
rect 15396 28218 15424 28358
rect 15384 28212 15436 28218
rect 15384 28154 15436 28160
rect 15384 27328 15436 27334
rect 15384 27270 15436 27276
rect 15396 26994 15424 27270
rect 15384 26988 15436 26994
rect 15384 26930 15436 26936
rect 15292 25696 15344 25702
rect 15292 25638 15344 25644
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15106 24712 15162 24721
rect 15106 24647 15162 24656
rect 15016 24608 15068 24614
rect 15016 24550 15068 24556
rect 15106 24576 15162 24585
rect 14740 24268 14792 24274
rect 14740 24210 14792 24216
rect 14648 24132 14700 24138
rect 14648 24074 14700 24080
rect 14660 23730 14688 24074
rect 14648 23724 14700 23730
rect 14648 23666 14700 23672
rect 14554 23488 14610 23497
rect 14554 23423 14610 23432
rect 14372 23248 14424 23254
rect 14372 23190 14424 23196
rect 14384 22642 14412 23190
rect 14464 23112 14516 23118
rect 14464 23054 14516 23060
rect 14372 22636 14424 22642
rect 14372 22578 14424 22584
rect 14188 22500 14240 22506
rect 14188 22442 14240 22448
rect 14200 21554 14228 22442
rect 14372 21956 14424 21962
rect 14372 21898 14424 21904
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 14384 20942 14412 21898
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14292 19145 14320 19994
rect 14384 19854 14412 20878
rect 14372 19848 14424 19854
rect 14372 19790 14424 19796
rect 14384 19689 14412 19790
rect 14370 19680 14426 19689
rect 14370 19615 14426 19624
rect 14372 19168 14424 19174
rect 14278 19136 14334 19145
rect 14372 19110 14424 19116
rect 14278 19071 14334 19080
rect 14188 18692 14240 18698
rect 14188 18634 14240 18640
rect 14094 18048 14150 18057
rect 14094 17983 14150 17992
rect 14096 17876 14148 17882
rect 14096 17818 14148 17824
rect 14004 17264 14056 17270
rect 14004 17206 14056 17212
rect 13912 16448 13964 16454
rect 13912 16390 13964 16396
rect 13924 16114 13952 16390
rect 14016 16250 14044 17206
rect 14108 17202 14136 17818
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 14004 16244 14056 16250
rect 14004 16186 14056 16192
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 14200 16046 14228 18634
rect 14292 18290 14320 19071
rect 14384 18766 14412 19110
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14476 18290 14504 23054
rect 14556 22636 14608 22642
rect 14556 22578 14608 22584
rect 14568 21457 14596 22578
rect 14554 21448 14610 21457
rect 14554 21383 14610 21392
rect 14568 19514 14596 21383
rect 14660 21350 14688 23666
rect 14924 23112 14976 23118
rect 14924 23054 14976 23060
rect 14936 22642 14964 23054
rect 14924 22636 14976 22642
rect 14924 22578 14976 22584
rect 14740 22500 14792 22506
rect 14740 22442 14792 22448
rect 14924 22500 14976 22506
rect 14924 22442 14976 22448
rect 14648 21344 14700 21350
rect 14648 21286 14700 21292
rect 14660 20942 14688 21286
rect 14648 20936 14700 20942
rect 14648 20878 14700 20884
rect 14648 19712 14700 19718
rect 14646 19680 14648 19689
rect 14752 19700 14780 22442
rect 14936 22166 14964 22442
rect 14924 22160 14976 22166
rect 14924 22102 14976 22108
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14844 21690 14872 21830
rect 14832 21684 14884 21690
rect 14832 21626 14884 21632
rect 14844 21457 14872 21626
rect 14936 21554 14964 22102
rect 14924 21548 14976 21554
rect 14924 21490 14976 21496
rect 14830 21448 14886 21457
rect 14830 21383 14886 21392
rect 14844 20874 14872 21383
rect 14832 20868 14884 20874
rect 14832 20810 14884 20816
rect 14700 19680 14780 19700
rect 14702 19672 14780 19680
rect 14832 19712 14884 19718
rect 14832 19654 14884 19660
rect 14646 19615 14702 19624
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14556 19304 14608 19310
rect 14556 19246 14608 19252
rect 14568 18630 14596 19246
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 14556 18624 14608 18630
rect 14556 18566 14608 18572
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14464 17196 14516 17202
rect 14568 17184 14596 18566
rect 14752 18154 14780 19110
rect 14740 18148 14792 18154
rect 14740 18090 14792 18096
rect 14648 18080 14700 18086
rect 14648 18022 14700 18028
rect 14660 17338 14688 18022
rect 14844 17678 14872 19654
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 14752 17338 14780 17614
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14516 17156 14596 17184
rect 14464 17138 14516 17144
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14370 16960 14426 16969
rect 14292 16250 14320 16934
rect 14370 16895 14426 16904
rect 14384 16590 14412 16895
rect 14476 16590 14504 17138
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14464 16584 14516 16590
rect 14464 16526 14516 16532
rect 14660 16522 14688 17274
rect 14844 17202 14872 17614
rect 14936 17270 14964 21490
rect 15028 19242 15056 24550
rect 15212 24562 15240 24754
rect 15162 24534 15240 24562
rect 15106 24511 15162 24520
rect 15384 24200 15436 24206
rect 15382 24168 15384 24177
rect 15436 24168 15438 24177
rect 15382 24103 15438 24112
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 15200 23112 15252 23118
rect 15200 23054 15252 23060
rect 15120 22506 15148 23054
rect 15108 22500 15160 22506
rect 15108 22442 15160 22448
rect 15108 21888 15160 21894
rect 15108 21830 15160 21836
rect 15120 21418 15148 21830
rect 15108 21412 15160 21418
rect 15108 21354 15160 21360
rect 15120 19854 15148 21354
rect 15212 20534 15240 23054
rect 15384 21956 15436 21962
rect 15384 21898 15436 21904
rect 15292 21548 15344 21554
rect 15292 21490 15344 21496
rect 15304 20942 15332 21490
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 15200 20528 15252 20534
rect 15200 20470 15252 20476
rect 15108 19848 15160 19854
rect 15108 19790 15160 19796
rect 15120 19514 15148 19790
rect 15108 19508 15160 19514
rect 15108 19450 15160 19456
rect 15292 19372 15344 19378
rect 15396 19360 15424 21898
rect 15488 20874 15516 31622
rect 15566 31512 15622 31521
rect 15566 31447 15568 31456
rect 15620 31447 15622 31456
rect 15568 31418 15620 31424
rect 15580 30433 15608 31418
rect 15566 30424 15622 30433
rect 15566 30359 15622 30368
rect 15660 30048 15712 30054
rect 15660 29990 15712 29996
rect 15672 29714 15700 29990
rect 15660 29708 15712 29714
rect 15660 29650 15712 29656
rect 15568 29504 15620 29510
rect 15568 29446 15620 29452
rect 15580 26586 15608 29446
rect 15672 27470 15700 29650
rect 15660 27464 15712 27470
rect 15660 27406 15712 27412
rect 15764 27130 15792 35430
rect 15856 35154 15884 35702
rect 16118 35592 16174 35601
rect 16118 35527 16174 35536
rect 16132 35494 16160 35527
rect 16120 35488 16172 35494
rect 16120 35430 16172 35436
rect 16488 35488 16540 35494
rect 16488 35430 16540 35436
rect 15844 35148 15896 35154
rect 15844 35090 15896 35096
rect 16132 34610 16160 35430
rect 16500 35068 16528 35430
rect 16776 35222 16804 36110
rect 17132 36032 17184 36038
rect 17132 35974 17184 35980
rect 16856 35624 16908 35630
rect 16856 35566 16908 35572
rect 16868 35290 16896 35566
rect 16856 35284 16908 35290
rect 16856 35226 16908 35232
rect 16764 35216 16816 35222
rect 16764 35158 16816 35164
rect 16776 35086 16804 35158
rect 16580 35080 16632 35086
rect 16500 35040 16580 35068
rect 16580 35022 16632 35028
rect 16764 35080 16816 35086
rect 16764 35022 16816 35028
rect 16672 35012 16724 35018
rect 16672 34954 16724 34960
rect 16856 35012 16908 35018
rect 16856 34954 16908 34960
rect 16684 34746 16712 34954
rect 16672 34740 16724 34746
rect 16672 34682 16724 34688
rect 16120 34604 16172 34610
rect 16120 34546 16172 34552
rect 16868 34474 16896 34954
rect 16856 34468 16908 34474
rect 16856 34410 16908 34416
rect 15936 33924 15988 33930
rect 15936 33866 15988 33872
rect 15948 33522 15976 33866
rect 17144 33658 17172 35974
rect 17696 35630 17724 37878
rect 17972 36786 18000 38354
rect 19444 38282 19472 38490
rect 21100 38350 21128 38490
rect 23204 38480 23256 38486
rect 23204 38422 23256 38428
rect 23216 38350 23244 38422
rect 21088 38344 21140 38350
rect 21088 38286 21140 38292
rect 23204 38344 23256 38350
rect 23204 38286 23256 38292
rect 19432 38276 19484 38282
rect 19432 38218 19484 38224
rect 19984 38276 20036 38282
rect 19984 38218 20036 38224
rect 22100 38276 22152 38282
rect 22100 38218 22152 38224
rect 19064 38208 19116 38214
rect 19064 38150 19116 38156
rect 19076 38010 19104 38150
rect 19064 38004 19116 38010
rect 19064 37946 19116 37952
rect 18052 37800 18104 37806
rect 18052 37742 18104 37748
rect 17960 36780 18012 36786
rect 17960 36722 18012 36728
rect 18064 35834 18092 37742
rect 19076 37126 19104 37946
rect 19340 37188 19392 37194
rect 19340 37130 19392 37136
rect 19064 37120 19116 37126
rect 19064 37062 19116 37068
rect 18420 36712 18472 36718
rect 18420 36654 18472 36660
rect 18432 36378 18460 36654
rect 18420 36372 18472 36378
rect 18420 36314 18472 36320
rect 18788 36236 18840 36242
rect 18788 36178 18840 36184
rect 18052 35828 18104 35834
rect 18052 35770 18104 35776
rect 18052 35692 18104 35698
rect 18052 35634 18104 35640
rect 17684 35624 17736 35630
rect 17684 35566 17736 35572
rect 17696 35494 17724 35566
rect 17868 35556 17920 35562
rect 17868 35498 17920 35504
rect 17684 35488 17736 35494
rect 17684 35430 17736 35436
rect 17880 35290 17908 35498
rect 18064 35290 18092 35634
rect 18800 35630 18828 36178
rect 19352 36009 19380 37130
rect 19444 36854 19472 38218
rect 19996 38010 20024 38218
rect 20720 38208 20772 38214
rect 20720 38150 20772 38156
rect 21456 38208 21508 38214
rect 21456 38150 21508 38156
rect 20732 38010 20760 38150
rect 19984 38004 20036 38010
rect 19984 37946 20036 37952
rect 20720 38004 20772 38010
rect 20720 37946 20772 37952
rect 19800 37800 19852 37806
rect 19800 37742 19852 37748
rect 20812 37800 20864 37806
rect 20812 37742 20864 37748
rect 19432 36848 19484 36854
rect 19432 36790 19484 36796
rect 19338 36000 19394 36009
rect 19338 35935 19394 35944
rect 18880 35692 18932 35698
rect 18880 35634 18932 35640
rect 18788 35624 18840 35630
rect 18788 35566 18840 35572
rect 18144 35488 18196 35494
rect 18144 35430 18196 35436
rect 17868 35284 17920 35290
rect 17868 35226 17920 35232
rect 18052 35284 18104 35290
rect 18052 35226 18104 35232
rect 17880 35086 17908 35226
rect 18156 35086 18184 35430
rect 18800 35222 18828 35566
rect 18788 35216 18840 35222
rect 18788 35158 18840 35164
rect 17868 35080 17920 35086
rect 17868 35022 17920 35028
rect 18144 35080 18196 35086
rect 18144 35022 18196 35028
rect 18236 35080 18288 35086
rect 18236 35022 18288 35028
rect 17868 34944 17920 34950
rect 17868 34886 17920 34892
rect 17880 34202 17908 34886
rect 18248 34678 18276 35022
rect 18236 34672 18288 34678
rect 18236 34614 18288 34620
rect 18236 34400 18288 34406
rect 18236 34342 18288 34348
rect 17868 34196 17920 34202
rect 17868 34138 17920 34144
rect 17880 33862 17908 34138
rect 18144 33992 18196 33998
rect 18144 33934 18196 33940
rect 17408 33856 17460 33862
rect 17408 33798 17460 33804
rect 17776 33856 17828 33862
rect 17776 33798 17828 33804
rect 17868 33856 17920 33862
rect 17868 33798 17920 33804
rect 17132 33652 17184 33658
rect 17132 33594 17184 33600
rect 15936 33516 15988 33522
rect 15936 33458 15988 33464
rect 16028 33516 16080 33522
rect 16028 33458 16080 33464
rect 15948 32892 15976 33458
rect 16040 33114 16068 33458
rect 17420 33454 17448 33798
rect 17684 33516 17736 33522
rect 17684 33458 17736 33464
rect 17408 33448 17460 33454
rect 17408 33390 17460 33396
rect 16028 33108 16080 33114
rect 16028 33050 16080 33056
rect 16304 32972 16356 32978
rect 16304 32914 16356 32920
rect 17040 32972 17092 32978
rect 17040 32914 17092 32920
rect 15948 32864 16160 32892
rect 15936 32768 15988 32774
rect 15936 32710 15988 32716
rect 16028 32768 16080 32774
rect 16028 32710 16080 32716
rect 15948 31754 15976 32710
rect 16040 32366 16068 32710
rect 16028 32360 16080 32366
rect 16028 32302 16080 32308
rect 15856 31726 15976 31754
rect 15856 31346 15884 31726
rect 16040 31396 16068 32302
rect 16132 31822 16160 32864
rect 16316 32774 16344 32914
rect 16304 32768 16356 32774
rect 16304 32710 16356 32716
rect 16488 32768 16540 32774
rect 16488 32710 16540 32716
rect 16500 31890 16528 32710
rect 16488 31884 16540 31890
rect 16488 31826 16540 31832
rect 16120 31816 16172 31822
rect 16120 31758 16172 31764
rect 16212 31816 16264 31822
rect 16212 31758 16264 31764
rect 15948 31368 16068 31396
rect 15844 31340 15896 31346
rect 15844 31282 15896 31288
rect 15948 31226 15976 31368
rect 16132 31328 16160 31758
rect 15856 31198 15976 31226
rect 16040 31300 16160 31328
rect 15856 29782 15884 31198
rect 16040 31142 16068 31300
rect 16224 31226 16252 31758
rect 16396 31680 16448 31686
rect 16396 31622 16448 31628
rect 16580 31680 16632 31686
rect 16580 31622 16632 31628
rect 16408 31482 16436 31622
rect 16396 31476 16448 31482
rect 16396 31418 16448 31424
rect 16592 31346 16620 31622
rect 17052 31346 17080 32914
rect 17420 32774 17448 33390
rect 17500 33108 17552 33114
rect 17500 33050 17552 33056
rect 17408 32768 17460 32774
rect 17408 32710 17460 32716
rect 17316 32564 17368 32570
rect 17316 32506 17368 32512
rect 16580 31340 16632 31346
rect 16580 31282 16632 31288
rect 16672 31340 16724 31346
rect 16672 31282 16724 31288
rect 17040 31340 17092 31346
rect 17040 31282 17092 31288
rect 16132 31198 16252 31226
rect 16304 31272 16356 31278
rect 16684 31249 16712 31282
rect 16304 31214 16356 31220
rect 16670 31240 16726 31249
rect 15936 31136 15988 31142
rect 15936 31078 15988 31084
rect 16028 31136 16080 31142
rect 16028 31078 16080 31084
rect 15948 30938 15976 31078
rect 15936 30932 15988 30938
rect 15936 30874 15988 30880
rect 16040 30802 16068 31078
rect 16132 30802 16160 31198
rect 16212 30932 16264 30938
rect 16212 30874 16264 30880
rect 15936 30796 15988 30802
rect 15936 30738 15988 30744
rect 16028 30796 16080 30802
rect 16028 30738 16080 30744
rect 16120 30796 16172 30802
rect 16120 30738 16172 30744
rect 15844 29776 15896 29782
rect 15844 29718 15896 29724
rect 15948 29714 15976 30738
rect 15936 29708 15988 29714
rect 15936 29650 15988 29656
rect 16120 29708 16172 29714
rect 16120 29650 16172 29656
rect 15844 29640 15896 29646
rect 15844 29582 15896 29588
rect 15856 29152 15884 29582
rect 15948 29306 15976 29650
rect 15936 29300 15988 29306
rect 16132 29288 16160 29650
rect 16224 29510 16252 30874
rect 16316 30802 16344 31214
rect 16580 31204 16632 31210
rect 16670 31175 16726 31184
rect 16580 31146 16632 31152
rect 16304 30796 16356 30802
rect 16304 30738 16356 30744
rect 16592 30734 16620 31146
rect 17224 31136 17276 31142
rect 17224 31078 17276 31084
rect 16580 30728 16632 30734
rect 16580 30670 16632 30676
rect 17236 29646 17264 31078
rect 17224 29640 17276 29646
rect 17224 29582 17276 29588
rect 16212 29504 16264 29510
rect 16212 29446 16264 29452
rect 15936 29242 15988 29248
rect 16040 29260 16160 29288
rect 15936 29164 15988 29170
rect 15856 29124 15936 29152
rect 15936 29106 15988 29112
rect 15948 28218 15976 29106
rect 15936 28212 15988 28218
rect 15936 28154 15988 28160
rect 15752 27124 15804 27130
rect 15752 27066 15804 27072
rect 16040 26602 16068 29260
rect 16120 29164 16172 29170
rect 16120 29106 16172 29112
rect 16132 28762 16160 29106
rect 17132 29028 17184 29034
rect 17132 28970 17184 28976
rect 16120 28756 16172 28762
rect 16120 28698 16172 28704
rect 16132 28082 16160 28698
rect 17144 28558 17172 28970
rect 17224 28688 17276 28694
rect 17224 28630 17276 28636
rect 17132 28552 17184 28558
rect 17132 28494 17184 28500
rect 16120 28076 16172 28082
rect 16120 28018 16172 28024
rect 17144 28014 17172 28494
rect 17132 28008 17184 28014
rect 17132 27950 17184 27956
rect 16396 27600 16448 27606
rect 16396 27542 16448 27548
rect 16408 26994 16436 27542
rect 16396 26988 16448 26994
rect 16396 26930 16448 26936
rect 16948 26988 17000 26994
rect 16948 26930 17000 26936
rect 16304 26784 16356 26790
rect 16304 26726 16356 26732
rect 15568 26580 15620 26586
rect 16040 26574 16160 26602
rect 15568 26522 15620 26528
rect 16028 26444 16080 26450
rect 16028 26386 16080 26392
rect 15568 25900 15620 25906
rect 15568 25842 15620 25848
rect 15580 25362 15608 25842
rect 15660 25696 15712 25702
rect 15660 25638 15712 25644
rect 15752 25696 15804 25702
rect 15752 25638 15804 25644
rect 15568 25356 15620 25362
rect 15568 25298 15620 25304
rect 15672 24886 15700 25638
rect 15660 24880 15712 24886
rect 15660 24822 15712 24828
rect 15764 23322 15792 25638
rect 16040 25294 16068 26386
rect 15844 25288 15896 25294
rect 15844 25230 15896 25236
rect 16028 25288 16080 25294
rect 16028 25230 16080 25236
rect 15856 24954 15884 25230
rect 15844 24948 15896 24954
rect 15844 24890 15896 24896
rect 16028 24200 16080 24206
rect 16028 24142 16080 24148
rect 15936 23656 15988 23662
rect 15936 23598 15988 23604
rect 15752 23316 15804 23322
rect 15752 23258 15804 23264
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15844 23112 15896 23118
rect 15844 23054 15896 23060
rect 15672 22778 15700 23054
rect 15660 22772 15712 22778
rect 15660 22714 15712 22720
rect 15752 22704 15804 22710
rect 15752 22646 15804 22652
rect 15764 22166 15792 22646
rect 15856 22438 15884 23054
rect 15948 22778 15976 23598
rect 16040 22982 16068 24142
rect 16132 23089 16160 26574
rect 16316 26382 16344 26726
rect 16960 26518 16988 26930
rect 16856 26512 16908 26518
rect 16854 26480 16856 26489
rect 16948 26512 17000 26518
rect 16908 26480 16910 26489
rect 16948 26454 17000 26460
rect 16854 26415 16910 26424
rect 16304 26376 16356 26382
rect 16224 26336 16304 26364
rect 16224 25974 16252 26336
rect 16304 26318 16356 26324
rect 17040 26376 17092 26382
rect 17040 26318 17092 26324
rect 16488 26308 16540 26314
rect 16488 26250 16540 26256
rect 16212 25968 16264 25974
rect 16396 25968 16448 25974
rect 16212 25910 16264 25916
rect 16394 25936 16396 25945
rect 16448 25936 16450 25945
rect 16394 25871 16450 25880
rect 16500 25838 16528 26250
rect 16580 25900 16632 25906
rect 16580 25842 16632 25848
rect 16488 25832 16540 25838
rect 16488 25774 16540 25780
rect 16212 25424 16264 25430
rect 16264 25384 16344 25412
rect 16212 25366 16264 25372
rect 16212 24880 16264 24886
rect 16212 24822 16264 24828
rect 16224 24410 16252 24822
rect 16212 24404 16264 24410
rect 16212 24346 16264 24352
rect 16118 23080 16174 23089
rect 16118 23015 16174 23024
rect 16028 22976 16080 22982
rect 16028 22918 16080 22924
rect 15936 22772 15988 22778
rect 15936 22714 15988 22720
rect 16028 22636 16080 22642
rect 16028 22578 16080 22584
rect 15844 22432 15896 22438
rect 15844 22374 15896 22380
rect 15752 22160 15804 22166
rect 15752 22102 15804 22108
rect 16040 22098 16068 22578
rect 16028 22092 16080 22098
rect 16028 22034 16080 22040
rect 16040 21690 16068 22034
rect 16028 21684 16080 21690
rect 16028 21626 16080 21632
rect 16040 21418 16068 21626
rect 16132 21418 16160 23015
rect 16212 22160 16264 22166
rect 16212 22102 16264 22108
rect 16028 21412 16080 21418
rect 16028 21354 16080 21360
rect 16120 21412 16172 21418
rect 16120 21354 16172 21360
rect 15476 20868 15528 20874
rect 15476 20810 15528 20816
rect 15568 20800 15620 20806
rect 15568 20742 15620 20748
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15344 19332 15424 19360
rect 15292 19314 15344 19320
rect 15016 19236 15068 19242
rect 15016 19178 15068 19184
rect 15396 18902 15424 19332
rect 15384 18896 15436 18902
rect 15384 18838 15436 18844
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 15304 18086 15332 18702
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15396 17898 15424 18838
rect 15304 17870 15424 17898
rect 14924 17264 14976 17270
rect 14924 17206 14976 17212
rect 14832 17196 14884 17202
rect 14832 17138 14884 17144
rect 15304 16640 15332 17870
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15396 16998 15424 17614
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15384 16652 15436 16658
rect 15304 16612 15384 16640
rect 15384 16594 15436 16600
rect 14648 16516 14700 16522
rect 14648 16458 14700 16464
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14280 16244 14332 16250
rect 14280 16186 14332 16192
rect 14464 16244 14516 16250
rect 14464 16186 14516 16192
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 14108 15638 14136 15982
rect 14096 15632 14148 15638
rect 14096 15574 14148 15580
rect 14200 15570 14228 15982
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14292 15502 14320 16050
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 13740 12406 13860 12434
rect 13634 11792 13690 11801
rect 13634 11727 13690 11736
rect 13452 11144 13504 11150
rect 13504 11104 13584 11132
rect 13452 11086 13504 11092
rect 13358 10704 13414 10713
rect 13358 10639 13414 10648
rect 13372 9674 13400 10639
rect 13556 10062 13584 11104
rect 13648 10606 13676 11727
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13372 9646 13492 9674
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13268 9444 13320 9450
rect 13268 9386 13320 9392
rect 13176 5296 13228 5302
rect 13176 5238 13228 5244
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 13096 4758 13124 5102
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 11980 4004 12032 4010
rect 11980 3946 12032 3952
rect 11520 3052 11572 3058
rect 11348 3012 11520 3040
rect 11520 2994 11572 3000
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 11532 2582 11560 2994
rect 11624 2650 11652 2994
rect 11992 2990 12020 3946
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12622 3904 12678 3913
rect 12176 3738 12204 3878
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 12268 3602 12296 3878
rect 12622 3839 12678 3848
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 12360 2530 12388 3334
rect 12452 3126 12480 3334
rect 12440 3120 12492 3126
rect 12440 3062 12492 3068
rect 12532 2848 12584 2854
rect 12532 2790 12584 2796
rect 8944 2508 8996 2514
rect 12360 2502 12480 2530
rect 8944 2450 8996 2456
rect 12452 2446 12480 2502
rect 12544 2446 12572 2790
rect 12636 2514 12664 3839
rect 12820 2922 12848 4082
rect 12808 2916 12860 2922
rect 12808 2858 12860 2864
rect 13280 2774 13308 9386
rect 13372 7868 13400 9522
rect 13464 8362 13492 9646
rect 13740 9568 13768 12406
rect 13818 11248 13874 11257
rect 13818 11183 13820 11192
rect 13872 11183 13874 11192
rect 13820 11154 13872 11160
rect 13820 11076 13872 11082
rect 13924 11064 13952 14554
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14186 13016 14242 13025
rect 14186 12951 14242 12960
rect 14004 11892 14056 11898
rect 14004 11834 14056 11840
rect 14016 11150 14044 11834
rect 14200 11830 14228 12951
rect 14292 12850 14320 14214
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14200 11234 14228 11766
rect 14292 11762 14320 12786
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 14108 11218 14228 11234
rect 14096 11212 14228 11218
rect 14148 11206 14228 11212
rect 14096 11154 14148 11160
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 13872 11036 13952 11064
rect 13820 11018 13872 11024
rect 13648 9540 13768 9568
rect 13542 9344 13598 9353
rect 13542 9279 13598 9288
rect 13556 8974 13584 9279
rect 13648 8974 13676 9540
rect 13726 9480 13782 9489
rect 13726 9415 13782 9424
rect 13740 8974 13768 9415
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13544 7880 13596 7886
rect 13372 7840 13544 7868
rect 13544 7822 13596 7828
rect 13556 6322 13584 7822
rect 13648 6390 13676 8910
rect 13832 8906 13860 11018
rect 14016 10674 14044 11086
rect 14096 11076 14148 11082
rect 14096 11018 14148 11024
rect 14108 10810 14136 11018
rect 14200 10810 14228 11086
rect 14292 11014 14320 11086
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 13912 9648 13964 9654
rect 13910 9616 13912 9625
rect 13964 9616 13966 9625
rect 13910 9551 13966 9560
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13464 5778 13492 6054
rect 13452 5772 13504 5778
rect 13452 5714 13504 5720
rect 13556 5302 13584 6258
rect 13832 6186 13860 8298
rect 13924 8090 13952 8910
rect 14108 8634 14136 10542
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14002 7304 14058 7313
rect 14002 7239 14058 7248
rect 13912 6384 13964 6390
rect 13912 6326 13964 6332
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13924 5710 13952 6326
rect 14016 6254 14044 7239
rect 14108 7206 14136 7686
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14108 6458 14136 6802
rect 14200 6798 14228 10406
rect 14292 9897 14320 10950
rect 14384 10674 14412 12582
rect 14476 11830 14504 16186
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 14556 15904 14608 15910
rect 14556 15846 14608 15852
rect 14568 15638 14596 15846
rect 14556 15632 14608 15638
rect 14556 15574 14608 15580
rect 14568 15026 14596 15574
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 14660 13938 14688 14418
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14568 13462 14596 13874
rect 14556 13456 14608 13462
rect 14556 13398 14608 13404
rect 14568 13161 14596 13398
rect 14554 13152 14610 13161
rect 14554 13087 14610 13096
rect 14660 12986 14688 13874
rect 14752 13462 14780 14010
rect 14844 13734 14872 15982
rect 14936 15638 14964 16390
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 14924 15632 14976 15638
rect 14924 15574 14976 15580
rect 14936 15026 14964 15574
rect 15396 15502 15424 16186
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15108 15428 15160 15434
rect 15108 15370 15160 15376
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14936 14074 14964 14214
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 14740 13456 14792 13462
rect 14740 13398 14792 13404
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 15028 12102 15056 14350
rect 15120 12646 15148 15370
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 15212 13530 15240 13670
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 15108 12164 15160 12170
rect 15108 12106 15160 12112
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 15016 11824 15068 11830
rect 15016 11766 15068 11772
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14464 11076 14516 11082
rect 14464 11018 14516 11024
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 14476 10985 14504 11018
rect 14462 10976 14518 10985
rect 14462 10911 14518 10920
rect 14568 10849 14596 11018
rect 14554 10840 14610 10849
rect 14476 10784 14554 10792
rect 14476 10775 14610 10784
rect 14476 10764 14596 10775
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14278 9888 14334 9897
rect 14278 9823 14334 9832
rect 14292 9450 14320 9823
rect 14280 9444 14332 9450
rect 14280 9386 14332 9392
rect 14292 8974 14320 9386
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14280 8560 14332 8566
rect 14280 8502 14332 8508
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 14292 6458 14320 8502
rect 14384 6798 14412 10610
rect 14476 10606 14504 10764
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14568 10062 14596 10610
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14476 8498 14504 9318
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 14004 6248 14056 6254
rect 14002 6216 14004 6225
rect 14056 6216 14058 6225
rect 14002 6151 14058 6160
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 13544 5296 13596 5302
rect 13464 5256 13544 5284
rect 13464 4214 13492 5256
rect 13544 5238 13596 5244
rect 14108 4758 14136 5510
rect 14096 4752 14148 4758
rect 14096 4694 14148 4700
rect 13452 4208 13504 4214
rect 13452 4150 13504 4156
rect 14370 4176 14426 4185
rect 13464 3534 13492 4150
rect 14370 4111 14426 4120
rect 14278 4040 14334 4049
rect 14278 3975 14334 3984
rect 14292 3534 14320 3975
rect 14384 3602 14412 4111
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 13912 3460 13964 3466
rect 13912 3402 13964 3408
rect 13924 3058 13952 3402
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 13924 2922 13952 2994
rect 13912 2916 13964 2922
rect 13912 2858 13964 2864
rect 13280 2746 13400 2774
rect 13372 2514 13400 2746
rect 14384 2514 14412 3538
rect 14476 3126 14504 8434
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14568 5574 14596 6598
rect 14660 5914 14688 11698
rect 15028 11529 15056 11766
rect 15014 11520 15070 11529
rect 15014 11455 15070 11464
rect 14922 11248 14978 11257
rect 14922 11183 14978 11192
rect 14936 11150 14964 11183
rect 14924 11144 14976 11150
rect 14924 11086 14976 11092
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14752 7868 14780 9998
rect 14936 9674 14964 11086
rect 14844 9646 14964 9674
rect 14844 8090 14872 9646
rect 14922 9208 14978 9217
rect 14922 9143 14978 9152
rect 14936 9110 14964 9143
rect 14924 9104 14976 9110
rect 14924 9046 14976 9052
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14832 7880 14884 7886
rect 14752 7840 14832 7868
rect 14752 7274 14780 7840
rect 14832 7822 14884 7828
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14740 7268 14792 7274
rect 14740 7210 14792 7216
rect 14752 7002 14780 7210
rect 14740 6996 14792 7002
rect 14740 6938 14792 6944
rect 14844 6730 14872 7278
rect 14832 6724 14884 6730
rect 14832 6666 14884 6672
rect 14740 6112 14792 6118
rect 14740 6054 14792 6060
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14568 5166 14596 5510
rect 14752 5166 14780 6054
rect 14832 5840 14884 5846
rect 14832 5782 14884 5788
rect 14556 5160 14608 5166
rect 14556 5102 14608 5108
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14844 5030 14872 5782
rect 14936 5778 14964 9046
rect 15028 8498 15056 11455
rect 15120 11354 15148 12106
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15212 11218 15240 11494
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 15120 8498 15148 10950
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15212 10577 15240 10610
rect 15198 10568 15254 10577
rect 15198 10503 15254 10512
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 15212 10062 15240 10202
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15304 10010 15332 14010
rect 15488 12832 15516 19654
rect 15580 18290 15608 20742
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15672 19854 15700 20402
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15752 19712 15804 19718
rect 15658 19680 15714 19689
rect 15752 19654 15804 19660
rect 15658 19615 15714 19624
rect 15672 19446 15700 19615
rect 15660 19440 15712 19446
rect 15660 19382 15712 19388
rect 15568 18284 15620 18290
rect 15568 18226 15620 18232
rect 15580 16794 15608 18226
rect 15660 18216 15712 18222
rect 15660 18158 15712 18164
rect 15672 17678 15700 18158
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15672 17202 15700 17614
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15660 16992 15712 16998
rect 15660 16934 15712 16940
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15672 16182 15700 16934
rect 15660 16176 15712 16182
rect 15660 16118 15712 16124
rect 15568 15972 15620 15978
rect 15568 15914 15620 15920
rect 15580 15434 15608 15914
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15568 15428 15620 15434
rect 15568 15370 15620 15376
rect 15580 14958 15608 15370
rect 15672 15026 15700 15846
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15396 12804 15516 12832
rect 15396 12481 15424 12804
rect 15580 12764 15608 14894
rect 15488 12736 15608 12764
rect 15382 12472 15438 12481
rect 15382 12407 15384 12416
rect 15436 12407 15438 12416
rect 15384 12378 15436 12384
rect 15382 12336 15438 12345
rect 15382 12271 15438 12280
rect 15396 10266 15424 12271
rect 15488 11762 15516 12736
rect 15672 12442 15700 14962
rect 15764 13394 15792 19654
rect 15856 18766 15884 20198
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15856 15978 15884 16526
rect 15936 16108 15988 16114
rect 16040 16096 16068 21354
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 16132 19854 16160 20402
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 16224 18902 16252 22102
rect 16316 22094 16344 25384
rect 16500 25226 16528 25774
rect 16592 25294 16620 25842
rect 17052 25294 17080 26318
rect 17132 25764 17184 25770
rect 17132 25706 17184 25712
rect 16580 25288 16632 25294
rect 16580 25230 16632 25236
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 16488 25220 16540 25226
rect 16488 25162 16540 25168
rect 17144 24886 17172 25706
rect 17132 24880 17184 24886
rect 17132 24822 17184 24828
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 16868 24274 16896 24754
rect 17132 24608 17184 24614
rect 17132 24550 17184 24556
rect 16856 24268 16908 24274
rect 16856 24210 16908 24216
rect 16396 24200 16448 24206
rect 16764 24200 16816 24206
rect 16396 24142 16448 24148
rect 16762 24168 16764 24177
rect 16816 24168 16818 24177
rect 16408 23866 16436 24142
rect 16762 24103 16818 24112
rect 16396 23860 16448 23866
rect 16396 23802 16448 23808
rect 16672 23520 16724 23526
rect 16672 23462 16724 23468
rect 16684 23322 16712 23462
rect 16776 23322 16804 24103
rect 17040 23724 17092 23730
rect 17040 23666 17092 23672
rect 17052 23322 17080 23666
rect 16672 23316 16724 23322
rect 16672 23258 16724 23264
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 17040 23316 17092 23322
rect 17040 23258 17092 23264
rect 17040 23112 17092 23118
rect 17040 23054 17092 23060
rect 16856 23044 16908 23050
rect 16856 22986 16908 22992
rect 16948 23044 17000 23050
rect 16948 22986 17000 22992
rect 16764 22568 16816 22574
rect 16764 22510 16816 22516
rect 16776 22234 16804 22510
rect 16868 22234 16896 22986
rect 16960 22778 16988 22986
rect 16948 22772 17000 22778
rect 16948 22714 17000 22720
rect 17052 22710 17080 23054
rect 17040 22704 17092 22710
rect 17040 22646 17092 22652
rect 17052 22506 17080 22646
rect 17040 22500 17092 22506
rect 17040 22442 17092 22448
rect 16764 22228 16816 22234
rect 16764 22170 16816 22176
rect 16856 22228 16908 22234
rect 16856 22170 16908 22176
rect 17038 22128 17094 22137
rect 16316 22066 16436 22094
rect 16304 20800 16356 20806
rect 16304 20742 16356 20748
rect 16316 19009 16344 20742
rect 16302 19000 16358 19009
rect 16302 18935 16358 18944
rect 16212 18896 16264 18902
rect 16212 18838 16264 18844
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 15988 16068 16068 16096
rect 15936 16050 15988 16056
rect 15844 15972 15896 15978
rect 15844 15914 15896 15920
rect 16040 15502 16068 16068
rect 15844 15496 15896 15502
rect 16028 15496 16080 15502
rect 15896 15456 15976 15484
rect 15844 15438 15896 15444
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15488 11014 15516 11698
rect 15580 11234 15608 12038
rect 15672 11665 15700 12174
rect 15658 11656 15714 11665
rect 15658 11591 15714 11600
rect 15672 11354 15700 11591
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15580 11206 15700 11234
rect 15568 11144 15620 11150
rect 15566 11112 15568 11121
rect 15620 11112 15622 11121
rect 15566 11047 15622 11056
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15488 10713 15516 10746
rect 15474 10704 15530 10713
rect 15474 10639 15530 10648
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15580 10010 15608 10610
rect 15212 9674 15240 9998
rect 15304 9982 15608 10010
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15212 9646 15332 9674
rect 15304 9586 15332 9646
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15396 9110 15424 9862
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 15016 8492 15068 8498
rect 15016 8434 15068 8440
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 15028 8022 15056 8230
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15016 8016 15068 8022
rect 15016 7958 15068 7964
rect 15120 6798 15148 8026
rect 15212 7886 15240 8910
rect 15396 8838 15424 9046
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15212 7342 15240 7822
rect 15292 7812 15344 7818
rect 15292 7754 15344 7760
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 15304 7274 15332 7754
rect 15396 7410 15424 8230
rect 15488 7886 15516 9982
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15580 9654 15608 9862
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15672 9586 15700 11206
rect 15764 10266 15792 13330
rect 15948 12442 15976 15456
rect 16028 15438 16080 15444
rect 16132 13938 16160 18566
rect 16316 18290 16344 18935
rect 16408 18329 16436 22066
rect 17038 22063 17040 22072
rect 17092 22063 17094 22072
rect 17040 22034 17092 22040
rect 17040 21956 17092 21962
rect 17040 21898 17092 21904
rect 17052 21865 17080 21898
rect 17038 21856 17094 21865
rect 17038 21791 17094 21800
rect 16672 21344 16724 21350
rect 16672 21286 16724 21292
rect 16684 21146 16712 21286
rect 16672 21140 16724 21146
rect 16672 21082 16724 21088
rect 17144 20466 17172 24550
rect 17236 22778 17264 28630
rect 17328 28626 17356 32506
rect 17512 30841 17540 33050
rect 17696 32910 17724 33458
rect 17788 32910 17816 33798
rect 18052 33448 18104 33454
rect 18052 33390 18104 33396
rect 17684 32904 17736 32910
rect 17684 32846 17736 32852
rect 17776 32904 17828 32910
rect 17960 32904 18012 32910
rect 17776 32846 17828 32852
rect 17880 32864 17960 32892
rect 17592 30864 17644 30870
rect 17498 30832 17554 30841
rect 17592 30806 17644 30812
rect 17498 30767 17554 30776
rect 17316 28620 17368 28626
rect 17316 28562 17368 28568
rect 17328 26518 17356 28562
rect 17500 27396 17552 27402
rect 17500 27338 17552 27344
rect 17512 27130 17540 27338
rect 17500 27124 17552 27130
rect 17500 27066 17552 27072
rect 17316 26512 17368 26518
rect 17604 26466 17632 30806
rect 17696 30326 17724 32846
rect 17880 32774 17908 32864
rect 17960 32846 18012 32852
rect 17868 32768 17920 32774
rect 17868 32710 17920 32716
rect 17960 32768 18012 32774
rect 17960 32710 18012 32716
rect 17880 32434 17908 32710
rect 17868 32428 17920 32434
rect 17868 32370 17920 32376
rect 17972 32366 18000 32710
rect 18064 32366 18092 33390
rect 18156 33114 18184 33934
rect 18144 33108 18196 33114
rect 18144 33050 18196 33056
rect 18156 32978 18184 33050
rect 18248 32978 18276 34342
rect 18328 33516 18380 33522
rect 18328 33458 18380 33464
rect 18144 32972 18196 32978
rect 18144 32914 18196 32920
rect 18236 32972 18288 32978
rect 18236 32914 18288 32920
rect 18248 32570 18276 32914
rect 18236 32564 18288 32570
rect 18236 32506 18288 32512
rect 17960 32360 18012 32366
rect 17960 32302 18012 32308
rect 18052 32360 18104 32366
rect 18052 32302 18104 32308
rect 18064 32230 18092 32302
rect 18052 32224 18104 32230
rect 18052 32166 18104 32172
rect 18340 31754 18368 33458
rect 18512 33312 18564 33318
rect 18512 33254 18564 33260
rect 18524 32910 18552 33254
rect 18512 32904 18564 32910
rect 18512 32846 18564 32852
rect 18788 32904 18840 32910
rect 18788 32846 18840 32852
rect 18800 32570 18828 32846
rect 18788 32564 18840 32570
rect 18788 32506 18840 32512
rect 18788 32428 18840 32434
rect 18788 32370 18840 32376
rect 18604 32360 18656 32366
rect 18604 32302 18656 32308
rect 18512 32224 18564 32230
rect 18512 32166 18564 32172
rect 18524 31890 18552 32166
rect 18512 31884 18564 31890
rect 18512 31826 18564 31832
rect 18248 31726 18368 31754
rect 18144 31408 18196 31414
rect 18144 31350 18196 31356
rect 17960 31136 18012 31142
rect 17960 31078 18012 31084
rect 17972 30666 18000 31078
rect 18156 30818 18184 31350
rect 18248 31346 18276 31726
rect 18616 31414 18644 32302
rect 18800 31754 18828 32370
rect 18788 31748 18840 31754
rect 18788 31690 18840 31696
rect 18604 31408 18656 31414
rect 18604 31350 18656 31356
rect 18236 31340 18288 31346
rect 18236 31282 18288 31288
rect 18604 31272 18656 31278
rect 18656 31220 18736 31226
rect 18604 31214 18736 31220
rect 18616 31198 18736 31214
rect 18604 31136 18656 31142
rect 18604 31078 18656 31084
rect 18616 30938 18644 31078
rect 18604 30932 18656 30938
rect 18604 30874 18656 30880
rect 18156 30790 18276 30818
rect 18248 30734 18276 30790
rect 18236 30728 18288 30734
rect 18236 30670 18288 30676
rect 17960 30660 18012 30666
rect 17960 30602 18012 30608
rect 17684 30320 17736 30326
rect 17684 30262 17736 30268
rect 17696 27470 17724 30262
rect 18144 29776 18196 29782
rect 18144 29718 18196 29724
rect 18156 29170 18184 29718
rect 17868 29164 17920 29170
rect 17868 29106 17920 29112
rect 17960 29164 18012 29170
rect 17960 29106 18012 29112
rect 18144 29164 18196 29170
rect 18144 29106 18196 29112
rect 17776 28620 17828 28626
rect 17776 28562 17828 28568
rect 17788 28218 17816 28562
rect 17880 28218 17908 29106
rect 17972 28422 18000 29106
rect 18052 28688 18104 28694
rect 18052 28630 18104 28636
rect 17960 28416 18012 28422
rect 17960 28358 18012 28364
rect 17776 28212 17828 28218
rect 17776 28154 17828 28160
rect 17868 28212 17920 28218
rect 17868 28154 17920 28160
rect 17972 28082 18000 28358
rect 17960 28076 18012 28082
rect 17960 28018 18012 28024
rect 17684 27464 17736 27470
rect 17684 27406 17736 27412
rect 17684 27328 17736 27334
rect 17684 27270 17736 27276
rect 17316 26454 17368 26460
rect 17328 25702 17356 26454
rect 17512 26438 17632 26466
rect 17512 26246 17540 26438
rect 17592 26376 17644 26382
rect 17592 26318 17644 26324
rect 17500 26240 17552 26246
rect 17500 26182 17552 26188
rect 17316 25696 17368 25702
rect 17316 25638 17368 25644
rect 17408 25696 17460 25702
rect 17408 25638 17460 25644
rect 17420 25498 17448 25638
rect 17408 25492 17460 25498
rect 17408 25434 17460 25440
rect 17316 25424 17368 25430
rect 17512 25378 17540 26182
rect 17604 25906 17632 26318
rect 17592 25900 17644 25906
rect 17592 25842 17644 25848
rect 17316 25366 17368 25372
rect 17328 24886 17356 25366
rect 17420 25350 17540 25378
rect 17316 24880 17368 24886
rect 17316 24822 17368 24828
rect 17420 24818 17448 25350
rect 17500 25288 17552 25294
rect 17498 25256 17500 25265
rect 17552 25256 17554 25265
rect 17498 25191 17554 25200
rect 17408 24812 17460 24818
rect 17408 24754 17460 24760
rect 17604 24342 17632 25842
rect 17592 24336 17644 24342
rect 17592 24278 17644 24284
rect 17592 23724 17644 23730
rect 17592 23666 17644 23672
rect 17604 23526 17632 23666
rect 17696 23662 17724 27270
rect 18064 27130 18092 28630
rect 18156 27946 18184 29106
rect 18144 27940 18196 27946
rect 18144 27882 18196 27888
rect 18052 27124 18104 27130
rect 18052 27066 18104 27072
rect 17776 26784 17828 26790
rect 17776 26726 17828 26732
rect 17684 23656 17736 23662
rect 17684 23598 17736 23604
rect 17592 23520 17644 23526
rect 17592 23462 17644 23468
rect 17316 23112 17368 23118
rect 17316 23054 17368 23060
rect 17408 23112 17460 23118
rect 17460 23072 17540 23100
rect 17408 23054 17460 23060
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 17328 22642 17356 23054
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 17316 22636 17368 22642
rect 17316 22578 17368 22584
rect 17224 22500 17276 22506
rect 17224 22442 17276 22448
rect 17236 20602 17264 22442
rect 17328 22098 17356 22578
rect 17316 22092 17368 22098
rect 17316 22034 17368 22040
rect 17328 21690 17356 22034
rect 17316 21684 17368 21690
rect 17316 21626 17368 21632
rect 17316 21480 17368 21486
rect 17316 21422 17368 21428
rect 17328 20806 17356 21422
rect 17316 20800 17368 20806
rect 17316 20742 17368 20748
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 16488 19848 16540 19854
rect 16486 19816 16488 19825
rect 16540 19816 16542 19825
rect 16486 19751 16542 19760
rect 16960 19689 16988 19858
rect 16946 19680 17002 19689
rect 16946 19615 17002 19624
rect 16672 19236 16724 19242
rect 16672 19178 16724 19184
rect 16684 18834 16712 19178
rect 16672 18828 16724 18834
rect 16724 18788 16804 18816
rect 16672 18770 16724 18776
rect 16394 18320 16450 18329
rect 16304 18284 16356 18290
rect 16394 18255 16450 18264
rect 16580 18284 16632 18290
rect 16304 18226 16356 18232
rect 16580 18226 16632 18232
rect 16302 18184 16358 18193
rect 16302 18119 16358 18128
rect 16212 17604 16264 17610
rect 16212 17546 16264 17552
rect 16224 16114 16252 17546
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16120 13932 16172 13938
rect 16172 13892 16252 13920
rect 16120 13874 16172 13880
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 16118 13424 16174 13433
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 15856 12322 15884 12378
rect 15856 12294 15976 12322
rect 15842 12200 15898 12209
rect 15842 12135 15844 12144
rect 15896 12135 15898 12144
rect 15844 12106 15896 12112
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15764 10130 15792 10202
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15672 9042 15700 9522
rect 15764 9466 15792 9862
rect 15856 9586 15884 12106
rect 15948 11694 15976 12294
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 16040 11354 16068 13398
rect 16118 13359 16120 13368
rect 16172 13359 16174 13368
rect 16120 13330 16172 13336
rect 16224 12918 16252 13892
rect 16212 12912 16264 12918
rect 16212 12854 16264 12860
rect 16316 12594 16344 18119
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16500 17610 16528 18022
rect 16592 17678 16620 18226
rect 16670 18048 16726 18057
rect 16670 17983 16726 17992
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16500 17270 16528 17546
rect 16488 17264 16540 17270
rect 16488 17206 16540 17212
rect 16486 17096 16542 17105
rect 16592 17082 16620 17614
rect 16542 17054 16620 17082
rect 16486 17031 16542 17040
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 16408 14074 16436 14894
rect 16488 14340 16540 14346
rect 16488 14282 16540 14288
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16500 13734 16528 14282
rect 16488 13728 16540 13734
rect 16488 13670 16540 13676
rect 16500 13326 16528 13670
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16316 12566 16436 12594
rect 16408 12442 16436 12566
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16120 12300 16172 12306
rect 16120 12242 16172 12248
rect 16132 11370 16160 12242
rect 16316 12220 16344 12378
rect 16488 12232 16540 12238
rect 16316 12192 16436 12220
rect 16408 11778 16436 12192
rect 16488 12174 16540 12180
rect 16500 12102 16528 12174
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16408 11750 16620 11778
rect 16302 11384 16358 11393
rect 16132 11354 16252 11370
rect 16028 11348 16080 11354
rect 16132 11348 16264 11354
rect 16132 11342 16212 11348
rect 16028 11290 16080 11296
rect 16302 11319 16358 11328
rect 16212 11290 16264 11296
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15948 9926 15976 10610
rect 15936 9920 15988 9926
rect 15936 9862 15988 9868
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15764 9438 15884 9466
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15292 7268 15344 7274
rect 15292 7210 15344 7216
rect 15488 6866 15516 7346
rect 15580 6882 15608 7754
rect 15672 7410 15700 8230
rect 15660 7404 15712 7410
rect 15660 7346 15712 7352
rect 15476 6860 15528 6866
rect 15580 6854 15700 6882
rect 15476 6802 15528 6808
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15488 6186 15516 6802
rect 15672 6798 15700 6854
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15476 6180 15528 6186
rect 15476 6122 15528 6128
rect 15580 5778 15608 6394
rect 14924 5772 14976 5778
rect 14924 5714 14976 5720
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15672 5710 15700 6734
rect 15764 6662 15792 8910
rect 15856 7886 15884 9438
rect 15948 9178 15976 9522
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 16040 7410 16068 11290
rect 16212 11212 16264 11218
rect 16316 11200 16344 11319
rect 16264 11172 16344 11200
rect 16212 11154 16264 11160
rect 16302 11112 16358 11121
rect 16302 11047 16358 11056
rect 16118 10840 16174 10849
rect 16174 10798 16252 10826
rect 16118 10775 16174 10784
rect 16224 10674 16252 10798
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16132 9704 16160 10610
rect 16132 9676 16252 9704
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 16132 8634 16160 9522
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16224 8430 16252 9676
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16224 7886 16252 8366
rect 16316 8294 16344 11047
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16316 7750 16344 7822
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16408 7410 16436 11750
rect 16592 11694 16620 11750
rect 16580 11688 16632 11694
rect 16580 11630 16632 11636
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 16500 9674 16528 11562
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16592 10470 16620 10950
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16684 9722 16712 17983
rect 16776 13394 16804 18788
rect 17040 18216 17092 18222
rect 17040 18158 17092 18164
rect 16856 18080 16908 18086
rect 16856 18022 16908 18028
rect 16868 17678 16896 18022
rect 17052 17746 17080 18158
rect 17040 17740 17092 17746
rect 17040 17682 17092 17688
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16868 17241 16896 17614
rect 17040 17604 17092 17610
rect 17040 17546 17092 17552
rect 16854 17232 16910 17241
rect 17052 17202 17080 17546
rect 16854 17167 16856 17176
rect 16908 17167 16910 17176
rect 17040 17196 17092 17202
rect 16856 17138 16908 17144
rect 17040 17138 17092 17144
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16960 16522 16988 16934
rect 17144 16674 17172 20402
rect 17420 19836 17448 22714
rect 17512 22030 17540 23072
rect 17604 22778 17632 23462
rect 17592 22772 17644 22778
rect 17592 22714 17644 22720
rect 17696 22658 17724 23598
rect 17604 22630 17724 22658
rect 17604 22506 17632 22630
rect 17788 22574 17816 26726
rect 18064 26382 18092 27066
rect 18052 26376 18104 26382
rect 18052 26318 18104 26324
rect 17868 26240 17920 26246
rect 17868 26182 17920 26188
rect 18052 26240 18104 26246
rect 18052 26182 18104 26188
rect 17880 24993 17908 26182
rect 17958 25800 18014 25809
rect 17958 25735 18014 25744
rect 17972 25498 18000 25735
rect 18064 25498 18092 26182
rect 17960 25492 18012 25498
rect 17960 25434 18012 25440
rect 18052 25492 18104 25498
rect 18052 25434 18104 25440
rect 18248 25378 18276 30670
rect 18602 30424 18658 30433
rect 18708 30410 18736 31198
rect 18658 30382 18736 30410
rect 18602 30359 18658 30368
rect 18512 28960 18564 28966
rect 18512 28902 18564 28908
rect 18524 28558 18552 28902
rect 18512 28552 18564 28558
rect 18512 28494 18564 28500
rect 18512 28076 18564 28082
rect 18512 28018 18564 28024
rect 18524 26926 18552 28018
rect 18696 27396 18748 27402
rect 18696 27338 18748 27344
rect 18512 26920 18564 26926
rect 18512 26862 18564 26868
rect 18326 26480 18382 26489
rect 18326 26415 18328 26424
rect 18380 26415 18382 26424
rect 18328 26386 18380 26392
rect 18524 26382 18552 26862
rect 18512 26376 18564 26382
rect 18512 26318 18564 26324
rect 17972 25350 18276 25378
rect 17866 24984 17922 24993
rect 17866 24919 17922 24928
rect 17868 24880 17920 24886
rect 17868 24822 17920 24828
rect 17776 22568 17828 22574
rect 17776 22510 17828 22516
rect 17592 22500 17644 22506
rect 17592 22442 17644 22448
rect 17776 22432 17828 22438
rect 17776 22374 17828 22380
rect 17788 22234 17816 22374
rect 17880 22234 17908 24822
rect 17776 22228 17828 22234
rect 17776 22170 17828 22176
rect 17868 22228 17920 22234
rect 17868 22170 17920 22176
rect 17774 22128 17830 22137
rect 17774 22063 17830 22072
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 17512 21690 17540 21966
rect 17684 21956 17736 21962
rect 17684 21898 17736 21904
rect 17696 21865 17724 21898
rect 17788 21894 17816 22063
rect 17868 22024 17920 22030
rect 17868 21966 17920 21972
rect 17776 21888 17828 21894
rect 17682 21856 17738 21865
rect 17776 21830 17828 21836
rect 17682 21791 17738 21800
rect 17500 21684 17552 21690
rect 17500 21626 17552 21632
rect 17880 21622 17908 21966
rect 17868 21616 17920 21622
rect 17868 21558 17920 21564
rect 17500 21548 17552 21554
rect 17500 21490 17552 21496
rect 17512 21457 17540 21490
rect 17498 21448 17554 21457
rect 17498 21383 17554 21392
rect 17512 21350 17540 21383
rect 17500 21344 17552 21350
rect 17500 21286 17552 21292
rect 17776 20460 17828 20466
rect 17776 20402 17828 20408
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 17592 20256 17644 20262
rect 17592 20198 17644 20204
rect 17512 19990 17540 20198
rect 17500 19984 17552 19990
rect 17500 19926 17552 19932
rect 17420 19808 17540 19836
rect 17224 19712 17276 19718
rect 17224 19654 17276 19660
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 17236 19514 17264 19654
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 17420 19310 17448 19654
rect 17408 19304 17460 19310
rect 17408 19246 17460 19252
rect 17512 17882 17540 19808
rect 17604 19446 17632 20198
rect 17788 19786 17816 20402
rect 17868 19984 17920 19990
rect 17868 19926 17920 19932
rect 17880 19854 17908 19926
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17776 19780 17828 19786
rect 17776 19722 17828 19728
rect 17592 19440 17644 19446
rect 17592 19382 17644 19388
rect 17592 18692 17644 18698
rect 17592 18634 17644 18640
rect 17500 17876 17552 17882
rect 17500 17818 17552 17824
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 17236 17270 17264 17614
rect 17224 17264 17276 17270
rect 17224 17206 17276 17212
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17512 16794 17540 16934
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17052 16646 17172 16674
rect 16948 16516 17000 16522
rect 16948 16458 17000 16464
rect 16948 15428 17000 15434
rect 16948 15370 17000 15376
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 16764 13388 16816 13394
rect 16764 13330 16816 13336
rect 16868 12646 16896 15098
rect 16960 14929 16988 15370
rect 16946 14920 17002 14929
rect 16946 14855 17002 14864
rect 16960 13462 16988 14855
rect 17052 14618 17080 16646
rect 17408 16584 17460 16590
rect 17408 16526 17460 16532
rect 17224 16516 17276 16522
rect 17224 16458 17276 16464
rect 17236 16114 17264 16458
rect 17224 16108 17276 16114
rect 17224 16050 17276 16056
rect 17236 15570 17264 16050
rect 17316 16040 17368 16046
rect 17316 15982 17368 15988
rect 17224 15564 17276 15570
rect 17224 15506 17276 15512
rect 17132 15428 17184 15434
rect 17132 15370 17184 15376
rect 17144 15026 17172 15370
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 16948 13456 17000 13462
rect 16948 13398 17000 13404
rect 16948 13252 17000 13258
rect 17052 13240 17080 13670
rect 17144 13326 17172 14962
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 17236 14550 17264 14826
rect 17224 14544 17276 14550
rect 17224 14486 17276 14492
rect 17328 14414 17356 15982
rect 17420 15502 17448 16526
rect 17512 16454 17540 16730
rect 17500 16448 17552 16454
rect 17500 16390 17552 16396
rect 17512 16114 17540 16390
rect 17604 16250 17632 18634
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 17788 17882 17816 18362
rect 17868 18216 17920 18222
rect 17868 18158 17920 18164
rect 17776 17876 17828 17882
rect 17776 17818 17828 17824
rect 17776 17672 17828 17678
rect 17776 17614 17828 17620
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 17512 15502 17540 16050
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17500 15496 17552 15502
rect 17500 15438 17552 15444
rect 17604 15314 17632 16186
rect 17420 15286 17632 15314
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17000 13212 17080 13240
rect 16948 13194 17000 13200
rect 16960 12889 16988 13194
rect 16946 12880 17002 12889
rect 16946 12815 17002 12824
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16868 12442 16896 12582
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 16868 12345 16896 12378
rect 16854 12336 16910 12345
rect 16854 12271 16910 12280
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16764 11348 16816 11354
rect 16764 11290 16816 11296
rect 16776 10742 16804 11290
rect 16764 10736 16816 10742
rect 16868 10713 16896 11494
rect 16764 10678 16816 10684
rect 16854 10704 16910 10713
rect 16854 10639 16910 10648
rect 16856 10600 16908 10606
rect 16960 10577 16988 12174
rect 17144 11558 17172 13262
rect 17328 13190 17356 13262
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17236 11082 17264 12174
rect 17328 11762 17356 12242
rect 17420 12102 17448 15286
rect 17498 15192 17554 15201
rect 17696 15162 17724 16390
rect 17788 15473 17816 17614
rect 17774 15464 17830 15473
rect 17774 15399 17830 15408
rect 17774 15192 17830 15201
rect 17684 15156 17736 15162
rect 17498 15127 17554 15136
rect 17512 14006 17540 15127
rect 17604 15116 17684 15144
rect 17500 14000 17552 14006
rect 17500 13942 17552 13948
rect 17604 13394 17632 15116
rect 17774 15127 17830 15136
rect 17684 15098 17736 15104
rect 17788 15026 17816 15127
rect 17776 15020 17828 15026
rect 17776 14962 17828 14968
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 17592 13388 17644 13394
rect 17592 13330 17644 13336
rect 17604 12374 17632 13330
rect 17592 12368 17644 12374
rect 17592 12310 17644 12316
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17316 11756 17368 11762
rect 17420 11744 17448 12038
rect 17696 11880 17724 14214
rect 17788 13954 17816 14962
rect 17880 14414 17908 18158
rect 17972 17252 18000 25350
rect 18052 25288 18104 25294
rect 18052 25230 18104 25236
rect 18144 25288 18196 25294
rect 18144 25230 18196 25236
rect 18064 24750 18092 25230
rect 18156 24818 18184 25230
rect 18524 25158 18552 26318
rect 18708 25498 18736 27338
rect 18788 26920 18840 26926
rect 18788 26862 18840 26868
rect 18800 25702 18828 26862
rect 18788 25696 18840 25702
rect 18788 25638 18840 25644
rect 18696 25492 18748 25498
rect 18696 25434 18748 25440
rect 18512 25152 18564 25158
rect 18512 25094 18564 25100
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 18052 24744 18104 24750
rect 18052 24686 18104 24692
rect 18524 24614 18552 25094
rect 18708 24886 18736 25434
rect 18696 24880 18748 24886
rect 18696 24822 18748 24828
rect 18800 24818 18828 25638
rect 18788 24812 18840 24818
rect 18788 24754 18840 24760
rect 18696 24744 18748 24750
rect 18696 24686 18748 24692
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18708 24206 18736 24686
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 18328 23520 18380 23526
rect 18328 23462 18380 23468
rect 18340 23186 18368 23462
rect 18892 23322 18920 35634
rect 19352 35154 19380 35935
rect 19340 35148 19392 35154
rect 19340 35090 19392 35096
rect 19064 34944 19116 34950
rect 19064 34886 19116 34892
rect 18970 34776 19026 34785
rect 18970 34711 19026 34720
rect 18984 32570 19012 34711
rect 19076 33114 19104 34886
rect 19444 34542 19472 36790
rect 19812 36242 19840 37742
rect 19984 37732 20036 37738
rect 19984 37674 20036 37680
rect 19996 37466 20024 37674
rect 19984 37460 20036 37466
rect 19984 37402 20036 37408
rect 20352 37460 20404 37466
rect 20352 37402 20404 37408
rect 20364 37346 20392 37402
rect 20180 37330 20392 37346
rect 20168 37324 20392 37330
rect 20220 37318 20392 37324
rect 20168 37266 20220 37272
rect 19892 37256 19944 37262
rect 19892 37198 19944 37204
rect 19800 36236 19852 36242
rect 19800 36178 19852 36184
rect 19616 36168 19668 36174
rect 19616 36110 19668 36116
rect 19628 35834 19656 36110
rect 19708 36032 19760 36038
rect 19708 35974 19760 35980
rect 19616 35828 19668 35834
rect 19616 35770 19668 35776
rect 19616 35488 19668 35494
rect 19616 35430 19668 35436
rect 19628 35154 19656 35430
rect 19720 35290 19748 35974
rect 19708 35284 19760 35290
rect 19708 35226 19760 35232
rect 19616 35148 19668 35154
rect 19616 35090 19668 35096
rect 19432 34536 19484 34542
rect 19432 34478 19484 34484
rect 19340 33516 19392 33522
rect 19340 33458 19392 33464
rect 19616 33516 19668 33522
rect 19616 33458 19668 33464
rect 19064 33108 19116 33114
rect 19064 33050 19116 33056
rect 19352 32910 19380 33458
rect 19432 33040 19484 33046
rect 19432 32982 19484 32988
rect 19340 32904 19392 32910
rect 19340 32846 19392 32852
rect 19248 32836 19300 32842
rect 19248 32778 19300 32784
rect 18972 32564 19024 32570
rect 18972 32506 19024 32512
rect 19260 32366 19288 32778
rect 19352 32434 19380 32846
rect 19340 32428 19392 32434
rect 19340 32370 19392 32376
rect 19064 32360 19116 32366
rect 19064 32302 19116 32308
rect 19156 32360 19208 32366
rect 19156 32302 19208 32308
rect 19248 32360 19300 32366
rect 19248 32302 19300 32308
rect 19076 32026 19104 32302
rect 19064 32020 19116 32026
rect 19064 31962 19116 31968
rect 19064 31816 19116 31822
rect 19064 31758 19116 31764
rect 19076 31482 19104 31758
rect 19064 31476 19116 31482
rect 19064 31418 19116 31424
rect 19064 31340 19116 31346
rect 19064 31282 19116 31288
rect 19076 30802 19104 31282
rect 19168 31210 19196 32302
rect 19352 31482 19380 32370
rect 19444 31754 19472 32982
rect 19628 32910 19656 33458
rect 19800 33312 19852 33318
rect 19800 33254 19852 33260
rect 19708 33108 19760 33114
rect 19708 33050 19760 33056
rect 19616 32904 19668 32910
rect 19616 32846 19668 32852
rect 19444 31726 19564 31754
rect 19340 31476 19392 31482
rect 19340 31418 19392 31424
rect 19156 31204 19208 31210
rect 19156 31146 19208 31152
rect 19064 30796 19116 30802
rect 19064 30738 19116 30744
rect 19536 29170 19564 31726
rect 19616 30252 19668 30258
rect 19616 30194 19668 30200
rect 19524 29164 19576 29170
rect 19524 29106 19576 29112
rect 19432 29028 19484 29034
rect 19432 28970 19484 28976
rect 18972 28484 19024 28490
rect 18972 28426 19024 28432
rect 19064 28484 19116 28490
rect 19064 28426 19116 28432
rect 18984 28014 19012 28426
rect 19076 28218 19104 28426
rect 19248 28416 19300 28422
rect 19248 28358 19300 28364
rect 19260 28218 19288 28358
rect 19064 28212 19116 28218
rect 19064 28154 19116 28160
rect 19248 28212 19300 28218
rect 19248 28154 19300 28160
rect 18972 28008 19024 28014
rect 18972 27950 19024 27956
rect 19340 27940 19392 27946
rect 19340 27882 19392 27888
rect 19352 27674 19380 27882
rect 19340 27668 19392 27674
rect 19340 27610 19392 27616
rect 19248 27396 19300 27402
rect 19248 27338 19300 27344
rect 19260 27130 19288 27338
rect 19444 27130 19472 28970
rect 19536 27606 19564 29106
rect 19524 27600 19576 27606
rect 19524 27542 19576 27548
rect 19524 27464 19576 27470
rect 19524 27406 19576 27412
rect 19248 27124 19300 27130
rect 19248 27066 19300 27072
rect 19432 27124 19484 27130
rect 19432 27066 19484 27072
rect 19444 26994 19472 27066
rect 19536 26994 19564 27406
rect 19628 26994 19656 30194
rect 19432 26988 19484 26994
rect 19432 26930 19484 26936
rect 19524 26988 19576 26994
rect 19524 26930 19576 26936
rect 19616 26988 19668 26994
rect 19616 26930 19668 26936
rect 19628 26874 19656 26930
rect 19536 26846 19656 26874
rect 19340 26580 19392 26586
rect 19340 26522 19392 26528
rect 19352 25906 19380 26522
rect 19248 25900 19300 25906
rect 19248 25842 19300 25848
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 19260 25786 19288 25842
rect 19260 25758 19380 25786
rect 18972 25696 19024 25702
rect 18972 25638 19024 25644
rect 18880 23316 18932 23322
rect 18880 23258 18932 23264
rect 18328 23180 18380 23186
rect 18328 23122 18380 23128
rect 18420 23112 18472 23118
rect 18248 23060 18420 23066
rect 18604 23112 18656 23118
rect 18248 23054 18472 23060
rect 18602 23080 18604 23089
rect 18696 23112 18748 23118
rect 18656 23080 18658 23089
rect 18248 23038 18460 23054
rect 18248 22982 18276 23038
rect 18696 23054 18748 23060
rect 18602 23015 18658 23024
rect 18236 22976 18288 22982
rect 18236 22918 18288 22924
rect 18328 22976 18380 22982
rect 18328 22918 18380 22924
rect 18144 22228 18196 22234
rect 18144 22170 18196 22176
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 18064 21350 18092 21966
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 18156 20466 18184 22170
rect 18248 21690 18276 22918
rect 18340 22574 18368 22918
rect 18420 22636 18472 22642
rect 18420 22578 18472 22584
rect 18328 22568 18380 22574
rect 18328 22510 18380 22516
rect 18432 22234 18460 22578
rect 18708 22506 18736 23054
rect 18696 22500 18748 22506
rect 18696 22442 18748 22448
rect 18420 22228 18472 22234
rect 18420 22170 18472 22176
rect 18236 21684 18288 21690
rect 18236 21626 18288 21632
rect 18144 20460 18196 20466
rect 18144 20402 18196 20408
rect 18604 20392 18656 20398
rect 18604 20334 18656 20340
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 18340 19446 18368 19722
rect 18418 19680 18474 19689
rect 18418 19615 18474 19624
rect 18328 19440 18380 19446
rect 18328 19382 18380 19388
rect 18340 18630 18368 19382
rect 18432 19242 18460 19615
rect 18420 19236 18472 19242
rect 18420 19178 18472 19184
rect 18432 18902 18460 19178
rect 18420 18896 18472 18902
rect 18420 18838 18472 18844
rect 18616 18766 18644 20334
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18420 18284 18472 18290
rect 18420 18226 18472 18232
rect 18052 17672 18104 17678
rect 18050 17640 18052 17649
rect 18236 17672 18288 17678
rect 18104 17640 18106 17649
rect 18236 17614 18288 17620
rect 18050 17575 18106 17584
rect 18144 17604 18196 17610
rect 18144 17546 18196 17552
rect 17972 17224 18092 17252
rect 17960 16720 18012 16726
rect 17960 16662 18012 16668
rect 17972 15502 18000 16662
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 17972 15026 18000 15098
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17972 14618 18000 14962
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17880 14278 17908 14350
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17788 13926 17908 13954
rect 17774 13832 17830 13841
rect 17774 13767 17776 13776
rect 17828 13767 17830 13776
rect 17776 13738 17828 13744
rect 17880 13258 17908 13926
rect 17868 13252 17920 13258
rect 17604 11852 17724 11880
rect 17788 13212 17868 13240
rect 17500 11756 17552 11762
rect 17420 11716 17500 11744
rect 17316 11698 17368 11704
rect 17500 11698 17552 11704
rect 17408 11620 17460 11626
rect 17408 11562 17460 11568
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17328 11150 17356 11494
rect 17420 11150 17448 11562
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17040 11076 17092 11082
rect 17040 11018 17092 11024
rect 17224 11076 17276 11082
rect 17224 11018 17276 11024
rect 17052 10810 17080 11018
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 16856 10542 16908 10548
rect 16946 10568 17002 10577
rect 16672 9716 16724 9722
rect 16500 9646 16620 9674
rect 16672 9658 16724 9664
rect 16486 9480 16542 9489
rect 16486 9415 16488 9424
rect 16540 9415 16542 9424
rect 16488 9386 16540 9392
rect 16488 8492 16540 8498
rect 16592 8480 16620 9646
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16540 8452 16620 8480
rect 16488 8434 16540 8440
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16488 7880 16540 7886
rect 16488 7822 16540 7828
rect 16500 7546 16528 7822
rect 16592 7546 16620 7890
rect 16488 7540 16540 7546
rect 16488 7482 16540 7488
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 16580 7268 16632 7274
rect 16580 7210 16632 7216
rect 16592 6934 16620 7210
rect 16580 6928 16632 6934
rect 16580 6870 16632 6876
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 16684 6322 16712 9522
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16776 8090 16804 9454
rect 16868 8294 16896 10542
rect 16946 10503 17002 10512
rect 16960 10198 16988 10503
rect 17052 10198 17080 10610
rect 16948 10192 17000 10198
rect 16948 10134 17000 10140
rect 17040 10192 17092 10198
rect 17040 10134 17092 10140
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16960 9897 16988 9998
rect 16946 9888 17002 9897
rect 16946 9823 17002 9832
rect 16960 9654 16988 9823
rect 17038 9752 17094 9761
rect 17038 9687 17094 9696
rect 16948 9648 17000 9654
rect 16948 9590 17000 9596
rect 17052 9450 17080 9687
rect 17040 9444 17092 9450
rect 17040 9386 17092 9392
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16868 7886 16896 8230
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16762 7712 16818 7721
rect 16762 7647 16818 7656
rect 16776 7478 16804 7647
rect 16764 7472 16816 7478
rect 16764 7414 16816 7420
rect 16868 6662 16896 7822
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16960 6458 16988 9318
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 17052 8401 17080 8434
rect 17038 8392 17094 8401
rect 17038 8327 17094 8336
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 17052 7410 17080 7958
rect 17144 7886 17172 10746
rect 17236 10742 17264 11018
rect 17328 10810 17356 11086
rect 17420 10810 17448 11086
rect 17500 11008 17552 11014
rect 17500 10950 17552 10956
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17408 10804 17460 10810
rect 17408 10746 17460 10752
rect 17224 10736 17276 10742
rect 17224 10678 17276 10684
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17224 10532 17276 10538
rect 17224 10474 17276 10480
rect 17132 7880 17184 7886
rect 17130 7848 17132 7857
rect 17184 7848 17186 7857
rect 17130 7783 17186 7792
rect 17144 7410 17172 7783
rect 17236 7449 17264 10474
rect 17328 10130 17356 10610
rect 17420 10418 17448 10610
rect 17512 10418 17540 10950
rect 17604 10538 17632 11852
rect 17788 11830 17816 13212
rect 17868 13194 17920 13200
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17592 10532 17644 10538
rect 17592 10474 17644 10480
rect 17420 10390 17632 10418
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17408 10056 17460 10062
rect 17406 10024 17408 10033
rect 17460 10024 17462 10033
rect 17316 9988 17368 9994
rect 17406 9959 17462 9968
rect 17316 9930 17368 9936
rect 17328 9674 17356 9930
rect 17328 9654 17540 9674
rect 17328 9648 17552 9654
rect 17328 9646 17500 9648
rect 17500 9590 17552 9596
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17316 9104 17368 9110
rect 17314 9072 17316 9081
rect 17368 9072 17370 9081
rect 17314 9007 17370 9016
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17328 7546 17356 8026
rect 17420 7585 17448 9522
rect 17500 9444 17552 9450
rect 17500 9386 17552 9392
rect 17406 7576 17462 7585
rect 17316 7540 17368 7546
rect 17406 7511 17462 7520
rect 17316 7482 17368 7488
rect 17222 7440 17278 7449
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 17132 7404 17184 7410
rect 17222 7375 17224 7384
rect 17132 7346 17184 7352
rect 17276 7375 17278 7384
rect 17224 7346 17276 7352
rect 17420 6458 17448 7511
rect 17512 7410 17540 9386
rect 17604 8430 17632 10390
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 17604 6798 17632 8366
rect 17696 7410 17724 11698
rect 17788 11150 17816 11766
rect 17776 11144 17828 11150
rect 17972 11098 18000 14350
rect 18064 12374 18092 17224
rect 18156 16522 18184 17546
rect 18144 16516 18196 16522
rect 18144 16458 18196 16464
rect 18156 14414 18184 16458
rect 18248 15026 18276 17614
rect 18432 16425 18460 18226
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 18524 17678 18552 18022
rect 18696 17876 18748 17882
rect 18696 17818 18748 17824
rect 18512 17672 18564 17678
rect 18512 17614 18564 17620
rect 18524 16794 18552 17614
rect 18708 17338 18736 17818
rect 18696 17332 18748 17338
rect 18696 17274 18748 17280
rect 18604 16992 18656 16998
rect 18604 16934 18656 16940
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18418 16416 18474 16425
rect 18418 16351 18474 16360
rect 18616 16114 18644 16934
rect 18696 16720 18748 16726
rect 18696 16662 18748 16668
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 18340 15026 18368 15982
rect 18420 15632 18472 15638
rect 18418 15600 18420 15609
rect 18472 15600 18474 15609
rect 18418 15535 18474 15544
rect 18420 15496 18472 15502
rect 18418 15464 18420 15473
rect 18604 15496 18656 15502
rect 18472 15464 18474 15473
rect 18604 15438 18656 15444
rect 18418 15399 18474 15408
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 18340 14498 18368 14962
rect 18432 14618 18460 14962
rect 18512 14816 18564 14822
rect 18512 14758 18564 14764
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 18340 14470 18460 14498
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 18144 13932 18196 13938
rect 18144 13874 18196 13880
rect 18236 13932 18288 13938
rect 18288 13892 18368 13920
rect 18236 13874 18288 13880
rect 18156 13530 18184 13874
rect 18340 13530 18368 13892
rect 18144 13524 18196 13530
rect 18144 13466 18196 13472
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 18236 13456 18288 13462
rect 18236 13398 18288 13404
rect 18248 13190 18276 13398
rect 18432 13326 18460 14470
rect 18524 13938 18552 14758
rect 18616 14346 18644 15438
rect 18708 15094 18736 16662
rect 18696 15088 18748 15094
rect 18696 15030 18748 15036
rect 18604 14340 18656 14346
rect 18604 14282 18656 14288
rect 18616 14006 18644 14282
rect 18708 14074 18736 15030
rect 18696 14068 18748 14074
rect 18696 14010 18748 14016
rect 18604 14000 18656 14006
rect 18604 13942 18656 13948
rect 18512 13932 18564 13938
rect 18512 13874 18564 13880
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18236 13184 18288 13190
rect 18236 13126 18288 13132
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 18340 12986 18368 13126
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18052 12368 18104 12374
rect 18052 12310 18104 12316
rect 18248 11830 18276 12718
rect 18326 12472 18382 12481
rect 18326 12407 18382 12416
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 17776 11086 17828 11092
rect 17880 11070 18000 11098
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17788 9722 17816 10406
rect 17880 10062 17908 11070
rect 17960 10668 18012 10674
rect 18064 10656 18092 11698
rect 18248 11665 18276 11766
rect 18234 11656 18290 11665
rect 18234 11591 18290 11600
rect 18248 11082 18276 11591
rect 18340 11218 18368 12407
rect 18616 12306 18644 13738
rect 18800 12782 18828 19314
rect 18984 19174 19012 25638
rect 19064 25424 19116 25430
rect 19062 25392 19064 25401
rect 19116 25392 19118 25401
rect 19062 25327 19118 25336
rect 19352 24818 19380 25758
rect 19536 25129 19564 26846
rect 19720 25974 19748 33050
rect 19812 32910 19840 33254
rect 19800 32904 19852 32910
rect 19800 32846 19852 32852
rect 19904 32756 19932 37198
rect 20364 35086 20392 37318
rect 20536 37256 20588 37262
rect 20536 37198 20588 37204
rect 20548 36145 20576 37198
rect 20824 36922 20852 37742
rect 21088 37460 21140 37466
rect 21088 37402 21140 37408
rect 20996 37256 21048 37262
rect 20996 37198 21048 37204
rect 20812 36916 20864 36922
rect 20812 36858 20864 36864
rect 20534 36136 20590 36145
rect 21008 36106 21036 37198
rect 21100 37194 21128 37402
rect 21088 37188 21140 37194
rect 21088 37130 21140 37136
rect 21272 36916 21324 36922
rect 21272 36858 21324 36864
rect 21284 36718 21312 36858
rect 21468 36854 21496 38150
rect 22112 38010 22140 38218
rect 22928 38208 22980 38214
rect 22928 38150 22980 38156
rect 22940 38010 22968 38150
rect 22100 38004 22152 38010
rect 22100 37946 22152 37952
rect 22928 38004 22980 38010
rect 22928 37946 22980 37952
rect 22836 37460 22888 37466
rect 22836 37402 22888 37408
rect 21548 37324 21600 37330
rect 21548 37266 21600 37272
rect 21560 37126 21588 37266
rect 22848 37194 22876 37402
rect 22940 37262 22968 37946
rect 23020 37800 23072 37806
rect 23020 37742 23072 37748
rect 22928 37256 22980 37262
rect 22928 37198 22980 37204
rect 22836 37188 22888 37194
rect 22836 37130 22888 37136
rect 21548 37120 21600 37126
rect 21548 37062 21600 37068
rect 21732 36916 21784 36922
rect 21732 36858 21784 36864
rect 21456 36848 21508 36854
rect 21456 36790 21508 36796
rect 21364 36780 21416 36786
rect 21364 36722 21416 36728
rect 21180 36712 21232 36718
rect 21180 36654 21232 36660
rect 21272 36712 21324 36718
rect 21272 36654 21324 36660
rect 21192 36378 21220 36654
rect 21272 36576 21324 36582
rect 21272 36518 21324 36524
rect 21180 36372 21232 36378
rect 21180 36314 21232 36320
rect 21284 36310 21312 36518
rect 21272 36304 21324 36310
rect 21272 36246 21324 36252
rect 20534 36071 20590 36080
rect 20996 36100 21048 36106
rect 20548 35154 20576 36071
rect 20996 36042 21048 36048
rect 20536 35148 20588 35154
rect 20536 35090 20588 35096
rect 20260 35080 20312 35086
rect 20260 35022 20312 35028
rect 20352 35080 20404 35086
rect 20352 35022 20404 35028
rect 21180 35080 21232 35086
rect 21180 35022 21232 35028
rect 20168 34944 20220 34950
rect 20168 34886 20220 34892
rect 19984 34604 20036 34610
rect 19984 34546 20036 34552
rect 19996 33114 20024 34546
rect 20076 33516 20128 33522
rect 20076 33458 20128 33464
rect 20088 33114 20116 33458
rect 20180 33402 20208 34886
rect 20272 34746 20300 35022
rect 20364 34746 20392 35022
rect 20996 34944 21048 34950
rect 20996 34886 21048 34892
rect 20260 34740 20312 34746
rect 20260 34682 20312 34688
rect 20352 34740 20404 34746
rect 20352 34682 20404 34688
rect 21008 33930 21036 34886
rect 21192 34746 21220 35022
rect 21272 34944 21324 34950
rect 21272 34886 21324 34892
rect 21180 34740 21232 34746
rect 21180 34682 21232 34688
rect 20996 33924 21048 33930
rect 20996 33866 21048 33872
rect 20180 33374 20300 33402
rect 19984 33108 20036 33114
rect 19984 33050 20036 33056
rect 20076 33108 20128 33114
rect 20076 33050 20128 33056
rect 19984 32904 20036 32910
rect 20036 32864 20208 32892
rect 19984 32846 20036 32852
rect 19904 32728 20024 32756
rect 19892 31952 19944 31958
rect 19892 31894 19944 31900
rect 19904 30122 19932 31894
rect 19892 30116 19944 30122
rect 19892 30058 19944 30064
rect 19904 29034 19932 30058
rect 19892 29028 19944 29034
rect 19892 28970 19944 28976
rect 19800 28688 19852 28694
rect 19800 28630 19852 28636
rect 19996 28642 20024 32728
rect 20076 32360 20128 32366
rect 20076 32302 20128 32308
rect 20088 30938 20116 32302
rect 20180 31686 20208 32864
rect 20168 31680 20220 31686
rect 20168 31622 20220 31628
rect 20180 31414 20208 31622
rect 20168 31408 20220 31414
rect 20168 31350 20220 31356
rect 20076 30932 20128 30938
rect 20076 30874 20128 30880
rect 20076 30796 20128 30802
rect 20076 30738 20128 30744
rect 20088 30258 20116 30738
rect 20180 30598 20208 31350
rect 20168 30592 20220 30598
rect 20168 30534 20220 30540
rect 20076 30252 20128 30258
rect 20076 30194 20128 30200
rect 19812 28558 19840 28630
rect 19996 28614 20116 28642
rect 19800 28552 19852 28558
rect 19800 28494 19852 28500
rect 19892 28552 19944 28558
rect 19892 28494 19944 28500
rect 19984 28552 20036 28558
rect 19984 28494 20036 28500
rect 19812 28064 19840 28494
rect 19904 28218 19932 28494
rect 19892 28212 19944 28218
rect 19892 28154 19944 28160
rect 19892 28076 19944 28082
rect 19812 28036 19892 28064
rect 19892 28018 19944 28024
rect 19996 28014 20024 28494
rect 19984 28008 20036 28014
rect 19984 27950 20036 27956
rect 19996 27674 20024 27950
rect 19984 27668 20036 27674
rect 19984 27610 20036 27616
rect 19892 27464 19944 27470
rect 19892 27406 19944 27412
rect 19800 26988 19852 26994
rect 19800 26930 19852 26936
rect 19812 26489 19840 26930
rect 19798 26480 19854 26489
rect 19798 26415 19854 26424
rect 19798 26344 19854 26353
rect 19904 26330 19932 27406
rect 20088 26926 20116 28614
rect 20076 26920 20128 26926
rect 20076 26862 20128 26868
rect 19854 26302 19932 26330
rect 19798 26279 19854 26288
rect 19708 25968 19760 25974
rect 19708 25910 19760 25916
rect 20088 25906 20116 26862
rect 20076 25900 20128 25906
rect 20076 25842 20128 25848
rect 20168 25900 20220 25906
rect 20168 25842 20220 25848
rect 19708 25764 19760 25770
rect 19708 25706 19760 25712
rect 19720 25498 19748 25706
rect 19984 25696 20036 25702
rect 19984 25638 20036 25644
rect 19708 25492 19760 25498
rect 19708 25434 19760 25440
rect 19996 25362 20024 25638
rect 19984 25356 20036 25362
rect 19984 25298 20036 25304
rect 19892 25288 19944 25294
rect 19890 25256 19892 25265
rect 19944 25256 19946 25265
rect 19890 25191 19946 25200
rect 19522 25120 19578 25129
rect 19522 25055 19578 25064
rect 19340 24812 19392 24818
rect 19340 24754 19392 24760
rect 19064 24404 19116 24410
rect 19064 24346 19116 24352
rect 19076 19854 19104 24346
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19444 21593 19472 22714
rect 19430 21584 19486 21593
rect 19430 21519 19432 21528
rect 19484 21519 19486 21528
rect 19432 21490 19484 21496
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19352 20534 19380 20878
rect 19432 20800 19484 20806
rect 19430 20768 19432 20777
rect 19484 20768 19486 20777
rect 19430 20703 19486 20712
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 19156 19984 19208 19990
rect 19156 19926 19208 19932
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 19076 19446 19104 19790
rect 19064 19440 19116 19446
rect 19064 19382 19116 19388
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 19064 18624 19116 18630
rect 19064 18566 19116 18572
rect 19076 18426 19104 18566
rect 19064 18420 19116 18426
rect 19064 18362 19116 18368
rect 19168 18193 19196 19926
rect 19352 19854 19380 20470
rect 19444 20466 19472 20703
rect 19536 20602 19564 25055
rect 20180 24818 20208 25842
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 19892 24608 19944 24614
rect 19892 24550 19944 24556
rect 19708 24404 19760 24410
rect 19708 24346 19760 24352
rect 19720 23186 19748 24346
rect 19708 23180 19760 23186
rect 19708 23122 19760 23128
rect 19616 22976 19668 22982
rect 19616 22918 19668 22924
rect 19524 20596 19576 20602
rect 19628 20584 19656 22918
rect 19720 22166 19748 23122
rect 19708 22160 19760 22166
rect 19708 22102 19760 22108
rect 19904 21865 19932 24550
rect 20168 24132 20220 24138
rect 20168 24074 20220 24080
rect 20076 23588 20128 23594
rect 20076 23530 20128 23536
rect 20088 23361 20116 23530
rect 20074 23352 20130 23361
rect 20180 23322 20208 24074
rect 20074 23287 20130 23296
rect 20168 23316 20220 23322
rect 20168 23258 20220 23264
rect 20180 22778 20208 23258
rect 20168 22772 20220 22778
rect 20168 22714 20220 22720
rect 20272 22438 20300 33374
rect 20812 33380 20864 33386
rect 20812 33322 20864 33328
rect 20444 32768 20496 32774
rect 20350 32736 20406 32745
rect 20444 32710 20496 32716
rect 20720 32768 20772 32774
rect 20720 32710 20772 32716
rect 20350 32671 20406 32680
rect 20364 32570 20392 32671
rect 20456 32570 20484 32710
rect 20352 32564 20404 32570
rect 20352 32506 20404 32512
rect 20444 32564 20496 32570
rect 20444 32506 20496 32512
rect 20534 32464 20590 32473
rect 20456 32434 20534 32450
rect 20444 32428 20534 32434
rect 20496 32422 20534 32428
rect 20534 32399 20590 32408
rect 20628 32428 20680 32434
rect 20444 32370 20496 32376
rect 20628 32370 20680 32376
rect 20640 31482 20668 32370
rect 20732 32026 20760 32710
rect 20720 32020 20772 32026
rect 20720 31962 20772 31968
rect 20628 31476 20680 31482
rect 20628 31418 20680 31424
rect 20352 30048 20404 30054
rect 20352 29990 20404 29996
rect 20720 30048 20772 30054
rect 20720 29990 20772 29996
rect 20364 29850 20392 29990
rect 20732 29850 20760 29990
rect 20352 29844 20404 29850
rect 20720 29844 20772 29850
rect 20404 29804 20484 29832
rect 20352 29786 20404 29792
rect 20456 29646 20484 29804
rect 20720 29786 20772 29792
rect 20444 29640 20496 29646
rect 20444 29582 20496 29588
rect 20824 29152 20852 33322
rect 21180 32972 21232 32978
rect 21180 32914 21232 32920
rect 21192 32298 21220 32914
rect 21180 32292 21232 32298
rect 21180 32234 21232 32240
rect 21284 31754 21312 34886
rect 21100 31726 21312 31754
rect 20996 30320 21048 30326
rect 20996 30262 21048 30268
rect 20904 29776 20956 29782
rect 20904 29718 20956 29724
rect 20916 29238 20944 29718
rect 21008 29646 21036 30262
rect 20996 29640 21048 29646
rect 20996 29582 21048 29588
rect 20996 29504 21048 29510
rect 20996 29446 21048 29452
rect 20904 29232 20956 29238
rect 20904 29174 20956 29180
rect 20732 29124 20852 29152
rect 20352 28416 20404 28422
rect 20352 28358 20404 28364
rect 20364 27674 20392 28358
rect 20352 27668 20404 27674
rect 20352 27610 20404 27616
rect 20732 27146 20760 29124
rect 20812 29028 20864 29034
rect 20812 28970 20864 28976
rect 20640 27118 20760 27146
rect 20640 26994 20668 27118
rect 20628 26988 20680 26994
rect 20628 26930 20680 26936
rect 20720 26988 20772 26994
rect 20720 26930 20772 26936
rect 20628 26580 20680 26586
rect 20628 26522 20680 26528
rect 20640 26042 20668 26522
rect 20732 26314 20760 26930
rect 20720 26308 20772 26314
rect 20720 26250 20772 26256
rect 20628 26036 20680 26042
rect 20628 25978 20680 25984
rect 20732 25809 20760 26250
rect 20718 25800 20774 25809
rect 20718 25735 20774 25744
rect 20536 25288 20588 25294
rect 20536 25230 20588 25236
rect 20548 24954 20576 25230
rect 20824 25226 20852 28970
rect 20812 25220 20864 25226
rect 20812 25162 20864 25168
rect 20536 24948 20588 24954
rect 20536 24890 20588 24896
rect 20718 24848 20774 24857
rect 20718 24783 20774 24792
rect 20732 24206 20760 24783
rect 20812 24744 20864 24750
rect 20812 24686 20864 24692
rect 20720 24200 20772 24206
rect 20720 24142 20772 24148
rect 20628 24064 20680 24070
rect 20628 24006 20680 24012
rect 20534 23896 20590 23905
rect 20534 23831 20590 23840
rect 20548 23662 20576 23831
rect 20640 23730 20668 24006
rect 20628 23724 20680 23730
rect 20628 23666 20680 23672
rect 20536 23656 20588 23662
rect 20536 23598 20588 23604
rect 20824 23186 20852 24686
rect 20916 23322 20944 29174
rect 21008 29034 21036 29446
rect 20996 29028 21048 29034
rect 20996 28970 21048 28976
rect 20996 26784 21048 26790
rect 20996 26726 21048 26732
rect 21008 26586 21036 26726
rect 20996 26580 21048 26586
rect 20996 26522 21048 26528
rect 20996 24268 21048 24274
rect 20996 24210 21048 24216
rect 21008 23730 21036 24210
rect 20996 23724 21048 23730
rect 20996 23666 21048 23672
rect 20904 23316 20956 23322
rect 20904 23258 20956 23264
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20824 22760 20852 23122
rect 20824 22732 20944 22760
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 20260 22432 20312 22438
rect 20260 22374 20312 22380
rect 20628 22228 20680 22234
rect 20628 22170 20680 22176
rect 20076 22160 20128 22166
rect 20076 22102 20128 22108
rect 19890 21856 19946 21865
rect 19890 21791 19946 21800
rect 19708 21548 19760 21554
rect 19708 21490 19760 21496
rect 19720 20942 19748 21490
rect 19800 21344 19852 21350
rect 19800 21286 19852 21292
rect 19708 20936 19760 20942
rect 19708 20878 19760 20884
rect 19628 20556 19748 20584
rect 19524 20538 19576 20544
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19248 19780 19300 19786
rect 19248 19722 19300 19728
rect 19260 19281 19288 19722
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19246 19272 19302 19281
rect 19246 19207 19302 19216
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19260 18329 19288 19110
rect 19352 18834 19380 19654
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19444 18714 19472 20198
rect 19536 19378 19564 20538
rect 19616 20460 19668 20466
rect 19616 20402 19668 20408
rect 19628 19786 19656 20402
rect 19616 19780 19668 19786
rect 19616 19722 19668 19728
rect 19614 19408 19670 19417
rect 19524 19372 19576 19378
rect 19720 19394 19748 20556
rect 19812 20466 19840 21286
rect 19800 20460 19852 20466
rect 19800 20402 19852 20408
rect 19812 20058 19840 20402
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19800 20052 19852 20058
rect 19800 19994 19852 20000
rect 19812 19786 19840 19994
rect 19996 19922 20024 20198
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 19800 19780 19852 19786
rect 19800 19722 19852 19728
rect 19670 19366 19748 19394
rect 19614 19343 19670 19352
rect 20088 19334 20116 22102
rect 20352 21888 20404 21894
rect 20352 21830 20404 21836
rect 20364 21554 20392 21830
rect 20640 21672 20668 22170
rect 20824 21690 20852 22578
rect 20916 22094 20944 22732
rect 21100 22658 21128 31726
rect 21180 29640 21232 29646
rect 21180 29582 21232 29588
rect 21192 28948 21220 29582
rect 21272 29572 21324 29578
rect 21272 29514 21324 29520
rect 21284 29238 21312 29514
rect 21272 29232 21324 29238
rect 21272 29174 21324 29180
rect 21376 28994 21404 36722
rect 21744 35154 21772 36858
rect 21916 36848 21968 36854
rect 21916 36790 21968 36796
rect 21928 36242 21956 36790
rect 22008 36576 22060 36582
rect 22060 36536 22140 36564
rect 22008 36518 22060 36524
rect 21916 36236 21968 36242
rect 21916 36178 21968 36184
rect 22112 36174 22140 36536
rect 22100 36168 22152 36174
rect 22100 36110 22152 36116
rect 22112 35766 22140 36110
rect 22848 36106 22876 37130
rect 22940 36786 22968 37198
rect 23032 36922 23060 37742
rect 23020 36916 23072 36922
rect 23020 36858 23072 36864
rect 22928 36780 22980 36786
rect 22928 36722 22980 36728
rect 22836 36100 22888 36106
rect 22888 36060 23060 36088
rect 22836 36042 22888 36048
rect 22100 35760 22152 35766
rect 22100 35702 22152 35708
rect 22744 35692 22796 35698
rect 22744 35634 22796 35640
rect 22468 35624 22520 35630
rect 22468 35566 22520 35572
rect 22480 35222 22508 35566
rect 22652 35488 22704 35494
rect 22652 35430 22704 35436
rect 22468 35216 22520 35222
rect 22468 35158 22520 35164
rect 21732 35148 21784 35154
rect 21732 35090 21784 35096
rect 22376 34944 22428 34950
rect 22376 34886 22428 34892
rect 22388 34746 22416 34886
rect 22480 34746 22508 35158
rect 22664 35086 22692 35430
rect 22756 35086 22784 35634
rect 22652 35080 22704 35086
rect 22652 35022 22704 35028
rect 22744 35080 22796 35086
rect 22744 35022 22796 35028
rect 22376 34740 22428 34746
rect 22376 34682 22428 34688
rect 22468 34740 22520 34746
rect 22468 34682 22520 34688
rect 21456 34536 21508 34542
rect 21456 34478 21508 34484
rect 21468 33930 21496 34478
rect 22480 34202 22508 34682
rect 22468 34196 22520 34202
rect 22468 34138 22520 34144
rect 22480 33998 22508 34138
rect 23032 34134 23060 36060
rect 23112 36032 23164 36038
rect 23112 35974 23164 35980
rect 23020 34128 23072 34134
rect 23020 34070 23072 34076
rect 22468 33992 22520 33998
rect 22468 33934 22520 33940
rect 23032 33930 23060 34070
rect 21456 33924 21508 33930
rect 21456 33866 21508 33872
rect 23020 33924 23072 33930
rect 23020 33866 23072 33872
rect 21640 33652 21692 33658
rect 21640 33594 21692 33600
rect 21456 32768 21508 32774
rect 21456 32710 21508 32716
rect 21468 32434 21496 32710
rect 21456 32428 21508 32434
rect 21456 32370 21508 32376
rect 21468 32298 21496 32370
rect 21456 32292 21508 32298
rect 21456 32234 21508 32240
rect 21456 29504 21508 29510
rect 21456 29446 21508 29452
rect 21468 29238 21496 29446
rect 21456 29232 21508 29238
rect 21456 29174 21508 29180
rect 21376 28966 21588 28994
rect 21272 28960 21324 28966
rect 21192 28920 21272 28948
rect 21272 28902 21324 28908
rect 21364 26376 21416 26382
rect 21364 26318 21416 26324
rect 21376 25498 21404 26318
rect 21364 25492 21416 25498
rect 21364 25434 21416 25440
rect 21180 24812 21232 24818
rect 21180 24754 21232 24760
rect 21192 23798 21220 24754
rect 21364 24676 21416 24682
rect 21364 24618 21416 24624
rect 21376 24206 21404 24618
rect 21364 24200 21416 24206
rect 21364 24142 21416 24148
rect 21376 23798 21404 24142
rect 21180 23792 21232 23798
rect 21180 23734 21232 23740
rect 21364 23792 21416 23798
rect 21364 23734 21416 23740
rect 21376 23662 21404 23734
rect 21364 23656 21416 23662
rect 21364 23598 21416 23604
rect 21364 23316 21416 23322
rect 21364 23258 21416 23264
rect 21376 23118 21404 23258
rect 21364 23112 21416 23118
rect 21362 23080 21364 23089
rect 21416 23080 21418 23089
rect 21272 23044 21324 23050
rect 21362 23015 21418 23024
rect 21272 22986 21324 22992
rect 21284 22681 21312 22986
rect 21008 22630 21128 22658
rect 21270 22672 21326 22681
rect 21008 22420 21036 22630
rect 21270 22607 21326 22616
rect 21088 22568 21140 22574
rect 21140 22528 21220 22556
rect 21088 22510 21140 22516
rect 21008 22392 21128 22420
rect 20996 22094 21048 22098
rect 20916 22092 21048 22094
rect 20916 22066 20996 22092
rect 20996 22034 21048 22040
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 20812 21684 20864 21690
rect 20640 21644 20760 21672
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20628 21548 20680 21554
rect 20628 21490 20680 21496
rect 20364 20913 20392 21490
rect 20640 21146 20668 21490
rect 20628 21140 20680 21146
rect 20628 21082 20680 21088
rect 20350 20904 20406 20913
rect 20350 20839 20406 20848
rect 20536 20596 20588 20602
rect 20536 20538 20588 20544
rect 19524 19314 19576 19320
rect 19352 18686 19472 18714
rect 19904 19306 20116 19334
rect 19352 18358 19380 18686
rect 19340 18352 19392 18358
rect 19246 18320 19302 18329
rect 19340 18294 19392 18300
rect 19246 18255 19302 18264
rect 19154 18184 19210 18193
rect 19154 18119 19210 18128
rect 18880 18080 18932 18086
rect 18880 18022 18932 18028
rect 18892 17796 18920 18022
rect 19156 17876 19208 17882
rect 19156 17818 19208 17824
rect 18972 17808 19024 17814
rect 18892 17768 18972 17796
rect 18892 17066 18920 17768
rect 18972 17750 19024 17756
rect 19168 17660 19196 17818
rect 19340 17672 19392 17678
rect 19168 17632 19340 17660
rect 18972 17604 19024 17610
rect 18972 17546 19024 17552
rect 18984 17202 19012 17546
rect 18972 17196 19024 17202
rect 18972 17138 19024 17144
rect 19168 17134 19196 17632
rect 19340 17614 19392 17620
rect 19156 17128 19208 17134
rect 19156 17070 19208 17076
rect 18880 17060 18932 17066
rect 18880 17002 18932 17008
rect 19168 16969 19196 17070
rect 19154 16960 19210 16969
rect 19154 16895 19210 16904
rect 18880 16788 18932 16794
rect 18880 16730 18932 16736
rect 18892 13802 18920 16730
rect 19338 16688 19394 16697
rect 19338 16623 19394 16632
rect 19352 16182 19380 16623
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19798 16552 19854 16561
rect 19340 16176 19392 16182
rect 19340 16118 19392 16124
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19246 15736 19302 15745
rect 19352 15706 19380 15982
rect 19246 15671 19302 15680
rect 19340 15700 19392 15706
rect 19064 15632 19116 15638
rect 19062 15600 19064 15609
rect 19116 15600 19118 15609
rect 19062 15535 19118 15544
rect 19154 14512 19210 14521
rect 19154 14447 19210 14456
rect 19064 13932 19116 13938
rect 19064 13874 19116 13880
rect 18880 13796 18932 13802
rect 18880 13738 18932 13744
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18604 12300 18656 12306
rect 18604 12242 18656 12248
rect 18696 12232 18748 12238
rect 18696 12174 18748 12180
rect 18788 12232 18840 12238
rect 18984 12220 19012 13194
rect 18788 12174 18840 12180
rect 18892 12192 19012 12220
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18524 11898 18552 12038
rect 18708 11898 18736 12174
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18420 11824 18472 11830
rect 18418 11792 18420 11801
rect 18472 11792 18474 11801
rect 18418 11727 18474 11736
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 18432 11354 18460 11630
rect 18604 11620 18656 11626
rect 18604 11562 18656 11568
rect 18512 11552 18564 11558
rect 18512 11494 18564 11500
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18328 11212 18380 11218
rect 18328 11154 18380 11160
rect 18420 11212 18472 11218
rect 18420 11154 18472 11160
rect 18236 11076 18288 11082
rect 18236 11018 18288 11024
rect 18012 10628 18092 10656
rect 18144 10668 18196 10674
rect 17960 10610 18012 10616
rect 18144 10610 18196 10616
rect 17960 10532 18012 10538
rect 17960 10474 18012 10480
rect 17972 10198 18000 10474
rect 18156 10266 18184 10610
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 17960 10192 18012 10198
rect 17960 10134 18012 10140
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 17960 9988 18012 9994
rect 17960 9930 18012 9936
rect 17776 9716 17828 9722
rect 17972 9674 18000 9930
rect 17776 9658 17828 9664
rect 17880 9646 18000 9674
rect 17880 9382 17908 9646
rect 18064 9586 18092 9998
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17960 9376 18012 9382
rect 18012 9336 18092 9364
rect 17960 9318 18012 9324
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17880 8634 17908 8910
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17972 8090 18000 8434
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17880 7410 17908 7822
rect 17960 7812 18012 7818
rect 17960 7754 18012 7760
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 17776 7404 17828 7410
rect 17776 7346 17828 7352
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17788 6934 17816 7346
rect 17880 7313 17908 7346
rect 17866 7304 17922 7313
rect 17866 7239 17922 7248
rect 17776 6928 17828 6934
rect 17776 6870 17828 6876
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17788 6458 17816 6870
rect 17972 6730 18000 7754
rect 18064 6798 18092 9336
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 16960 6186 16988 6394
rect 18064 6322 18092 6734
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 16948 6180 17000 6186
rect 16948 6122 17000 6128
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15016 5160 15068 5166
rect 15016 5102 15068 5108
rect 14832 5024 14884 5030
rect 14832 4966 14884 4972
rect 15028 4758 15056 5102
rect 15212 4758 15240 5510
rect 15672 5166 15700 5646
rect 16960 5642 16988 6122
rect 17052 5642 17080 6190
rect 17420 5846 17448 6258
rect 17408 5840 17460 5846
rect 17408 5782 17460 5788
rect 17420 5710 17448 5782
rect 17604 5710 17632 6258
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 16948 5636 17000 5642
rect 16948 5578 17000 5584
rect 17040 5636 17092 5642
rect 17040 5578 17092 5584
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 17052 4758 17080 5578
rect 17788 5574 17816 6258
rect 18156 6254 18184 10202
rect 18340 9674 18368 11154
rect 18432 10810 18460 11154
rect 18524 11150 18552 11494
rect 18616 11393 18644 11562
rect 18602 11384 18658 11393
rect 18602 11319 18658 11328
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18616 10810 18644 11086
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18604 10804 18656 10810
rect 18800 10792 18828 12174
rect 18892 11694 18920 12192
rect 18972 11756 19024 11762
rect 18972 11698 19024 11704
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18892 11014 18920 11630
rect 18984 11218 19012 11698
rect 18972 11212 19024 11218
rect 18972 11154 19024 11160
rect 18880 11008 18932 11014
rect 18880 10950 18932 10956
rect 18984 10849 19012 11154
rect 18970 10840 19026 10849
rect 18604 10746 18656 10752
rect 18708 10764 18828 10792
rect 18880 10804 18932 10810
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 18604 10668 18656 10674
rect 18604 10610 18656 10616
rect 18524 9722 18552 10610
rect 18248 9646 18368 9674
rect 18512 9716 18564 9722
rect 18512 9658 18564 9664
rect 18248 9081 18276 9646
rect 18510 9616 18566 9625
rect 18510 9551 18566 9560
rect 18524 9110 18552 9551
rect 18512 9104 18564 9110
rect 18234 9072 18290 9081
rect 18512 9046 18564 9052
rect 18234 9007 18290 9016
rect 18248 8090 18276 9007
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 18340 8838 18368 8910
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 18236 7948 18288 7954
rect 18236 7890 18288 7896
rect 18248 7002 18276 7890
rect 18236 6996 18288 7002
rect 18236 6938 18288 6944
rect 18340 6882 18368 8774
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18432 7750 18460 8570
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18432 7410 18460 7686
rect 18524 7546 18552 7822
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18420 7404 18472 7410
rect 18420 7346 18472 7352
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18432 6934 18460 7142
rect 18248 6866 18368 6882
rect 18420 6928 18472 6934
rect 18420 6870 18472 6876
rect 18236 6860 18368 6866
rect 18288 6854 18368 6860
rect 18236 6802 18288 6808
rect 18328 6792 18380 6798
rect 18616 6780 18644 10610
rect 18708 9110 18736 10764
rect 18970 10775 19026 10784
rect 19076 10792 19104 13874
rect 19168 11354 19196 14447
rect 19260 14414 19288 15671
rect 19340 15642 19392 15648
rect 19444 15638 19472 16526
rect 19616 16516 19668 16522
rect 19798 16487 19854 16496
rect 19616 16458 19668 16464
rect 19628 16250 19656 16458
rect 19616 16244 19668 16250
rect 19616 16186 19668 16192
rect 19708 16244 19760 16250
rect 19708 16186 19760 16192
rect 19628 16114 19656 16186
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 19616 16108 19668 16114
rect 19616 16050 19668 16056
rect 19432 15632 19484 15638
rect 19432 15574 19484 15580
rect 19536 15094 19564 16050
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 19628 15502 19656 15846
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19524 15088 19576 15094
rect 19524 15030 19576 15036
rect 19628 15026 19656 15302
rect 19720 15162 19748 16186
rect 19812 15910 19840 16487
rect 19904 16046 19932 19306
rect 20548 18834 20576 20538
rect 20640 19854 20668 21082
rect 20732 20806 20760 21644
rect 20812 21626 20864 21632
rect 20812 21548 20864 21554
rect 20812 21490 20864 21496
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20732 19990 20760 20334
rect 20720 19984 20772 19990
rect 20720 19926 20772 19932
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20732 18970 20760 19926
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 20536 18828 20588 18834
rect 20536 18770 20588 18776
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19996 18426 20024 18634
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 20444 18284 20496 18290
rect 20444 18226 20496 18232
rect 20352 17740 20404 17746
rect 20352 17682 20404 17688
rect 20364 17202 20392 17682
rect 20456 17542 20484 18226
rect 20824 18057 20852 21490
rect 20916 21078 20944 21966
rect 20904 21072 20956 21078
rect 20902 21040 20904 21049
rect 20956 21040 20958 21049
rect 20902 20975 20958 20984
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 20916 20058 20944 20334
rect 20904 20052 20956 20058
rect 20904 19994 20956 20000
rect 20916 19174 20944 19994
rect 21008 19990 21036 22034
rect 21100 21894 21128 22392
rect 21088 21888 21140 21894
rect 21088 21830 21140 21836
rect 21192 21690 21220 22528
rect 21180 21684 21232 21690
rect 21180 21626 21232 21632
rect 21088 21412 21140 21418
rect 21088 21354 21140 21360
rect 21100 20942 21128 21354
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 20996 19984 21048 19990
rect 20996 19926 21048 19932
rect 21192 19938 21220 21626
rect 21272 21140 21324 21146
rect 21272 21082 21324 21088
rect 21284 20602 21312 21082
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21468 20602 21496 20742
rect 21272 20596 21324 20602
rect 21272 20538 21324 20544
rect 21456 20596 21508 20602
rect 21456 20538 21508 20544
rect 21560 20262 21588 28966
rect 21652 24614 21680 33594
rect 21732 33108 21784 33114
rect 21732 33050 21784 33056
rect 21744 32910 21772 33050
rect 22744 33040 22796 33046
rect 22744 32982 22796 32988
rect 21732 32904 21784 32910
rect 21732 32846 21784 32852
rect 22008 32904 22060 32910
rect 22008 32846 22060 32852
rect 21744 31958 21772 32846
rect 21824 32836 21876 32842
rect 21824 32778 21876 32784
rect 21836 32745 21864 32778
rect 22020 32745 22048 32846
rect 22376 32836 22428 32842
rect 22376 32778 22428 32784
rect 22284 32768 22336 32774
rect 21822 32736 21878 32745
rect 21822 32671 21878 32680
rect 22006 32736 22062 32745
rect 22284 32710 22336 32716
rect 22006 32671 22062 32680
rect 22296 32570 22324 32710
rect 22388 32570 22416 32778
rect 21824 32564 21876 32570
rect 21824 32506 21876 32512
rect 22284 32564 22336 32570
rect 22284 32506 22336 32512
rect 22376 32564 22428 32570
rect 22376 32506 22428 32512
rect 21836 32026 21864 32506
rect 22284 32360 22336 32366
rect 22284 32302 22336 32308
rect 22008 32224 22060 32230
rect 22008 32166 22060 32172
rect 21824 32020 21876 32026
rect 21824 31962 21876 31968
rect 21732 31952 21784 31958
rect 21732 31894 21784 31900
rect 22020 31890 22048 32166
rect 22008 31884 22060 31890
rect 22008 31826 22060 31832
rect 22192 31680 22244 31686
rect 22192 31622 22244 31628
rect 22204 31346 22232 31622
rect 22296 31521 22324 32302
rect 22282 31512 22338 31521
rect 22282 31447 22338 31456
rect 22192 31340 22244 31346
rect 22192 31282 22244 31288
rect 21916 31204 21968 31210
rect 21916 31146 21968 31152
rect 21824 31136 21876 31142
rect 21824 31078 21876 31084
rect 21732 29164 21784 29170
rect 21732 29106 21784 29112
rect 21744 28762 21772 29106
rect 21732 28756 21784 28762
rect 21732 28698 21784 28704
rect 21640 24608 21692 24614
rect 21640 24550 21692 24556
rect 21836 24426 21864 31078
rect 21928 30326 21956 31146
rect 22388 30802 22416 32506
rect 22652 32496 22704 32502
rect 22650 32464 22652 32473
rect 22704 32464 22706 32473
rect 22650 32399 22706 32408
rect 22468 32224 22520 32230
rect 22468 32166 22520 32172
rect 22480 31754 22508 32166
rect 22756 31890 22784 32982
rect 23020 32904 23072 32910
rect 23020 32846 23072 32852
rect 23032 32434 23060 32846
rect 23020 32428 23072 32434
rect 23020 32370 23072 32376
rect 23020 32224 23072 32230
rect 23020 32166 23072 32172
rect 23032 32026 23060 32166
rect 23020 32020 23072 32026
rect 23020 31962 23072 31968
rect 22744 31884 22796 31890
rect 22744 31826 22796 31832
rect 22468 31748 22520 31754
rect 22468 31690 22520 31696
rect 22480 31482 22508 31690
rect 22468 31476 22520 31482
rect 22468 31418 22520 31424
rect 22376 30796 22428 30802
rect 22376 30738 22428 30744
rect 22756 30326 22784 31826
rect 23124 31754 23152 35974
rect 23400 35290 23428 38898
rect 23480 38480 23532 38486
rect 23480 38422 23532 38428
rect 23492 38282 23520 38422
rect 23480 38276 23532 38282
rect 23480 38218 23532 38224
rect 23756 37800 23808 37806
rect 23756 37742 23808 37748
rect 23664 36780 23716 36786
rect 23664 36722 23716 36728
rect 23388 35284 23440 35290
rect 23388 35226 23440 35232
rect 23296 34536 23348 34542
rect 23296 34478 23348 34484
rect 23572 34536 23624 34542
rect 23572 34478 23624 34484
rect 23308 34066 23336 34478
rect 23584 34202 23612 34478
rect 23572 34196 23624 34202
rect 23572 34138 23624 34144
rect 23296 34060 23348 34066
rect 23296 34002 23348 34008
rect 23296 33856 23348 33862
rect 23296 33798 23348 33804
rect 23204 32428 23256 32434
rect 23204 32370 23256 32376
rect 23216 32026 23244 32370
rect 23204 32020 23256 32026
rect 23204 31962 23256 31968
rect 23124 31726 23244 31754
rect 21916 30320 21968 30326
rect 21916 30262 21968 30268
rect 22744 30320 22796 30326
rect 22744 30262 22796 30268
rect 22192 29776 22244 29782
rect 22192 29718 22244 29724
rect 22006 29200 22062 29209
rect 21928 29158 22006 29186
rect 21928 29102 21956 29158
rect 22006 29135 22062 29144
rect 21916 29096 21968 29102
rect 21916 29038 21968 29044
rect 22100 29028 22152 29034
rect 22100 28970 22152 28976
rect 22112 28694 22140 28970
rect 22204 28762 22232 29718
rect 22284 28960 22336 28966
rect 22284 28902 22336 28908
rect 22192 28756 22244 28762
rect 22192 28698 22244 28704
rect 22100 28688 22152 28694
rect 22100 28630 22152 28636
rect 22204 28490 22232 28698
rect 22296 28626 22324 28902
rect 22284 28620 22336 28626
rect 22284 28562 22336 28568
rect 22192 28484 22244 28490
rect 22192 28426 22244 28432
rect 23020 28484 23072 28490
rect 23020 28426 23072 28432
rect 22468 28416 22520 28422
rect 22468 28358 22520 28364
rect 22836 28416 22888 28422
rect 22836 28358 22888 28364
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22192 27464 22244 27470
rect 22192 27406 22244 27412
rect 22204 26314 22232 27406
rect 22296 27334 22324 28018
rect 22480 28014 22508 28358
rect 22848 28082 22876 28358
rect 22836 28076 22888 28082
rect 22836 28018 22888 28024
rect 22468 28008 22520 28014
rect 22468 27950 22520 27956
rect 22480 27878 22508 27950
rect 22376 27872 22428 27878
rect 22376 27814 22428 27820
rect 22468 27872 22520 27878
rect 22468 27814 22520 27820
rect 22744 27872 22796 27878
rect 22744 27814 22796 27820
rect 22388 27674 22416 27814
rect 22376 27668 22428 27674
rect 22376 27610 22428 27616
rect 22756 27470 22784 27814
rect 23032 27606 23060 28426
rect 23112 27872 23164 27878
rect 23112 27814 23164 27820
rect 23124 27606 23152 27814
rect 23020 27600 23072 27606
rect 23020 27542 23072 27548
rect 23112 27600 23164 27606
rect 23112 27542 23164 27548
rect 22744 27464 22796 27470
rect 22744 27406 22796 27412
rect 22836 27464 22888 27470
rect 22836 27406 22888 27412
rect 22284 27328 22336 27334
rect 22848 27282 22876 27406
rect 22284 27270 22336 27276
rect 22664 27254 22876 27282
rect 22560 27124 22612 27130
rect 22560 27066 22612 27072
rect 22376 26376 22428 26382
rect 22376 26318 22428 26324
rect 22192 26308 22244 26314
rect 22192 26250 22244 26256
rect 22388 25906 22416 26318
rect 22376 25900 22428 25906
rect 22376 25842 22428 25848
rect 22192 25424 22244 25430
rect 22192 25366 22244 25372
rect 21916 25356 21968 25362
rect 21916 25298 21968 25304
rect 21744 24398 21864 24426
rect 21744 24154 21772 24398
rect 21824 24336 21876 24342
rect 21824 24278 21876 24284
rect 21652 24126 21772 24154
rect 21652 24070 21680 24126
rect 21640 24064 21692 24070
rect 21640 24006 21692 24012
rect 21640 23588 21692 23594
rect 21640 23530 21692 23536
rect 21652 20942 21680 23530
rect 21836 22094 21864 24278
rect 21744 22066 21864 22094
rect 21640 20936 21692 20942
rect 21640 20878 21692 20884
rect 21548 20256 21600 20262
rect 21548 20198 21600 20204
rect 21192 19910 21312 19938
rect 21178 19816 21234 19825
rect 21178 19751 21180 19760
rect 21232 19751 21234 19760
rect 21180 19722 21232 19728
rect 21284 19334 21312 19910
rect 21546 19408 21602 19417
rect 21546 19343 21602 19352
rect 21192 19306 21312 19334
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 21088 18896 21140 18902
rect 21088 18838 21140 18844
rect 20902 18320 20958 18329
rect 20902 18255 20958 18264
rect 20916 18222 20944 18255
rect 20904 18216 20956 18222
rect 20904 18158 20956 18164
rect 21100 18086 21128 18838
rect 21088 18080 21140 18086
rect 20810 18048 20866 18057
rect 21088 18022 21140 18028
rect 20810 17983 20866 17992
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20444 17536 20496 17542
rect 20444 17478 20496 17484
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 20456 16998 20484 17478
rect 20444 16992 20496 16998
rect 20444 16934 20496 16940
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 19892 16040 19944 16046
rect 19892 15982 19944 15988
rect 19800 15904 19852 15910
rect 19800 15846 19852 15852
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19708 15156 19760 15162
rect 19708 15098 19760 15104
rect 19812 15026 19840 15302
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19616 15020 19668 15026
rect 19616 14962 19668 14968
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19444 14822 19472 14962
rect 19708 14884 19760 14890
rect 19708 14826 19760 14832
rect 19432 14816 19484 14822
rect 19720 14793 19748 14826
rect 19432 14758 19484 14764
rect 19706 14784 19762 14793
rect 19706 14719 19762 14728
rect 19248 14408 19300 14414
rect 19248 14350 19300 14356
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19156 11348 19208 11354
rect 19156 11290 19208 11296
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 19076 10764 19196 10792
rect 18880 10746 18932 10752
rect 18892 10690 18920 10746
rect 18800 10662 18920 10690
rect 19064 10668 19116 10674
rect 18696 9104 18748 9110
rect 18696 9046 18748 9052
rect 18694 8256 18750 8265
rect 18694 8191 18750 8200
rect 18708 8090 18736 8191
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18696 7812 18748 7818
rect 18696 7754 18748 7760
rect 18708 7002 18736 7754
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 18696 6792 18748 6798
rect 18616 6752 18696 6780
rect 18328 6734 18380 6740
rect 18696 6734 18748 6740
rect 18340 6458 18368 6734
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18510 6216 18566 6225
rect 17960 6180 18012 6186
rect 17880 6140 17960 6168
rect 17880 5846 17908 6140
rect 18510 6151 18566 6160
rect 17960 6122 18012 6128
rect 18524 5846 18552 6151
rect 17868 5840 17920 5846
rect 17868 5782 17920 5788
rect 18512 5840 18564 5846
rect 18512 5782 18564 5788
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 15016 4752 15068 4758
rect 15016 4694 15068 4700
rect 15200 4752 15252 4758
rect 15200 4694 15252 4700
rect 17040 4752 17092 4758
rect 17040 4694 17092 4700
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 14556 4004 14608 4010
rect 14556 3946 14608 3952
rect 14568 3738 14596 3946
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14660 3534 14688 3878
rect 15856 3641 15884 4422
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 16120 4208 16172 4214
rect 16120 4150 16172 4156
rect 15842 3632 15898 3641
rect 15842 3567 15844 3576
rect 15896 3567 15898 3576
rect 15844 3538 15896 3544
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 15568 3392 15620 3398
rect 15568 3334 15620 3340
rect 14660 3194 14688 3334
rect 14752 3194 14780 3334
rect 14936 3194 14964 3334
rect 14648 3188 14700 3194
rect 14648 3130 14700 3136
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 15580 2990 15608 3334
rect 16132 3126 16160 4150
rect 16120 3120 16172 3126
rect 16120 3062 16172 3068
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 16224 2514 16252 4218
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16316 3738 16344 4082
rect 16684 4078 16712 4422
rect 16672 4072 16724 4078
rect 16672 4014 16724 4020
rect 17590 4040 17646 4049
rect 17590 3975 17646 3984
rect 17500 3936 17552 3942
rect 17500 3878 17552 3884
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 17512 3398 17540 3878
rect 17604 3398 17632 3975
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 16316 2854 16344 3334
rect 16960 3194 16988 3334
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17696 3126 17724 5170
rect 18800 3720 18828 10662
rect 18984 10628 19064 10656
rect 18880 10600 18932 10606
rect 18878 10568 18880 10577
rect 18932 10568 18934 10577
rect 18878 10503 18934 10512
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18892 10033 18920 10066
rect 18878 10024 18934 10033
rect 18878 9959 18934 9968
rect 18984 9674 19012 10628
rect 19064 10610 19116 10616
rect 19168 10554 19196 10764
rect 19260 10674 19288 10950
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 19076 10526 19196 10554
rect 19076 9926 19104 10526
rect 19352 10266 19380 14350
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19444 12986 19472 13126
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19616 12776 19668 12782
rect 19720 12764 19748 13126
rect 19668 12736 19748 12764
rect 19616 12718 19668 12724
rect 19524 12708 19576 12714
rect 19524 12650 19576 12656
rect 19536 12374 19564 12650
rect 19524 12368 19576 12374
rect 19524 12310 19576 12316
rect 19708 12300 19760 12306
rect 19708 12242 19760 12248
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19340 10260 19392 10266
rect 19340 10202 19392 10208
rect 19064 9920 19116 9926
rect 19064 9862 19116 9868
rect 19156 9920 19208 9926
rect 19156 9862 19208 9868
rect 18892 9646 19012 9674
rect 19076 9654 19104 9862
rect 19064 9648 19116 9654
rect 18892 5370 18920 9646
rect 19064 9590 19116 9596
rect 19168 8566 19196 9862
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19246 9072 19302 9081
rect 19246 9007 19302 9016
rect 19260 8906 19288 9007
rect 19248 8900 19300 8906
rect 19248 8842 19300 8848
rect 19156 8560 19208 8566
rect 19156 8502 19208 8508
rect 19062 8392 19118 8401
rect 19062 8327 19118 8336
rect 18970 7848 19026 7857
rect 18970 7783 19026 7792
rect 18984 7410 19012 7783
rect 19076 7750 19104 8327
rect 19064 7744 19116 7750
rect 19064 7686 19116 7692
rect 19154 7712 19210 7721
rect 19154 7647 19210 7656
rect 19168 7478 19196 7647
rect 19156 7472 19208 7478
rect 19156 7414 19208 7420
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 19062 7304 19118 7313
rect 19062 7239 19118 7248
rect 19076 7206 19104 7239
rect 18972 7200 19024 7206
rect 18972 7142 19024 7148
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 18984 6866 19012 7142
rect 18972 6860 19024 6866
rect 18972 6802 19024 6808
rect 19248 5568 19300 5574
rect 19248 5510 19300 5516
rect 18880 5364 18932 5370
rect 18880 5306 18932 5312
rect 19260 5166 19288 5510
rect 19248 5160 19300 5166
rect 19248 5102 19300 5108
rect 19352 4826 19380 9522
rect 19444 7342 19472 11086
rect 19720 11082 19748 12242
rect 19708 11076 19760 11082
rect 19708 11018 19760 11024
rect 19524 10600 19576 10606
rect 19524 10542 19576 10548
rect 19536 10062 19564 10542
rect 19614 10160 19670 10169
rect 19614 10095 19670 10104
rect 19628 10062 19656 10095
rect 19524 10056 19576 10062
rect 19524 9998 19576 10004
rect 19616 10056 19668 10062
rect 19616 9998 19668 10004
rect 19524 9920 19576 9926
rect 19524 9862 19576 9868
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 19444 6497 19472 7278
rect 19430 6488 19486 6497
rect 19430 6423 19486 6432
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19444 4622 19472 5646
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 18708 3692 18828 3720
rect 17960 3664 18012 3670
rect 17960 3606 18012 3612
rect 17972 3194 18000 3606
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 18248 2990 18276 3130
rect 18616 2990 18644 3470
rect 18236 2984 18288 2990
rect 18236 2926 18288 2932
rect 18604 2984 18656 2990
rect 18604 2926 18656 2932
rect 18708 2922 18736 3692
rect 18878 3632 18934 3641
rect 18788 3596 18840 3602
rect 18878 3567 18934 3576
rect 18788 3538 18840 3544
rect 18800 3505 18828 3538
rect 18892 3534 18920 3567
rect 18880 3528 18932 3534
rect 18786 3496 18842 3505
rect 18880 3470 18932 3476
rect 18786 3431 18842 3440
rect 19352 2990 19380 4082
rect 19536 3194 19564 9862
rect 19614 9208 19670 9217
rect 19614 9143 19670 9152
rect 19628 9110 19656 9143
rect 19616 9104 19668 9110
rect 19616 9046 19668 9052
rect 19616 8968 19668 8974
rect 19614 8936 19616 8945
rect 19668 8936 19670 8945
rect 19614 8871 19670 8880
rect 19614 8528 19670 8537
rect 19614 8463 19616 8472
rect 19668 8463 19670 8472
rect 19616 8434 19668 8440
rect 19616 8288 19668 8294
rect 19616 8230 19668 8236
rect 19628 7274 19656 8230
rect 19720 7528 19748 11018
rect 19812 9382 19840 14962
rect 19904 14618 19932 15438
rect 19892 14612 19944 14618
rect 19892 14554 19944 14560
rect 19904 14482 19932 14554
rect 19892 14476 19944 14482
rect 19892 14418 19944 14424
rect 19996 14414 20024 16594
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20076 15972 20128 15978
rect 20076 15914 20128 15920
rect 20088 15638 20116 15914
rect 20076 15632 20128 15638
rect 20076 15574 20128 15580
rect 20548 15570 20576 16050
rect 20536 15564 20588 15570
rect 20536 15506 20588 15512
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20076 15428 20128 15434
rect 20076 15370 20128 15376
rect 19984 14408 20036 14414
rect 19982 14376 19984 14385
rect 20036 14376 20038 14385
rect 19982 14311 20038 14320
rect 20088 11914 20116 15370
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 20180 14482 20208 14962
rect 20272 14657 20300 15438
rect 20536 15428 20588 15434
rect 20536 15370 20588 15376
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20258 14648 20314 14657
rect 20258 14583 20314 14592
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 20168 14000 20220 14006
rect 20220 13960 20300 13988
rect 20168 13942 20220 13948
rect 20166 13424 20222 13433
rect 20166 13359 20168 13368
rect 20220 13359 20222 13368
rect 20168 13330 20220 13336
rect 20180 13025 20208 13330
rect 20272 13161 20300 13960
rect 20258 13152 20314 13161
rect 20258 13087 20314 13096
rect 20166 13016 20222 13025
rect 20166 12951 20222 12960
rect 19904 11886 20116 11914
rect 19904 10985 19932 11886
rect 20074 11792 20130 11801
rect 20074 11727 20130 11736
rect 20088 11286 20116 11727
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20076 11280 20128 11286
rect 20076 11222 20128 11228
rect 19890 10976 19946 10985
rect 19946 10934 20024 10962
rect 19890 10911 19946 10920
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19800 9376 19852 9382
rect 19800 9318 19852 9324
rect 19800 9104 19852 9110
rect 19800 9046 19852 9052
rect 19812 8634 19840 9046
rect 19800 8628 19852 8634
rect 19800 8570 19852 8576
rect 19904 8362 19932 9998
rect 19892 8356 19944 8362
rect 19892 8298 19944 8304
rect 19800 7540 19852 7546
rect 19720 7500 19800 7528
rect 19800 7482 19852 7488
rect 19616 7268 19668 7274
rect 19616 7210 19668 7216
rect 19812 6662 19840 7482
rect 19904 7410 19932 8298
rect 19996 7546 20024 10934
rect 20180 9722 20208 11290
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 20088 8566 20116 9522
rect 20180 9110 20208 9658
rect 20272 9518 20300 13087
rect 20364 10044 20392 15098
rect 20548 15026 20576 15370
rect 20640 15201 20668 16050
rect 20732 15434 20760 17818
rect 21100 17678 21128 18022
rect 21192 17678 21220 19306
rect 21560 18766 21588 19343
rect 21548 18760 21600 18766
rect 21548 18702 21600 18708
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 21284 18086 21312 18566
rect 21744 18442 21772 22066
rect 21928 21622 21956 25298
rect 22008 25152 22060 25158
rect 22006 25120 22008 25129
rect 22100 25152 22152 25158
rect 22060 25120 22062 25129
rect 22100 25094 22152 25100
rect 22006 25055 22062 25064
rect 22008 24812 22060 24818
rect 22008 24754 22060 24760
rect 22020 24614 22048 24754
rect 22008 24608 22060 24614
rect 22008 24550 22060 24556
rect 22112 24342 22140 25094
rect 22204 24954 22232 25366
rect 22192 24948 22244 24954
rect 22192 24890 22244 24896
rect 22100 24336 22152 24342
rect 22100 24278 22152 24284
rect 22572 24274 22600 27066
rect 22560 24268 22612 24274
rect 22560 24210 22612 24216
rect 22284 24200 22336 24206
rect 22284 24142 22336 24148
rect 22296 23633 22324 24142
rect 22468 24064 22520 24070
rect 22468 24006 22520 24012
rect 22282 23624 22338 23633
rect 22282 23559 22338 23568
rect 22480 23497 22508 24006
rect 22466 23488 22522 23497
rect 22466 23423 22522 23432
rect 22100 23316 22152 23322
rect 22100 23258 22152 23264
rect 22112 22710 22140 23258
rect 22100 22704 22152 22710
rect 22100 22646 22152 22652
rect 22008 22636 22060 22642
rect 22008 22578 22060 22584
rect 22020 22098 22048 22578
rect 22008 22092 22060 22098
rect 22008 22034 22060 22040
rect 22112 22030 22140 22646
rect 22284 22636 22336 22642
rect 22204 22596 22284 22624
rect 22204 22166 22232 22596
rect 22284 22578 22336 22584
rect 22284 22500 22336 22506
rect 22284 22442 22336 22448
rect 22376 22500 22428 22506
rect 22376 22442 22428 22448
rect 22192 22160 22244 22166
rect 22192 22102 22244 22108
rect 22204 22030 22232 22102
rect 22100 22024 22152 22030
rect 22192 22024 22244 22030
rect 22100 21966 22152 21972
rect 22190 21992 22192 22001
rect 22244 21992 22246 22001
rect 22190 21927 22246 21936
rect 21916 21616 21968 21622
rect 21916 21558 21968 21564
rect 22296 20262 22324 22442
rect 22388 21962 22416 22442
rect 22376 21956 22428 21962
rect 22376 21898 22428 21904
rect 22572 21146 22600 24210
rect 22560 21140 22612 21146
rect 22560 21082 22612 21088
rect 22560 20800 22612 20806
rect 22560 20742 22612 20748
rect 22572 20466 22600 20742
rect 22560 20460 22612 20466
rect 22560 20402 22612 20408
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 22284 20256 22336 20262
rect 22284 20198 22336 20204
rect 21824 19848 21876 19854
rect 21824 19790 21876 19796
rect 21836 19514 21864 19790
rect 22204 19514 22232 20198
rect 21824 19508 21876 19514
rect 21824 19450 21876 19456
rect 22192 19508 22244 19514
rect 22192 19450 22244 19456
rect 22572 19417 22600 20402
rect 22558 19408 22614 19417
rect 22100 19372 22152 19378
rect 22558 19343 22614 19352
rect 22100 19314 22152 19320
rect 22112 18970 22140 19314
rect 22284 19236 22336 19242
rect 22284 19178 22336 19184
rect 22100 18964 22152 18970
rect 22100 18906 22152 18912
rect 22112 18766 22140 18906
rect 22296 18766 22324 19178
rect 22664 18834 22692 27254
rect 23032 26994 23060 27542
rect 23112 27396 23164 27402
rect 23112 27338 23164 27344
rect 22928 26988 22980 26994
rect 22928 26930 22980 26936
rect 23020 26988 23072 26994
rect 23020 26930 23072 26936
rect 22940 26586 22968 26930
rect 22928 26580 22980 26586
rect 22928 26522 22980 26528
rect 22836 24948 22888 24954
rect 22836 24890 22888 24896
rect 22848 24138 22876 24890
rect 22928 24812 22980 24818
rect 22928 24754 22980 24760
rect 23032 24800 23060 26930
rect 23124 26858 23152 27338
rect 23112 26852 23164 26858
rect 23112 26794 23164 26800
rect 23216 25974 23244 31726
rect 23308 26518 23336 33798
rect 23480 32768 23532 32774
rect 23480 32710 23532 32716
rect 23388 32360 23440 32366
rect 23388 32302 23440 32308
rect 23400 31822 23428 32302
rect 23492 32230 23520 32710
rect 23572 32428 23624 32434
rect 23572 32370 23624 32376
rect 23584 32230 23612 32370
rect 23480 32224 23532 32230
rect 23480 32166 23532 32172
rect 23572 32224 23624 32230
rect 23572 32166 23624 32172
rect 23388 31816 23440 31822
rect 23440 31776 23520 31804
rect 23388 31758 23440 31764
rect 23388 30320 23440 30326
rect 23388 30262 23440 30268
rect 23400 29850 23428 30262
rect 23492 30258 23520 31776
rect 23572 30592 23624 30598
rect 23572 30534 23624 30540
rect 23480 30252 23532 30258
rect 23480 30194 23532 30200
rect 23584 30190 23612 30534
rect 23676 30433 23704 36722
rect 23768 35154 23796 37742
rect 23756 35148 23808 35154
rect 23756 35090 23808 35096
rect 23768 34406 23796 35090
rect 23756 34400 23808 34406
rect 23756 34342 23808 34348
rect 23848 33108 23900 33114
rect 23848 33050 23900 33056
rect 23860 32502 23888 33050
rect 23848 32496 23900 32502
rect 23848 32438 23900 32444
rect 23756 32292 23808 32298
rect 23756 32234 23808 32240
rect 23768 31958 23796 32234
rect 23756 31952 23808 31958
rect 23756 31894 23808 31900
rect 23768 31822 23796 31894
rect 23756 31816 23808 31822
rect 23756 31758 23808 31764
rect 23662 30424 23718 30433
rect 23662 30359 23718 30368
rect 23768 30258 23796 31758
rect 23756 30252 23808 30258
rect 23756 30194 23808 30200
rect 23572 30184 23624 30190
rect 23572 30126 23624 30132
rect 23480 30116 23532 30122
rect 23480 30058 23532 30064
rect 23388 29844 23440 29850
rect 23388 29786 23440 29792
rect 23492 29646 23520 30058
rect 23480 29640 23532 29646
rect 23480 29582 23532 29588
rect 23388 29028 23440 29034
rect 23388 28970 23440 28976
rect 23584 28994 23612 30126
rect 23768 29646 23796 30194
rect 23848 30184 23900 30190
rect 23848 30126 23900 30132
rect 23756 29640 23808 29646
rect 23756 29582 23808 29588
rect 23860 29510 23888 30126
rect 23848 29504 23900 29510
rect 23848 29446 23900 29452
rect 23296 26512 23348 26518
rect 23296 26454 23348 26460
rect 23204 25968 23256 25974
rect 23204 25910 23256 25916
rect 23204 25220 23256 25226
rect 23204 25162 23256 25168
rect 23112 24812 23164 24818
rect 23032 24772 23112 24800
rect 22940 24206 22968 24754
rect 23032 24342 23060 24772
rect 23112 24754 23164 24760
rect 23112 24608 23164 24614
rect 23112 24550 23164 24556
rect 23020 24336 23072 24342
rect 23020 24278 23072 24284
rect 22928 24200 22980 24206
rect 22928 24142 22980 24148
rect 22836 24132 22888 24138
rect 22836 24074 22888 24080
rect 23032 23066 23060 24278
rect 22848 23038 23060 23066
rect 22744 22976 22796 22982
rect 22744 22918 22796 22924
rect 22756 22817 22784 22918
rect 22742 22808 22798 22817
rect 22742 22743 22798 22752
rect 22744 22704 22796 22710
rect 22744 22646 22796 22652
rect 22756 21554 22784 22646
rect 22848 22094 22876 23038
rect 23020 22636 23072 22642
rect 23020 22578 23072 22584
rect 23032 22234 23060 22578
rect 23020 22228 23072 22234
rect 23020 22170 23072 22176
rect 22848 22066 22968 22094
rect 22744 21548 22796 21554
rect 22744 21490 22796 21496
rect 22652 18828 22704 18834
rect 22652 18770 22704 18776
rect 22100 18760 22152 18766
rect 22100 18702 22152 18708
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 22376 18760 22428 18766
rect 22376 18702 22428 18708
rect 22468 18760 22520 18766
rect 22468 18702 22520 18708
rect 21822 18456 21878 18465
rect 21744 18414 21822 18442
rect 21822 18391 21878 18400
rect 21364 18284 21416 18290
rect 21364 18226 21416 18232
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21272 18080 21324 18086
rect 21272 18022 21324 18028
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 21088 17672 21140 17678
rect 21088 17614 21140 17620
rect 21180 17672 21232 17678
rect 21180 17614 21232 17620
rect 20824 17338 20852 17614
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 21192 17338 21220 17478
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 21180 17332 21232 17338
rect 21180 17274 21232 17280
rect 20812 16720 20864 16726
rect 20812 16662 20864 16668
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20626 15192 20682 15201
rect 20626 15127 20628 15136
rect 20680 15127 20682 15136
rect 20628 15098 20680 15104
rect 20824 15094 20852 16662
rect 20904 16516 20956 16522
rect 20904 16458 20956 16464
rect 20916 16114 20944 16458
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20904 15904 20956 15910
rect 20904 15846 20956 15852
rect 20916 15366 20944 15846
rect 21284 15502 21312 18022
rect 21376 16114 21404 18226
rect 21548 17196 21600 17202
rect 21548 17138 21600 17144
rect 21364 16108 21416 16114
rect 21364 16050 21416 16056
rect 21376 15638 21404 16050
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21468 15706 21496 15846
rect 21560 15745 21588 17138
rect 21640 16176 21692 16182
rect 21640 16118 21692 16124
rect 21546 15736 21602 15745
rect 21456 15700 21508 15706
rect 21546 15671 21602 15680
rect 21456 15642 21508 15648
rect 21364 15632 21416 15638
rect 21364 15574 21416 15580
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 20904 15360 20956 15366
rect 20904 15302 20956 15308
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20628 15020 20680 15026
rect 20628 14962 20680 14968
rect 20640 14793 20668 14962
rect 20720 14884 20772 14890
rect 20720 14826 20772 14832
rect 20626 14784 20682 14793
rect 20626 14719 20682 14728
rect 20536 14544 20588 14550
rect 20456 14492 20536 14498
rect 20456 14486 20588 14492
rect 20456 14470 20576 14486
rect 20456 14346 20484 14470
rect 20732 14414 20760 14826
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 20536 14340 20588 14346
rect 20536 14282 20588 14288
rect 20456 14006 20484 14282
rect 20444 14000 20496 14006
rect 20444 13942 20496 13948
rect 20548 13870 20576 14282
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20732 12170 20760 13466
rect 20824 13190 20852 15030
rect 20916 14278 20944 15302
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 21008 14618 21036 15098
rect 21284 14958 21312 15438
rect 21180 14952 21232 14958
rect 21180 14894 21232 14900
rect 21272 14952 21324 14958
rect 21272 14894 21324 14900
rect 21192 14770 21220 14894
rect 21192 14742 21312 14770
rect 20996 14612 21048 14618
rect 20996 14554 21048 14560
rect 21284 14346 21312 14742
rect 21180 14340 21232 14346
rect 21180 14282 21232 14288
rect 21272 14340 21324 14346
rect 21272 14282 21324 14288
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 21192 13988 21220 14282
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 21192 13960 21312 13988
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 21088 13932 21140 13938
rect 21140 13892 21220 13920
rect 21088 13874 21140 13880
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 20824 12306 20852 13126
rect 20916 12434 20944 13874
rect 21192 12442 21220 13892
rect 21180 12436 21232 12442
rect 20916 12406 21036 12434
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20720 12164 20772 12170
rect 20720 12106 20772 12112
rect 20904 12164 20956 12170
rect 20904 12106 20956 12112
rect 20732 11218 20760 12106
rect 20916 11830 20944 12106
rect 20904 11824 20956 11830
rect 20904 11766 20956 11772
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20720 11212 20772 11218
rect 20640 11172 20720 11200
rect 20536 10804 20588 10810
rect 20536 10746 20588 10752
rect 20548 10538 20576 10746
rect 20536 10532 20588 10538
rect 20536 10474 20588 10480
rect 20444 10056 20496 10062
rect 20364 10016 20444 10044
rect 20260 9512 20312 9518
rect 20260 9454 20312 9460
rect 20364 9330 20392 10016
rect 20444 9998 20496 10004
rect 20444 9920 20496 9926
rect 20444 9862 20496 9868
rect 20456 9518 20484 9862
rect 20444 9512 20496 9518
rect 20640 9466 20668 11172
rect 20720 11154 20772 11160
rect 20824 10742 20852 11494
rect 20916 11218 20944 11766
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 20904 11076 20956 11082
rect 20904 11018 20956 11024
rect 20916 10810 20944 11018
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 20812 10736 20864 10742
rect 20812 10678 20864 10684
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 20444 9454 20496 9460
rect 20272 9302 20392 9330
rect 20548 9438 20668 9466
rect 20168 9104 20220 9110
rect 20168 9046 20220 9052
rect 20076 8560 20128 8566
rect 20076 8502 20128 8508
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 20088 7274 20116 8502
rect 20272 8498 20300 9302
rect 20548 9194 20576 9438
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20456 9178 20576 9194
rect 20444 9172 20576 9178
rect 20496 9166 20576 9172
rect 20444 9114 20496 9120
rect 20456 8838 20484 9114
rect 20536 9104 20588 9110
rect 20534 9072 20536 9081
rect 20588 9072 20590 9081
rect 20534 9007 20590 9016
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 20444 8832 20496 8838
rect 20444 8774 20496 8780
rect 20442 8664 20498 8673
rect 20442 8599 20498 8608
rect 20352 8560 20404 8566
rect 20352 8502 20404 8508
rect 20260 8492 20312 8498
rect 20260 8434 20312 8440
rect 20168 8356 20220 8362
rect 20168 8298 20220 8304
rect 20180 8022 20208 8298
rect 20168 8016 20220 8022
rect 20168 7958 20220 7964
rect 20076 7268 20128 7274
rect 20076 7210 20128 7216
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 19800 6656 19852 6662
rect 19800 6598 19852 6604
rect 20088 6458 20116 6734
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 19616 5568 19668 5574
rect 19616 5510 19668 5516
rect 19628 5370 19656 5510
rect 19616 5364 19668 5370
rect 19616 5306 19668 5312
rect 19892 5024 19944 5030
rect 19892 4966 19944 4972
rect 19904 4690 19932 4966
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 20180 4622 20208 7958
rect 20272 7206 20300 8434
rect 20364 7206 20392 8502
rect 20456 7886 20484 8599
rect 20548 8090 20576 8910
rect 20536 8084 20588 8090
rect 20536 8026 20588 8032
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20548 7546 20576 7822
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20640 7426 20668 9318
rect 20732 7585 20760 10610
rect 21008 10146 21036 12406
rect 21180 12378 21232 12384
rect 21192 12170 21220 12378
rect 21284 12238 21312 13960
rect 21376 13938 21404 14214
rect 21364 13932 21416 13938
rect 21364 13874 21416 13880
rect 21376 13258 21404 13874
rect 21364 13252 21416 13258
rect 21364 13194 21416 13200
rect 21376 12986 21404 13194
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21272 12232 21324 12238
rect 21324 12192 21496 12220
rect 21272 12174 21324 12180
rect 21180 12164 21232 12170
rect 21180 12106 21232 12112
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 21100 10266 21128 10610
rect 21088 10260 21140 10266
rect 21088 10202 21140 10208
rect 21008 10118 21128 10146
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20824 8945 20852 9318
rect 20810 8936 20866 8945
rect 20810 8871 20812 8880
rect 20864 8871 20866 8880
rect 20812 8842 20864 8848
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 20824 7800 20852 8570
rect 20916 8537 20944 9658
rect 20994 9208 21050 9217
rect 20994 9143 20996 9152
rect 21048 9143 21050 9152
rect 20996 9114 21048 9120
rect 20902 8528 20958 8537
rect 20902 8463 20904 8472
rect 20956 8463 20958 8472
rect 20904 8434 20956 8440
rect 20904 7812 20956 7818
rect 20824 7772 20904 7800
rect 20904 7754 20956 7760
rect 20718 7576 20774 7585
rect 20718 7511 20774 7520
rect 20720 7472 20772 7478
rect 20640 7420 20720 7426
rect 20640 7414 20772 7420
rect 20536 7404 20588 7410
rect 20640 7398 20760 7414
rect 20536 7346 20588 7352
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 20272 6866 20300 7142
rect 20260 6860 20312 6866
rect 20260 6802 20312 6808
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 19708 4480 19760 4486
rect 19708 4422 19760 4428
rect 19720 3398 19748 4422
rect 20364 4010 20392 7142
rect 20548 7002 20576 7346
rect 20536 6996 20588 7002
rect 20536 6938 20588 6944
rect 20916 6730 20944 7754
rect 20628 6724 20680 6730
rect 20628 6666 20680 6672
rect 20904 6724 20956 6730
rect 20904 6666 20956 6672
rect 20352 4004 20404 4010
rect 20352 3946 20404 3952
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 19812 3602 19840 3878
rect 19800 3596 19852 3602
rect 19800 3538 19852 3544
rect 20640 3534 20668 6666
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 20732 4622 20760 4966
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 21008 4214 21036 9114
rect 21100 8634 21128 10118
rect 21192 9081 21220 12106
rect 21272 11144 21324 11150
rect 21468 11121 21496 12192
rect 21560 11830 21588 15671
rect 21548 11824 21600 11830
rect 21548 11766 21600 11772
rect 21652 11286 21680 16118
rect 21836 15706 21864 18226
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22204 17660 22232 18022
rect 22284 17672 22336 17678
rect 22204 17632 22284 17660
rect 22204 17134 22232 17632
rect 22284 17614 22336 17620
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 22192 17128 22244 17134
rect 22192 17070 22244 17076
rect 22100 16584 22152 16590
rect 22204 16572 22232 17070
rect 22296 16590 22324 17206
rect 22152 16544 22232 16572
rect 22284 16584 22336 16590
rect 22100 16526 22152 16532
rect 22284 16526 22336 16532
rect 22388 16250 22416 18702
rect 22480 18426 22508 18702
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 22940 18222 22968 22066
rect 23020 18624 23072 18630
rect 23020 18566 23072 18572
rect 22928 18216 22980 18222
rect 22928 18158 22980 18164
rect 22940 17921 22968 18158
rect 22926 17912 22982 17921
rect 22926 17847 22982 17856
rect 23032 17796 23060 18566
rect 23124 18170 23152 24550
rect 23216 24206 23244 25162
rect 23400 24886 23428 28970
rect 23584 28966 23888 28994
rect 23480 28688 23532 28694
rect 23480 28630 23532 28636
rect 23492 26450 23520 28630
rect 23860 28558 23888 28966
rect 23848 28552 23900 28558
rect 23848 28494 23900 28500
rect 23860 26518 23888 28494
rect 23952 27962 23980 38966
rect 25228 38956 25280 38962
rect 25228 38898 25280 38904
rect 27252 38956 27304 38962
rect 27252 38898 27304 38904
rect 33600 38956 33652 38962
rect 33600 38898 33652 38904
rect 24032 38344 24084 38350
rect 24032 38286 24084 38292
rect 24044 38010 24072 38286
rect 24124 38276 24176 38282
rect 24124 38218 24176 38224
rect 24032 38004 24084 38010
rect 24032 37946 24084 37952
rect 24136 34678 24164 38218
rect 25044 38208 25096 38214
rect 25044 38150 25096 38156
rect 25056 38010 25084 38150
rect 25240 38010 25268 38898
rect 26056 38208 26108 38214
rect 26056 38150 26108 38156
rect 25044 38004 25096 38010
rect 25044 37946 25096 37952
rect 25228 38004 25280 38010
rect 25228 37946 25280 37952
rect 24860 37800 24912 37806
rect 24860 37742 24912 37748
rect 24676 37392 24728 37398
rect 24676 37334 24728 37340
rect 24400 34944 24452 34950
rect 24400 34886 24452 34892
rect 24124 34672 24176 34678
rect 24124 34614 24176 34620
rect 24412 33998 24440 34886
rect 24400 33992 24452 33998
rect 24400 33934 24452 33940
rect 24124 33856 24176 33862
rect 24124 33798 24176 33804
rect 24136 32502 24164 33798
rect 24688 33658 24716 37334
rect 24872 36378 24900 37742
rect 24952 37664 25004 37670
rect 24952 37606 25004 37612
rect 24860 36372 24912 36378
rect 24860 36314 24912 36320
rect 24964 36145 24992 37606
rect 25056 37210 25084 37946
rect 25596 37868 25648 37874
rect 25596 37810 25648 37816
rect 25688 37868 25740 37874
rect 25688 37810 25740 37816
rect 25056 37194 25176 37210
rect 25056 37188 25188 37194
rect 25056 37182 25136 37188
rect 25136 37130 25188 37136
rect 25136 36780 25188 36786
rect 25136 36722 25188 36728
rect 24950 36136 25006 36145
rect 24950 36071 25006 36080
rect 24676 33652 24728 33658
rect 24676 33594 24728 33600
rect 24216 32768 24268 32774
rect 24216 32710 24268 32716
rect 24308 32768 24360 32774
rect 24308 32710 24360 32716
rect 24124 32496 24176 32502
rect 24124 32438 24176 32444
rect 24228 32230 24256 32710
rect 24124 32224 24176 32230
rect 24124 32166 24176 32172
rect 24216 32224 24268 32230
rect 24216 32166 24268 32172
rect 24136 31346 24164 32166
rect 24124 31340 24176 31346
rect 24124 31282 24176 31288
rect 24032 30048 24084 30054
rect 24032 29990 24084 29996
rect 24124 30048 24176 30054
rect 24124 29990 24176 29996
rect 24044 29850 24072 29990
rect 24032 29844 24084 29850
rect 24032 29786 24084 29792
rect 24136 29102 24164 29990
rect 24124 29096 24176 29102
rect 24124 29038 24176 29044
rect 23952 27934 24072 27962
rect 23940 27872 23992 27878
rect 23940 27814 23992 27820
rect 23848 26512 23900 26518
rect 23848 26454 23900 26460
rect 23480 26444 23532 26450
rect 23480 26386 23532 26392
rect 23492 25906 23520 26386
rect 23848 26376 23900 26382
rect 23848 26318 23900 26324
rect 23860 26042 23888 26318
rect 23848 26036 23900 26042
rect 23848 25978 23900 25984
rect 23480 25900 23532 25906
rect 23480 25842 23532 25848
rect 23756 25288 23808 25294
rect 23756 25230 23808 25236
rect 23388 24880 23440 24886
rect 23388 24822 23440 24828
rect 23768 24818 23796 25230
rect 23848 24880 23900 24886
rect 23848 24822 23900 24828
rect 23572 24812 23624 24818
rect 23572 24754 23624 24760
rect 23756 24812 23808 24818
rect 23756 24754 23808 24760
rect 23388 24744 23440 24750
rect 23388 24686 23440 24692
rect 23204 24200 23256 24206
rect 23204 24142 23256 24148
rect 23400 23769 23428 24686
rect 23480 24608 23532 24614
rect 23480 24550 23532 24556
rect 23386 23760 23442 23769
rect 23386 23695 23442 23704
rect 23388 23180 23440 23186
rect 23388 23122 23440 23128
rect 23296 23112 23348 23118
rect 23296 23054 23348 23060
rect 23308 22642 23336 23054
rect 23400 22642 23428 23122
rect 23296 22636 23348 22642
rect 23296 22578 23348 22584
rect 23388 22636 23440 22642
rect 23388 22578 23440 22584
rect 23204 22432 23256 22438
rect 23204 22374 23256 22380
rect 23216 21690 23244 22374
rect 23308 22166 23336 22578
rect 23296 22160 23348 22166
rect 23296 22102 23348 22108
rect 23204 21684 23256 21690
rect 23204 21626 23256 21632
rect 23308 21554 23336 22102
rect 23388 22092 23440 22098
rect 23388 22034 23440 22040
rect 23400 21690 23428 22034
rect 23388 21684 23440 21690
rect 23388 21626 23440 21632
rect 23296 21548 23348 21554
rect 23296 21490 23348 21496
rect 23492 20806 23520 24550
rect 23584 23730 23612 24754
rect 23664 24336 23716 24342
rect 23664 24278 23716 24284
rect 23572 23724 23624 23730
rect 23572 23666 23624 23672
rect 23676 23633 23704 24278
rect 23860 23798 23888 24822
rect 23952 23905 23980 27814
rect 24044 24818 24072 27934
rect 24228 26874 24256 32166
rect 24320 28218 24348 32710
rect 24400 32428 24452 32434
rect 24400 32370 24452 32376
rect 24584 32428 24636 32434
rect 24584 32370 24636 32376
rect 24412 32065 24440 32370
rect 24596 32212 24624 32370
rect 24504 32184 24624 32212
rect 24398 32056 24454 32065
rect 24398 31991 24454 32000
rect 24400 31680 24452 31686
rect 24400 31622 24452 31628
rect 24412 31482 24440 31622
rect 24400 31476 24452 31482
rect 24400 31418 24452 31424
rect 24504 31346 24532 32184
rect 24584 31884 24636 31890
rect 24584 31826 24636 31832
rect 24492 31340 24544 31346
rect 24492 31282 24544 31288
rect 24400 28416 24452 28422
rect 24400 28358 24452 28364
rect 24412 28218 24440 28358
rect 24308 28212 24360 28218
rect 24308 28154 24360 28160
rect 24400 28212 24452 28218
rect 24400 28154 24452 28160
rect 24400 27600 24452 27606
rect 24400 27542 24452 27548
rect 24228 26846 24348 26874
rect 24124 26784 24176 26790
rect 24124 26726 24176 26732
rect 24136 26194 24164 26726
rect 24214 26344 24270 26353
rect 24214 26279 24216 26288
rect 24268 26279 24270 26288
rect 24216 26250 24268 26256
rect 24136 26166 24256 26194
rect 24124 25696 24176 25702
rect 24124 25638 24176 25644
rect 24136 24993 24164 25638
rect 24122 24984 24178 24993
rect 24122 24919 24178 24928
rect 24032 24812 24084 24818
rect 24032 24754 24084 24760
rect 24124 24812 24176 24818
rect 24124 24754 24176 24760
rect 23938 23896 23994 23905
rect 24044 23866 24072 24754
rect 24136 24721 24164 24754
rect 24122 24712 24178 24721
rect 24122 24647 24178 24656
rect 24136 23905 24164 24647
rect 24228 24206 24256 26166
rect 24216 24200 24268 24206
rect 24216 24142 24268 24148
rect 24122 23896 24178 23905
rect 23938 23831 23994 23840
rect 24032 23860 24084 23866
rect 23848 23792 23900 23798
rect 23848 23734 23900 23740
rect 23756 23724 23808 23730
rect 23756 23666 23808 23672
rect 23662 23624 23718 23633
rect 23662 23559 23718 23568
rect 23768 23497 23796 23666
rect 23754 23488 23810 23497
rect 23754 23423 23810 23432
rect 23848 23112 23900 23118
rect 23848 23054 23900 23060
rect 23860 22778 23888 23054
rect 23848 22772 23900 22778
rect 23848 22714 23900 22720
rect 23572 22636 23624 22642
rect 23572 22578 23624 22584
rect 23584 21962 23612 22578
rect 23572 21956 23624 21962
rect 23572 21898 23624 21904
rect 23480 20800 23532 20806
rect 23480 20742 23532 20748
rect 23952 20602 23980 23831
rect 24122 23831 24178 23840
rect 24032 23802 24084 23808
rect 24228 23798 24256 24142
rect 24216 23792 24268 23798
rect 24216 23734 24268 23740
rect 24216 23520 24268 23526
rect 24216 23462 24268 23468
rect 24124 22636 24176 22642
rect 24124 22578 24176 22584
rect 24136 22030 24164 22578
rect 24124 22024 24176 22030
rect 24124 21966 24176 21972
rect 24136 21486 24164 21966
rect 24124 21480 24176 21486
rect 24124 21422 24176 21428
rect 24032 20936 24084 20942
rect 24032 20878 24084 20884
rect 24044 20602 24072 20878
rect 24228 20806 24256 23462
rect 24216 20800 24268 20806
rect 24216 20742 24268 20748
rect 23940 20596 23992 20602
rect 23940 20538 23992 20544
rect 24032 20596 24084 20602
rect 24032 20538 24084 20544
rect 24216 20392 24268 20398
rect 24216 20334 24268 20340
rect 24228 20058 24256 20334
rect 24216 20052 24268 20058
rect 24216 19994 24268 20000
rect 24032 19780 24084 19786
rect 24032 19722 24084 19728
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 23676 19378 23704 19654
rect 23664 19372 23716 19378
rect 23664 19314 23716 19320
rect 23480 18216 23532 18222
rect 23124 18142 23336 18170
rect 23480 18158 23532 18164
rect 22940 17768 23060 17796
rect 22940 17649 22968 17768
rect 23020 17672 23072 17678
rect 22926 17640 22982 17649
rect 22744 17604 22796 17610
rect 22664 17564 22744 17592
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 22192 16108 22244 16114
rect 22192 16050 22244 16056
rect 21824 15700 21876 15706
rect 21824 15642 21876 15648
rect 21732 15020 21784 15026
rect 21732 14962 21784 14968
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 21744 14770 21772 14962
rect 21928 14929 21956 14962
rect 21914 14920 21970 14929
rect 21914 14855 21970 14864
rect 21744 14742 21864 14770
rect 21732 14612 21784 14618
rect 21732 14554 21784 14560
rect 21744 14074 21772 14554
rect 21732 14068 21784 14074
rect 21732 14010 21784 14016
rect 21836 11370 21864 14742
rect 21916 14408 21968 14414
rect 21916 14350 21968 14356
rect 21928 14074 21956 14350
rect 22112 14346 22140 16050
rect 22204 15706 22232 16050
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22376 15700 22428 15706
rect 22376 15642 22428 15648
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 22296 15026 22324 15438
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22192 14816 22244 14822
rect 22192 14758 22244 14764
rect 22204 14414 22232 14758
rect 22192 14408 22244 14414
rect 22192 14350 22244 14356
rect 22100 14340 22152 14346
rect 22100 14282 22152 14288
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 22296 13938 22324 14962
rect 21916 13932 21968 13938
rect 21916 13874 21968 13880
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 21928 11665 21956 13874
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 22192 12640 22244 12646
rect 22296 12617 22324 12786
rect 22192 12582 22244 12588
rect 22282 12608 22338 12617
rect 22204 12458 22232 12582
rect 22282 12543 22338 12552
rect 22388 12458 22416 15642
rect 22480 14822 22508 17478
rect 22572 17202 22600 17478
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22572 16590 22600 17138
rect 22664 16658 22692 17564
rect 23020 17614 23072 17620
rect 22926 17575 22928 17584
rect 22744 17546 22796 17552
rect 22980 17575 22982 17584
rect 22928 17546 22980 17552
rect 22836 17060 22888 17066
rect 22836 17002 22888 17008
rect 22652 16652 22704 16658
rect 22652 16594 22704 16600
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 22664 16454 22692 16594
rect 22848 16590 22876 17002
rect 22836 16584 22888 16590
rect 22836 16526 22888 16532
rect 22652 16448 22704 16454
rect 22652 16390 22704 16396
rect 22744 16448 22796 16454
rect 22744 16390 22796 16396
rect 22558 15600 22614 15609
rect 22558 15535 22560 15544
rect 22612 15535 22614 15544
rect 22560 15506 22612 15512
rect 22468 14816 22520 14822
rect 22520 14776 22600 14804
rect 22468 14758 22520 14764
rect 22468 14408 22520 14414
rect 22468 14350 22520 14356
rect 22480 14074 22508 14350
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 22468 13932 22520 13938
rect 22468 13874 22520 13880
rect 22204 12430 22416 12458
rect 22192 12164 22244 12170
rect 22192 12106 22244 12112
rect 22098 11928 22154 11937
rect 22098 11863 22154 11872
rect 22112 11830 22140 11863
rect 22204 11830 22232 12106
rect 22296 11830 22324 12430
rect 22376 12232 22428 12238
rect 22374 12200 22376 12209
rect 22428 12200 22430 12209
rect 22374 12135 22430 12144
rect 22480 11898 22508 13874
rect 22572 12889 22600 14776
rect 22652 13932 22704 13938
rect 22652 13874 22704 13880
rect 22664 13326 22692 13874
rect 22652 13320 22704 13326
rect 22652 13262 22704 13268
rect 22558 12880 22614 12889
rect 22558 12815 22614 12824
rect 22560 12232 22612 12238
rect 22560 12174 22612 12180
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22100 11824 22152 11830
rect 22100 11766 22152 11772
rect 22192 11824 22244 11830
rect 22192 11766 22244 11772
rect 22284 11824 22336 11830
rect 22284 11766 22336 11772
rect 21914 11656 21970 11665
rect 21914 11591 21970 11600
rect 21744 11342 21864 11370
rect 21640 11280 21692 11286
rect 21640 11222 21692 11228
rect 21272 11086 21324 11092
rect 21454 11112 21510 11121
rect 21284 10849 21312 11086
rect 21454 11047 21510 11056
rect 21270 10840 21326 10849
rect 21270 10775 21326 10784
rect 21284 9761 21312 10775
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 21270 9752 21326 9761
rect 21376 9722 21404 10610
rect 21270 9687 21326 9696
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 21178 9072 21234 9081
rect 21178 9007 21234 9016
rect 21192 8974 21220 9007
rect 21180 8968 21232 8974
rect 21284 8945 21312 9590
rect 21180 8910 21232 8916
rect 21270 8936 21326 8945
rect 21270 8871 21326 8880
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 21088 8628 21140 8634
rect 21088 8570 21140 8576
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 21100 7886 21128 8434
rect 21192 8412 21220 8774
rect 21284 8566 21312 8871
rect 21272 8560 21324 8566
rect 21272 8502 21324 8508
rect 21192 8384 21312 8412
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 21088 7880 21140 7886
rect 21088 7822 21140 7828
rect 21100 7206 21128 7822
rect 21192 7546 21220 8230
rect 21284 7834 21312 8384
rect 21376 7954 21404 9658
rect 21468 8634 21496 11047
rect 21548 10736 21600 10742
rect 21548 10678 21600 10684
rect 21560 10198 21588 10678
rect 21548 10192 21600 10198
rect 21548 10134 21600 10140
rect 21560 10033 21588 10134
rect 21652 10062 21680 11222
rect 21744 10674 21772 11342
rect 21824 11280 21876 11286
rect 21822 11248 21824 11257
rect 21876 11248 21878 11257
rect 21822 11183 21878 11192
rect 21824 11144 21876 11150
rect 21824 11086 21876 11092
rect 21732 10668 21784 10674
rect 21732 10610 21784 10616
rect 21640 10056 21692 10062
rect 21546 10024 21602 10033
rect 21640 9998 21692 10004
rect 21546 9959 21602 9968
rect 21744 9897 21772 10610
rect 21730 9888 21786 9897
rect 21730 9823 21786 9832
rect 21548 9716 21600 9722
rect 21548 9658 21600 9664
rect 21560 8974 21588 9658
rect 21640 9172 21692 9178
rect 21640 9114 21692 9120
rect 21548 8968 21600 8974
rect 21548 8910 21600 8916
rect 21456 8628 21508 8634
rect 21456 8570 21508 8576
rect 21454 8528 21510 8537
rect 21454 8463 21456 8472
rect 21508 8463 21510 8472
rect 21456 8434 21508 8440
rect 21454 8256 21510 8265
rect 21454 8191 21510 8200
rect 21364 7948 21416 7954
rect 21364 7890 21416 7896
rect 21284 7806 21404 7834
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21284 7410 21312 7686
rect 21272 7404 21324 7410
rect 21272 7346 21324 7352
rect 21088 7200 21140 7206
rect 21088 7142 21140 7148
rect 21100 6866 21128 7142
rect 21088 6860 21140 6866
rect 21088 6802 21140 6808
rect 21376 6780 21404 7806
rect 21468 7410 21496 8191
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21560 6934 21588 8910
rect 21652 8498 21680 9114
rect 21640 8492 21692 8498
rect 21640 8434 21692 8440
rect 21548 6928 21600 6934
rect 21548 6870 21600 6876
rect 21640 6928 21692 6934
rect 21640 6870 21692 6876
rect 21376 6752 21588 6780
rect 21652 6769 21680 6870
rect 21744 6780 21772 9823
rect 21836 9586 21864 11086
rect 21824 9580 21876 9586
rect 21824 9522 21876 9528
rect 21836 9042 21864 9522
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 21928 8974 21956 11591
rect 22100 11552 22152 11558
rect 22100 11494 22152 11500
rect 22112 11121 22140 11494
rect 22204 11150 22232 11766
rect 22192 11144 22244 11150
rect 22098 11112 22154 11121
rect 22192 11086 22244 11092
rect 22098 11047 22154 11056
rect 22098 10976 22154 10985
rect 22098 10911 22154 10920
rect 22112 10266 22140 10911
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 22100 10056 22152 10062
rect 22100 9998 22152 10004
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 22112 8922 22140 9998
rect 22296 9382 22324 11766
rect 22480 10742 22508 11834
rect 22572 11150 22600 12174
rect 22560 11144 22612 11150
rect 22560 11086 22612 11092
rect 22468 10736 22520 10742
rect 22572 10713 22600 11086
rect 22468 10678 22520 10684
rect 22558 10704 22614 10713
rect 22480 10470 22508 10678
rect 22558 10639 22614 10648
rect 22468 10464 22520 10470
rect 22468 10406 22520 10412
rect 22560 10056 22612 10062
rect 22560 9998 22612 10004
rect 22468 9920 22520 9926
rect 22468 9862 22520 9868
rect 22480 9382 22508 9862
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 22468 9376 22520 9382
rect 22468 9318 22520 9324
rect 21824 8900 21876 8906
rect 22112 8894 22416 8922
rect 22572 8906 22600 9998
rect 22664 9722 22692 13262
rect 22756 10810 22784 16390
rect 22834 15600 22890 15609
rect 22834 15535 22890 15544
rect 22848 15434 22876 15535
rect 22836 15428 22888 15434
rect 22836 15370 22888 15376
rect 22848 11082 22876 15370
rect 22940 13530 22968 17546
rect 23032 17270 23060 17614
rect 23020 17264 23072 17270
rect 23020 17206 23072 17212
rect 23308 17218 23336 18142
rect 23492 17678 23520 18158
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 23032 16590 23060 17206
rect 23308 17190 23520 17218
rect 23204 17128 23256 17134
rect 23204 17070 23256 17076
rect 23216 16998 23244 17070
rect 23204 16992 23256 16998
rect 23204 16934 23256 16940
rect 23216 16590 23244 16934
rect 23386 16824 23442 16833
rect 23492 16794 23520 17190
rect 23572 17128 23624 17134
rect 23572 17070 23624 17076
rect 23386 16759 23442 16768
rect 23480 16788 23532 16794
rect 23020 16584 23072 16590
rect 23020 16526 23072 16532
rect 23204 16584 23256 16590
rect 23204 16526 23256 16532
rect 23400 15570 23428 16759
rect 23480 16730 23532 16736
rect 23388 15564 23440 15570
rect 23388 15506 23440 15512
rect 23296 15428 23348 15434
rect 23296 15370 23348 15376
rect 23204 14816 23256 14822
rect 23204 14758 23256 14764
rect 23216 14482 23244 14758
rect 23204 14476 23256 14482
rect 23204 14418 23256 14424
rect 23204 14340 23256 14346
rect 23308 14328 23336 15370
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 23256 14300 23336 14328
rect 23204 14282 23256 14288
rect 22928 13524 22980 13530
rect 22928 13466 22980 13472
rect 23216 12918 23244 14282
rect 23400 14074 23428 14962
rect 23492 14074 23520 16730
rect 23584 15473 23612 17070
rect 23570 15464 23626 15473
rect 23570 15399 23626 15408
rect 23584 14958 23612 15399
rect 23572 14952 23624 14958
rect 23572 14894 23624 14900
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23480 13796 23532 13802
rect 23480 13738 23532 13744
rect 23492 13705 23520 13738
rect 23478 13696 23534 13705
rect 23478 13631 23534 13640
rect 23204 12912 23256 12918
rect 23204 12854 23256 12860
rect 23388 12640 23440 12646
rect 23388 12582 23440 12588
rect 22928 12368 22980 12374
rect 22928 12310 22980 12316
rect 22940 11286 22968 12310
rect 23296 12096 23348 12102
rect 23296 12038 23348 12044
rect 23308 11762 23336 12038
rect 23296 11756 23348 11762
rect 23296 11698 23348 11704
rect 23112 11552 23164 11558
rect 23112 11494 23164 11500
rect 22928 11280 22980 11286
rect 22928 11222 22980 11228
rect 22836 11076 22888 11082
rect 22836 11018 22888 11024
rect 22940 10810 22968 11222
rect 22744 10804 22796 10810
rect 22744 10746 22796 10752
rect 22928 10804 22980 10810
rect 22980 10764 23060 10792
rect 22928 10746 22980 10752
rect 22836 10668 22888 10674
rect 22836 10610 22888 10616
rect 22928 10668 22980 10674
rect 22928 10610 22980 10616
rect 22742 10296 22798 10305
rect 22848 10266 22876 10610
rect 22742 10231 22798 10240
rect 22836 10260 22888 10266
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22650 9616 22706 9625
rect 22650 9551 22706 9560
rect 21824 8842 21876 8848
rect 21836 8090 21864 8842
rect 22284 8832 22336 8838
rect 22284 8774 22336 8780
rect 22296 8566 22324 8774
rect 21916 8560 21968 8566
rect 22284 8560 22336 8566
rect 21968 8520 22048 8548
rect 21916 8502 21968 8508
rect 21916 8424 21968 8430
rect 21916 8366 21968 8372
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21836 7410 21864 8026
rect 21928 7818 21956 8366
rect 21916 7812 21968 7818
rect 22020 7800 22048 8520
rect 22284 8502 22336 8508
rect 22388 8514 22416 8894
rect 22468 8900 22520 8906
rect 22468 8842 22520 8848
rect 22560 8900 22612 8906
rect 22560 8842 22612 8848
rect 22480 8634 22508 8842
rect 22664 8634 22692 9551
rect 22468 8628 22520 8634
rect 22468 8570 22520 8576
rect 22652 8628 22704 8634
rect 22652 8570 22704 8576
rect 22388 8486 22692 8514
rect 22756 8498 22784 10231
rect 22836 10202 22888 10208
rect 22940 10198 22968 10610
rect 22928 10192 22980 10198
rect 22926 10160 22928 10169
rect 22980 10160 22982 10169
rect 22926 10095 22982 10104
rect 22836 9580 22888 9586
rect 22836 9522 22888 9528
rect 22848 9110 22876 9522
rect 22928 9444 22980 9450
rect 22928 9386 22980 9392
rect 22836 9104 22888 9110
rect 22836 9046 22888 9052
rect 22940 8974 22968 9386
rect 22928 8968 22980 8974
rect 22928 8910 22980 8916
rect 23032 8673 23060 10764
rect 23124 10690 23152 11494
rect 23296 11144 23348 11150
rect 23296 11086 23348 11092
rect 23308 10810 23336 11086
rect 23296 10804 23348 10810
rect 23296 10746 23348 10752
rect 23124 10662 23336 10690
rect 23204 10464 23256 10470
rect 23204 10406 23256 10412
rect 23216 9654 23244 10406
rect 23204 9648 23256 9654
rect 23204 9590 23256 9596
rect 23112 9172 23164 9178
rect 23112 9114 23164 9120
rect 23018 8664 23074 8673
rect 23018 8599 23074 8608
rect 23124 8498 23152 9114
rect 22664 8362 22692 8486
rect 22744 8492 22796 8498
rect 22744 8434 22796 8440
rect 22836 8492 22888 8498
rect 22836 8434 22888 8440
rect 23112 8492 23164 8498
rect 23216 8480 23244 9590
rect 23308 8616 23336 10662
rect 23400 10130 23428 12582
rect 23676 12434 23704 19314
rect 23848 18760 23900 18766
rect 23848 18702 23900 18708
rect 23860 18290 23888 18702
rect 23848 18284 23900 18290
rect 23848 18226 23900 18232
rect 23756 18080 23808 18086
rect 23756 18022 23808 18028
rect 23768 16114 23796 18022
rect 23860 17814 23888 18226
rect 23848 17808 23900 17814
rect 23848 17750 23900 17756
rect 23940 17740 23992 17746
rect 23940 17682 23992 17688
rect 23848 17536 23900 17542
rect 23848 17478 23900 17484
rect 23860 16998 23888 17478
rect 23952 17134 23980 17682
rect 24044 17649 24072 19722
rect 24030 17640 24086 17649
rect 24030 17575 24086 17584
rect 24124 17604 24176 17610
rect 23940 17128 23992 17134
rect 23940 17070 23992 17076
rect 23848 16992 23900 16998
rect 23848 16934 23900 16940
rect 23756 16108 23808 16114
rect 23756 16050 23808 16056
rect 24044 15434 24072 17575
rect 24124 17546 24176 17552
rect 24136 17066 24164 17546
rect 24320 17218 24348 26846
rect 24412 26586 24440 27542
rect 24400 26580 24452 26586
rect 24400 26522 24452 26528
rect 24412 24818 24440 26522
rect 24400 24812 24452 24818
rect 24400 24754 24452 24760
rect 24400 24608 24452 24614
rect 24400 24550 24452 24556
rect 24412 23050 24440 24550
rect 24400 23044 24452 23050
rect 24400 22986 24452 22992
rect 24400 20596 24452 20602
rect 24400 20538 24452 20544
rect 24412 20058 24440 20538
rect 24400 20052 24452 20058
rect 24400 19994 24452 20000
rect 24504 18970 24532 31282
rect 24596 29646 24624 31826
rect 24584 29640 24636 29646
rect 24584 29582 24636 29588
rect 24584 27328 24636 27334
rect 24584 27270 24636 27276
rect 24596 26994 24624 27270
rect 24584 26988 24636 26994
rect 24584 26930 24636 26936
rect 24688 25294 24716 33594
rect 24860 32224 24912 32230
rect 24860 32166 24912 32172
rect 24872 32026 24900 32166
rect 24860 32020 24912 32026
rect 24860 31962 24912 31968
rect 24964 31346 24992 36071
rect 25148 35834 25176 36722
rect 25412 36712 25464 36718
rect 25412 36654 25464 36660
rect 25320 36576 25372 36582
rect 25320 36518 25372 36524
rect 25332 36378 25360 36518
rect 25320 36372 25372 36378
rect 25320 36314 25372 36320
rect 25424 36242 25452 36654
rect 25412 36236 25464 36242
rect 25412 36178 25464 36184
rect 25228 36032 25280 36038
rect 25228 35974 25280 35980
rect 25136 35828 25188 35834
rect 25136 35770 25188 35776
rect 25136 35692 25188 35698
rect 25136 35634 25188 35640
rect 25148 35086 25176 35634
rect 25136 35080 25188 35086
rect 25136 35022 25188 35028
rect 25148 34746 25176 35022
rect 25136 34740 25188 34746
rect 25136 34682 25188 34688
rect 25148 33998 25176 34682
rect 25136 33992 25188 33998
rect 25136 33934 25188 33940
rect 25240 33946 25268 35974
rect 25424 35154 25452 36178
rect 25608 36009 25636 37810
rect 25700 37466 25728 37810
rect 25780 37800 25832 37806
rect 25780 37742 25832 37748
rect 25688 37460 25740 37466
rect 25688 37402 25740 37408
rect 25688 36168 25740 36174
rect 25688 36110 25740 36116
rect 25594 36000 25650 36009
rect 25594 35935 25650 35944
rect 25608 35578 25636 35935
rect 25700 35766 25728 36110
rect 25688 35760 25740 35766
rect 25688 35702 25740 35708
rect 25608 35550 25728 35578
rect 25504 35488 25556 35494
rect 25504 35430 25556 35436
rect 25516 35290 25544 35430
rect 25504 35284 25556 35290
rect 25504 35226 25556 35232
rect 25412 35148 25464 35154
rect 25412 35090 25464 35096
rect 25596 34944 25648 34950
rect 25596 34886 25648 34892
rect 25608 34649 25636 34886
rect 25594 34640 25650 34649
rect 25594 34575 25650 34584
rect 25700 34490 25728 35550
rect 25608 34462 25728 34490
rect 25240 33918 25544 33946
rect 25044 33856 25096 33862
rect 25044 33798 25096 33804
rect 25056 31498 25084 33798
rect 25136 32428 25188 32434
rect 25136 32370 25188 32376
rect 25148 31754 25176 32370
rect 25148 31726 25268 31754
rect 25056 31470 25176 31498
rect 25044 31408 25096 31414
rect 25044 31350 25096 31356
rect 24952 31340 25004 31346
rect 24952 31282 25004 31288
rect 24860 30252 24912 30258
rect 24860 30194 24912 30200
rect 24768 29504 24820 29510
rect 24768 29446 24820 29452
rect 24780 28558 24808 29446
rect 24872 28762 24900 30194
rect 24860 28756 24912 28762
rect 24860 28698 24912 28704
rect 24768 28552 24820 28558
rect 24768 28494 24820 28500
rect 24872 28082 24900 28698
rect 24964 28694 24992 31282
rect 24952 28688 25004 28694
rect 24952 28630 25004 28636
rect 24860 28076 24912 28082
rect 24860 28018 24912 28024
rect 24952 28076 25004 28082
rect 24952 28018 25004 28024
rect 24872 27112 24900 28018
rect 24780 27084 24900 27112
rect 24780 26994 24808 27084
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24768 26512 24820 26518
rect 24768 26454 24820 26460
rect 24676 25288 24728 25294
rect 24676 25230 24728 25236
rect 24676 24744 24728 24750
rect 24676 24686 24728 24692
rect 24584 23316 24636 23322
rect 24584 23258 24636 23264
rect 24596 22778 24624 23258
rect 24584 22772 24636 22778
rect 24584 22714 24636 22720
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 24596 21690 24624 21966
rect 24584 21684 24636 21690
rect 24584 21626 24636 21632
rect 24688 20618 24716 24686
rect 24780 22681 24808 26454
rect 24860 25832 24912 25838
rect 24860 25774 24912 25780
rect 24872 24818 24900 25774
rect 24860 24812 24912 24818
rect 24860 24754 24912 24760
rect 24872 24070 24900 24754
rect 24860 24064 24912 24070
rect 24860 24006 24912 24012
rect 24860 23248 24912 23254
rect 24964 23236 24992 28018
rect 25056 26382 25084 31350
rect 25148 31346 25176 31470
rect 25136 31340 25188 31346
rect 25136 31282 25188 31288
rect 25240 30870 25268 31726
rect 25228 30864 25280 30870
rect 25228 30806 25280 30812
rect 25412 28960 25464 28966
rect 25412 28902 25464 28908
rect 25424 27946 25452 28902
rect 25412 27940 25464 27946
rect 25412 27882 25464 27888
rect 25136 27872 25188 27878
rect 25136 27814 25188 27820
rect 25148 27470 25176 27814
rect 25424 27674 25452 27882
rect 25412 27668 25464 27674
rect 25412 27610 25464 27616
rect 25136 27464 25188 27470
rect 25136 27406 25188 27412
rect 25228 27396 25280 27402
rect 25228 27338 25280 27344
rect 25240 27130 25268 27338
rect 25136 27124 25188 27130
rect 25136 27066 25188 27072
rect 25228 27124 25280 27130
rect 25228 27066 25280 27072
rect 25148 26994 25176 27066
rect 25136 26988 25188 26994
rect 25136 26930 25188 26936
rect 25228 26988 25280 26994
rect 25280 26948 25360 26976
rect 25228 26930 25280 26936
rect 25136 26852 25188 26858
rect 25136 26794 25188 26800
rect 25044 26376 25096 26382
rect 25044 26318 25096 26324
rect 25044 25288 25096 25294
rect 25044 25230 25096 25236
rect 25056 24206 25084 25230
rect 25148 24614 25176 26794
rect 25228 26784 25280 26790
rect 25228 26726 25280 26732
rect 25136 24608 25188 24614
rect 25136 24550 25188 24556
rect 25044 24200 25096 24206
rect 25044 24142 25096 24148
rect 25240 23882 25268 26726
rect 25332 26382 25360 26948
rect 25516 26586 25544 33918
rect 25608 31414 25636 34462
rect 25792 33980 25820 37742
rect 25964 36576 26016 36582
rect 25964 36518 26016 36524
rect 25976 36378 26004 36518
rect 25964 36372 26016 36378
rect 25964 36314 26016 36320
rect 26068 36174 26096 38150
rect 27264 38010 27292 38898
rect 27252 38004 27304 38010
rect 27252 37946 27304 37952
rect 26148 37868 26200 37874
rect 26148 37810 26200 37816
rect 27252 37868 27304 37874
rect 27252 37810 27304 37816
rect 26160 37466 26188 37810
rect 26148 37460 26200 37466
rect 26148 37402 26200 37408
rect 26056 36168 26108 36174
rect 26056 36110 26108 36116
rect 25872 36032 25924 36038
rect 25872 35974 25924 35980
rect 25884 35766 25912 35974
rect 25872 35760 25924 35766
rect 25872 35702 25924 35708
rect 26068 35494 26096 36110
rect 26056 35488 26108 35494
rect 26056 35430 26108 35436
rect 26608 34740 26660 34746
rect 26608 34682 26660 34688
rect 26424 34060 26476 34066
rect 26424 34002 26476 34008
rect 25792 33952 26096 33980
rect 25872 33516 25924 33522
rect 25872 33458 25924 33464
rect 25688 33312 25740 33318
rect 25688 33254 25740 33260
rect 25700 32910 25728 33254
rect 25688 32904 25740 32910
rect 25688 32846 25740 32852
rect 25688 31680 25740 31686
rect 25688 31622 25740 31628
rect 25780 31680 25832 31686
rect 25780 31622 25832 31628
rect 25596 31408 25648 31414
rect 25596 31350 25648 31356
rect 25700 30870 25728 31622
rect 25688 30864 25740 30870
rect 25688 30806 25740 30812
rect 25792 30666 25820 31622
rect 25780 30660 25832 30666
rect 25780 30602 25832 30608
rect 25596 28076 25648 28082
rect 25596 28018 25648 28024
rect 25608 27130 25636 28018
rect 25792 27946 25820 30602
rect 25884 28082 25912 33458
rect 26068 32298 26096 33952
rect 26332 33856 26384 33862
rect 26332 33798 26384 33804
rect 26344 33522 26372 33798
rect 26436 33658 26464 34002
rect 26620 33998 26648 34682
rect 26792 34196 26844 34202
rect 26792 34138 26844 34144
rect 26608 33992 26660 33998
rect 26608 33934 26660 33940
rect 26424 33652 26476 33658
rect 26424 33594 26476 33600
rect 26332 33516 26384 33522
rect 26332 33458 26384 33464
rect 26516 33516 26568 33522
rect 26516 33458 26568 33464
rect 26528 33114 26556 33458
rect 26608 33448 26660 33454
rect 26608 33390 26660 33396
rect 26620 33114 26648 33390
rect 26516 33108 26568 33114
rect 26516 33050 26568 33056
rect 26608 33108 26660 33114
rect 26608 33050 26660 33056
rect 26804 33046 26832 34138
rect 27264 33862 27292 37810
rect 33612 36922 33640 38898
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 35594 38108 35902 38117
rect 35594 38106 35600 38108
rect 35656 38106 35680 38108
rect 35736 38106 35760 38108
rect 35816 38106 35840 38108
rect 35896 38106 35902 38108
rect 35656 38054 35658 38106
rect 35838 38054 35840 38106
rect 35594 38052 35600 38054
rect 35656 38052 35680 38054
rect 35736 38052 35760 38054
rect 35816 38052 35840 38054
rect 35896 38052 35902 38054
rect 35594 38043 35902 38052
rect 37648 37868 37700 37874
rect 37648 37810 37700 37816
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 37660 36922 37688 37810
rect 37832 37664 37884 37670
rect 37832 37606 37884 37612
rect 37844 37505 37872 37606
rect 37830 37496 37886 37505
rect 37830 37431 37886 37440
rect 33600 36916 33652 36922
rect 33600 36858 33652 36864
rect 37648 36916 37700 36922
rect 37648 36858 37700 36864
rect 28448 36780 28500 36786
rect 28448 36722 28500 36728
rect 37372 36780 37424 36786
rect 37372 36722 37424 36728
rect 28460 36378 28488 36722
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 37384 36378 37412 36722
rect 28448 36372 28500 36378
rect 28448 36314 28500 36320
rect 37372 36372 37424 36378
rect 37372 36314 37424 36320
rect 27804 36168 27856 36174
rect 27804 36110 27856 36116
rect 28632 36168 28684 36174
rect 28632 36110 28684 36116
rect 27528 34740 27580 34746
rect 27528 34682 27580 34688
rect 27540 34202 27568 34682
rect 27528 34196 27580 34202
rect 27528 34138 27580 34144
rect 27344 34128 27396 34134
rect 27396 34088 27476 34116
rect 27344 34070 27396 34076
rect 27448 34082 27476 34088
rect 27448 34054 27568 34082
rect 27540 33998 27568 34054
rect 27528 33992 27580 33998
rect 27528 33934 27580 33940
rect 27068 33856 27120 33862
rect 27068 33798 27120 33804
rect 27252 33856 27304 33862
rect 27252 33798 27304 33804
rect 27080 33658 27108 33798
rect 27068 33652 27120 33658
rect 27068 33594 27120 33600
rect 27264 33386 27292 33798
rect 27528 33516 27580 33522
rect 27528 33458 27580 33464
rect 27252 33380 27304 33386
rect 27252 33322 27304 33328
rect 27436 33380 27488 33386
rect 27436 33322 27488 33328
rect 26792 33040 26844 33046
rect 26792 32982 26844 32988
rect 27160 32904 27212 32910
rect 27160 32846 27212 32852
rect 26516 32836 26568 32842
rect 26516 32778 26568 32784
rect 26056 32292 26108 32298
rect 26056 32234 26108 32240
rect 26068 31754 26096 32234
rect 25976 31726 26096 31754
rect 25872 28076 25924 28082
rect 25872 28018 25924 28024
rect 25780 27940 25832 27946
rect 25780 27882 25832 27888
rect 25596 27124 25648 27130
rect 25596 27066 25648 27072
rect 25504 26580 25556 26586
rect 25504 26522 25556 26528
rect 25412 26444 25464 26450
rect 25412 26386 25464 26392
rect 25320 26376 25372 26382
rect 25320 26318 25372 26324
rect 25320 25152 25372 25158
rect 25320 25094 25372 25100
rect 25332 24206 25360 25094
rect 25320 24200 25372 24206
rect 25320 24142 25372 24148
rect 24912 23208 24992 23236
rect 25056 23854 25268 23882
rect 24860 23190 24912 23196
rect 24872 22982 24900 23190
rect 24860 22976 24912 22982
rect 24860 22918 24912 22924
rect 24766 22672 24822 22681
rect 24766 22607 24822 22616
rect 24860 22636 24912 22642
rect 24780 22574 24808 22607
rect 24860 22578 24912 22584
rect 24768 22568 24820 22574
rect 24768 22510 24820 22516
rect 24872 21554 24900 22578
rect 25056 22234 25084 23854
rect 25332 23769 25360 24142
rect 25318 23760 25374 23769
rect 25318 23695 25374 23704
rect 25424 23662 25452 26386
rect 25688 26308 25740 26314
rect 25688 26250 25740 26256
rect 25596 24200 25648 24206
rect 25516 24160 25596 24188
rect 25412 23656 25464 23662
rect 25332 23616 25412 23644
rect 25332 23474 25360 23616
rect 25412 23598 25464 23604
rect 25148 23446 25360 23474
rect 25044 22228 25096 22234
rect 25044 22170 25096 22176
rect 25148 22094 25176 23446
rect 25412 23112 25464 23118
rect 25412 23054 25464 23060
rect 25424 22574 25452 23054
rect 25412 22568 25464 22574
rect 25412 22510 25464 22516
rect 25516 22094 25544 24160
rect 25596 24142 25648 24148
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25608 23361 25636 23666
rect 25594 23352 25650 23361
rect 25594 23287 25650 23296
rect 25596 22976 25648 22982
rect 25596 22918 25648 22924
rect 25608 22710 25636 22918
rect 25596 22704 25648 22710
rect 25596 22646 25648 22652
rect 25056 22066 25176 22094
rect 25240 22066 25544 22094
rect 24860 21548 24912 21554
rect 24860 21490 24912 21496
rect 25056 21434 25084 22066
rect 25136 21616 25188 21622
rect 25136 21558 25188 21564
rect 24872 21406 25084 21434
rect 24768 20868 24820 20874
rect 24768 20810 24820 20816
rect 24596 20590 24716 20618
rect 24780 20602 24808 20810
rect 24768 20596 24820 20602
rect 24596 20346 24624 20590
rect 24768 20538 24820 20544
rect 24766 20496 24822 20505
rect 24688 20466 24766 20482
rect 24676 20460 24766 20466
rect 24728 20454 24766 20460
rect 24872 20466 24900 21406
rect 25148 21010 25176 21558
rect 25240 21010 25268 22066
rect 25608 21622 25636 22646
rect 25596 21616 25648 21622
rect 25410 21584 25466 21593
rect 25596 21558 25648 21564
rect 25410 21519 25466 21528
rect 25424 21146 25452 21519
rect 25596 21344 25648 21350
rect 25596 21286 25648 21292
rect 25412 21140 25464 21146
rect 25412 21082 25464 21088
rect 25608 21078 25636 21286
rect 25596 21072 25648 21078
rect 25596 21014 25648 21020
rect 25136 21004 25188 21010
rect 25136 20946 25188 20952
rect 25228 21004 25280 21010
rect 25228 20946 25280 20952
rect 25504 20800 25556 20806
rect 25504 20742 25556 20748
rect 24766 20431 24822 20440
rect 24860 20460 24912 20466
rect 24676 20402 24728 20408
rect 24860 20402 24912 20408
rect 24596 20318 24716 20346
rect 24584 19916 24636 19922
rect 24584 19858 24636 19864
rect 24596 19310 24624 19858
rect 24584 19304 24636 19310
rect 24584 19246 24636 19252
rect 24596 19174 24624 19246
rect 24584 19168 24636 19174
rect 24584 19110 24636 19116
rect 24688 18970 24716 20318
rect 24872 19854 24900 20402
rect 24860 19848 24912 19854
rect 24860 19790 24912 19796
rect 25228 19848 25280 19854
rect 25228 19790 25280 19796
rect 24952 19780 25004 19786
rect 24952 19722 25004 19728
rect 25044 19780 25096 19786
rect 25044 19722 25096 19728
rect 24492 18964 24544 18970
rect 24492 18906 24544 18912
rect 24676 18964 24728 18970
rect 24676 18906 24728 18912
rect 24676 18760 24728 18766
rect 24676 18702 24728 18708
rect 24688 18426 24716 18702
rect 24676 18420 24728 18426
rect 24676 18362 24728 18368
rect 24676 18148 24728 18154
rect 24676 18090 24728 18096
rect 24584 17536 24636 17542
rect 24584 17478 24636 17484
rect 24596 17338 24624 17478
rect 24688 17338 24716 18090
rect 24860 17876 24912 17882
rect 24860 17818 24912 17824
rect 24584 17332 24636 17338
rect 24584 17274 24636 17280
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 24228 17190 24348 17218
rect 24400 17196 24452 17202
rect 24124 17060 24176 17066
rect 24124 17002 24176 17008
rect 24136 16658 24164 17002
rect 24124 16652 24176 16658
rect 24124 16594 24176 16600
rect 24124 16516 24176 16522
rect 24124 16458 24176 16464
rect 24136 16250 24164 16458
rect 24124 16244 24176 16250
rect 24124 16186 24176 16192
rect 24136 15978 24164 16186
rect 24124 15972 24176 15978
rect 24124 15914 24176 15920
rect 24032 15428 24084 15434
rect 24032 15370 24084 15376
rect 23848 15360 23900 15366
rect 23848 15302 23900 15308
rect 23584 12406 23704 12434
rect 23480 11824 23532 11830
rect 23480 11766 23532 11772
rect 23492 11694 23520 11766
rect 23480 11688 23532 11694
rect 23480 11630 23532 11636
rect 23492 11529 23520 11630
rect 23478 11520 23534 11529
rect 23478 11455 23534 11464
rect 23480 11076 23532 11082
rect 23480 11018 23532 11024
rect 23492 10849 23520 11018
rect 23478 10840 23534 10849
rect 23478 10775 23534 10784
rect 23480 10600 23532 10606
rect 23480 10542 23532 10548
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 23492 10062 23520 10542
rect 23480 10056 23532 10062
rect 23480 9998 23532 10004
rect 23492 9466 23520 9998
rect 23584 9586 23612 12406
rect 23664 11280 23716 11286
rect 23664 11222 23716 11228
rect 23676 10577 23704 11222
rect 23756 11144 23808 11150
rect 23756 11086 23808 11092
rect 23662 10568 23718 10577
rect 23662 10503 23718 10512
rect 23664 9988 23716 9994
rect 23664 9930 23716 9936
rect 23676 9586 23704 9930
rect 23768 9586 23796 11086
rect 23860 10305 23888 15302
rect 23938 14648 23994 14657
rect 23938 14583 23994 14592
rect 23952 14550 23980 14583
rect 23940 14544 23992 14550
rect 23940 14486 23992 14492
rect 23952 12374 23980 14486
rect 24124 14000 24176 14006
rect 24124 13942 24176 13948
rect 23940 12368 23992 12374
rect 24136 12322 24164 13942
rect 23940 12310 23992 12316
rect 24044 12294 24164 12322
rect 23940 12164 23992 12170
rect 23940 12106 23992 12112
rect 23952 11558 23980 12106
rect 23940 11552 23992 11558
rect 23940 11494 23992 11500
rect 24044 11506 24072 12294
rect 24124 12232 24176 12238
rect 24124 12174 24176 12180
rect 24136 11830 24164 12174
rect 24124 11824 24176 11830
rect 24122 11792 24124 11801
rect 24176 11792 24178 11801
rect 24122 11727 24178 11736
rect 23952 11150 23980 11494
rect 24044 11478 24164 11506
rect 23940 11144 23992 11150
rect 23940 11086 23992 11092
rect 24032 11076 24084 11082
rect 24032 11018 24084 11024
rect 24044 10538 24072 11018
rect 24136 10606 24164 11478
rect 24228 11286 24256 17190
rect 24400 17138 24452 17144
rect 24412 16250 24440 17138
rect 24768 16992 24820 16998
rect 24768 16934 24820 16940
rect 24780 16794 24808 16934
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 24490 16552 24546 16561
rect 24490 16487 24546 16496
rect 24400 16244 24452 16250
rect 24400 16186 24452 16192
rect 24306 16144 24362 16153
rect 24306 16079 24362 16088
rect 24320 15978 24348 16079
rect 24308 15972 24360 15978
rect 24308 15914 24360 15920
rect 24412 15178 24440 16186
rect 24504 16114 24532 16487
rect 24676 16176 24728 16182
rect 24676 16118 24728 16124
rect 24492 16108 24544 16114
rect 24492 16050 24544 16056
rect 24320 15162 24440 15178
rect 24320 15156 24452 15162
rect 24320 15150 24400 15156
rect 24320 14618 24348 15150
rect 24400 15098 24452 15104
rect 24400 15020 24452 15026
rect 24400 14962 24452 14968
rect 24584 15020 24636 15026
rect 24584 14962 24636 14968
rect 24308 14612 24360 14618
rect 24308 14554 24360 14560
rect 24320 14074 24348 14554
rect 24308 14068 24360 14074
rect 24308 14010 24360 14016
rect 24306 13832 24362 13841
rect 24306 13767 24308 13776
rect 24360 13767 24362 13776
rect 24308 13738 24360 13744
rect 24320 12986 24348 13738
rect 24308 12980 24360 12986
rect 24308 12922 24360 12928
rect 24308 12776 24360 12782
rect 24306 12744 24308 12753
rect 24360 12744 24362 12753
rect 24306 12679 24362 12688
rect 24308 12300 24360 12306
rect 24308 12242 24360 12248
rect 24320 11558 24348 12242
rect 24412 11665 24440 14962
rect 24492 13388 24544 13394
rect 24492 13330 24544 13336
rect 24504 12238 24532 13330
rect 24492 12232 24544 12238
rect 24492 12174 24544 12180
rect 24596 12170 24624 14962
rect 24688 14482 24716 16118
rect 24768 15360 24820 15366
rect 24768 15302 24820 15308
rect 24780 15162 24808 15302
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24780 14498 24808 15098
rect 24872 14600 24900 17818
rect 24964 17610 24992 19722
rect 25056 19514 25084 19722
rect 25136 19712 25188 19718
rect 25136 19654 25188 19660
rect 25044 19508 25096 19514
rect 25044 19450 25096 19456
rect 25148 19378 25176 19654
rect 25240 19514 25268 19790
rect 25228 19508 25280 19514
rect 25228 19450 25280 19456
rect 25136 19372 25188 19378
rect 25136 19314 25188 19320
rect 25320 19168 25372 19174
rect 25320 19110 25372 19116
rect 25136 18828 25188 18834
rect 25136 18770 25188 18776
rect 25044 18760 25096 18766
rect 25044 18702 25096 18708
rect 24952 17604 25004 17610
rect 24952 17546 25004 17552
rect 24964 16794 24992 17546
rect 24952 16788 25004 16794
rect 24952 16730 25004 16736
rect 25056 16250 25084 18702
rect 25148 18290 25176 18770
rect 25332 18766 25360 19110
rect 25320 18760 25372 18766
rect 25320 18702 25372 18708
rect 25136 18284 25188 18290
rect 25136 18226 25188 18232
rect 25228 18284 25280 18290
rect 25228 18226 25280 18232
rect 25240 17882 25268 18226
rect 25228 17876 25280 17882
rect 25228 17818 25280 17824
rect 25516 17814 25544 20742
rect 25700 19174 25728 26250
rect 25792 24070 25820 27882
rect 25884 27062 25912 28018
rect 25976 27606 26004 31726
rect 26332 31680 26384 31686
rect 26332 31622 26384 31628
rect 26344 31482 26372 31622
rect 26332 31476 26384 31482
rect 26332 31418 26384 31424
rect 26424 30252 26476 30258
rect 26424 30194 26476 30200
rect 26056 29776 26108 29782
rect 26056 29718 26108 29724
rect 26068 29306 26096 29718
rect 26436 29646 26464 30194
rect 26424 29640 26476 29646
rect 26330 29608 26386 29617
rect 26160 29566 26330 29594
rect 26056 29300 26108 29306
rect 26056 29242 26108 29248
rect 26160 29170 26188 29566
rect 26424 29582 26476 29588
rect 26330 29543 26386 29552
rect 26240 29504 26292 29510
rect 26240 29446 26292 29452
rect 26148 29164 26200 29170
rect 26148 29106 26200 29112
rect 26160 28762 26188 29106
rect 26252 29102 26280 29446
rect 26424 29232 26476 29238
rect 26528 29220 26556 32778
rect 27172 32026 27200 32846
rect 27160 32020 27212 32026
rect 27160 31962 27212 31968
rect 27172 31346 27200 31962
rect 27160 31340 27212 31346
rect 27160 31282 27212 31288
rect 26976 31272 27028 31278
rect 26976 31214 27028 31220
rect 27252 31272 27304 31278
rect 27252 31214 27304 31220
rect 26988 30938 27016 31214
rect 26976 30932 27028 30938
rect 26976 30874 27028 30880
rect 26700 30660 26752 30666
rect 26700 30602 26752 30608
rect 26608 29844 26660 29850
rect 26608 29786 26660 29792
rect 26620 29646 26648 29786
rect 26608 29640 26660 29646
rect 26608 29582 26660 29588
rect 26712 29458 26740 30602
rect 27160 29844 27212 29850
rect 27160 29786 27212 29792
rect 26976 29640 27028 29646
rect 26976 29582 27028 29588
rect 26988 29458 27016 29582
rect 26476 29192 26556 29220
rect 26620 29430 27016 29458
rect 26424 29174 26476 29180
rect 26240 29096 26292 29102
rect 26240 29038 26292 29044
rect 26148 28756 26200 28762
rect 26148 28698 26200 28704
rect 26056 28416 26108 28422
rect 26056 28358 26108 28364
rect 25964 27600 26016 27606
rect 25964 27542 26016 27548
rect 25872 27056 25924 27062
rect 25872 26998 25924 27004
rect 25964 26988 26016 26994
rect 25964 26930 26016 26936
rect 25872 26784 25924 26790
rect 25976 26772 26004 26930
rect 25924 26744 26004 26772
rect 25872 26726 25924 26732
rect 25884 24818 25912 26726
rect 25962 24848 26018 24857
rect 25872 24812 25924 24818
rect 25962 24783 26018 24792
rect 25872 24754 25924 24760
rect 25884 24410 25912 24754
rect 25872 24404 25924 24410
rect 25872 24346 25924 24352
rect 25780 24064 25832 24070
rect 25780 24006 25832 24012
rect 25976 23662 26004 24783
rect 25964 23656 26016 23662
rect 25964 23598 26016 23604
rect 25780 23112 25832 23118
rect 25780 23054 25832 23060
rect 25792 22642 25820 23054
rect 26068 22778 26096 28358
rect 26148 26784 26200 26790
rect 26148 26726 26200 26732
rect 26160 26382 26188 26726
rect 26332 26512 26384 26518
rect 26332 26454 26384 26460
rect 26148 26376 26200 26382
rect 26148 26318 26200 26324
rect 26160 25906 26188 26318
rect 26344 26042 26372 26454
rect 26332 26036 26384 26042
rect 26332 25978 26384 25984
rect 26148 25900 26200 25906
rect 26148 25842 26200 25848
rect 26344 25498 26372 25978
rect 26332 25492 26384 25498
rect 26332 25434 26384 25440
rect 26436 24886 26464 29174
rect 26620 28082 26648 29430
rect 26792 29300 26844 29306
rect 26792 29242 26844 29248
rect 26804 28558 26832 29242
rect 26884 29164 26936 29170
rect 26884 29106 26936 29112
rect 26700 28552 26752 28558
rect 26700 28494 26752 28500
rect 26792 28552 26844 28558
rect 26792 28494 26844 28500
rect 26608 28076 26660 28082
rect 26608 28018 26660 28024
rect 26608 26988 26660 26994
rect 26608 26930 26660 26936
rect 26424 24880 26476 24886
rect 26424 24822 26476 24828
rect 26436 24750 26464 24822
rect 26240 24744 26292 24750
rect 26240 24686 26292 24692
rect 26424 24744 26476 24750
rect 26424 24686 26476 24692
rect 26148 24200 26200 24206
rect 26148 24142 26200 24148
rect 26160 23594 26188 24142
rect 26148 23588 26200 23594
rect 26148 23530 26200 23536
rect 26252 23526 26280 24686
rect 26620 24410 26648 26930
rect 26712 26353 26740 28494
rect 26792 28076 26844 28082
rect 26792 28018 26844 28024
rect 26804 27878 26832 28018
rect 26792 27872 26844 27878
rect 26792 27814 26844 27820
rect 26804 26994 26832 27814
rect 26792 26988 26844 26994
rect 26792 26930 26844 26936
rect 26896 26518 26924 29106
rect 26976 28552 27028 28558
rect 26976 28494 27028 28500
rect 26884 26512 26936 26518
rect 26884 26454 26936 26460
rect 26896 26382 26924 26454
rect 26884 26376 26936 26382
rect 26698 26344 26754 26353
rect 26884 26318 26936 26324
rect 26698 26279 26754 26288
rect 26712 25378 26740 26279
rect 26712 25350 26832 25378
rect 26700 25288 26752 25294
rect 26700 25230 26752 25236
rect 26608 24404 26660 24410
rect 26608 24346 26660 24352
rect 26240 23520 26292 23526
rect 26240 23462 26292 23468
rect 26516 23112 26568 23118
rect 26516 23054 26568 23060
rect 26240 23044 26292 23050
rect 26240 22986 26292 22992
rect 26056 22772 26108 22778
rect 26056 22714 26108 22720
rect 26252 22658 26280 22986
rect 26332 22976 26384 22982
rect 26332 22918 26384 22924
rect 26344 22817 26372 22918
rect 26330 22808 26386 22817
rect 26528 22778 26556 23054
rect 26330 22743 26332 22752
rect 26384 22743 26386 22752
rect 26516 22772 26568 22778
rect 26332 22714 26384 22720
rect 26516 22714 26568 22720
rect 25780 22636 25832 22642
rect 26252 22630 26372 22658
rect 25780 22578 25832 22584
rect 25792 22438 25820 22578
rect 25780 22432 25832 22438
rect 25780 22374 25832 22380
rect 25792 22030 25820 22374
rect 25780 22024 25832 22030
rect 25780 21966 25832 21972
rect 26240 22024 26292 22030
rect 26240 21966 26292 21972
rect 25780 21888 25832 21894
rect 25780 21830 25832 21836
rect 25792 21690 25820 21830
rect 25780 21684 25832 21690
rect 25780 21626 25832 21632
rect 25792 21570 25820 21626
rect 25792 21554 25912 21570
rect 25792 21548 25924 21554
rect 25792 21542 25872 21548
rect 25872 21490 25924 21496
rect 26252 21486 26280 21966
rect 26344 21486 26372 22630
rect 26712 22094 26740 25230
rect 26804 22166 26832 25350
rect 26988 24818 27016 28494
rect 27172 28082 27200 29786
rect 27264 28150 27292 31214
rect 27344 29504 27396 29510
rect 27344 29446 27396 29452
rect 27356 28218 27384 29446
rect 27448 28762 27476 33322
rect 27540 31362 27568 33458
rect 27620 32972 27672 32978
rect 27620 32914 27672 32920
rect 27632 31482 27660 32914
rect 27816 32230 27844 36110
rect 27896 33856 27948 33862
rect 27896 33798 27948 33804
rect 27908 33454 27936 33798
rect 28172 33516 28224 33522
rect 28172 33458 28224 33464
rect 27896 33448 27948 33454
rect 27896 33390 27948 33396
rect 28080 33380 28132 33386
rect 28080 33322 28132 33328
rect 27804 32224 27856 32230
rect 27804 32166 27856 32172
rect 27804 31952 27856 31958
rect 27804 31894 27856 31900
rect 27620 31476 27672 31482
rect 27620 31418 27672 31424
rect 27540 31334 27660 31362
rect 27528 29300 27580 29306
rect 27528 29242 27580 29248
rect 27540 29170 27568 29242
rect 27632 29170 27660 31334
rect 27712 30728 27764 30734
rect 27712 30670 27764 30676
rect 27724 30326 27752 30670
rect 27712 30320 27764 30326
rect 27712 30262 27764 30268
rect 27528 29164 27580 29170
rect 27528 29106 27580 29112
rect 27620 29164 27672 29170
rect 27620 29106 27672 29112
rect 27528 29028 27580 29034
rect 27528 28970 27580 28976
rect 27436 28756 27488 28762
rect 27436 28698 27488 28704
rect 27344 28212 27396 28218
rect 27344 28154 27396 28160
rect 27252 28144 27304 28150
rect 27252 28086 27304 28092
rect 27160 28076 27212 28082
rect 27080 28036 27160 28064
rect 27080 27130 27108 28036
rect 27160 28018 27212 28024
rect 27160 27464 27212 27470
rect 27160 27406 27212 27412
rect 27068 27124 27120 27130
rect 27068 27066 27120 27072
rect 27172 27010 27200 27406
rect 27264 27130 27292 28086
rect 27540 27606 27568 28970
rect 27816 28558 27844 31894
rect 28092 31822 28120 33322
rect 28184 33046 28212 33458
rect 28172 33040 28224 33046
rect 28172 32982 28224 32988
rect 28644 32745 28672 36110
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 37648 35692 37700 35698
rect 37648 35634 37700 35640
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 37660 35290 37688 35634
rect 37832 35488 37884 35494
rect 37830 35456 37832 35465
rect 37884 35456 37886 35465
rect 37830 35391 37886 35400
rect 37648 35284 37700 35290
rect 37648 35226 37700 35232
rect 37372 35080 37424 35086
rect 37372 35022 37424 35028
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 29380 34610 29868 34626
rect 29368 34604 29880 34610
rect 29420 34598 29828 34604
rect 29368 34546 29420 34552
rect 29828 34546 29880 34552
rect 28908 34536 28960 34542
rect 28908 34478 28960 34484
rect 28816 32768 28868 32774
rect 28630 32736 28686 32745
rect 28816 32710 28868 32716
rect 28630 32671 28686 32680
rect 27896 31816 27948 31822
rect 27896 31758 27948 31764
rect 28080 31816 28132 31822
rect 28080 31758 28132 31764
rect 27908 29306 27936 31758
rect 28356 31340 28408 31346
rect 28356 31282 28408 31288
rect 28540 31340 28592 31346
rect 28540 31282 28592 31288
rect 28172 30796 28224 30802
rect 28172 30738 28224 30744
rect 28080 30388 28132 30394
rect 28080 30330 28132 30336
rect 28092 29646 28120 30330
rect 28184 30326 28212 30738
rect 28264 30728 28316 30734
rect 28264 30670 28316 30676
rect 28172 30320 28224 30326
rect 28172 30262 28224 30268
rect 28276 30258 28304 30670
rect 28264 30252 28316 30258
rect 28264 30194 28316 30200
rect 28172 30048 28224 30054
rect 28172 29990 28224 29996
rect 28080 29640 28132 29646
rect 28080 29582 28132 29588
rect 28080 29504 28132 29510
rect 28080 29446 28132 29452
rect 28092 29345 28120 29446
rect 28078 29336 28134 29345
rect 27896 29300 27948 29306
rect 28078 29271 28134 29280
rect 27896 29242 27948 29248
rect 28078 29064 28134 29073
rect 28078 28999 28134 29008
rect 28092 28966 28120 28999
rect 28080 28960 28132 28966
rect 28080 28902 28132 28908
rect 28184 28762 28212 29990
rect 28276 29306 28304 30194
rect 28264 29300 28316 29306
rect 28264 29242 28316 29248
rect 28276 29034 28304 29242
rect 28264 29028 28316 29034
rect 28264 28970 28316 28976
rect 28172 28756 28224 28762
rect 28172 28698 28224 28704
rect 27804 28552 27856 28558
rect 27804 28494 27856 28500
rect 27528 27600 27580 27606
rect 27528 27542 27580 27548
rect 27804 27600 27856 27606
rect 27804 27542 27856 27548
rect 27436 27464 27488 27470
rect 27436 27406 27488 27412
rect 27448 27130 27476 27406
rect 27252 27124 27304 27130
rect 27252 27066 27304 27072
rect 27436 27124 27488 27130
rect 27436 27066 27488 27072
rect 27080 26982 27200 27010
rect 27252 26988 27304 26994
rect 27080 25702 27108 26982
rect 27252 26930 27304 26936
rect 27712 26988 27764 26994
rect 27712 26930 27764 26936
rect 27160 26852 27212 26858
rect 27160 26794 27212 26800
rect 27172 26382 27200 26794
rect 27160 26376 27212 26382
rect 27160 26318 27212 26324
rect 27264 26246 27292 26930
rect 27436 26784 27488 26790
rect 27436 26726 27488 26732
rect 27448 26382 27476 26726
rect 27724 26586 27752 26930
rect 27712 26580 27764 26586
rect 27712 26522 27764 26528
rect 27344 26376 27396 26382
rect 27344 26318 27396 26324
rect 27436 26376 27488 26382
rect 27436 26318 27488 26324
rect 27252 26240 27304 26246
rect 27252 26182 27304 26188
rect 27068 25696 27120 25702
rect 27068 25638 27120 25644
rect 26976 24812 27028 24818
rect 26976 24754 27028 24760
rect 27080 24614 27108 25638
rect 27264 25294 27292 26182
rect 27356 25294 27384 26318
rect 27252 25288 27304 25294
rect 27252 25230 27304 25236
rect 27344 25288 27396 25294
rect 27344 25230 27396 25236
rect 27448 25106 27476 26318
rect 27356 25078 27476 25106
rect 27620 25152 27672 25158
rect 27620 25094 27672 25100
rect 27160 24812 27212 24818
rect 27160 24754 27212 24760
rect 27068 24608 27120 24614
rect 27068 24550 27120 24556
rect 26792 22160 26844 22166
rect 26792 22102 26844 22108
rect 26620 22066 26740 22094
rect 26422 21856 26478 21865
rect 26422 21791 26478 21800
rect 26240 21480 26292 21486
rect 26332 21480 26384 21486
rect 26240 21422 26292 21428
rect 26330 21448 26332 21457
rect 26384 21448 26386 21457
rect 26330 21383 26386 21392
rect 25780 20868 25832 20874
rect 25780 20810 25832 20816
rect 25792 20534 25820 20810
rect 25780 20528 25832 20534
rect 25780 20470 25832 20476
rect 26056 20528 26108 20534
rect 26056 20470 26108 20476
rect 26068 19174 26096 20470
rect 26240 19916 26292 19922
rect 26240 19858 26292 19864
rect 26252 19394 26280 19858
rect 26332 19712 26384 19718
rect 26332 19654 26384 19660
rect 26160 19378 26280 19394
rect 26148 19372 26280 19378
rect 26200 19366 26280 19372
rect 26148 19314 26200 19320
rect 26344 19310 26372 19654
rect 26436 19310 26464 21791
rect 26620 21690 26648 22066
rect 27172 21690 27200 24754
rect 27250 23896 27306 23905
rect 27356 23866 27384 25078
rect 27436 24812 27488 24818
rect 27436 24754 27488 24760
rect 27528 24812 27580 24818
rect 27528 24754 27580 24760
rect 27448 24410 27476 24754
rect 27540 24410 27568 24754
rect 27436 24404 27488 24410
rect 27436 24346 27488 24352
rect 27528 24404 27580 24410
rect 27528 24346 27580 24352
rect 27632 24342 27660 25094
rect 27620 24336 27672 24342
rect 27620 24278 27672 24284
rect 27816 24206 27844 27542
rect 28368 27130 28396 31282
rect 28448 31272 28500 31278
rect 28448 31214 28500 31220
rect 28460 30666 28488 31214
rect 28448 30660 28500 30666
rect 28448 30602 28500 30608
rect 28460 28558 28488 30602
rect 28552 30394 28580 31282
rect 28632 31136 28684 31142
rect 28632 31078 28684 31084
rect 28724 31136 28776 31142
rect 28724 31078 28776 31084
rect 28644 30394 28672 31078
rect 28736 30802 28764 31078
rect 28724 30796 28776 30802
rect 28724 30738 28776 30744
rect 28828 30734 28856 32710
rect 28920 31346 28948 34478
rect 29736 33992 29788 33998
rect 29736 33934 29788 33940
rect 29092 33924 29144 33930
rect 29092 33866 29144 33872
rect 29104 33658 29132 33866
rect 29748 33658 29776 33934
rect 29092 33652 29144 33658
rect 29092 33594 29144 33600
rect 29736 33652 29788 33658
rect 29736 33594 29788 33600
rect 29184 33516 29236 33522
rect 29184 33458 29236 33464
rect 29276 33516 29328 33522
rect 29276 33458 29328 33464
rect 29196 33114 29224 33458
rect 29288 33114 29316 33458
rect 29644 33312 29696 33318
rect 29644 33254 29696 33260
rect 29184 33108 29236 33114
rect 29184 33050 29236 33056
rect 29276 33108 29328 33114
rect 29276 33050 29328 33056
rect 29196 32502 29224 33050
rect 29656 32978 29684 33254
rect 29736 33040 29788 33046
rect 29736 32982 29788 32988
rect 29644 32972 29696 32978
rect 29644 32914 29696 32920
rect 29552 32768 29604 32774
rect 29552 32710 29604 32716
rect 29564 32570 29592 32710
rect 29552 32564 29604 32570
rect 29552 32506 29604 32512
rect 29184 32496 29236 32502
rect 29184 32438 29236 32444
rect 29748 32230 29776 32982
rect 29736 32224 29788 32230
rect 29736 32166 29788 32172
rect 29748 31890 29776 32166
rect 29736 31884 29788 31890
rect 29736 31826 29788 31832
rect 29840 31754 29868 34546
rect 30104 34400 30156 34406
rect 30104 34342 30156 34348
rect 30116 34066 30144 34342
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 30104 34060 30156 34066
rect 30104 34002 30156 34008
rect 31392 34060 31444 34066
rect 31392 34002 31444 34008
rect 30472 33856 30524 33862
rect 30472 33798 30524 33804
rect 30564 33856 30616 33862
rect 30564 33798 30616 33804
rect 30484 33454 30512 33798
rect 30576 33658 30604 33798
rect 30564 33652 30616 33658
rect 30564 33594 30616 33600
rect 30288 33448 30340 33454
rect 30288 33390 30340 33396
rect 30472 33448 30524 33454
rect 30472 33390 30524 33396
rect 31208 33448 31260 33454
rect 31208 33390 31260 33396
rect 30104 33380 30156 33386
rect 30104 33322 30156 33328
rect 30012 33108 30064 33114
rect 30012 33050 30064 33056
rect 30024 32570 30052 33050
rect 30116 32994 30144 33322
rect 30116 32966 30236 32994
rect 30104 32904 30156 32910
rect 30104 32846 30156 32852
rect 30012 32564 30064 32570
rect 30012 32506 30064 32512
rect 29840 31726 29960 31754
rect 29932 31346 29960 31726
rect 30012 31748 30064 31754
rect 30012 31690 30064 31696
rect 30024 31346 30052 31690
rect 30116 31482 30144 32846
rect 30208 32570 30236 32966
rect 30300 32842 30328 33390
rect 31220 32910 31248 33390
rect 31404 33386 31432 34002
rect 31760 33992 31812 33998
rect 31760 33934 31812 33940
rect 31772 33658 31800 33934
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 31760 33652 31812 33658
rect 31760 33594 31812 33600
rect 31484 33516 31536 33522
rect 31852 33516 31904 33522
rect 31536 33476 31852 33504
rect 31484 33458 31536 33464
rect 31852 33458 31904 33464
rect 32312 33516 32364 33522
rect 32312 33458 32364 33464
rect 32036 33448 32088 33454
rect 32036 33390 32088 33396
rect 31392 33380 31444 33386
rect 31392 33322 31444 33328
rect 31484 33380 31536 33386
rect 31484 33322 31536 33328
rect 31208 32904 31260 32910
rect 31208 32846 31260 32852
rect 30288 32836 30340 32842
rect 30288 32778 30340 32784
rect 30196 32564 30248 32570
rect 30196 32506 30248 32512
rect 30208 31754 30236 32506
rect 30208 31726 30328 31754
rect 30104 31476 30156 31482
rect 30104 31418 30156 31424
rect 28908 31340 28960 31346
rect 28908 31282 28960 31288
rect 29920 31340 29972 31346
rect 29920 31282 29972 31288
rect 30012 31340 30064 31346
rect 30196 31340 30248 31346
rect 30064 31300 30144 31328
rect 30012 31282 30064 31288
rect 29092 31204 29144 31210
rect 29092 31146 29144 31152
rect 29104 30734 29132 31146
rect 28816 30728 28868 30734
rect 28816 30670 28868 30676
rect 29092 30728 29144 30734
rect 29092 30670 29144 30676
rect 28540 30388 28592 30394
rect 28540 30330 28592 30336
rect 28632 30388 28684 30394
rect 28632 30330 28684 30336
rect 28540 29776 28592 29782
rect 28540 29718 28592 29724
rect 28552 29646 28580 29718
rect 28828 29714 28856 30670
rect 28908 29776 28960 29782
rect 28908 29718 28960 29724
rect 28816 29708 28868 29714
rect 28816 29650 28868 29656
rect 28920 29646 28948 29718
rect 28540 29640 28592 29646
rect 28724 29640 28776 29646
rect 28540 29582 28592 29588
rect 28722 29608 28724 29617
rect 28908 29640 28960 29646
rect 28776 29608 28778 29617
rect 28908 29582 28960 29588
rect 28722 29543 28778 29552
rect 28632 29164 28684 29170
rect 28632 29106 28684 29112
rect 28540 29028 28592 29034
rect 28644 29016 28672 29106
rect 28592 28988 28672 29016
rect 28540 28970 28592 28976
rect 28816 28960 28868 28966
rect 28816 28902 28868 28908
rect 28828 28762 28856 28902
rect 28816 28756 28868 28762
rect 28816 28698 28868 28704
rect 28448 28552 28500 28558
rect 28448 28494 28500 28500
rect 28356 27124 28408 27130
rect 28356 27066 28408 27072
rect 27896 26988 27948 26994
rect 27896 26930 27948 26936
rect 27988 26988 28040 26994
rect 27988 26930 28040 26936
rect 27908 26586 27936 26930
rect 28000 26858 28028 26930
rect 27988 26852 28040 26858
rect 27988 26794 28040 26800
rect 27896 26580 27948 26586
rect 27896 26522 27948 26528
rect 27896 26308 27948 26314
rect 27896 26250 27948 26256
rect 27908 24274 27936 26250
rect 28000 25786 28028 26794
rect 28172 26376 28224 26382
rect 28172 26318 28224 26324
rect 28184 26042 28212 26318
rect 28172 26036 28224 26042
rect 28172 25978 28224 25984
rect 28000 25758 28120 25786
rect 28092 24886 28120 25758
rect 28172 24948 28224 24954
rect 28172 24890 28224 24896
rect 28080 24880 28132 24886
rect 28080 24822 28132 24828
rect 27896 24268 27948 24274
rect 27896 24210 27948 24216
rect 27804 24200 27856 24206
rect 27804 24142 27856 24148
rect 27436 24064 27488 24070
rect 27436 24006 27488 24012
rect 27620 24064 27672 24070
rect 27620 24006 27672 24012
rect 27250 23831 27252 23840
rect 27304 23831 27306 23840
rect 27344 23860 27396 23866
rect 27252 23802 27304 23808
rect 27344 23802 27396 23808
rect 27252 22976 27304 22982
rect 27252 22918 27304 22924
rect 27264 22030 27292 22918
rect 27356 22710 27384 23802
rect 27448 23118 27476 24006
rect 27632 23322 27660 24006
rect 27712 23656 27764 23662
rect 27712 23598 27764 23604
rect 27620 23316 27672 23322
rect 27620 23258 27672 23264
rect 27436 23112 27488 23118
rect 27436 23054 27488 23060
rect 27620 23112 27672 23118
rect 27620 23054 27672 23060
rect 27632 22710 27660 23054
rect 27344 22704 27396 22710
rect 27344 22646 27396 22652
rect 27620 22704 27672 22710
rect 27620 22646 27672 22652
rect 27724 22094 27752 23598
rect 27804 23112 27856 23118
rect 27908 23100 27936 24210
rect 27988 24200 28040 24206
rect 27988 24142 28040 24148
rect 27856 23072 27936 23100
rect 27804 23054 27856 23060
rect 27816 22642 27844 23054
rect 28000 22642 28028 24142
rect 28092 23662 28120 24822
rect 28184 24206 28212 24890
rect 28460 24834 28488 28494
rect 28632 28416 28684 28422
rect 28632 28358 28684 28364
rect 28540 28076 28592 28082
rect 28540 28018 28592 28024
rect 28552 26450 28580 28018
rect 28540 26444 28592 26450
rect 28540 26386 28592 26392
rect 28540 26240 28592 26246
rect 28540 26182 28592 26188
rect 28552 25906 28580 26182
rect 28540 25900 28592 25906
rect 28540 25842 28592 25848
rect 28552 24954 28580 25842
rect 28540 24948 28592 24954
rect 28540 24890 28592 24896
rect 28460 24806 28580 24834
rect 28172 24200 28224 24206
rect 28172 24142 28224 24148
rect 28172 23724 28224 23730
rect 28172 23666 28224 23672
rect 28080 23656 28132 23662
rect 28080 23598 28132 23604
rect 27804 22636 27856 22642
rect 27804 22578 27856 22584
rect 27988 22636 28040 22642
rect 27988 22578 28040 22584
rect 27540 22066 27752 22094
rect 27252 22024 27304 22030
rect 27252 21966 27304 21972
rect 26516 21684 26568 21690
rect 26516 21626 26568 21632
rect 26608 21684 26660 21690
rect 26608 21626 26660 21632
rect 27160 21684 27212 21690
rect 27160 21626 27212 21632
rect 26528 21486 26556 21626
rect 27264 21554 27292 21966
rect 27540 21894 27568 22066
rect 27528 21888 27580 21894
rect 27528 21830 27580 21836
rect 27712 21888 27764 21894
rect 27712 21830 27764 21836
rect 27620 21684 27672 21690
rect 27620 21626 27672 21632
rect 27252 21548 27304 21554
rect 27252 21490 27304 21496
rect 26516 21480 26568 21486
rect 26516 21422 26568 21428
rect 27632 21418 27660 21626
rect 27620 21412 27672 21418
rect 27620 21354 27672 21360
rect 27344 21344 27396 21350
rect 27344 21286 27396 21292
rect 27356 21078 27384 21286
rect 27344 21072 27396 21078
rect 27620 21072 27672 21078
rect 27344 21014 27396 21020
rect 27540 21020 27620 21026
rect 27540 21014 27672 21020
rect 27540 20998 27660 21014
rect 26792 20800 26844 20806
rect 26790 20768 26792 20777
rect 27540 20777 27568 20998
rect 27724 20942 27752 21830
rect 28000 21554 28028 22578
rect 27988 21548 28040 21554
rect 27988 21490 28040 21496
rect 27894 21448 27950 21457
rect 28000 21434 28028 21490
rect 27950 21406 28028 21434
rect 27894 21383 27950 21392
rect 27712 20936 27764 20942
rect 27712 20878 27764 20884
rect 26844 20768 26846 20777
rect 26790 20703 26846 20712
rect 27526 20768 27582 20777
rect 27526 20703 27582 20712
rect 27804 20596 27856 20602
rect 27804 20538 27856 20544
rect 26976 20460 27028 20466
rect 26976 20402 27028 20408
rect 26516 19984 26568 19990
rect 26516 19926 26568 19932
rect 26332 19304 26384 19310
rect 26332 19246 26384 19252
rect 26424 19304 26476 19310
rect 26424 19246 26476 19252
rect 25688 19168 25740 19174
rect 25688 19110 25740 19116
rect 26056 19168 26108 19174
rect 26056 19110 26108 19116
rect 26240 19168 26292 19174
rect 26528 19156 26556 19926
rect 26988 19514 27016 20402
rect 27068 20256 27120 20262
rect 27068 20198 27120 20204
rect 26976 19508 27028 19514
rect 26976 19450 27028 19456
rect 27080 19394 27108 20198
rect 27252 20052 27304 20058
rect 27252 19994 27304 20000
rect 27264 19854 27292 19994
rect 27816 19854 27844 20538
rect 28184 19922 28212 23666
rect 28264 22636 28316 22642
rect 28264 22578 28316 22584
rect 28276 22030 28304 22578
rect 28552 22234 28580 24806
rect 28644 24410 28672 28358
rect 28724 27464 28776 27470
rect 28724 27406 28776 27412
rect 28736 27062 28764 27406
rect 28920 27334 28948 29582
rect 28998 29336 29054 29345
rect 28998 29271 29054 29280
rect 29012 29170 29040 29271
rect 29000 29164 29052 29170
rect 29000 29106 29052 29112
rect 29104 28762 29132 30670
rect 29932 30258 29960 31282
rect 29920 30252 29972 30258
rect 29920 30194 29972 30200
rect 29644 30184 29696 30190
rect 29696 30132 29960 30138
rect 29644 30126 29960 30132
rect 29656 30110 29960 30126
rect 29932 30054 29960 30110
rect 29460 30048 29512 30054
rect 29460 29990 29512 29996
rect 29644 30048 29696 30054
rect 29644 29990 29696 29996
rect 29920 30048 29972 30054
rect 29920 29990 29972 29996
rect 29092 28756 29144 28762
rect 29092 28698 29144 28704
rect 29472 27606 29500 29990
rect 29656 29170 29684 29990
rect 29644 29164 29696 29170
rect 29644 29106 29696 29112
rect 29736 28552 29788 28558
rect 29736 28494 29788 28500
rect 29460 27600 29512 27606
rect 29460 27542 29512 27548
rect 29748 27538 29776 28494
rect 29736 27532 29788 27538
rect 29736 27474 29788 27480
rect 29932 27470 29960 29990
rect 30012 29572 30064 29578
rect 30012 29514 30064 29520
rect 30024 29170 30052 29514
rect 30116 29170 30144 31300
rect 30196 31282 30248 31288
rect 30208 30326 30236 31282
rect 30196 30320 30248 30326
rect 30196 30262 30248 30268
rect 30012 29164 30064 29170
rect 30012 29106 30064 29112
rect 30104 29164 30156 29170
rect 30104 29106 30156 29112
rect 30116 28626 30144 29106
rect 30104 28620 30156 28626
rect 30104 28562 30156 28568
rect 29368 27464 29420 27470
rect 29368 27406 29420 27412
rect 29920 27464 29972 27470
rect 29920 27406 29972 27412
rect 28908 27328 28960 27334
rect 28908 27270 28960 27276
rect 28724 27056 28776 27062
rect 28724 26998 28776 27004
rect 29184 26988 29236 26994
rect 29184 26930 29236 26936
rect 29196 26586 29224 26930
rect 29184 26580 29236 26586
rect 29184 26522 29236 26528
rect 28724 26444 28776 26450
rect 28776 26404 28856 26432
rect 28724 26386 28776 26392
rect 28828 26330 28856 26404
rect 28908 26376 28960 26382
rect 28828 26324 28908 26330
rect 28828 26318 28960 26324
rect 28828 26302 28948 26318
rect 29380 26314 29408 27406
rect 29644 27396 29696 27402
rect 29644 27338 29696 27344
rect 30012 27396 30064 27402
rect 30012 27338 30064 27344
rect 29552 27328 29604 27334
rect 29552 27270 29604 27276
rect 29564 26314 29592 27270
rect 29656 26586 29684 27338
rect 30024 27062 30052 27338
rect 30300 27112 30328 31726
rect 31024 31272 31076 31278
rect 31024 31214 31076 31220
rect 31300 31272 31352 31278
rect 31300 31214 31352 31220
rect 30380 31204 30432 31210
rect 30380 31146 30432 31152
rect 30392 30802 30420 31146
rect 30380 30796 30432 30802
rect 30380 30738 30432 30744
rect 30932 30592 30984 30598
rect 30932 30534 30984 30540
rect 30380 30252 30432 30258
rect 30380 30194 30432 30200
rect 30392 29646 30420 30194
rect 30944 30190 30972 30534
rect 30932 30184 30984 30190
rect 30932 30126 30984 30132
rect 31036 29850 31064 31214
rect 31024 29844 31076 29850
rect 31024 29786 31076 29792
rect 30380 29640 30432 29646
rect 30380 29582 30432 29588
rect 30840 29640 30892 29646
rect 30840 29582 30892 29588
rect 30852 28626 30880 29582
rect 31024 29028 31076 29034
rect 31024 28970 31076 28976
rect 30840 28620 30892 28626
rect 30840 28562 30892 28568
rect 30656 28552 30708 28558
rect 30656 28494 30708 28500
rect 30748 28552 30800 28558
rect 30748 28494 30800 28500
rect 30380 27464 30432 27470
rect 30380 27406 30432 27412
rect 30116 27084 30328 27112
rect 30012 27056 30064 27062
rect 30012 26998 30064 27004
rect 29644 26580 29696 26586
rect 29644 26522 29696 26528
rect 29368 26308 29420 26314
rect 29368 26250 29420 26256
rect 29552 26308 29604 26314
rect 29552 26250 29604 26256
rect 29184 26240 29236 26246
rect 29184 26182 29236 26188
rect 29092 26036 29144 26042
rect 29092 25978 29144 25984
rect 29104 25838 29132 25978
rect 29196 25974 29224 26182
rect 29184 25968 29236 25974
rect 29184 25910 29236 25916
rect 29092 25832 29144 25838
rect 29092 25774 29144 25780
rect 29000 24948 29052 24954
rect 29000 24890 29052 24896
rect 28724 24744 28776 24750
rect 28724 24686 28776 24692
rect 28632 24404 28684 24410
rect 28632 24346 28684 24352
rect 28736 24206 28764 24686
rect 29012 24410 29040 24890
rect 29000 24404 29052 24410
rect 29000 24346 29052 24352
rect 28816 24268 28868 24274
rect 28816 24210 28868 24216
rect 28724 24200 28776 24206
rect 28724 24142 28776 24148
rect 28828 23730 28856 24210
rect 28908 24200 28960 24206
rect 28960 24148 29040 24154
rect 28908 24142 29040 24148
rect 28920 24126 29040 24142
rect 28908 24064 28960 24070
rect 28908 24006 28960 24012
rect 28816 23724 28868 23730
rect 28816 23666 28868 23672
rect 28828 23322 28856 23666
rect 28816 23316 28868 23322
rect 28816 23258 28868 23264
rect 28724 23180 28776 23186
rect 28724 23122 28776 23128
rect 28736 22438 28764 23122
rect 28828 23118 28856 23258
rect 28816 23112 28868 23118
rect 28816 23054 28868 23060
rect 28724 22432 28776 22438
rect 28724 22374 28776 22380
rect 28448 22228 28500 22234
rect 28448 22170 28500 22176
rect 28540 22228 28592 22234
rect 28540 22170 28592 22176
rect 28264 22024 28316 22030
rect 28264 21966 28316 21972
rect 28276 21690 28304 21966
rect 28264 21684 28316 21690
rect 28264 21626 28316 21632
rect 28460 21350 28488 22170
rect 28552 22098 28580 22170
rect 28920 22098 28948 24006
rect 29012 23866 29040 24126
rect 29000 23860 29052 23866
rect 29000 23802 29052 23808
rect 29000 22160 29052 22166
rect 29000 22102 29052 22108
rect 28540 22092 28592 22098
rect 28540 22034 28592 22040
rect 28908 22092 28960 22098
rect 28908 22034 28960 22040
rect 29012 21554 29040 22102
rect 28724 21548 28776 21554
rect 28724 21490 28776 21496
rect 29000 21548 29052 21554
rect 29000 21490 29052 21496
rect 28632 21480 28684 21486
rect 28632 21422 28684 21428
rect 28448 21344 28500 21350
rect 28448 21286 28500 21292
rect 28644 20602 28672 21422
rect 28736 21146 28764 21490
rect 28816 21480 28868 21486
rect 28816 21422 28868 21428
rect 28724 21140 28776 21146
rect 28724 21082 28776 21088
rect 28828 21078 28856 21422
rect 28816 21072 28868 21078
rect 28816 21014 28868 21020
rect 28632 20596 28684 20602
rect 28632 20538 28684 20544
rect 29104 19990 29132 25774
rect 29196 24750 29224 25910
rect 29276 24812 29328 24818
rect 29276 24754 29328 24760
rect 29184 24744 29236 24750
rect 29184 24686 29236 24692
rect 29196 23186 29224 24686
rect 29288 23798 29316 24754
rect 29276 23792 29328 23798
rect 29276 23734 29328 23740
rect 29276 23656 29328 23662
rect 29276 23598 29328 23604
rect 29184 23180 29236 23186
rect 29184 23122 29236 23128
rect 29288 23050 29316 23598
rect 29184 23044 29236 23050
rect 29184 22986 29236 22992
rect 29276 23044 29328 23050
rect 29276 22986 29328 22992
rect 29196 22778 29224 22986
rect 29184 22772 29236 22778
rect 29184 22714 29236 22720
rect 29196 20058 29224 22714
rect 29288 22030 29316 22986
rect 29276 22024 29328 22030
rect 29276 21966 29328 21972
rect 29184 20052 29236 20058
rect 29184 19994 29236 20000
rect 29092 19984 29144 19990
rect 29092 19926 29144 19932
rect 28172 19916 28224 19922
rect 28172 19858 28224 19864
rect 27252 19848 27304 19854
rect 27252 19790 27304 19796
rect 27344 19848 27396 19854
rect 27344 19790 27396 19796
rect 27804 19848 27856 19854
rect 27804 19790 27856 19796
rect 28632 19848 28684 19854
rect 28632 19790 28684 19796
rect 27252 19712 27304 19718
rect 27252 19654 27304 19660
rect 27160 19440 27212 19446
rect 27080 19388 27160 19394
rect 27080 19382 27212 19388
rect 27080 19366 27200 19382
rect 26700 19304 26752 19310
rect 26700 19246 26752 19252
rect 26292 19128 26556 19156
rect 26240 19110 26292 19116
rect 26068 18426 26096 19110
rect 26056 18420 26108 18426
rect 26056 18362 26108 18368
rect 26056 18080 26108 18086
rect 26056 18022 26108 18028
rect 25504 17808 25556 17814
rect 25504 17750 25556 17756
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 25148 17338 25176 17682
rect 25504 17672 25556 17678
rect 25504 17614 25556 17620
rect 25228 17604 25280 17610
rect 25228 17546 25280 17552
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 25044 16244 25096 16250
rect 25044 16186 25096 16192
rect 25240 16153 25268 17546
rect 25412 17196 25464 17202
rect 25412 17138 25464 17144
rect 25226 16144 25282 16153
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 25136 16108 25188 16114
rect 25226 16079 25282 16088
rect 25136 16050 25188 16056
rect 24952 16040 25004 16046
rect 24952 15982 25004 15988
rect 24964 14890 24992 15982
rect 25056 15910 25084 16050
rect 25044 15904 25096 15910
rect 25044 15846 25096 15852
rect 25148 15570 25176 16050
rect 25136 15564 25188 15570
rect 25136 15506 25188 15512
rect 25044 15428 25096 15434
rect 25044 15370 25096 15376
rect 24952 14884 25004 14890
rect 24952 14826 25004 14832
rect 24872 14572 24992 14600
rect 24676 14476 24728 14482
rect 24780 14470 24900 14498
rect 24676 14418 24728 14424
rect 24768 14340 24820 14346
rect 24768 14282 24820 14288
rect 24676 13728 24728 13734
rect 24676 13670 24728 13676
rect 24688 12850 24716 13670
rect 24676 12844 24728 12850
rect 24676 12786 24728 12792
rect 24688 12374 24716 12786
rect 24676 12368 24728 12374
rect 24676 12310 24728 12316
rect 24780 12186 24808 14282
rect 24872 14278 24900 14470
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24964 13802 24992 14572
rect 24952 13796 25004 13802
rect 24952 13738 25004 13744
rect 24872 13258 24992 13274
rect 24860 13252 24992 13258
rect 24912 13246 24992 13252
rect 24860 13194 24912 13200
rect 24858 13152 24914 13161
rect 24858 13087 24914 13096
rect 24872 12238 24900 13087
rect 24584 12164 24636 12170
rect 24584 12106 24636 12112
rect 24688 12158 24808 12186
rect 24860 12232 24912 12238
rect 24860 12174 24912 12180
rect 24688 12102 24716 12158
rect 24676 12096 24728 12102
rect 24596 12044 24676 12050
rect 24596 12038 24728 12044
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24596 12022 24716 12038
rect 24398 11656 24454 11665
rect 24398 11591 24454 11600
rect 24308 11552 24360 11558
rect 24308 11494 24360 11500
rect 24492 11552 24544 11558
rect 24492 11494 24544 11500
rect 24504 11370 24532 11494
rect 24320 11354 24532 11370
rect 24320 11348 24544 11354
rect 24320 11342 24492 11348
rect 24216 11280 24268 11286
rect 24216 11222 24268 11228
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 24032 10532 24084 10538
rect 24032 10474 24084 10480
rect 23846 10296 23902 10305
rect 23846 10231 23848 10240
rect 23900 10231 23902 10240
rect 23848 10202 23900 10208
rect 24044 10146 24072 10474
rect 24124 10260 24176 10266
rect 24124 10202 24176 10208
rect 23860 10118 24072 10146
rect 23860 10062 23888 10118
rect 23848 10056 23900 10062
rect 23848 9998 23900 10004
rect 23952 9654 23980 10118
rect 24032 10056 24084 10062
rect 24136 10044 24164 10202
rect 24084 10016 24164 10044
rect 24032 9998 24084 10004
rect 24216 9716 24268 9722
rect 24216 9658 24268 9664
rect 23940 9648 23992 9654
rect 23940 9590 23992 9596
rect 23572 9580 23624 9586
rect 23572 9522 23624 9528
rect 23664 9580 23716 9586
rect 23664 9522 23716 9528
rect 23756 9580 23808 9586
rect 23756 9522 23808 9528
rect 23492 9438 23612 9466
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 23308 8588 23428 8616
rect 23296 8492 23348 8498
rect 23216 8452 23296 8480
rect 23112 8434 23164 8440
rect 23296 8434 23348 8440
rect 22560 8356 22612 8362
rect 22560 8298 22612 8304
rect 22652 8356 22704 8362
rect 22652 8298 22704 8304
rect 22468 7812 22520 7818
rect 22020 7772 22468 7800
rect 21916 7754 21968 7760
rect 22468 7754 22520 7760
rect 22376 7540 22428 7546
rect 22376 7482 22428 7488
rect 21914 7440 21970 7449
rect 21824 7404 21876 7410
rect 21914 7375 21916 7384
rect 21824 7346 21876 7352
rect 21968 7375 21970 7384
rect 22192 7404 22244 7410
rect 21916 7346 21968 7352
rect 22192 7346 22244 7352
rect 22204 7206 22232 7346
rect 22284 7336 22336 7342
rect 22284 7278 22336 7284
rect 22192 7200 22244 7206
rect 22192 7142 22244 7148
rect 22296 7002 22324 7278
rect 22284 6996 22336 7002
rect 22284 6938 22336 6944
rect 22008 6792 22060 6798
rect 21456 6384 21508 6390
rect 21456 6326 21508 6332
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 21376 5574 21404 6258
rect 21468 5710 21496 6326
rect 21560 6254 21588 6752
rect 21638 6760 21694 6769
rect 21744 6752 22008 6780
rect 22192 6792 22244 6798
rect 22008 6734 22060 6740
rect 22112 6740 22192 6746
rect 22112 6734 22244 6740
rect 21638 6695 21694 6704
rect 22112 6718 22232 6734
rect 21652 6662 21680 6695
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 22112 6458 22140 6718
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 22284 6656 22336 6662
rect 22284 6598 22336 6604
rect 22204 6458 22232 6598
rect 22296 6458 22324 6598
rect 22388 6458 22416 7482
rect 22480 7410 22508 7754
rect 22572 7546 22600 8298
rect 22560 7540 22612 7546
rect 22560 7482 22612 7488
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22100 6452 22152 6458
rect 22100 6394 22152 6400
rect 22192 6452 22244 6458
rect 22192 6394 22244 6400
rect 22284 6452 22336 6458
rect 22284 6394 22336 6400
rect 22376 6452 22428 6458
rect 22376 6394 22428 6400
rect 21914 6352 21970 6361
rect 22480 6338 22508 7346
rect 22664 6882 22692 8298
rect 22756 8022 22784 8434
rect 22744 8016 22796 8022
rect 22744 7958 22796 7964
rect 22848 7002 22876 8434
rect 23400 8022 23428 8588
rect 23492 8566 23520 9318
rect 23480 8560 23532 8566
rect 23480 8502 23532 8508
rect 23388 8016 23440 8022
rect 23388 7958 23440 7964
rect 23112 7948 23164 7954
rect 23112 7890 23164 7896
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 23032 7410 23060 7482
rect 23124 7410 23152 7890
rect 23204 7540 23256 7546
rect 23204 7482 23256 7488
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 23112 7404 23164 7410
rect 23112 7346 23164 7352
rect 23032 7018 23060 7346
rect 22836 6996 22888 7002
rect 23032 6990 23152 7018
rect 22836 6938 22888 6944
rect 22664 6854 22876 6882
rect 22560 6724 22612 6730
rect 22560 6666 22612 6672
rect 22572 6361 22600 6666
rect 21914 6287 21916 6296
rect 21968 6287 21970 6296
rect 22008 6316 22060 6322
rect 21916 6258 21968 6264
rect 22008 6258 22060 6264
rect 22296 6310 22508 6338
rect 22558 6352 22614 6361
rect 21548 6248 21600 6254
rect 21548 6190 21600 6196
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 21364 5568 21416 5574
rect 21364 5510 21416 5516
rect 21364 4548 21416 4554
rect 21364 4490 21416 4496
rect 21376 4282 21404 4490
rect 21364 4276 21416 4282
rect 21364 4218 21416 4224
rect 20996 4208 21048 4214
rect 20996 4150 21048 4156
rect 21560 4146 21588 6190
rect 22020 5642 22048 6258
rect 22296 6186 22324 6310
rect 22558 6287 22614 6296
rect 22848 6254 22876 6854
rect 22928 6792 22980 6798
rect 22928 6734 22980 6740
rect 23020 6792 23072 6798
rect 23124 6780 23152 6990
rect 23072 6752 23152 6780
rect 23020 6734 23072 6740
rect 22940 6497 22968 6734
rect 23124 6662 23152 6752
rect 23020 6656 23072 6662
rect 23020 6598 23072 6604
rect 23112 6656 23164 6662
rect 23112 6598 23164 6604
rect 22926 6488 22982 6497
rect 23032 6458 23060 6598
rect 22926 6423 22982 6432
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 23216 6322 23244 7482
rect 23294 7032 23350 7041
rect 23492 6984 23520 8502
rect 23584 8498 23612 9438
rect 23664 9172 23716 9178
rect 23664 9114 23716 9120
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23584 8294 23612 8434
rect 23572 8288 23624 8294
rect 23572 8230 23624 8236
rect 23294 6967 23350 6976
rect 23308 6866 23336 6967
rect 23400 6956 23520 6984
rect 23296 6860 23348 6866
rect 23296 6802 23348 6808
rect 23296 6724 23348 6730
rect 23400 6712 23428 6956
rect 23478 6896 23534 6905
rect 23478 6831 23534 6840
rect 23348 6684 23428 6712
rect 23296 6666 23348 6672
rect 23492 6458 23520 6831
rect 23676 6798 23704 9114
rect 23768 8945 23796 9522
rect 24032 9444 24084 9450
rect 24032 9386 24084 9392
rect 23754 8936 23810 8945
rect 23754 8871 23810 8880
rect 24044 8498 24072 9386
rect 23848 8492 23900 8498
rect 23848 8434 23900 8440
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 23756 8288 23808 8294
rect 23756 8230 23808 8236
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23664 6792 23716 6798
rect 23664 6734 23716 6740
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23204 6316 23256 6322
rect 23204 6258 23256 6264
rect 22836 6248 22888 6254
rect 22836 6190 22888 6196
rect 22284 6180 22336 6186
rect 22284 6122 22336 6128
rect 22008 5636 22060 5642
rect 22008 5578 22060 5584
rect 22192 5296 22244 5302
rect 22192 5238 22244 5244
rect 21916 5024 21968 5030
rect 21916 4966 21968 4972
rect 21928 4146 21956 4966
rect 22204 4282 22232 5238
rect 22296 5234 22324 6122
rect 23388 5840 23440 5846
rect 23388 5782 23440 5788
rect 22560 5772 22612 5778
rect 22560 5714 22612 5720
rect 22572 5370 22600 5714
rect 23294 5536 23350 5545
rect 23294 5471 23350 5480
rect 22560 5364 22612 5370
rect 22560 5306 22612 5312
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 22572 5166 22600 5306
rect 23308 5302 23336 5471
rect 23400 5302 23428 5782
rect 23296 5296 23348 5302
rect 23296 5238 23348 5244
rect 23388 5296 23440 5302
rect 23388 5238 23440 5244
rect 22836 5228 22888 5234
rect 22836 5170 22888 5176
rect 22560 5160 22612 5166
rect 22560 5102 22612 5108
rect 22744 5024 22796 5030
rect 22744 4966 22796 4972
rect 22652 4548 22704 4554
rect 22652 4490 22704 4496
rect 22664 4282 22692 4490
rect 22756 4486 22784 4966
rect 22848 4826 22876 5170
rect 22836 4820 22888 4826
rect 22836 4762 22888 4768
rect 23308 4486 23336 5238
rect 23400 4690 23428 5238
rect 23388 4684 23440 4690
rect 23388 4626 23440 4632
rect 23584 4622 23612 6734
rect 23768 6474 23796 8230
rect 23860 8090 23888 8434
rect 23848 8084 23900 8090
rect 23848 8026 23900 8032
rect 23846 7576 23902 7585
rect 23846 7511 23902 7520
rect 23676 6446 23796 6474
rect 23860 6458 23888 7511
rect 23952 6662 23980 8434
rect 24228 7410 24256 9658
rect 24320 8537 24348 11342
rect 24492 11290 24544 11296
rect 24492 10804 24544 10810
rect 24492 10746 24544 10752
rect 24504 9330 24532 10746
rect 24596 9450 24624 12022
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24780 10985 24808 11630
rect 24766 10976 24822 10985
rect 24766 10911 24822 10920
rect 24768 10600 24820 10606
rect 24768 10542 24820 10548
rect 24676 9648 24728 9654
rect 24674 9616 24676 9625
rect 24728 9616 24730 9625
rect 24674 9551 24730 9560
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 24584 9444 24636 9450
rect 24584 9386 24636 9392
rect 24688 9330 24716 9454
rect 24504 9302 24716 9330
rect 24398 9208 24454 9217
rect 24398 9143 24454 9152
rect 24412 9042 24440 9143
rect 24400 9036 24452 9042
rect 24400 8978 24452 8984
rect 24306 8528 24362 8537
rect 24306 8463 24362 8472
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 24308 7200 24360 7206
rect 24308 7142 24360 7148
rect 23940 6656 23992 6662
rect 23940 6598 23992 6604
rect 23848 6452 23900 6458
rect 23676 5914 23704 6446
rect 23848 6394 23900 6400
rect 23664 5908 23716 5914
rect 23664 5850 23716 5856
rect 23676 5166 23704 5850
rect 23952 5250 23980 6598
rect 24320 6390 24348 7142
rect 24504 6458 24532 9302
rect 24584 8968 24636 8974
rect 24584 8910 24636 8916
rect 24596 8090 24624 8910
rect 24584 8084 24636 8090
rect 24584 8026 24636 8032
rect 24676 7404 24728 7410
rect 24676 7346 24728 7352
rect 24688 7206 24716 7346
rect 24676 7200 24728 7206
rect 24676 7142 24728 7148
rect 24492 6452 24544 6458
rect 24492 6394 24544 6400
rect 24308 6384 24360 6390
rect 24308 6326 24360 6332
rect 24504 5574 24532 6394
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 24596 5642 24624 6258
rect 24584 5636 24636 5642
rect 24584 5578 24636 5584
rect 24492 5568 24544 5574
rect 24492 5510 24544 5516
rect 23952 5234 24348 5250
rect 23940 5228 24348 5234
rect 23992 5222 24348 5228
rect 23940 5170 23992 5176
rect 23664 5160 23716 5166
rect 23664 5102 23716 5108
rect 24216 5024 24268 5030
rect 24216 4966 24268 4972
rect 24228 4826 24256 4966
rect 24320 4826 24348 5222
rect 24216 4820 24268 4826
rect 24216 4762 24268 4768
rect 24308 4820 24360 4826
rect 24308 4762 24360 4768
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 22744 4480 22796 4486
rect 22744 4422 22796 4428
rect 22928 4480 22980 4486
rect 22928 4422 22980 4428
rect 23296 4480 23348 4486
rect 23296 4422 23348 4428
rect 22192 4276 22244 4282
rect 22192 4218 22244 4224
rect 22652 4276 22704 4282
rect 22652 4218 22704 4224
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 21916 4140 21968 4146
rect 21916 4082 21968 4088
rect 22940 3534 22968 4422
rect 23388 4276 23440 4282
rect 23388 4218 23440 4224
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 22928 3528 22980 3534
rect 22928 3470 22980 3476
rect 19708 3392 19760 3398
rect 19708 3334 19760 3340
rect 20352 3392 20404 3398
rect 20352 3334 20404 3340
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 20364 3126 20392 3334
rect 20352 3120 20404 3126
rect 20352 3062 20404 3068
rect 20640 2990 20668 3470
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 22192 3392 22244 3398
rect 22192 3334 22244 3340
rect 20916 3194 20944 3334
rect 22020 3194 22048 3334
rect 22204 3194 22232 3334
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 23400 3126 23428 4218
rect 23584 3194 23612 4558
rect 24584 3596 24636 3602
rect 24584 3538 24636 3544
rect 24596 3505 24624 3538
rect 24582 3496 24638 3505
rect 24688 3466 24716 7142
rect 24780 5098 24808 10542
rect 24872 10033 24900 12038
rect 24964 11150 24992 13246
rect 25056 13002 25084 15370
rect 25136 15360 25188 15366
rect 25136 15302 25188 15308
rect 25148 13161 25176 15302
rect 25240 15162 25268 16079
rect 25320 15904 25372 15910
rect 25320 15846 25372 15852
rect 25332 15706 25360 15846
rect 25320 15700 25372 15706
rect 25320 15642 25372 15648
rect 25320 15564 25372 15570
rect 25320 15506 25372 15512
rect 25228 15156 25280 15162
rect 25228 15098 25280 15104
rect 25228 13320 25280 13326
rect 25332 13308 25360 15506
rect 25424 14385 25452 17138
rect 25516 16454 25544 17614
rect 25964 17536 26016 17542
rect 25964 17478 26016 17484
rect 25976 17338 26004 17478
rect 25872 17332 25924 17338
rect 25872 17274 25924 17280
rect 25964 17332 26016 17338
rect 25964 17274 26016 17280
rect 25688 16516 25740 16522
rect 25688 16458 25740 16464
rect 25504 16448 25556 16454
rect 25504 16390 25556 16396
rect 25516 15366 25544 16390
rect 25596 15496 25648 15502
rect 25596 15438 25648 15444
rect 25504 15360 25556 15366
rect 25502 15328 25504 15337
rect 25556 15328 25558 15337
rect 25502 15263 25558 15272
rect 25504 15020 25556 15026
rect 25504 14962 25556 14968
rect 25410 14376 25466 14385
rect 25410 14311 25466 14320
rect 25424 13546 25452 14311
rect 25516 14074 25544 14962
rect 25608 14890 25636 15438
rect 25700 15162 25728 16458
rect 25884 16454 25912 17274
rect 25872 16448 25924 16454
rect 25872 16390 25924 16396
rect 25778 16144 25834 16153
rect 25778 16079 25780 16088
rect 25832 16079 25834 16088
rect 25964 16108 26016 16114
rect 25780 16050 25832 16056
rect 25964 16050 26016 16056
rect 25872 15972 25924 15978
rect 25872 15914 25924 15920
rect 25778 15464 25834 15473
rect 25778 15399 25780 15408
rect 25832 15399 25834 15408
rect 25780 15370 25832 15376
rect 25778 15328 25834 15337
rect 25778 15263 25834 15272
rect 25688 15156 25740 15162
rect 25688 15098 25740 15104
rect 25596 14884 25648 14890
rect 25596 14826 25648 14832
rect 25688 14476 25740 14482
rect 25688 14418 25740 14424
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25424 13518 25544 13546
rect 25412 13456 25464 13462
rect 25412 13398 25464 13404
rect 25280 13280 25360 13308
rect 25228 13262 25280 13268
rect 25134 13152 25190 13161
rect 25134 13087 25190 13096
rect 25056 12974 25176 13002
rect 25042 12880 25098 12889
rect 25042 12815 25044 12824
rect 25096 12815 25098 12824
rect 25044 12786 25096 12792
rect 25044 12708 25096 12714
rect 25044 12650 25096 12656
rect 25056 12374 25084 12650
rect 25044 12368 25096 12374
rect 25044 12310 25096 12316
rect 25044 12096 25096 12102
rect 25148 12084 25176 12974
rect 25096 12056 25176 12084
rect 25044 12038 25096 12044
rect 25056 11937 25084 12038
rect 25042 11928 25098 11937
rect 25042 11863 25098 11872
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 24952 11008 25004 11014
rect 24952 10950 25004 10956
rect 24964 10180 24992 10950
rect 25056 10282 25084 11863
rect 25136 11824 25188 11830
rect 25136 11766 25188 11772
rect 25148 11150 25176 11766
rect 25136 11144 25188 11150
rect 25136 11086 25188 11092
rect 25148 10470 25176 11086
rect 25240 10674 25268 13262
rect 25318 13016 25374 13025
rect 25424 12986 25452 13398
rect 25516 13258 25544 13518
rect 25700 13462 25728 14418
rect 25596 13456 25648 13462
rect 25596 13398 25648 13404
rect 25688 13456 25740 13462
rect 25688 13398 25740 13404
rect 25504 13252 25556 13258
rect 25504 13194 25556 13200
rect 25318 12951 25320 12960
rect 25372 12951 25374 12960
rect 25412 12980 25464 12986
rect 25320 12922 25372 12928
rect 25412 12922 25464 12928
rect 25516 12866 25544 13194
rect 25332 12838 25544 12866
rect 25332 11830 25360 12838
rect 25608 12646 25636 13398
rect 25688 13320 25740 13326
rect 25792 13297 25820 15263
rect 25688 13262 25740 13268
rect 25778 13288 25834 13297
rect 25700 12646 25728 13262
rect 25884 13258 25912 15914
rect 25976 15745 26004 16050
rect 25962 15736 26018 15745
rect 26068 15706 26096 18022
rect 26148 17060 26200 17066
rect 26148 17002 26200 17008
rect 25962 15671 26018 15680
rect 26056 15700 26108 15706
rect 25976 15638 26004 15671
rect 26056 15642 26108 15648
rect 25964 15632 26016 15638
rect 25964 15574 26016 15580
rect 26056 15496 26108 15502
rect 26160 15473 26188 17002
rect 26056 15438 26108 15444
rect 26146 15464 26202 15473
rect 25964 15360 26016 15366
rect 25964 15302 26016 15308
rect 25976 14618 26004 15302
rect 25964 14612 26016 14618
rect 25964 14554 26016 14560
rect 25964 13456 26016 13462
rect 25964 13398 26016 13404
rect 25778 13223 25834 13232
rect 25872 13252 25924 13258
rect 25872 13194 25924 13200
rect 25780 13184 25832 13190
rect 25780 13126 25832 13132
rect 25792 12782 25820 13126
rect 25780 12776 25832 12782
rect 25780 12718 25832 12724
rect 25596 12640 25648 12646
rect 25410 12608 25466 12617
rect 25596 12582 25648 12588
rect 25688 12640 25740 12646
rect 25688 12582 25740 12588
rect 25410 12543 25466 12552
rect 25424 12170 25452 12543
rect 25502 12472 25558 12481
rect 25558 12416 25636 12434
rect 25502 12407 25636 12416
rect 25516 12406 25636 12407
rect 25412 12164 25464 12170
rect 25412 12106 25464 12112
rect 25504 12096 25556 12102
rect 25424 12044 25504 12050
rect 25424 12038 25556 12044
rect 25424 12022 25544 12038
rect 25320 11824 25372 11830
rect 25320 11766 25372 11772
rect 25424 10810 25452 12022
rect 25504 11688 25556 11694
rect 25502 11656 25504 11665
rect 25556 11656 25558 11665
rect 25502 11591 25558 11600
rect 25504 11144 25556 11150
rect 25502 11112 25504 11121
rect 25556 11112 25558 11121
rect 25502 11047 25558 11056
rect 25502 10840 25558 10849
rect 25412 10804 25464 10810
rect 25502 10775 25558 10784
rect 25412 10746 25464 10752
rect 25228 10668 25280 10674
rect 25228 10610 25280 10616
rect 25136 10464 25188 10470
rect 25136 10406 25188 10412
rect 25056 10254 25176 10282
rect 24964 10152 25084 10180
rect 24952 10056 25004 10062
rect 24858 10024 24914 10033
rect 24952 9998 25004 10004
rect 24858 9959 24914 9968
rect 24872 9654 24900 9959
rect 24964 9722 24992 9998
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 24860 9648 24912 9654
rect 24860 9590 24912 9596
rect 25056 9042 25084 10152
rect 25148 9625 25176 10254
rect 25134 9616 25190 9625
rect 25134 9551 25190 9560
rect 25044 9036 25096 9042
rect 25044 8978 25096 8984
rect 25044 8424 25096 8430
rect 25044 8366 25096 8372
rect 24952 7880 25004 7886
rect 24952 7822 25004 7828
rect 24964 7546 24992 7822
rect 24952 7540 25004 7546
rect 24952 7482 25004 7488
rect 24860 6724 24912 6730
rect 24860 6666 24912 6672
rect 24872 6458 24900 6666
rect 25056 6662 25084 8366
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 24860 6452 24912 6458
rect 24860 6394 24912 6400
rect 24952 6112 25004 6118
rect 24952 6054 25004 6060
rect 24964 5914 24992 6054
rect 24952 5908 25004 5914
rect 24952 5850 25004 5856
rect 25148 5778 25176 9551
rect 25240 9178 25268 10610
rect 25516 10606 25544 10775
rect 25504 10600 25556 10606
rect 25504 10542 25556 10548
rect 25412 10532 25464 10538
rect 25412 10474 25464 10480
rect 25424 10441 25452 10474
rect 25410 10432 25466 10441
rect 25410 10367 25466 10376
rect 25320 9444 25372 9450
rect 25320 9386 25372 9392
rect 25332 9178 25360 9386
rect 25228 9172 25280 9178
rect 25228 9114 25280 9120
rect 25320 9172 25372 9178
rect 25320 9114 25372 9120
rect 25412 7880 25464 7886
rect 25412 7822 25464 7828
rect 25424 7546 25452 7822
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 25516 7528 25544 10542
rect 25608 10248 25636 12406
rect 25700 12374 25728 12582
rect 25884 12442 25912 13194
rect 25872 12436 25924 12442
rect 25872 12378 25924 12384
rect 25688 12368 25740 12374
rect 25688 12310 25740 12316
rect 25780 11144 25832 11150
rect 25780 11086 25832 11092
rect 25872 11144 25924 11150
rect 25872 11086 25924 11092
rect 25688 11008 25740 11014
rect 25688 10950 25740 10956
rect 25700 10674 25728 10950
rect 25688 10668 25740 10674
rect 25688 10610 25740 10616
rect 25608 10220 25728 10248
rect 25594 10160 25650 10169
rect 25594 10095 25650 10104
rect 25608 9926 25636 10095
rect 25700 10062 25728 10220
rect 25688 10056 25740 10062
rect 25688 9998 25740 10004
rect 25596 9920 25648 9926
rect 25596 9862 25648 9868
rect 25700 9761 25728 9998
rect 25686 9752 25742 9761
rect 25686 9687 25742 9696
rect 25792 9450 25820 11086
rect 25884 10266 25912 11086
rect 25976 10849 26004 13398
rect 26068 12850 26096 15438
rect 26146 15399 26202 15408
rect 26148 15156 26200 15162
rect 26148 15098 26200 15104
rect 26160 13258 26188 15098
rect 26148 13252 26200 13258
rect 26148 13194 26200 13200
rect 26056 12844 26108 12850
rect 26056 12786 26108 12792
rect 25962 10840 26018 10849
rect 25962 10775 26018 10784
rect 25964 10668 26016 10674
rect 25964 10610 26016 10616
rect 25872 10260 25924 10266
rect 25872 10202 25924 10208
rect 25976 9994 26004 10610
rect 25964 9988 26016 9994
rect 25964 9930 26016 9936
rect 26068 9897 26096 12786
rect 26160 10674 26188 13194
rect 26252 12866 26280 19110
rect 26608 18352 26660 18358
rect 26608 18294 26660 18300
rect 26332 17536 26384 17542
rect 26332 17478 26384 17484
rect 26344 17270 26372 17478
rect 26332 17264 26384 17270
rect 26332 17206 26384 17212
rect 26332 16584 26384 16590
rect 26330 16552 26332 16561
rect 26384 16552 26386 16561
rect 26330 16487 26386 16496
rect 26424 16516 26476 16522
rect 26424 16458 26476 16464
rect 26332 16448 26384 16454
rect 26332 16390 26384 16396
rect 26344 16182 26372 16390
rect 26332 16176 26384 16182
rect 26332 16118 26384 16124
rect 26332 15972 26384 15978
rect 26332 15914 26384 15920
rect 26344 15609 26372 15914
rect 26436 15706 26464 16458
rect 26620 16046 26648 18294
rect 26608 16040 26660 16046
rect 26608 15982 26660 15988
rect 26424 15700 26476 15706
rect 26424 15642 26476 15648
rect 26330 15600 26386 15609
rect 26330 15535 26386 15544
rect 26344 15502 26372 15535
rect 26620 15502 26648 15982
rect 26712 15502 26740 19246
rect 26976 18284 27028 18290
rect 26976 18226 27028 18232
rect 26988 17338 27016 18226
rect 26976 17332 27028 17338
rect 26976 17274 27028 17280
rect 27080 16794 27108 19366
rect 27264 18086 27292 19654
rect 27160 18080 27212 18086
rect 27160 18022 27212 18028
rect 27252 18080 27304 18086
rect 27252 18022 27304 18028
rect 27172 17746 27200 18022
rect 27160 17740 27212 17746
rect 27160 17682 27212 17688
rect 27068 16788 27120 16794
rect 27068 16730 27120 16736
rect 27160 16584 27212 16590
rect 26882 16552 26938 16561
rect 26792 16516 26844 16522
rect 27160 16526 27212 16532
rect 26882 16487 26938 16496
rect 26792 16458 26844 16464
rect 26804 16250 26832 16458
rect 26792 16244 26844 16250
rect 26792 16186 26844 16192
rect 26790 15736 26846 15745
rect 26896 15706 26924 16487
rect 26790 15671 26846 15680
rect 26884 15700 26936 15706
rect 26804 15570 26832 15671
rect 26884 15642 26936 15648
rect 26896 15609 26924 15642
rect 26882 15600 26938 15609
rect 26792 15564 26844 15570
rect 26882 15535 26938 15544
rect 26792 15506 26844 15512
rect 26332 15496 26384 15502
rect 26332 15438 26384 15444
rect 26424 15496 26476 15502
rect 26424 15438 26476 15444
rect 26608 15496 26660 15502
rect 26608 15438 26660 15444
rect 26700 15496 26752 15502
rect 26700 15438 26752 15444
rect 27068 15496 27120 15502
rect 27068 15438 27120 15444
rect 26344 14006 26372 15438
rect 26436 15162 26464 15438
rect 26424 15156 26476 15162
rect 26424 15098 26476 15104
rect 26424 14952 26476 14958
rect 26424 14894 26476 14900
rect 26436 14550 26464 14894
rect 26516 14612 26568 14618
rect 26516 14554 26568 14560
rect 26424 14544 26476 14550
rect 26424 14486 26476 14492
rect 26332 14000 26384 14006
rect 26332 13942 26384 13948
rect 26424 13184 26476 13190
rect 26424 13126 26476 13132
rect 26436 13025 26464 13126
rect 26422 13016 26478 13025
rect 26422 12951 26478 12960
rect 26528 12918 26556 14554
rect 26712 14006 26740 15438
rect 26700 14000 26752 14006
rect 26700 13942 26752 13948
rect 26792 13728 26844 13734
rect 26792 13670 26844 13676
rect 26608 13252 26660 13258
rect 26608 13194 26660 13200
rect 26516 12912 26568 12918
rect 26251 12838 26280 12866
rect 26422 12880 26478 12889
rect 26251 12730 26279 12838
rect 26516 12854 26568 12860
rect 26422 12815 26478 12824
rect 26251 12714 26280 12730
rect 26240 12708 26292 12714
rect 26240 12650 26292 12656
rect 26436 12594 26464 12815
rect 26344 12566 26464 12594
rect 26344 11121 26372 12566
rect 26528 12345 26556 12854
rect 26620 12714 26648 13194
rect 26804 12850 26832 13670
rect 26974 13016 27030 13025
rect 26974 12951 26976 12960
rect 27028 12951 27030 12960
rect 26976 12922 27028 12928
rect 26792 12844 26844 12850
rect 26792 12786 26844 12792
rect 26976 12844 27028 12850
rect 26976 12786 27028 12792
rect 26608 12708 26660 12714
rect 26608 12650 26660 12656
rect 26792 12708 26844 12714
rect 26792 12650 26844 12656
rect 26884 12708 26936 12714
rect 26884 12650 26936 12656
rect 26620 12374 26648 12650
rect 26700 12436 26752 12442
rect 26700 12378 26752 12384
rect 26608 12368 26660 12374
rect 26514 12336 26570 12345
rect 26608 12310 26660 12316
rect 26514 12271 26570 12280
rect 26424 11144 26476 11150
rect 26330 11112 26386 11121
rect 26424 11086 26476 11092
rect 26516 11144 26568 11150
rect 26516 11086 26568 11092
rect 26608 11144 26660 11150
rect 26608 11086 26660 11092
rect 26330 11047 26386 11056
rect 26148 10668 26200 10674
rect 26148 10610 26200 10616
rect 26240 10192 26292 10198
rect 26240 10134 26292 10140
rect 26054 9888 26110 9897
rect 26054 9823 26110 9832
rect 26068 9602 26096 9823
rect 25884 9586 26096 9602
rect 25872 9580 26096 9586
rect 25924 9574 26096 9580
rect 26146 9616 26202 9625
rect 26252 9586 26280 10134
rect 26146 9551 26148 9560
rect 25872 9522 25924 9528
rect 26200 9551 26202 9560
rect 26240 9580 26292 9586
rect 26148 9522 26200 9528
rect 26240 9522 26292 9528
rect 25780 9444 25832 9450
rect 25780 9386 25832 9392
rect 26240 9036 26292 9042
rect 26240 8978 26292 8984
rect 25780 8968 25832 8974
rect 25780 8910 25832 8916
rect 25872 8968 25924 8974
rect 26252 8922 26280 8978
rect 25872 8910 25924 8916
rect 25792 8566 25820 8910
rect 25780 8560 25832 8566
rect 25780 8502 25832 8508
rect 25884 8412 25912 8910
rect 26068 8894 26280 8922
rect 26068 8634 26096 8894
rect 26148 8832 26200 8838
rect 26148 8774 26200 8780
rect 26160 8634 26188 8774
rect 26056 8628 26108 8634
rect 26056 8570 26108 8576
rect 26148 8628 26200 8634
rect 26148 8570 26200 8576
rect 26344 8498 26372 11047
rect 26436 11014 26464 11086
rect 26424 11008 26476 11014
rect 26424 10950 26476 10956
rect 26436 9042 26464 10950
rect 26528 9450 26556 11086
rect 26620 10810 26648 11086
rect 26608 10804 26660 10810
rect 26608 10746 26660 10752
rect 26712 9654 26740 12378
rect 26804 11762 26832 12650
rect 26896 12170 26924 12650
rect 26884 12164 26936 12170
rect 26884 12106 26936 12112
rect 26792 11756 26844 11762
rect 26792 11698 26844 11704
rect 26884 10464 26936 10470
rect 26884 10406 26936 10412
rect 26700 9648 26752 9654
rect 26700 9590 26752 9596
rect 26790 9616 26846 9625
rect 26608 9580 26660 9586
rect 26790 9551 26846 9560
rect 26608 9522 26660 9528
rect 26620 9466 26648 9522
rect 26516 9444 26568 9450
rect 26620 9438 26740 9466
rect 26516 9386 26568 9392
rect 26424 9036 26476 9042
rect 26424 8978 26476 8984
rect 25964 8492 26016 8498
rect 25964 8434 26016 8440
rect 26332 8492 26384 8498
rect 26332 8434 26384 8440
rect 25792 8384 25912 8412
rect 25792 7954 25820 8384
rect 25780 7948 25832 7954
rect 25780 7890 25832 7896
rect 25516 7500 25728 7528
rect 25226 7440 25282 7449
rect 25516 7410 25544 7500
rect 25226 7375 25282 7384
rect 25504 7404 25556 7410
rect 25240 6866 25268 7375
rect 25504 7346 25556 7352
rect 25596 7404 25648 7410
rect 25596 7346 25648 7352
rect 25410 7168 25466 7177
rect 25410 7103 25466 7112
rect 25228 6860 25280 6866
rect 25228 6802 25280 6808
rect 25424 6730 25452 7103
rect 25502 6760 25558 6769
rect 25412 6724 25464 6730
rect 25608 6730 25636 7346
rect 25700 6934 25728 7500
rect 25688 6928 25740 6934
rect 25688 6870 25740 6876
rect 25792 6882 25820 7890
rect 25872 7404 25924 7410
rect 25872 7346 25924 7352
rect 25884 7177 25912 7346
rect 25976 7274 26004 8434
rect 26148 7744 26200 7750
rect 26148 7686 26200 7692
rect 26056 7404 26108 7410
rect 26056 7346 26108 7352
rect 25964 7268 26016 7274
rect 25964 7210 26016 7216
rect 25870 7168 25926 7177
rect 25870 7103 25926 7112
rect 26068 7002 26096 7346
rect 26160 7274 26188 7686
rect 26332 7540 26384 7546
rect 26332 7482 26384 7488
rect 26148 7268 26200 7274
rect 26148 7210 26200 7216
rect 26056 6996 26108 7002
rect 26056 6938 26108 6944
rect 26160 6934 26188 7210
rect 26240 7200 26292 7206
rect 26240 7142 26292 7148
rect 26148 6928 26200 6934
rect 25700 6780 25728 6870
rect 25792 6854 25907 6882
rect 26148 6870 26200 6876
rect 25879 6848 25907 6854
rect 25879 6820 25912 6848
rect 25780 6792 25832 6798
rect 25700 6752 25780 6780
rect 25884 6780 25912 6820
rect 26252 6798 26280 7142
rect 26148 6792 26200 6798
rect 25884 6752 26004 6780
rect 25780 6734 25832 6740
rect 25502 6695 25504 6704
rect 25412 6666 25464 6672
rect 25556 6695 25558 6704
rect 25596 6724 25648 6730
rect 25504 6666 25556 6672
rect 25596 6666 25648 6672
rect 25320 6656 25372 6662
rect 25320 6598 25372 6604
rect 25332 6118 25360 6598
rect 25608 6458 25636 6666
rect 25870 6488 25926 6497
rect 25596 6452 25648 6458
rect 25870 6423 25926 6432
rect 25596 6394 25648 6400
rect 25594 6352 25650 6361
rect 25884 6322 25912 6423
rect 25976 6322 26004 6752
rect 26148 6734 26200 6740
rect 26240 6792 26292 6798
rect 26240 6734 26292 6740
rect 26160 6322 26188 6734
rect 25594 6287 25596 6296
rect 25648 6287 25650 6296
rect 25872 6316 25924 6322
rect 25596 6258 25648 6264
rect 25872 6258 25924 6264
rect 25964 6316 26016 6322
rect 25964 6258 26016 6264
rect 26148 6316 26200 6322
rect 26148 6258 26200 6264
rect 26344 6186 26372 7482
rect 26516 7404 26568 7410
rect 26516 7346 26568 7352
rect 26608 7404 26660 7410
rect 26608 7346 26660 7352
rect 26528 7041 26556 7346
rect 26514 7032 26570 7041
rect 26514 6967 26570 6976
rect 26528 6798 26556 6967
rect 26424 6792 26476 6798
rect 26424 6734 26476 6740
rect 26516 6792 26568 6798
rect 26516 6734 26568 6740
rect 26436 6458 26464 6734
rect 26620 6730 26648 7346
rect 26608 6724 26660 6730
rect 26608 6666 26660 6672
rect 26424 6452 26476 6458
rect 26424 6394 26476 6400
rect 26332 6180 26384 6186
rect 26332 6122 26384 6128
rect 25320 6112 25372 6118
rect 25320 6054 25372 6060
rect 26436 5846 26464 6394
rect 26424 5840 26476 5846
rect 26424 5782 26476 5788
rect 25136 5772 25188 5778
rect 25136 5714 25188 5720
rect 26516 5160 26568 5166
rect 26516 5102 26568 5108
rect 24768 5092 24820 5098
rect 24768 5034 24820 5040
rect 26528 4690 26556 5102
rect 26516 4684 26568 4690
rect 26516 4626 26568 4632
rect 25780 4616 25832 4622
rect 25780 4558 25832 4564
rect 25792 4282 25820 4558
rect 25780 4276 25832 4282
rect 25780 4218 25832 4224
rect 25320 4208 25372 4214
rect 25320 4150 25372 4156
rect 24768 4140 24820 4146
rect 24768 4082 24820 4088
rect 24780 3602 24808 4082
rect 25226 3904 25282 3913
rect 25226 3839 25282 3848
rect 25240 3602 25268 3839
rect 25332 3602 25360 4150
rect 24768 3596 24820 3602
rect 24768 3538 24820 3544
rect 25228 3596 25280 3602
rect 25228 3538 25280 3544
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 24582 3431 24638 3440
rect 24676 3460 24728 3466
rect 24676 3402 24728 3408
rect 24032 3392 24084 3398
rect 24032 3334 24084 3340
rect 24860 3392 24912 3398
rect 24860 3334 24912 3340
rect 25228 3392 25280 3398
rect 25688 3392 25740 3398
rect 25280 3352 25360 3380
rect 25228 3334 25280 3340
rect 24044 3194 24072 3334
rect 24872 3194 24900 3334
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 24032 3188 24084 3194
rect 24032 3130 24084 3136
rect 24860 3188 24912 3194
rect 24860 3130 24912 3136
rect 23388 3120 23440 3126
rect 23388 3062 23440 3068
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 18696 2916 18748 2922
rect 18696 2858 18748 2864
rect 16304 2848 16356 2854
rect 16304 2790 16356 2796
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 19720 2514 19748 2790
rect 19812 2650 19840 2790
rect 24674 2680 24730 2689
rect 19800 2644 19852 2650
rect 25148 2650 25176 2926
rect 25332 2774 25360 3352
rect 25688 3334 25740 3340
rect 25700 3058 25728 3334
rect 25688 3052 25740 3058
rect 25688 2994 25740 3000
rect 25792 2990 25820 4218
rect 26332 3664 26384 3670
rect 26332 3606 26384 3612
rect 25780 2984 25832 2990
rect 25780 2926 25832 2932
rect 26344 2922 26372 3606
rect 26516 3392 26568 3398
rect 26620 3380 26648 6666
rect 26712 6254 26740 9438
rect 26804 8566 26832 9551
rect 26792 8560 26844 8566
rect 26792 8502 26844 8508
rect 26792 6656 26844 6662
rect 26792 6598 26844 6604
rect 26700 6248 26752 6254
rect 26700 6190 26752 6196
rect 26804 6186 26832 6598
rect 26896 6390 26924 10406
rect 26988 9586 27016 12786
rect 27080 12170 27108 15438
rect 27172 13190 27200 16526
rect 27252 15904 27304 15910
rect 27252 15846 27304 15852
rect 27264 15366 27292 15846
rect 27252 15360 27304 15366
rect 27252 15302 27304 15308
rect 27264 13734 27292 15302
rect 27252 13728 27304 13734
rect 27252 13670 27304 13676
rect 27356 13530 27384 19790
rect 27816 19446 27844 19790
rect 27804 19440 27856 19446
rect 27804 19382 27856 19388
rect 28644 19378 28672 19790
rect 27436 19372 27488 19378
rect 27436 19314 27488 19320
rect 28632 19372 28684 19378
rect 28632 19314 28684 19320
rect 27448 18630 27476 19314
rect 27436 18624 27488 18630
rect 27436 18566 27488 18572
rect 27448 17542 27476 18566
rect 28644 18154 28672 19314
rect 28816 18760 28868 18766
rect 28816 18702 28868 18708
rect 28724 18624 28776 18630
rect 28724 18566 28776 18572
rect 28736 18329 28764 18566
rect 28722 18320 28778 18329
rect 28722 18255 28778 18264
rect 28632 18148 28684 18154
rect 28632 18090 28684 18096
rect 27526 17640 27582 17649
rect 27582 17584 27660 17592
rect 27526 17575 27528 17584
rect 27580 17564 27660 17584
rect 27528 17546 27580 17552
rect 27436 17536 27488 17542
rect 27436 17478 27488 17484
rect 27448 16250 27476 17478
rect 27528 17128 27580 17134
rect 27528 17070 27580 17076
rect 27540 16697 27568 17070
rect 27526 16688 27582 16697
rect 27632 16658 27660 17564
rect 28540 17536 28592 17542
rect 28540 17478 28592 17484
rect 28552 17338 28580 17478
rect 28172 17332 28224 17338
rect 28172 17274 28224 17280
rect 28540 17332 28592 17338
rect 28540 17274 28592 17280
rect 27988 17196 28040 17202
rect 27988 17138 28040 17144
rect 27526 16623 27582 16632
rect 27620 16652 27672 16658
rect 27620 16594 27672 16600
rect 27896 16448 27948 16454
rect 27896 16390 27948 16396
rect 27436 16244 27488 16250
rect 27436 16186 27488 16192
rect 27344 13524 27396 13530
rect 27344 13466 27396 13472
rect 27344 13388 27396 13394
rect 27344 13330 27396 13336
rect 27160 13184 27212 13190
rect 27160 13126 27212 13132
rect 27068 12164 27120 12170
rect 27068 12106 27120 12112
rect 27080 11898 27108 12106
rect 27068 11892 27120 11898
rect 27068 11834 27120 11840
rect 27080 11626 27108 11834
rect 27068 11620 27120 11626
rect 27068 11562 27120 11568
rect 27066 10976 27122 10985
rect 27066 10911 27122 10920
rect 26976 9580 27028 9586
rect 26976 9522 27028 9528
rect 27080 6644 27108 10911
rect 27172 9586 27200 13126
rect 27252 12844 27304 12850
rect 27252 12786 27304 12792
rect 27264 12442 27292 12786
rect 27356 12714 27384 13330
rect 27344 12708 27396 12714
rect 27344 12650 27396 12656
rect 27252 12436 27304 12442
rect 27252 12378 27304 12384
rect 27344 12232 27396 12238
rect 27344 12174 27396 12180
rect 27356 11694 27384 12174
rect 27344 11688 27396 11694
rect 27344 11630 27396 11636
rect 27356 10305 27384 11630
rect 27342 10296 27398 10305
rect 27342 10231 27398 10240
rect 27252 10192 27304 10198
rect 27252 10134 27304 10140
rect 27160 9580 27212 9586
rect 27160 9522 27212 9528
rect 27264 9450 27292 10134
rect 27448 10010 27476 16186
rect 27908 15502 27936 16390
rect 28000 16046 28028 17138
rect 28078 16144 28134 16153
rect 28078 16079 28134 16088
rect 28092 16046 28120 16079
rect 27988 16040 28040 16046
rect 27988 15982 28040 15988
rect 28080 16040 28132 16046
rect 28080 15982 28132 15988
rect 28184 15502 28212 17274
rect 28540 16176 28592 16182
rect 28540 16118 28592 16124
rect 28356 15972 28408 15978
rect 28356 15914 28408 15920
rect 28264 15904 28316 15910
rect 28264 15846 28316 15852
rect 28276 15638 28304 15846
rect 28368 15706 28396 15914
rect 28552 15706 28580 16118
rect 28644 16114 28672 18090
rect 28736 16697 28764 18255
rect 28828 17678 28856 18702
rect 28908 18624 28960 18630
rect 28908 18566 28960 18572
rect 29276 18624 29328 18630
rect 29276 18566 29328 18572
rect 28920 18426 28948 18566
rect 28908 18420 28960 18426
rect 28908 18362 28960 18368
rect 29000 18216 29052 18222
rect 29000 18158 29052 18164
rect 29012 17882 29040 18158
rect 29288 17882 29316 18566
rect 29000 17876 29052 17882
rect 29000 17818 29052 17824
rect 29276 17876 29328 17882
rect 29276 17818 29328 17824
rect 28816 17672 28868 17678
rect 28816 17614 28868 17620
rect 28722 16688 28778 16697
rect 28722 16623 28778 16632
rect 29184 16516 29236 16522
rect 29184 16458 29236 16464
rect 28632 16108 28684 16114
rect 28632 16050 28684 16056
rect 29092 16108 29144 16114
rect 29092 16050 29144 16056
rect 28632 15904 28684 15910
rect 28632 15846 28684 15852
rect 28356 15700 28408 15706
rect 28356 15642 28408 15648
rect 28540 15700 28592 15706
rect 28540 15642 28592 15648
rect 28264 15632 28316 15638
rect 28264 15574 28316 15580
rect 27896 15496 27948 15502
rect 27896 15438 27948 15444
rect 28172 15496 28224 15502
rect 28172 15438 28224 15444
rect 28264 15496 28316 15502
rect 28264 15438 28316 15444
rect 28080 15428 28132 15434
rect 28080 15370 28132 15376
rect 27528 15360 27580 15366
rect 27580 15320 27660 15348
rect 27528 15302 27580 15308
rect 27528 14476 27580 14482
rect 27528 14418 27580 14424
rect 27540 11354 27568 14418
rect 27632 11694 27660 15320
rect 28092 15144 28120 15370
rect 27908 15116 28120 15144
rect 27908 14929 27936 15116
rect 28276 15042 28304 15438
rect 28000 15014 28304 15042
rect 28368 15026 28396 15642
rect 28448 15428 28500 15434
rect 28448 15370 28500 15376
rect 28356 15020 28408 15026
rect 27894 14920 27950 14929
rect 27894 14855 27950 14864
rect 27712 14408 27764 14414
rect 27712 14350 27764 14356
rect 27620 11688 27672 11694
rect 27620 11630 27672 11636
rect 27724 11558 27752 14350
rect 28000 14346 28028 15014
rect 28356 14962 28408 14968
rect 28172 14952 28224 14958
rect 28172 14894 28224 14900
rect 27988 14340 28040 14346
rect 27988 14282 28040 14288
rect 27988 14000 28040 14006
rect 27988 13942 28040 13948
rect 27804 13728 27856 13734
rect 27804 13670 27856 13676
rect 27816 13326 27844 13670
rect 27804 13320 27856 13326
rect 27804 13262 27856 13268
rect 27896 13320 27948 13326
rect 27896 13262 27948 13268
rect 27908 12986 27936 13262
rect 27896 12980 27948 12986
rect 27896 12922 27948 12928
rect 27804 12844 27856 12850
rect 27804 12786 27856 12792
rect 27712 11552 27764 11558
rect 27712 11494 27764 11500
rect 27816 11370 27844 12786
rect 27896 12640 27948 12646
rect 27896 12582 27948 12588
rect 27908 12170 27936 12582
rect 28000 12374 28028 13942
rect 27988 12368 28040 12374
rect 27988 12310 28040 12316
rect 28184 12209 28212 14894
rect 28264 14408 28316 14414
rect 28264 14350 28316 14356
rect 28276 13977 28304 14350
rect 28262 13968 28318 13977
rect 28262 13903 28318 13912
rect 28264 13864 28316 13870
rect 28264 13806 28316 13812
rect 28170 12200 28226 12209
rect 27896 12164 27948 12170
rect 28170 12135 28226 12144
rect 27896 12106 27948 12112
rect 27528 11348 27580 11354
rect 27528 11290 27580 11296
rect 27632 11342 27844 11370
rect 27632 11286 27660 11342
rect 27620 11280 27672 11286
rect 27620 11222 27672 11228
rect 27632 10130 27660 11222
rect 27804 11144 27856 11150
rect 27804 11086 27856 11092
rect 27816 10810 27844 11086
rect 27804 10804 27856 10810
rect 27804 10746 27856 10752
rect 27712 10668 27764 10674
rect 27908 10656 27936 12106
rect 27988 11756 28040 11762
rect 27988 11698 28040 11704
rect 27764 10628 27936 10656
rect 27712 10610 27764 10616
rect 27620 10124 27672 10130
rect 27620 10066 27672 10072
rect 27448 9982 27660 10010
rect 27632 9926 27660 9982
rect 27620 9920 27672 9926
rect 27620 9862 27672 9868
rect 27252 9444 27304 9450
rect 27252 9386 27304 9392
rect 27436 8968 27488 8974
rect 27436 8910 27488 8916
rect 27448 8498 27476 8910
rect 27436 8492 27488 8498
rect 27436 8434 27488 8440
rect 27252 8016 27304 8022
rect 27252 7958 27304 7964
rect 27264 6798 27292 7958
rect 27252 6792 27304 6798
rect 27252 6734 27304 6740
rect 27160 6656 27212 6662
rect 27080 6616 27160 6644
rect 27160 6598 27212 6604
rect 27172 6390 27200 6598
rect 26884 6384 26936 6390
rect 26884 6326 26936 6332
rect 27160 6384 27212 6390
rect 27160 6326 27212 6332
rect 27264 6322 27292 6734
rect 27252 6316 27304 6322
rect 27252 6258 27304 6264
rect 26792 6180 26844 6186
rect 26792 6122 26844 6128
rect 27068 6180 27120 6186
rect 27068 6122 27120 6128
rect 26976 5228 27028 5234
rect 26976 5170 27028 5176
rect 26790 4992 26846 5001
rect 26790 4927 26846 4936
rect 26804 4486 26832 4927
rect 26792 4480 26844 4486
rect 26792 4422 26844 4428
rect 26804 4282 26832 4422
rect 26988 4282 27016 5170
rect 27080 4622 27108 6122
rect 27344 5364 27396 5370
rect 27344 5306 27396 5312
rect 27252 5228 27304 5234
rect 27252 5170 27304 5176
rect 27160 5024 27212 5030
rect 27160 4966 27212 4972
rect 27068 4616 27120 4622
rect 27068 4558 27120 4564
rect 27080 4282 27108 4558
rect 27172 4486 27200 4966
rect 27264 4826 27292 5170
rect 27356 4826 27384 5306
rect 27252 4820 27304 4826
rect 27252 4762 27304 4768
rect 27344 4820 27396 4826
rect 27344 4762 27396 4768
rect 27448 4706 27476 8434
rect 27632 5166 27660 9862
rect 27724 9081 27752 10610
rect 27896 10464 27948 10470
rect 27896 10406 27948 10412
rect 27908 10169 27936 10406
rect 27894 10160 27950 10169
rect 27804 10124 27856 10130
rect 27894 10095 27950 10104
rect 27804 10066 27856 10072
rect 27710 9072 27766 9081
rect 27710 9007 27766 9016
rect 27724 8498 27752 9007
rect 27712 8492 27764 8498
rect 27712 8434 27764 8440
rect 27710 7984 27766 7993
rect 27710 7919 27766 7928
rect 27620 5160 27672 5166
rect 27620 5102 27672 5108
rect 27528 5024 27580 5030
rect 27528 4966 27580 4972
rect 27356 4678 27476 4706
rect 27160 4480 27212 4486
rect 27160 4422 27212 4428
rect 26792 4276 26844 4282
rect 26792 4218 26844 4224
rect 26976 4276 27028 4282
rect 26976 4218 27028 4224
rect 27068 4276 27120 4282
rect 27068 4218 27120 4224
rect 26804 3602 26832 4218
rect 26792 3596 26844 3602
rect 26792 3538 26844 3544
rect 26568 3352 26648 3380
rect 26700 3392 26752 3398
rect 26516 3334 26568 3340
rect 26700 3334 26752 3340
rect 27160 3392 27212 3398
rect 27160 3334 27212 3340
rect 26528 2922 26556 3334
rect 26712 3058 26740 3334
rect 27172 3126 27200 3334
rect 27356 3194 27384 4678
rect 27436 4616 27488 4622
rect 27540 4570 27568 4966
rect 27488 4564 27568 4570
rect 27436 4558 27568 4564
rect 27448 4542 27568 4558
rect 27632 4554 27660 5102
rect 27620 4548 27672 4554
rect 27620 4490 27672 4496
rect 27724 3534 27752 7919
rect 27816 7886 27844 10066
rect 28000 10062 28028 11698
rect 28276 11150 28304 13806
rect 28356 13796 28408 13802
rect 28356 13738 28408 13744
rect 28368 11354 28396 13738
rect 28460 13326 28488 15370
rect 28540 15156 28592 15162
rect 28644 15144 28672 15846
rect 29104 15706 29132 16050
rect 29092 15700 29144 15706
rect 29092 15642 29144 15648
rect 28724 15496 28776 15502
rect 28724 15438 28776 15444
rect 28816 15496 28868 15502
rect 28816 15438 28868 15444
rect 28908 15496 28960 15502
rect 28908 15438 28960 15444
rect 28736 15162 28764 15438
rect 28592 15116 28672 15144
rect 28540 15098 28592 15104
rect 28540 15020 28592 15026
rect 28540 14962 28592 14968
rect 28448 13320 28500 13326
rect 28448 13262 28500 13268
rect 28460 12288 28488 13262
rect 28552 12918 28580 14962
rect 28644 14056 28672 15116
rect 28724 15156 28776 15162
rect 28724 15098 28776 15104
rect 28828 15026 28856 15438
rect 28816 15020 28868 15026
rect 28816 14962 28868 14968
rect 28828 14618 28856 14962
rect 28920 14890 28948 15438
rect 29092 15428 29144 15434
rect 29092 15370 29144 15376
rect 28908 14884 28960 14890
rect 28908 14826 28960 14832
rect 28816 14612 28868 14618
rect 28816 14554 28868 14560
rect 29104 14278 29132 15370
rect 29092 14272 29144 14278
rect 29092 14214 29144 14220
rect 28644 14028 28948 14056
rect 28816 13932 28868 13938
rect 28816 13874 28868 13880
rect 28828 13530 28856 13874
rect 28816 13524 28868 13530
rect 28816 13466 28868 13472
rect 28724 13252 28776 13258
rect 28724 13194 28776 13200
rect 28736 12986 28764 13194
rect 28724 12980 28776 12986
rect 28724 12922 28776 12928
rect 28540 12912 28592 12918
rect 28540 12854 28592 12860
rect 28552 12646 28580 12854
rect 28540 12640 28592 12646
rect 28540 12582 28592 12588
rect 28460 12260 28764 12288
rect 28630 12200 28686 12209
rect 28630 12135 28686 12144
rect 28448 11892 28500 11898
rect 28448 11834 28500 11840
rect 28460 11354 28488 11834
rect 28540 11688 28592 11694
rect 28540 11630 28592 11636
rect 28552 11354 28580 11630
rect 28356 11348 28408 11354
rect 28356 11290 28408 11296
rect 28448 11348 28500 11354
rect 28448 11290 28500 11296
rect 28540 11348 28592 11354
rect 28540 11290 28592 11296
rect 28264 11144 28316 11150
rect 28264 11086 28316 11092
rect 28172 11008 28224 11014
rect 28172 10950 28224 10956
rect 28184 10742 28212 10950
rect 28172 10736 28224 10742
rect 28172 10678 28224 10684
rect 28080 10600 28132 10606
rect 28080 10542 28132 10548
rect 28092 10266 28120 10542
rect 28172 10464 28224 10470
rect 28172 10406 28224 10412
rect 28080 10260 28132 10266
rect 28080 10202 28132 10208
rect 28184 10198 28212 10406
rect 28172 10192 28224 10198
rect 28172 10134 28224 10140
rect 27988 10056 28040 10062
rect 27988 9998 28040 10004
rect 28172 9988 28224 9994
rect 28172 9930 28224 9936
rect 28184 9722 28212 9930
rect 28172 9716 28224 9722
rect 28172 9658 28224 9664
rect 28080 9648 28132 9654
rect 28080 9590 28132 9596
rect 27896 8900 27948 8906
rect 27896 8842 27948 8848
rect 27908 8566 27936 8842
rect 27896 8560 27948 8566
rect 27896 8502 27948 8508
rect 27988 8492 28040 8498
rect 27988 8434 28040 8440
rect 28000 8090 28028 8434
rect 27988 8084 28040 8090
rect 27988 8026 28040 8032
rect 27804 7880 27856 7886
rect 27804 7822 27856 7828
rect 27804 7744 27856 7750
rect 27804 7686 27856 7692
rect 27896 7744 27948 7750
rect 27896 7686 27948 7692
rect 27816 6304 27844 7686
rect 27908 7206 27936 7686
rect 27896 7200 27948 7206
rect 27896 7142 27948 7148
rect 27908 6458 27936 7142
rect 28092 6882 28120 9590
rect 28276 9330 28304 11086
rect 28356 10668 28408 10674
rect 28356 10610 28408 10616
rect 28368 9518 28396 10610
rect 28540 10600 28592 10606
rect 28460 10560 28540 10588
rect 28460 10130 28488 10560
rect 28644 10588 28672 12135
rect 28736 10674 28764 12260
rect 28828 10849 28856 13466
rect 28920 13326 28948 14028
rect 28908 13320 28960 13326
rect 28908 13262 28960 13268
rect 28920 12986 28948 13262
rect 29000 13252 29052 13258
rect 29000 13194 29052 13200
rect 28908 12980 28960 12986
rect 28908 12922 28960 12928
rect 28920 12434 28948 12922
rect 29012 12918 29040 13194
rect 29000 12912 29052 12918
rect 29000 12854 29052 12860
rect 28998 12744 29054 12753
rect 28998 12679 29000 12688
rect 29052 12679 29054 12688
rect 29000 12650 29052 12656
rect 28920 12406 29040 12434
rect 28814 10840 28870 10849
rect 28814 10775 28870 10784
rect 28816 10736 28868 10742
rect 28816 10678 28868 10684
rect 28724 10668 28776 10674
rect 28724 10610 28776 10616
rect 28592 10560 28672 10588
rect 28540 10542 28592 10548
rect 28632 10464 28684 10470
rect 28632 10406 28684 10412
rect 28538 10296 28594 10305
rect 28538 10231 28540 10240
rect 28592 10231 28594 10240
rect 28540 10202 28592 10208
rect 28448 10124 28500 10130
rect 28448 10066 28500 10072
rect 28446 10024 28502 10033
rect 28446 9959 28502 9968
rect 28460 9722 28488 9959
rect 28448 9716 28500 9722
rect 28448 9658 28500 9664
rect 28356 9512 28408 9518
rect 28356 9454 28408 9460
rect 28184 9302 28304 9330
rect 28184 8974 28212 9302
rect 28264 9172 28316 9178
rect 28264 9114 28316 9120
rect 28172 8968 28224 8974
rect 28172 8910 28224 8916
rect 28276 8498 28304 9114
rect 28172 8492 28224 8498
rect 28172 8434 28224 8440
rect 28264 8492 28316 8498
rect 28264 8434 28316 8440
rect 28000 6854 28120 6882
rect 28000 6662 28028 6854
rect 28184 6798 28212 8434
rect 28356 8356 28408 8362
rect 28356 8298 28408 8304
rect 28368 6934 28396 8298
rect 28552 7002 28580 10202
rect 28644 10169 28672 10406
rect 28630 10160 28686 10169
rect 28630 10095 28686 10104
rect 28736 9110 28764 10610
rect 28828 10062 28856 10678
rect 29012 10674 29040 12406
rect 29000 10668 29052 10674
rect 29000 10610 29052 10616
rect 28906 10568 28962 10577
rect 28906 10503 28962 10512
rect 28816 10056 28868 10062
rect 28816 9998 28868 10004
rect 28816 9920 28868 9926
rect 28816 9862 28868 9868
rect 28828 9722 28856 9862
rect 28816 9716 28868 9722
rect 28816 9658 28868 9664
rect 28816 9172 28868 9178
rect 28816 9114 28868 9120
rect 28724 9104 28776 9110
rect 28724 9046 28776 9052
rect 28736 8566 28764 9046
rect 28724 8560 28776 8566
rect 28724 8502 28776 8508
rect 28632 8492 28684 8498
rect 28632 8434 28684 8440
rect 28644 7274 28672 8434
rect 28828 8090 28856 9114
rect 28920 9042 28948 10503
rect 29012 10130 29040 10610
rect 29000 10124 29052 10130
rect 29000 10066 29052 10072
rect 28998 9616 29054 9625
rect 28998 9551 29054 9560
rect 29012 9178 29040 9551
rect 29000 9172 29052 9178
rect 29000 9114 29052 9120
rect 28908 9036 28960 9042
rect 28908 8978 28960 8984
rect 28908 8560 28960 8566
rect 28908 8502 28960 8508
rect 28816 8084 28868 8090
rect 28816 8026 28868 8032
rect 28920 7954 28948 8502
rect 28908 7948 28960 7954
rect 28908 7890 28960 7896
rect 28724 7540 28776 7546
rect 28724 7482 28776 7488
rect 28632 7268 28684 7274
rect 28632 7210 28684 7216
rect 28540 6996 28592 7002
rect 28540 6938 28592 6944
rect 28736 6934 28764 7482
rect 29000 7472 29052 7478
rect 29104 7460 29132 14214
rect 29196 14074 29224 16458
rect 29276 15904 29328 15910
rect 29276 15846 29328 15852
rect 29288 15706 29316 15846
rect 29276 15700 29328 15706
rect 29276 15642 29328 15648
rect 29276 14544 29328 14550
rect 29276 14486 29328 14492
rect 29184 14068 29236 14074
rect 29184 14010 29236 14016
rect 29196 13938 29224 14010
rect 29288 13938 29316 14486
rect 29380 14414 29408 26250
rect 29564 25945 29592 26250
rect 29550 25936 29606 25945
rect 29550 25871 29606 25880
rect 29564 25838 29592 25871
rect 29552 25832 29604 25838
rect 29552 25774 29604 25780
rect 29920 24608 29972 24614
rect 29920 24550 29972 24556
rect 29736 24336 29788 24342
rect 29736 24278 29788 24284
rect 29644 24132 29696 24138
rect 29644 24074 29696 24080
rect 29460 23792 29512 23798
rect 29460 23734 29512 23740
rect 29472 22094 29500 23734
rect 29656 23662 29684 24074
rect 29644 23656 29696 23662
rect 29644 23598 29696 23604
rect 29644 23044 29696 23050
rect 29644 22986 29696 22992
rect 29472 22066 29592 22094
rect 29564 20482 29592 22066
rect 29656 21690 29684 22986
rect 29748 22982 29776 24278
rect 29828 24064 29880 24070
rect 29828 24006 29880 24012
rect 29736 22976 29788 22982
rect 29736 22918 29788 22924
rect 29748 22642 29776 22918
rect 29840 22710 29868 24006
rect 29932 23594 29960 24550
rect 30116 24206 30144 27084
rect 30392 27010 30420 27406
rect 30196 26988 30248 26994
rect 30196 26930 30248 26936
rect 30300 26982 30420 27010
rect 30472 26988 30524 26994
rect 30208 26042 30236 26930
rect 30300 26926 30328 26982
rect 30472 26930 30524 26936
rect 30288 26920 30340 26926
rect 30288 26862 30340 26868
rect 30300 26586 30328 26862
rect 30380 26784 30432 26790
rect 30380 26726 30432 26732
rect 30288 26580 30340 26586
rect 30288 26522 30340 26528
rect 30196 26036 30248 26042
rect 30196 25978 30248 25984
rect 30288 25968 30340 25974
rect 30288 25910 30340 25916
rect 30300 25498 30328 25910
rect 30392 25906 30420 26726
rect 30380 25900 30432 25906
rect 30380 25842 30432 25848
rect 30288 25492 30340 25498
rect 30288 25434 30340 25440
rect 30300 24954 30328 25434
rect 30484 25378 30512 26930
rect 30564 26784 30616 26790
rect 30564 26726 30616 26732
rect 30576 25838 30604 26726
rect 30564 25832 30616 25838
rect 30564 25774 30616 25780
rect 30392 25350 30512 25378
rect 30392 25226 30420 25350
rect 30472 25288 30524 25294
rect 30472 25230 30524 25236
rect 30380 25220 30432 25226
rect 30380 25162 30432 25168
rect 30288 24948 30340 24954
rect 30288 24890 30340 24896
rect 30484 24206 30512 25230
rect 30576 24886 30604 25774
rect 30564 24880 30616 24886
rect 30564 24822 30616 24828
rect 30104 24200 30156 24206
rect 30472 24200 30524 24206
rect 30156 24160 30236 24188
rect 30104 24142 30156 24148
rect 30012 23656 30064 23662
rect 30012 23598 30064 23604
rect 29920 23588 29972 23594
rect 29920 23530 29972 23536
rect 29828 22704 29880 22710
rect 29828 22646 29880 22652
rect 29736 22636 29788 22642
rect 29736 22578 29788 22584
rect 29932 22556 29960 23530
rect 30024 22710 30052 23598
rect 30104 23112 30156 23118
rect 30104 23054 30156 23060
rect 30012 22704 30064 22710
rect 30012 22646 30064 22652
rect 29932 22528 30052 22556
rect 29736 22432 29788 22438
rect 29736 22374 29788 22380
rect 29748 22166 29776 22374
rect 29736 22160 29788 22166
rect 29736 22102 29788 22108
rect 29920 22024 29972 22030
rect 29920 21966 29972 21972
rect 29828 21956 29880 21962
rect 29828 21898 29880 21904
rect 29644 21684 29696 21690
rect 29644 21626 29696 21632
rect 29644 21548 29696 21554
rect 29644 21490 29696 21496
rect 29656 20942 29684 21490
rect 29840 21010 29868 21898
rect 29932 21690 29960 21966
rect 29920 21684 29972 21690
rect 29920 21626 29972 21632
rect 29828 21004 29880 21010
rect 29828 20946 29880 20952
rect 29644 20936 29696 20942
rect 29644 20878 29696 20884
rect 30024 20618 30052 22528
rect 30116 22166 30144 23054
rect 30208 22710 30236 24160
rect 30472 24142 30524 24148
rect 30484 23594 30512 24142
rect 30564 24132 30616 24138
rect 30564 24074 30616 24080
rect 30668 24120 30696 28494
rect 30760 28218 30788 28494
rect 30932 28416 30984 28422
rect 30932 28358 30984 28364
rect 30748 28212 30800 28218
rect 30748 28154 30800 28160
rect 30760 26858 30788 28154
rect 30944 27334 30972 28358
rect 30932 27328 30984 27334
rect 30932 27270 30984 27276
rect 30944 26994 30972 27270
rect 30932 26988 30984 26994
rect 30932 26930 30984 26936
rect 30748 26852 30800 26858
rect 30748 26794 30800 26800
rect 30840 25900 30892 25906
rect 30840 25842 30892 25848
rect 30852 25294 30880 25842
rect 30748 25288 30800 25294
rect 30748 25230 30800 25236
rect 30840 25288 30892 25294
rect 30840 25230 30892 25236
rect 30760 24682 30788 25230
rect 30748 24676 30800 24682
rect 30748 24618 30800 24624
rect 30840 24200 30892 24206
rect 30840 24142 30892 24148
rect 30748 24132 30800 24138
rect 30668 24092 30748 24120
rect 30472 23588 30524 23594
rect 30472 23530 30524 23536
rect 30484 23186 30512 23530
rect 30472 23180 30524 23186
rect 30472 23122 30524 23128
rect 30288 23112 30340 23118
rect 30288 23054 30340 23060
rect 30300 22778 30328 23054
rect 30472 22976 30524 22982
rect 30472 22918 30524 22924
rect 30484 22778 30512 22918
rect 30288 22772 30340 22778
rect 30288 22714 30340 22720
rect 30472 22772 30524 22778
rect 30472 22714 30524 22720
rect 30196 22704 30248 22710
rect 30196 22646 30248 22652
rect 30576 22506 30604 24074
rect 30668 22658 30696 24092
rect 30748 24074 30800 24080
rect 30852 23730 30880 24142
rect 30840 23724 30892 23730
rect 30840 23666 30892 23672
rect 30748 23248 30800 23254
rect 30748 23190 30800 23196
rect 30760 22778 30788 23190
rect 30748 22772 30800 22778
rect 30748 22714 30800 22720
rect 30668 22630 30788 22658
rect 30564 22500 30616 22506
rect 30564 22442 30616 22448
rect 30656 22500 30708 22506
rect 30656 22442 30708 22448
rect 30104 22160 30156 22166
rect 30104 22102 30156 22108
rect 30104 21888 30156 21894
rect 30104 21830 30156 21836
rect 30116 21418 30144 21830
rect 30104 21412 30156 21418
rect 30104 21354 30156 21360
rect 30668 21146 30696 22442
rect 30656 21140 30708 21146
rect 30656 21082 30708 21088
rect 30288 21072 30340 21078
rect 30288 21014 30340 21020
rect 30196 21004 30248 21010
rect 30196 20946 30248 20952
rect 30024 20602 30144 20618
rect 30208 20602 30236 20946
rect 30012 20596 30144 20602
rect 30064 20590 30144 20596
rect 30012 20538 30064 20544
rect 29564 20466 29684 20482
rect 30116 20466 30144 20590
rect 30196 20596 30248 20602
rect 30196 20538 30248 20544
rect 29460 20460 29512 20466
rect 29564 20460 29696 20466
rect 29564 20454 29644 20460
rect 29460 20402 29512 20408
rect 29644 20402 29696 20408
rect 30012 20460 30064 20466
rect 30012 20402 30064 20408
rect 30104 20460 30156 20466
rect 30104 20402 30156 20408
rect 29472 19854 29500 20402
rect 29460 19848 29512 19854
rect 29460 19790 29512 19796
rect 29368 14408 29420 14414
rect 29368 14350 29420 14356
rect 29184 13932 29236 13938
rect 29184 13874 29236 13880
rect 29276 13932 29328 13938
rect 29276 13874 29328 13880
rect 29196 10810 29224 13874
rect 29288 12306 29316 13874
rect 29368 13320 29420 13326
rect 29368 13262 29420 13268
rect 29380 12850 29408 13262
rect 29368 12844 29420 12850
rect 29368 12786 29420 12792
rect 29276 12300 29328 12306
rect 29276 12242 29328 12248
rect 29366 11928 29422 11937
rect 29366 11863 29422 11872
rect 29380 11830 29408 11863
rect 29368 11824 29420 11830
rect 29368 11766 29420 11772
rect 29184 10804 29236 10810
rect 29184 10746 29236 10752
rect 29184 10056 29236 10062
rect 29184 9998 29236 10004
rect 29052 7432 29132 7460
rect 29000 7414 29052 7420
rect 29092 7268 29144 7274
rect 29092 7210 29144 7216
rect 28356 6928 28408 6934
rect 28356 6870 28408 6876
rect 28724 6928 28776 6934
rect 28724 6870 28776 6876
rect 28080 6792 28132 6798
rect 28080 6734 28132 6740
rect 28172 6792 28224 6798
rect 28172 6734 28224 6740
rect 28724 6792 28776 6798
rect 28724 6734 28776 6740
rect 28092 6662 28120 6734
rect 27988 6656 28040 6662
rect 27988 6598 28040 6604
rect 28080 6656 28132 6662
rect 28080 6598 28132 6604
rect 27896 6452 27948 6458
rect 27896 6394 27948 6400
rect 27896 6316 27948 6322
rect 27816 6276 27896 6304
rect 27896 6258 27948 6264
rect 28092 6254 28120 6598
rect 28736 6458 28764 6734
rect 28724 6452 28776 6458
rect 28724 6394 28776 6400
rect 28080 6248 28132 6254
rect 28080 6190 28132 6196
rect 28080 5364 28132 5370
rect 28080 5306 28132 5312
rect 27896 5228 27948 5234
rect 27896 5170 27948 5176
rect 27908 5098 27936 5170
rect 27896 5092 27948 5098
rect 27896 5034 27948 5040
rect 27804 5024 27856 5030
rect 27804 4966 27856 4972
rect 27816 4078 27844 4966
rect 28092 4078 28120 5306
rect 28264 5228 28316 5234
rect 28264 5170 28316 5176
rect 27804 4072 27856 4078
rect 27804 4014 27856 4020
rect 28080 4072 28132 4078
rect 28080 4014 28132 4020
rect 28276 3534 28304 5170
rect 29104 4758 29132 7210
rect 29196 6798 29224 9998
rect 29380 9654 29408 11766
rect 29472 11354 29500 19790
rect 29552 16788 29604 16794
rect 29552 16730 29604 16736
rect 29564 15978 29592 16730
rect 29552 15972 29604 15978
rect 29552 15914 29604 15920
rect 29656 14482 29684 20402
rect 30024 19786 30052 20402
rect 30208 19922 30236 20538
rect 30300 20466 30328 21014
rect 30564 20868 30616 20874
rect 30564 20810 30616 20816
rect 30380 20800 30432 20806
rect 30380 20742 30432 20748
rect 30288 20460 30340 20466
rect 30288 20402 30340 20408
rect 30300 20369 30328 20402
rect 30286 20360 30342 20369
rect 30286 20295 30342 20304
rect 30392 20058 30420 20742
rect 30472 20460 30524 20466
rect 30472 20402 30524 20408
rect 30288 20052 30340 20058
rect 30288 19994 30340 20000
rect 30380 20052 30432 20058
rect 30380 19994 30432 20000
rect 30196 19916 30248 19922
rect 30196 19858 30248 19864
rect 30104 19848 30156 19854
rect 30104 19790 30156 19796
rect 30012 19780 30064 19786
rect 30012 19722 30064 19728
rect 29736 18964 29788 18970
rect 29736 18906 29788 18912
rect 29644 14476 29696 14482
rect 29644 14418 29696 14424
rect 29552 13728 29604 13734
rect 29552 13670 29604 13676
rect 29564 13462 29592 13670
rect 29552 13456 29604 13462
rect 29552 13398 29604 13404
rect 29644 13252 29696 13258
rect 29644 13194 29696 13200
rect 29656 12442 29684 13194
rect 29644 12436 29696 12442
rect 29644 12378 29696 12384
rect 29644 12300 29696 12306
rect 29644 12242 29696 12248
rect 29460 11348 29512 11354
rect 29460 11290 29512 11296
rect 29656 10674 29684 12242
rect 29748 12186 29776 18906
rect 29920 18760 29972 18766
rect 29920 18702 29972 18708
rect 29826 16280 29882 16289
rect 29826 16215 29828 16224
rect 29880 16215 29882 16224
rect 29828 16186 29880 16192
rect 29828 16108 29880 16114
rect 29828 16050 29880 16056
rect 29840 14822 29868 16050
rect 29828 14816 29880 14822
rect 29828 14758 29880 14764
rect 29828 13932 29880 13938
rect 29828 13874 29880 13880
rect 29840 12753 29868 13874
rect 29826 12744 29882 12753
rect 29826 12679 29882 12688
rect 29748 12158 29868 12186
rect 29840 11762 29868 12158
rect 29932 11762 29960 18702
rect 30024 11898 30052 19722
rect 30116 18834 30144 19790
rect 30300 19786 30328 19994
rect 30288 19780 30340 19786
rect 30288 19722 30340 19728
rect 30196 19440 30248 19446
rect 30300 19428 30328 19722
rect 30380 19508 30432 19514
rect 30380 19450 30432 19456
rect 30248 19400 30328 19428
rect 30196 19382 30248 19388
rect 30104 18828 30156 18834
rect 30104 18770 30156 18776
rect 30104 16516 30156 16522
rect 30104 16458 30156 16464
rect 30116 16182 30144 16458
rect 30208 16454 30236 19382
rect 30392 18290 30420 19450
rect 30484 19360 30512 20402
rect 30576 20058 30604 20810
rect 30656 20460 30708 20466
rect 30656 20402 30708 20408
rect 30668 20262 30696 20402
rect 30656 20256 30708 20262
rect 30656 20198 30708 20204
rect 30564 20052 30616 20058
rect 30564 19994 30616 20000
rect 30760 19990 30788 22630
rect 30852 21622 30880 23666
rect 30840 21616 30892 21622
rect 30840 21558 30892 21564
rect 30944 20398 30972 26930
rect 31036 25974 31064 28970
rect 31116 28552 31168 28558
rect 31116 28494 31168 28500
rect 31128 28218 31156 28494
rect 31116 28212 31168 28218
rect 31116 28154 31168 28160
rect 31312 27130 31340 31214
rect 31404 30326 31432 33322
rect 31496 32570 31524 33322
rect 31760 33312 31812 33318
rect 31760 33254 31812 33260
rect 31576 32904 31628 32910
rect 31576 32846 31628 32852
rect 31484 32564 31536 32570
rect 31484 32506 31536 32512
rect 31588 32502 31616 32846
rect 31772 32774 31800 33254
rect 31852 33040 31904 33046
rect 31852 32982 31904 32988
rect 31760 32768 31812 32774
rect 31760 32710 31812 32716
rect 31576 32496 31628 32502
rect 31576 32438 31628 32444
rect 31576 31884 31628 31890
rect 31576 31826 31628 31832
rect 31484 31816 31536 31822
rect 31484 31758 31536 31764
rect 31496 31346 31524 31758
rect 31484 31340 31536 31346
rect 31484 31282 31536 31288
rect 31392 30320 31444 30326
rect 31392 30262 31444 30268
rect 31484 29572 31536 29578
rect 31484 29514 31536 29520
rect 31496 29345 31524 29514
rect 31482 29336 31538 29345
rect 31482 29271 31538 29280
rect 31588 28762 31616 31826
rect 31668 29708 31720 29714
rect 31668 29650 31720 29656
rect 31680 29102 31708 29650
rect 31668 29096 31720 29102
rect 31668 29038 31720 29044
rect 31576 28756 31628 28762
rect 31576 28698 31628 28704
rect 31300 27124 31352 27130
rect 31300 27066 31352 27072
rect 31576 26988 31628 26994
rect 31576 26930 31628 26936
rect 31116 26444 31168 26450
rect 31116 26386 31168 26392
rect 31024 25968 31076 25974
rect 31024 25910 31076 25916
rect 31036 24614 31064 25910
rect 31128 25294 31156 26386
rect 31208 26240 31260 26246
rect 31208 26182 31260 26188
rect 31220 25906 31248 26182
rect 31208 25900 31260 25906
rect 31208 25842 31260 25848
rect 31392 25900 31444 25906
rect 31392 25842 31444 25848
rect 31484 25900 31536 25906
rect 31484 25842 31536 25848
rect 31300 25764 31352 25770
rect 31300 25706 31352 25712
rect 31116 25288 31168 25294
rect 31116 25230 31168 25236
rect 31312 24614 31340 25706
rect 31404 25498 31432 25842
rect 31392 25492 31444 25498
rect 31392 25434 31444 25440
rect 31496 25158 31524 25842
rect 31484 25152 31536 25158
rect 31484 25094 31536 25100
rect 31392 24676 31444 24682
rect 31392 24618 31444 24624
rect 31024 24608 31076 24614
rect 31024 24550 31076 24556
rect 31300 24608 31352 24614
rect 31300 24550 31352 24556
rect 31404 24274 31432 24618
rect 31588 24410 31616 26930
rect 31772 24954 31800 32710
rect 31760 24948 31812 24954
rect 31760 24890 31812 24896
rect 31576 24404 31628 24410
rect 31576 24346 31628 24352
rect 31392 24268 31444 24274
rect 31392 24210 31444 24216
rect 31208 23520 31260 23526
rect 31208 23462 31260 23468
rect 31024 22976 31076 22982
rect 31024 22918 31076 22924
rect 31036 22642 31064 22918
rect 31220 22778 31248 23462
rect 31300 23316 31352 23322
rect 31300 23258 31352 23264
rect 31312 22778 31340 23258
rect 31208 22772 31260 22778
rect 31208 22714 31260 22720
rect 31300 22772 31352 22778
rect 31300 22714 31352 22720
rect 31024 22636 31076 22642
rect 31024 22578 31076 22584
rect 31208 22636 31260 22642
rect 31208 22578 31260 22584
rect 31036 20942 31064 22578
rect 31024 20936 31076 20942
rect 31024 20878 31076 20884
rect 31116 20936 31168 20942
rect 31116 20878 31168 20884
rect 30932 20392 30984 20398
rect 30932 20334 30984 20340
rect 30932 20256 30984 20262
rect 30932 20198 30984 20204
rect 30748 19984 30800 19990
rect 30748 19926 30800 19932
rect 30944 19922 30972 20198
rect 31128 20058 31156 20878
rect 31220 20466 31248 22578
rect 31300 21956 31352 21962
rect 31300 21898 31352 21904
rect 31312 20942 31340 21898
rect 31300 20936 31352 20942
rect 31300 20878 31352 20884
rect 31404 20534 31432 24210
rect 31668 23180 31720 23186
rect 31668 23122 31720 23128
rect 31484 23044 31536 23050
rect 31484 22986 31536 22992
rect 31496 22642 31524 22986
rect 31484 22636 31536 22642
rect 31484 22578 31536 22584
rect 31680 22098 31708 23122
rect 31668 22092 31720 22098
rect 31864 22094 31892 32982
rect 31944 32904 31996 32910
rect 31944 32846 31996 32852
rect 31956 30734 31984 32846
rect 31944 30728 31996 30734
rect 31944 30670 31996 30676
rect 32048 29646 32076 33390
rect 32128 32428 32180 32434
rect 32128 32370 32180 32376
rect 32140 31958 32168 32370
rect 32128 31952 32180 31958
rect 32128 31894 32180 31900
rect 32324 31890 32352 33458
rect 33140 33380 33192 33386
rect 33140 33322 33192 33328
rect 34152 33380 34204 33386
rect 34152 33322 34204 33328
rect 33048 33108 33100 33114
rect 33048 33050 33100 33056
rect 32404 32836 32456 32842
rect 32404 32778 32456 32784
rect 32416 32434 32444 32778
rect 32404 32428 32456 32434
rect 32404 32370 32456 32376
rect 32864 32428 32916 32434
rect 32864 32370 32916 32376
rect 32312 31884 32364 31890
rect 32312 31826 32364 31832
rect 32324 31482 32352 31826
rect 32312 31476 32364 31482
rect 32312 31418 32364 31424
rect 32876 31346 32904 32370
rect 33060 31414 33088 33050
rect 33152 32910 33180 33322
rect 34060 33312 34112 33318
rect 34060 33254 34112 33260
rect 33324 33108 33376 33114
rect 33324 33050 33376 33056
rect 33140 32904 33192 32910
rect 33140 32846 33192 32852
rect 33336 32230 33364 33050
rect 34072 32910 34100 33254
rect 34164 33046 34192 33322
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34152 33040 34204 33046
rect 34152 32982 34204 32988
rect 35164 33040 35216 33046
rect 35216 32988 35480 32994
rect 35164 32982 35480 32988
rect 35176 32966 35480 32982
rect 34060 32904 34112 32910
rect 34060 32846 34112 32852
rect 34980 32904 35032 32910
rect 34980 32846 35032 32852
rect 33692 32836 33744 32842
rect 33692 32778 33744 32784
rect 33600 32768 33652 32774
rect 33600 32710 33652 32716
rect 33612 32502 33640 32710
rect 33600 32496 33652 32502
rect 33600 32438 33652 32444
rect 33704 32434 33732 32778
rect 34992 32774 35020 32846
rect 34980 32768 35032 32774
rect 34980 32710 35032 32716
rect 33692 32428 33744 32434
rect 33692 32370 33744 32376
rect 33416 32360 33468 32366
rect 33416 32302 33468 32308
rect 34336 32360 34388 32366
rect 34336 32302 34388 32308
rect 34612 32360 34664 32366
rect 34612 32302 34664 32308
rect 34704 32360 34756 32366
rect 34704 32302 34756 32308
rect 35348 32360 35400 32366
rect 35348 32302 35400 32308
rect 33324 32224 33376 32230
rect 33324 32166 33376 32172
rect 33048 31408 33100 31414
rect 33048 31350 33100 31356
rect 32864 31340 32916 31346
rect 33336 31328 33364 32166
rect 33428 31482 33456 32302
rect 34348 31890 34376 32302
rect 34152 31884 34204 31890
rect 34152 31826 34204 31832
rect 34336 31884 34388 31890
rect 34336 31826 34388 31832
rect 33416 31476 33468 31482
rect 33416 31418 33468 31424
rect 34164 31346 34192 31826
rect 34244 31680 34296 31686
rect 34244 31622 34296 31628
rect 34336 31680 34388 31686
rect 34336 31622 34388 31628
rect 33416 31340 33468 31346
rect 33336 31300 33416 31328
rect 32864 31282 32916 31288
rect 33416 31282 33468 31288
rect 33600 31340 33652 31346
rect 33600 31282 33652 31288
rect 34152 31340 34204 31346
rect 34152 31282 34204 31288
rect 32496 31272 32548 31278
rect 32496 31214 32548 31220
rect 32508 31142 32536 31214
rect 32496 31136 32548 31142
rect 32496 31078 32548 31084
rect 32036 29640 32088 29646
rect 32036 29582 32088 29588
rect 31944 29504 31996 29510
rect 31944 29446 31996 29452
rect 31956 29170 31984 29446
rect 31944 29164 31996 29170
rect 31944 29106 31996 29112
rect 32048 28966 32076 29582
rect 32508 28994 32536 31078
rect 32772 30796 32824 30802
rect 32772 30738 32824 30744
rect 32784 30258 32812 30738
rect 32772 30252 32824 30258
rect 32772 30194 32824 30200
rect 32680 30184 32732 30190
rect 32680 30126 32732 30132
rect 32416 28966 32536 28994
rect 32036 28960 32088 28966
rect 32036 28902 32088 28908
rect 32048 28762 32076 28902
rect 32036 28756 32088 28762
rect 32036 28698 32088 28704
rect 32416 28082 32444 28966
rect 32496 28756 32548 28762
rect 32496 28698 32548 28704
rect 32508 28558 32536 28698
rect 32496 28552 32548 28558
rect 32496 28494 32548 28500
rect 32128 28076 32180 28082
rect 32128 28018 32180 28024
rect 32404 28076 32456 28082
rect 32404 28018 32456 28024
rect 32140 27130 32168 28018
rect 32128 27124 32180 27130
rect 32128 27066 32180 27072
rect 32416 26994 32444 28018
rect 32508 27878 32536 28494
rect 32588 28008 32640 28014
rect 32588 27950 32640 27956
rect 32496 27872 32548 27878
rect 32496 27814 32548 27820
rect 32404 26988 32456 26994
rect 32404 26930 32456 26936
rect 32508 26450 32536 27814
rect 32496 26444 32548 26450
rect 32496 26386 32548 26392
rect 32220 26376 32272 26382
rect 32220 26318 32272 26324
rect 32232 26042 32260 26318
rect 32312 26308 32364 26314
rect 32312 26250 32364 26256
rect 32220 26036 32272 26042
rect 32220 25978 32272 25984
rect 32218 25936 32274 25945
rect 32324 25906 32352 26250
rect 32600 26042 32628 27950
rect 32588 26036 32640 26042
rect 32588 25978 32640 25984
rect 32218 25871 32220 25880
rect 32272 25871 32274 25880
rect 32312 25900 32364 25906
rect 32220 25842 32272 25848
rect 32312 25842 32364 25848
rect 32496 25832 32548 25838
rect 32496 25774 32548 25780
rect 31944 25764 31996 25770
rect 31944 25706 31996 25712
rect 31956 24070 31984 25706
rect 32128 25220 32180 25226
rect 32128 25162 32180 25168
rect 32036 24812 32088 24818
rect 32036 24754 32088 24760
rect 32048 24206 32076 24754
rect 32140 24206 32168 25162
rect 32508 25158 32536 25774
rect 32588 25288 32640 25294
rect 32588 25230 32640 25236
rect 32496 25152 32548 25158
rect 32496 25094 32548 25100
rect 32220 24948 32272 24954
rect 32220 24890 32272 24896
rect 32232 24342 32260 24890
rect 32220 24336 32272 24342
rect 32220 24278 32272 24284
rect 32036 24200 32088 24206
rect 32036 24142 32088 24148
rect 32128 24200 32180 24206
rect 32128 24142 32180 24148
rect 31944 24064 31996 24070
rect 31944 24006 31996 24012
rect 31956 23866 31984 24006
rect 31944 23860 31996 23866
rect 31944 23802 31996 23808
rect 31944 22772 31996 22778
rect 31944 22714 31996 22720
rect 31956 22574 31984 22714
rect 32048 22642 32076 24142
rect 32232 23746 32260 24278
rect 32404 24064 32456 24070
rect 32404 24006 32456 24012
rect 32416 23866 32444 24006
rect 32404 23860 32456 23866
rect 32404 23802 32456 23808
rect 32140 23730 32260 23746
rect 32600 23730 32628 25230
rect 32128 23724 32260 23730
rect 32180 23718 32260 23724
rect 32312 23724 32364 23730
rect 32128 23666 32180 23672
rect 32312 23666 32364 23672
rect 32404 23724 32456 23730
rect 32404 23666 32456 23672
rect 32588 23724 32640 23730
rect 32588 23666 32640 23672
rect 32140 23254 32168 23666
rect 32128 23248 32180 23254
rect 32128 23190 32180 23196
rect 32220 23044 32272 23050
rect 32220 22986 32272 22992
rect 32232 22642 32260 22986
rect 32324 22710 32352 23666
rect 32312 22704 32364 22710
rect 32312 22646 32364 22652
rect 32416 22642 32444 23666
rect 32600 22778 32628 23666
rect 32692 23322 32720 30126
rect 32772 29504 32824 29510
rect 32772 29446 32824 29452
rect 32784 28626 32812 29446
rect 32772 28620 32824 28626
rect 32772 28562 32824 28568
rect 32784 28082 32812 28562
rect 32772 28076 32824 28082
rect 32772 28018 32824 28024
rect 32876 27538 32904 31282
rect 32956 31136 33008 31142
rect 32956 31078 33008 31084
rect 32968 30938 32996 31078
rect 32956 30932 33008 30938
rect 32956 30874 33008 30880
rect 33508 30660 33560 30666
rect 33508 30602 33560 30608
rect 33048 29300 33100 29306
rect 33048 29242 33100 29248
rect 33060 28762 33088 29242
rect 33520 29170 33548 30602
rect 33140 29164 33192 29170
rect 33140 29106 33192 29112
rect 33508 29164 33560 29170
rect 33508 29106 33560 29112
rect 33048 28756 33100 28762
rect 33048 28698 33100 28704
rect 33152 28694 33180 29106
rect 33140 28688 33192 28694
rect 33140 28630 33192 28636
rect 33048 28552 33100 28558
rect 33048 28494 33100 28500
rect 32956 28076 33008 28082
rect 32956 28018 33008 28024
rect 32864 27532 32916 27538
rect 32864 27474 32916 27480
rect 32968 27418 32996 28018
rect 32876 27390 32996 27418
rect 32772 26920 32824 26926
rect 32772 26862 32824 26868
rect 32784 24070 32812 26862
rect 32876 25838 32904 27390
rect 32956 26920 33008 26926
rect 32956 26862 33008 26868
rect 32968 26586 32996 26862
rect 32956 26580 33008 26586
rect 32956 26522 33008 26528
rect 32956 26376 33008 26382
rect 32956 26318 33008 26324
rect 32968 26042 32996 26318
rect 32956 26036 33008 26042
rect 32956 25978 33008 25984
rect 32864 25832 32916 25838
rect 32864 25774 32916 25780
rect 32876 25430 32904 25774
rect 32864 25424 32916 25430
rect 32864 25366 32916 25372
rect 32968 25294 32996 25978
rect 33060 25498 33088 28494
rect 33324 28484 33376 28490
rect 33324 28426 33376 28432
rect 33336 28082 33364 28426
rect 33612 28082 33640 31282
rect 33968 31136 34020 31142
rect 33968 31078 34020 31084
rect 33980 29646 34008 31078
rect 34164 30682 34192 31282
rect 34256 31210 34284 31622
rect 34348 31346 34376 31622
rect 34624 31346 34652 32302
rect 34716 32026 34744 32302
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34704 32020 34756 32026
rect 34704 31962 34756 31968
rect 35360 31414 35388 32302
rect 35452 31482 35480 32966
rect 36636 32904 36688 32910
rect 36636 32846 36688 32852
rect 35992 32768 36044 32774
rect 35992 32710 36044 32716
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 36004 31482 36032 32710
rect 35440 31476 35492 31482
rect 35440 31418 35492 31424
rect 35992 31476 36044 31482
rect 35992 31418 36044 31424
rect 35348 31408 35400 31414
rect 35348 31350 35400 31356
rect 34336 31340 34388 31346
rect 34336 31282 34388 31288
rect 34612 31340 34664 31346
rect 34612 31282 34664 31288
rect 34796 31340 34848 31346
rect 34796 31282 34848 31288
rect 34244 31204 34296 31210
rect 34244 31146 34296 31152
rect 34072 30666 34192 30682
rect 34348 30666 34376 31282
rect 34624 30938 34652 31282
rect 34612 30932 34664 30938
rect 34612 30874 34664 30880
rect 34612 30796 34664 30802
rect 34612 30738 34664 30744
rect 34060 30660 34192 30666
rect 34112 30654 34192 30660
rect 34336 30660 34388 30666
rect 34060 30602 34112 30608
rect 34336 30602 34388 30608
rect 33784 29640 33836 29646
rect 33784 29582 33836 29588
rect 33968 29640 34020 29646
rect 33968 29582 34020 29588
rect 33796 28218 33824 29582
rect 33784 28212 33836 28218
rect 33784 28154 33836 28160
rect 33324 28076 33376 28082
rect 33324 28018 33376 28024
rect 33600 28076 33652 28082
rect 33600 28018 33652 28024
rect 33876 28076 33928 28082
rect 33876 28018 33928 28024
rect 33232 26988 33284 26994
rect 33232 26930 33284 26936
rect 33140 26784 33192 26790
rect 33140 26726 33192 26732
rect 33152 26382 33180 26726
rect 33244 26450 33272 26930
rect 33232 26444 33284 26450
rect 33232 26386 33284 26392
rect 33140 26376 33192 26382
rect 33336 26330 33364 28018
rect 33784 26988 33836 26994
rect 33784 26930 33836 26936
rect 33416 26784 33468 26790
rect 33416 26726 33468 26732
rect 33428 26586 33456 26726
rect 33416 26580 33468 26586
rect 33416 26522 33468 26528
rect 33140 26318 33192 26324
rect 33244 26302 33364 26330
rect 33416 26376 33468 26382
rect 33796 26353 33824 26930
rect 33416 26318 33468 26324
rect 33782 26344 33838 26353
rect 33244 25838 33272 26302
rect 33232 25832 33284 25838
rect 33232 25774 33284 25780
rect 33048 25492 33100 25498
rect 33048 25434 33100 25440
rect 32956 25288 33008 25294
rect 32956 25230 33008 25236
rect 33244 25226 33272 25774
rect 33324 25288 33376 25294
rect 33324 25230 33376 25236
rect 33232 25220 33284 25226
rect 33232 25162 33284 25168
rect 33048 24608 33100 24614
rect 33048 24550 33100 24556
rect 33232 24608 33284 24614
rect 33232 24550 33284 24556
rect 32864 24200 32916 24206
rect 32864 24142 32916 24148
rect 32772 24064 32824 24070
rect 32772 24006 32824 24012
rect 32772 23792 32824 23798
rect 32772 23734 32824 23740
rect 32680 23316 32732 23322
rect 32680 23258 32732 23264
rect 32680 23044 32732 23050
rect 32680 22986 32732 22992
rect 32588 22772 32640 22778
rect 32588 22714 32640 22720
rect 32036 22636 32088 22642
rect 32036 22578 32088 22584
rect 32128 22636 32180 22642
rect 32128 22578 32180 22584
rect 32220 22636 32272 22642
rect 32220 22578 32272 22584
rect 32404 22636 32456 22642
rect 32404 22578 32456 22584
rect 32496 22636 32548 22642
rect 32496 22578 32548 22584
rect 31944 22568 31996 22574
rect 31944 22510 31996 22516
rect 31668 22034 31720 22040
rect 31772 22066 31892 22094
rect 31484 21548 31536 21554
rect 31484 21490 31536 21496
rect 31496 20874 31524 21490
rect 31576 21344 31628 21350
rect 31576 21286 31628 21292
rect 31588 21078 31616 21286
rect 31772 21078 31800 22066
rect 32048 22030 32076 22578
rect 32140 22234 32168 22578
rect 32128 22228 32180 22234
rect 32128 22170 32180 22176
rect 32036 22024 32088 22030
rect 32036 21966 32088 21972
rect 32404 21956 32456 21962
rect 32404 21898 32456 21904
rect 32416 21146 32444 21898
rect 32508 21894 32536 22578
rect 32692 22234 32720 22986
rect 32784 22642 32812 23734
rect 32772 22636 32824 22642
rect 32772 22578 32824 22584
rect 32680 22228 32732 22234
rect 32680 22170 32732 22176
rect 32496 21888 32548 21894
rect 32496 21830 32548 21836
rect 31852 21140 31904 21146
rect 31852 21082 31904 21088
rect 32404 21140 32456 21146
rect 32404 21082 32456 21088
rect 31576 21072 31628 21078
rect 31576 21014 31628 21020
rect 31760 21072 31812 21078
rect 31760 21014 31812 21020
rect 31484 20868 31536 20874
rect 31484 20810 31536 20816
rect 31576 20868 31628 20874
rect 31576 20810 31628 20816
rect 31588 20602 31616 20810
rect 31576 20596 31628 20602
rect 31576 20538 31628 20544
rect 31392 20528 31444 20534
rect 31392 20470 31444 20476
rect 31208 20460 31260 20466
rect 31208 20402 31260 20408
rect 31300 20392 31352 20398
rect 31206 20360 31262 20369
rect 31300 20334 31352 20340
rect 31206 20295 31208 20304
rect 31260 20295 31262 20304
rect 31208 20266 31260 20272
rect 31116 20052 31168 20058
rect 31116 19994 31168 20000
rect 31220 19922 31248 20266
rect 30932 19916 30984 19922
rect 30932 19858 30984 19864
rect 31208 19916 31260 19922
rect 31208 19858 31260 19864
rect 30656 19712 30708 19718
rect 30656 19654 30708 19660
rect 30668 19514 30696 19654
rect 31220 19514 31248 19858
rect 31312 19854 31340 20334
rect 31772 19990 31800 21014
rect 31864 20398 31892 21082
rect 32876 20942 32904 24142
rect 33060 24138 33088 24550
rect 33140 24404 33192 24410
rect 33140 24346 33192 24352
rect 33048 24132 33100 24138
rect 33048 24074 33100 24080
rect 33152 23730 33180 24346
rect 33244 23866 33272 24550
rect 33336 24138 33364 25230
rect 33428 24682 33456 26318
rect 33782 26279 33838 26288
rect 33692 25288 33744 25294
rect 33692 25230 33744 25236
rect 33508 25152 33560 25158
rect 33508 25094 33560 25100
rect 33416 24676 33468 24682
rect 33416 24618 33468 24624
rect 33324 24132 33376 24138
rect 33324 24074 33376 24080
rect 33428 24018 33456 24618
rect 33336 23990 33456 24018
rect 33232 23860 33284 23866
rect 33232 23802 33284 23808
rect 33140 23724 33192 23730
rect 33140 23666 33192 23672
rect 32956 22432 33008 22438
rect 32956 22374 33008 22380
rect 32968 22030 32996 22374
rect 32956 22024 33008 22030
rect 32956 21966 33008 21972
rect 33336 21010 33364 23990
rect 33520 22234 33548 25094
rect 33704 24954 33732 25230
rect 33784 25152 33836 25158
rect 33784 25094 33836 25100
rect 33692 24948 33744 24954
rect 33692 24890 33744 24896
rect 33796 24614 33824 25094
rect 33784 24608 33836 24614
rect 33784 24550 33836 24556
rect 33796 24206 33824 24550
rect 33784 24200 33836 24206
rect 33784 24142 33836 24148
rect 33600 22500 33652 22506
rect 33600 22442 33652 22448
rect 33508 22228 33560 22234
rect 33508 22170 33560 22176
rect 33508 22024 33560 22030
rect 33612 22012 33640 22442
rect 33560 21984 33640 22012
rect 33692 22024 33744 22030
rect 33508 21966 33560 21972
rect 33692 21966 33744 21972
rect 33324 21004 33376 21010
rect 33324 20946 33376 20952
rect 32864 20936 32916 20942
rect 32864 20878 32916 20884
rect 33232 20936 33284 20942
rect 33232 20878 33284 20884
rect 32402 20496 32458 20505
rect 32402 20431 32458 20440
rect 31852 20392 31904 20398
rect 31852 20334 31904 20340
rect 31760 19984 31812 19990
rect 31760 19926 31812 19932
rect 31300 19848 31352 19854
rect 31300 19790 31352 19796
rect 30656 19508 30708 19514
rect 30656 19450 30708 19456
rect 31208 19508 31260 19514
rect 31208 19450 31260 19456
rect 31312 19378 31340 19790
rect 31668 19780 31720 19786
rect 31668 19722 31720 19728
rect 31680 19378 31708 19722
rect 30748 19372 30800 19378
rect 30484 19332 30748 19360
rect 30748 19314 30800 19320
rect 31300 19372 31352 19378
rect 31300 19314 31352 19320
rect 31668 19372 31720 19378
rect 31668 19314 31720 19320
rect 30656 18896 30708 18902
rect 30656 18838 30708 18844
rect 30380 18284 30432 18290
rect 30380 18226 30432 18232
rect 30472 18080 30524 18086
rect 30472 18022 30524 18028
rect 30484 17746 30512 18022
rect 30472 17740 30524 17746
rect 30472 17682 30524 17688
rect 30564 17672 30616 17678
rect 30564 17614 30616 17620
rect 30472 17264 30524 17270
rect 30472 17206 30524 17212
rect 30196 16448 30248 16454
rect 30196 16390 30248 16396
rect 30208 16182 30236 16390
rect 30104 16176 30156 16182
rect 30104 16118 30156 16124
rect 30196 16176 30248 16182
rect 30196 16118 30248 16124
rect 30380 16108 30432 16114
rect 30380 16050 30432 16056
rect 30392 15638 30420 16050
rect 30380 15632 30432 15638
rect 30380 15574 30432 15580
rect 30196 15496 30248 15502
rect 30196 15438 30248 15444
rect 30102 15056 30158 15065
rect 30102 14991 30158 15000
rect 30116 14958 30144 14991
rect 30104 14952 30156 14958
rect 30104 14894 30156 14900
rect 30208 14550 30236 15438
rect 30484 15026 30512 17206
rect 30576 16833 30604 17614
rect 30562 16824 30618 16833
rect 30562 16759 30618 16768
rect 30668 16046 30696 18838
rect 30760 16794 30788 19314
rect 32416 18766 32444 20431
rect 33244 20398 33272 20878
rect 33336 20534 33364 20946
rect 33416 20936 33468 20942
rect 33416 20878 33468 20884
rect 33428 20534 33456 20878
rect 33520 20602 33548 21966
rect 33704 21146 33732 21966
rect 33692 21140 33744 21146
rect 33692 21082 33744 21088
rect 33796 20602 33824 24142
rect 33888 23186 33916 28018
rect 34072 26994 34100 30602
rect 34348 29782 34376 30602
rect 34624 30326 34652 30738
rect 34612 30320 34664 30326
rect 34612 30262 34664 30268
rect 34336 29776 34388 29782
rect 34336 29718 34388 29724
rect 34152 29164 34204 29170
rect 34152 29106 34204 29112
rect 34164 29073 34192 29106
rect 34348 29102 34376 29718
rect 34428 29640 34480 29646
rect 34428 29582 34480 29588
rect 34440 29170 34468 29582
rect 34428 29164 34480 29170
rect 34428 29106 34480 29112
rect 34336 29096 34388 29102
rect 34150 29064 34206 29073
rect 34336 29038 34388 29044
rect 34150 28999 34206 29008
rect 34164 28218 34192 28999
rect 34428 28960 34480 28966
rect 34428 28902 34480 28908
rect 34440 28490 34468 28902
rect 34428 28484 34480 28490
rect 34428 28426 34480 28432
rect 34152 28212 34204 28218
rect 34152 28154 34204 28160
rect 34428 28076 34480 28082
rect 34428 28018 34480 28024
rect 34440 27402 34468 28018
rect 34520 27464 34572 27470
rect 34520 27406 34572 27412
rect 34428 27396 34480 27402
rect 34428 27338 34480 27344
rect 34336 27328 34388 27334
rect 34336 27270 34388 27276
rect 34060 26988 34112 26994
rect 34060 26930 34112 26936
rect 34348 26382 34376 27270
rect 34440 27062 34468 27338
rect 34428 27056 34480 27062
rect 34428 26998 34480 27004
rect 34336 26376 34388 26382
rect 34336 26318 34388 26324
rect 34244 26308 34296 26314
rect 34244 26250 34296 26256
rect 33968 24812 34020 24818
rect 33968 24754 34020 24760
rect 33980 23474 34008 24754
rect 34256 24614 34284 26250
rect 34336 26240 34388 26246
rect 34532 26228 34560 27406
rect 34624 26466 34652 30262
rect 34808 29850 34836 31282
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34796 29844 34848 29850
rect 34796 29786 34848 29792
rect 34980 29504 35032 29510
rect 34980 29446 35032 29452
rect 34992 29238 35020 29446
rect 35162 29336 35218 29345
rect 35162 29271 35218 29280
rect 34980 29232 35032 29238
rect 34980 29174 35032 29180
rect 35176 29170 35204 29271
rect 34796 29164 34848 29170
rect 34796 29106 34848 29112
rect 35164 29164 35216 29170
rect 35164 29106 35216 29112
rect 34704 28076 34756 28082
rect 34704 28018 34756 28024
rect 34716 26994 34744 28018
rect 34808 27470 34836 29106
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35256 28484 35308 28490
rect 35256 28426 35308 28432
rect 35268 28082 35296 28426
rect 35256 28076 35308 28082
rect 35256 28018 35308 28024
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34796 27464 34848 27470
rect 34796 27406 34848 27412
rect 34888 27464 34940 27470
rect 34888 27406 34940 27412
rect 34900 27130 34928 27406
rect 34888 27124 34940 27130
rect 34888 27066 34940 27072
rect 35360 26994 35388 31350
rect 35440 31340 35492 31346
rect 35440 31282 35492 31288
rect 35716 31340 35768 31346
rect 35716 31282 35768 31288
rect 36084 31340 36136 31346
rect 36084 31282 36136 31288
rect 36268 31340 36320 31346
rect 36268 31282 36320 31288
rect 36360 31340 36412 31346
rect 36360 31282 36412 31288
rect 36544 31340 36596 31346
rect 36544 31282 36596 31288
rect 35452 30734 35480 31282
rect 35728 30802 35756 31282
rect 35716 30796 35768 30802
rect 35716 30738 35768 30744
rect 35992 30796 36044 30802
rect 35992 30738 36044 30744
rect 35440 30728 35492 30734
rect 35440 30670 35492 30676
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 36004 29170 36032 30738
rect 36096 30734 36124 31282
rect 36084 30728 36136 30734
rect 36136 30688 36216 30716
rect 36084 30670 36136 30676
rect 36188 29170 36216 30688
rect 35532 29164 35584 29170
rect 35532 29106 35584 29112
rect 35992 29164 36044 29170
rect 35992 29106 36044 29112
rect 36176 29164 36228 29170
rect 36176 29106 36228 29112
rect 35440 29028 35492 29034
rect 35440 28970 35492 28976
rect 35452 28694 35480 28970
rect 35544 28694 35572 29106
rect 35808 28960 35860 28966
rect 35808 28902 35860 28908
rect 35624 28756 35676 28762
rect 35624 28698 35676 28704
rect 35440 28688 35492 28694
rect 35440 28630 35492 28636
rect 35532 28688 35584 28694
rect 35532 28630 35584 28636
rect 35452 28014 35480 28630
rect 35636 28490 35664 28698
rect 35820 28558 35848 28902
rect 36188 28608 36216 29106
rect 36280 28762 36308 31282
rect 36372 30938 36400 31282
rect 36360 30932 36412 30938
rect 36360 30874 36412 30880
rect 36452 29708 36504 29714
rect 36452 29650 36504 29656
rect 36360 29640 36412 29646
rect 36360 29582 36412 29588
rect 36372 29306 36400 29582
rect 36360 29300 36412 29306
rect 36360 29242 36412 29248
rect 36360 29164 36412 29170
rect 36360 29106 36412 29112
rect 36372 28762 36400 29106
rect 36268 28756 36320 28762
rect 36268 28698 36320 28704
rect 36360 28756 36412 28762
rect 36360 28698 36412 28704
rect 36268 28620 36320 28626
rect 36188 28580 36268 28608
rect 36268 28562 36320 28568
rect 35808 28552 35860 28558
rect 35808 28494 35860 28500
rect 35900 28552 35952 28558
rect 35900 28494 35952 28500
rect 35992 28552 36044 28558
rect 36464 28529 36492 29650
rect 35992 28494 36044 28500
rect 36450 28520 36506 28529
rect 35624 28484 35676 28490
rect 35624 28426 35676 28432
rect 35912 28422 35940 28494
rect 35900 28416 35952 28422
rect 35900 28358 35952 28364
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 36004 28218 36032 28494
rect 36450 28455 36506 28464
rect 36452 28416 36504 28422
rect 36452 28358 36504 28364
rect 35992 28212 36044 28218
rect 35992 28154 36044 28160
rect 35440 28008 35492 28014
rect 35440 27950 35492 27956
rect 36464 27470 36492 28358
rect 36452 27464 36504 27470
rect 36452 27406 36504 27412
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 36176 27056 36228 27062
rect 36176 26998 36228 27004
rect 34704 26988 34756 26994
rect 34704 26930 34756 26936
rect 35348 26988 35400 26994
rect 35348 26930 35400 26936
rect 35440 26988 35492 26994
rect 35440 26930 35492 26936
rect 34716 26586 34744 26930
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34704 26580 34756 26586
rect 34704 26522 34756 26528
rect 34624 26438 34744 26466
rect 34388 26200 34560 26228
rect 34336 26182 34388 26188
rect 34244 24608 34296 24614
rect 34244 24550 34296 24556
rect 33980 23446 34284 23474
rect 33876 23180 33928 23186
rect 33928 23140 34008 23168
rect 33876 23122 33928 23128
rect 33874 23080 33930 23089
rect 33874 23015 33930 23024
rect 33888 22982 33916 23015
rect 33876 22976 33928 22982
rect 33876 22918 33928 22924
rect 33888 22642 33916 22918
rect 33980 22778 34008 23140
rect 33968 22772 34020 22778
rect 33968 22714 34020 22720
rect 33876 22636 33928 22642
rect 33876 22578 33928 22584
rect 34060 22568 34112 22574
rect 34060 22510 34112 22516
rect 34072 22030 34100 22510
rect 34060 22024 34112 22030
rect 34060 21966 34112 21972
rect 33876 21004 33928 21010
rect 33876 20946 33928 20952
rect 33508 20596 33560 20602
rect 33508 20538 33560 20544
rect 33784 20596 33836 20602
rect 33784 20538 33836 20544
rect 33324 20528 33376 20534
rect 33324 20470 33376 20476
rect 33416 20528 33468 20534
rect 33416 20470 33468 20476
rect 33232 20392 33284 20398
rect 33232 20334 33284 20340
rect 33140 20256 33192 20262
rect 33140 20198 33192 20204
rect 33232 20256 33284 20262
rect 33232 20198 33284 20204
rect 32404 18760 32456 18766
rect 32404 18702 32456 18708
rect 33152 18306 33180 20198
rect 33244 19990 33272 20198
rect 33232 19984 33284 19990
rect 33232 19926 33284 19932
rect 33428 19718 33456 20470
rect 33888 20398 33916 20946
rect 34072 20602 34100 21966
rect 34152 21344 34204 21350
rect 34152 21286 34204 21292
rect 34164 20942 34192 21286
rect 34256 21078 34284 23446
rect 34348 22642 34376 26182
rect 34428 24812 34480 24818
rect 34428 24754 34480 24760
rect 34440 24206 34468 24754
rect 34428 24200 34480 24206
rect 34428 24142 34480 24148
rect 34612 24200 34664 24206
rect 34612 24142 34664 24148
rect 34426 23896 34482 23905
rect 34426 23831 34482 23840
rect 34440 22760 34468 23831
rect 34624 23798 34652 24142
rect 34612 23792 34664 23798
rect 34612 23734 34664 23740
rect 34520 23520 34572 23526
rect 34520 23462 34572 23468
rect 34532 23186 34560 23462
rect 34520 23180 34572 23186
rect 34520 23122 34572 23128
rect 34612 22772 34664 22778
rect 34440 22732 34612 22760
rect 34612 22714 34664 22720
rect 34716 22658 34744 26438
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34888 24200 34940 24206
rect 34888 24142 34940 24148
rect 35164 24200 35216 24206
rect 35164 24142 35216 24148
rect 34900 23866 34928 24142
rect 34888 23860 34940 23866
rect 34888 23802 34940 23808
rect 34796 23656 34848 23662
rect 34796 23598 34848 23604
rect 35176 23610 35204 24142
rect 35256 24064 35308 24070
rect 35256 24006 35308 24012
rect 35268 23730 35296 24006
rect 35256 23724 35308 23730
rect 35256 23666 35308 23672
rect 35360 23662 35388 26930
rect 35452 26586 35480 26930
rect 35992 26920 36044 26926
rect 35992 26862 36044 26868
rect 35440 26580 35492 26586
rect 35440 26522 35492 26528
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 36004 23866 36032 26862
rect 36188 24818 36216 26998
rect 36464 25362 36492 27406
rect 36556 27130 36584 31282
rect 36544 27124 36596 27130
rect 36544 27066 36596 27072
rect 36648 27062 36676 32846
rect 37188 30048 37240 30054
rect 37188 29990 37240 29996
rect 37200 29646 37228 29990
rect 37188 29640 37240 29646
rect 37188 29582 37240 29588
rect 36820 29504 36872 29510
rect 36820 29446 36872 29452
rect 36832 29209 36860 29446
rect 36818 29200 36874 29209
rect 36818 29135 36874 29144
rect 36728 29096 36780 29102
rect 36728 29038 36780 29044
rect 36740 28966 36768 29038
rect 36728 28960 36780 28966
rect 36728 28902 36780 28908
rect 36740 28762 36768 28902
rect 36728 28756 36780 28762
rect 36728 28698 36780 28704
rect 36728 28620 36780 28626
rect 36728 28562 36780 28568
rect 36740 28218 36768 28562
rect 37096 28552 37148 28558
rect 37096 28494 37148 28500
rect 37278 28520 37334 28529
rect 36728 28212 36780 28218
rect 36728 28154 36780 28160
rect 36728 27940 36780 27946
rect 36728 27882 36780 27888
rect 36740 27452 36768 27882
rect 37108 27538 37136 28494
rect 37278 28455 37334 28464
rect 37096 27532 37148 27538
rect 37096 27474 37148 27480
rect 36820 27464 36872 27470
rect 36740 27424 36820 27452
rect 36740 27062 36768 27424
rect 36820 27406 36872 27412
rect 36636 27056 36688 27062
rect 36636 26998 36688 27004
rect 36728 27056 36780 27062
rect 36728 26998 36780 27004
rect 36740 26518 36768 26998
rect 36820 26988 36872 26994
rect 36820 26930 36872 26936
rect 36832 26586 36860 26930
rect 37004 26784 37056 26790
rect 37004 26726 37056 26732
rect 37016 26586 37044 26726
rect 36820 26580 36872 26586
rect 36820 26522 36872 26528
rect 37004 26580 37056 26586
rect 37004 26522 37056 26528
rect 36728 26512 36780 26518
rect 36728 26454 36780 26460
rect 36728 26376 36780 26382
rect 36728 26318 36780 26324
rect 36740 25498 36768 26318
rect 36728 25492 36780 25498
rect 36728 25434 36780 25440
rect 36452 25356 36504 25362
rect 36452 25298 36504 25304
rect 37004 25288 37056 25294
rect 37004 25230 37056 25236
rect 36636 25152 36688 25158
rect 36636 25094 36688 25100
rect 36728 25152 36780 25158
rect 36728 25094 36780 25100
rect 36176 24812 36228 24818
rect 36176 24754 36228 24760
rect 36648 24614 36676 25094
rect 36740 24750 36768 25094
rect 36728 24744 36780 24750
rect 36728 24686 36780 24692
rect 36912 24744 36964 24750
rect 36912 24686 36964 24692
rect 36636 24608 36688 24614
rect 36636 24550 36688 24556
rect 36268 24336 36320 24342
rect 36268 24278 36320 24284
rect 36084 24200 36136 24206
rect 36084 24142 36136 24148
rect 35992 23860 36044 23866
rect 35992 23802 36044 23808
rect 36096 23746 36124 24142
rect 36280 23866 36308 24278
rect 36648 23866 36676 24550
rect 36268 23860 36320 23866
rect 36268 23802 36320 23808
rect 36636 23860 36688 23866
rect 36636 23802 36688 23808
rect 35440 23724 35492 23730
rect 35440 23666 35492 23672
rect 36004 23718 36124 23746
rect 35348 23656 35400 23662
rect 34336 22636 34388 22642
rect 34336 22578 34388 22584
rect 34624 22630 34744 22658
rect 34808 22642 34836 23598
rect 35176 23582 35296 23610
rect 35348 23598 35400 23604
rect 35268 23474 35296 23582
rect 35268 23446 35301 23474
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35273 23338 35301 23446
rect 35268 23310 35301 23338
rect 34796 22636 34848 22642
rect 34428 22568 34480 22574
rect 34428 22510 34480 22516
rect 34440 22030 34468 22510
rect 34624 22098 34652 22630
rect 34796 22578 34848 22584
rect 34704 22500 34756 22506
rect 34704 22442 34756 22448
rect 34612 22092 34664 22098
rect 34612 22034 34664 22040
rect 34428 22024 34480 22030
rect 34428 21966 34480 21972
rect 34440 21078 34468 21966
rect 34716 21894 34744 22442
rect 34808 22094 34836 22578
rect 34888 22568 34940 22574
rect 34886 22536 34888 22545
rect 34940 22536 34942 22545
rect 34886 22471 34942 22480
rect 35268 22386 35296 23310
rect 35360 22778 35388 23598
rect 35348 22772 35400 22778
rect 35452 22760 35480 23666
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 36004 22778 36032 23718
rect 36268 23656 36320 23662
rect 36268 23598 36320 23604
rect 36084 23520 36136 23526
rect 36084 23462 36136 23468
rect 35900 22772 35952 22778
rect 35452 22732 35664 22760
rect 35348 22714 35400 22720
rect 35636 22642 35664 22732
rect 35900 22714 35952 22720
rect 35992 22772 36044 22778
rect 35992 22714 36044 22720
rect 35532 22636 35584 22642
rect 35532 22578 35584 22584
rect 35624 22636 35676 22642
rect 35624 22578 35676 22584
rect 35716 22636 35768 22642
rect 35716 22578 35768 22584
rect 35268 22358 35301 22386
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35273 22250 35301 22358
rect 35268 22234 35301 22250
rect 35544 22234 35572 22578
rect 35256 22228 35308 22234
rect 35256 22170 35308 22176
rect 35532 22228 35584 22234
rect 35532 22170 35584 22176
rect 35268 22094 35296 22170
rect 35728 22166 35756 22578
rect 35912 22234 35940 22714
rect 36004 22438 36032 22714
rect 35992 22432 36044 22438
rect 35992 22374 36044 22380
rect 35900 22228 35952 22234
rect 35900 22170 35952 22176
rect 35716 22160 35768 22166
rect 35716 22102 35768 22108
rect 34808 22066 34928 22094
rect 34704 21888 34756 21894
rect 34704 21830 34756 21836
rect 34796 21888 34848 21894
rect 34796 21830 34848 21836
rect 34520 21548 34572 21554
rect 34520 21490 34572 21496
rect 34244 21072 34296 21078
rect 34244 21014 34296 21020
rect 34428 21072 34480 21078
rect 34428 21014 34480 21020
rect 34152 20936 34204 20942
rect 34152 20878 34204 20884
rect 34060 20596 34112 20602
rect 34060 20538 34112 20544
rect 33968 20460 34020 20466
rect 33968 20402 34020 20408
rect 33784 20392 33836 20398
rect 33784 20334 33836 20340
rect 33876 20392 33928 20398
rect 33876 20334 33928 20340
rect 33416 19712 33468 19718
rect 33416 19654 33468 19660
rect 33428 19378 33456 19654
rect 33416 19372 33468 19378
rect 33416 19314 33468 19320
rect 33428 18970 33456 19314
rect 33416 18964 33468 18970
rect 33416 18906 33468 18912
rect 33796 18902 33824 20334
rect 33980 20058 34008 20402
rect 33968 20052 34020 20058
rect 33968 19994 34020 20000
rect 33876 19916 33928 19922
rect 33876 19858 33928 19864
rect 33888 19378 33916 19858
rect 34256 19825 34284 21014
rect 34532 21010 34560 21490
rect 34716 21146 34744 21830
rect 34704 21140 34756 21146
rect 34704 21082 34756 21088
rect 34520 21004 34572 21010
rect 34520 20946 34572 20952
rect 34428 20936 34480 20942
rect 34428 20878 34480 20884
rect 34242 19816 34298 19825
rect 34242 19751 34298 19760
rect 34440 19378 34468 20878
rect 34532 19922 34560 20946
rect 34612 20868 34664 20874
rect 34612 20810 34664 20816
rect 34520 19916 34572 19922
rect 34520 19858 34572 19864
rect 34624 19378 34652 20810
rect 34808 20058 34836 21830
rect 34900 21690 34928 22066
rect 35176 22066 35296 22094
rect 35176 22030 35204 22066
rect 35164 22024 35216 22030
rect 35164 21966 35216 21972
rect 35164 21888 35216 21894
rect 35164 21830 35216 21836
rect 35176 21690 35204 21830
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 34888 21684 34940 21690
rect 34888 21626 34940 21632
rect 35164 21684 35216 21690
rect 35164 21626 35216 21632
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 36004 20942 36032 22374
rect 35992 20936 36044 20942
rect 35992 20878 36044 20884
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 36096 20058 36124 23462
rect 36280 23322 36308 23598
rect 36268 23316 36320 23322
rect 36268 23258 36320 23264
rect 36266 22672 36322 22681
rect 36266 22607 36268 22616
rect 36320 22607 36322 22616
rect 36268 22578 36320 22584
rect 36266 22536 36322 22545
rect 36266 22471 36268 22480
rect 36320 22471 36322 22480
rect 36268 22442 36320 22448
rect 36544 20256 36596 20262
rect 36544 20198 36596 20204
rect 36556 20058 36584 20198
rect 36648 20058 36676 23802
rect 36740 23662 36768 24686
rect 36820 24608 36872 24614
rect 36820 24550 36872 24556
rect 36832 23866 36860 24550
rect 36924 24138 36952 24686
rect 37016 24206 37044 25230
rect 37004 24200 37056 24206
rect 37004 24142 37056 24148
rect 36912 24132 36964 24138
rect 36912 24074 36964 24080
rect 36820 23860 36872 23866
rect 36820 23802 36872 23808
rect 36924 23798 36952 24074
rect 37108 24052 37136 27474
rect 37188 26240 37240 26246
rect 37188 26182 37240 26188
rect 37200 25498 37228 26182
rect 37188 25492 37240 25498
rect 37188 25434 37240 25440
rect 37188 25152 37240 25158
rect 37188 25094 37240 25100
rect 37200 24206 37228 25094
rect 37188 24200 37240 24206
rect 37188 24142 37240 24148
rect 37016 24024 37136 24052
rect 36912 23792 36964 23798
rect 36912 23734 36964 23740
rect 36728 23656 36780 23662
rect 36728 23598 36780 23604
rect 36820 23112 36872 23118
rect 36820 23054 36872 23060
rect 36728 22976 36780 22982
rect 36728 22918 36780 22924
rect 36740 22710 36768 22918
rect 36728 22704 36780 22710
rect 36728 22646 36780 22652
rect 36832 22642 36860 23054
rect 36820 22636 36872 22642
rect 36820 22578 36872 22584
rect 36832 21690 36860 22578
rect 36820 21684 36872 21690
rect 36820 21626 36872 21632
rect 36912 21548 36964 21554
rect 37016 21536 37044 24024
rect 36964 21508 37044 21536
rect 37096 21548 37148 21554
rect 36912 21490 36964 21496
rect 37096 21490 37148 21496
rect 36924 21078 36952 21490
rect 36912 21072 36964 21078
rect 36912 21014 36964 21020
rect 36820 21004 36872 21010
rect 36820 20946 36872 20952
rect 36832 20534 36860 20946
rect 36912 20936 36964 20942
rect 36912 20878 36964 20884
rect 36924 20534 36952 20878
rect 37108 20602 37136 21490
rect 37200 21146 37228 24142
rect 37292 22438 37320 28455
rect 37280 22432 37332 22438
rect 37280 22374 37332 22380
rect 37384 22094 37412 35022
rect 38292 32904 38344 32910
rect 38292 32846 38344 32852
rect 37740 32768 37792 32774
rect 38304 32745 38332 32846
rect 37740 32710 37792 32716
rect 38290 32736 38346 32745
rect 37752 32366 37780 32710
rect 38290 32671 38346 32680
rect 37740 32360 37792 32366
rect 37740 32302 37792 32308
rect 37556 30388 37608 30394
rect 37556 30330 37608 30336
rect 37292 22066 37412 22094
rect 37188 21140 37240 21146
rect 37188 21082 37240 21088
rect 37188 20936 37240 20942
rect 37188 20878 37240 20884
rect 37096 20596 37148 20602
rect 37096 20538 37148 20544
rect 36820 20528 36872 20534
rect 36820 20470 36872 20476
rect 36912 20528 36964 20534
rect 36912 20470 36964 20476
rect 37200 20262 37228 20878
rect 37188 20256 37240 20262
rect 37188 20198 37240 20204
rect 34796 20052 34848 20058
rect 34796 19994 34848 20000
rect 35348 20052 35400 20058
rect 35348 19994 35400 20000
rect 36084 20052 36136 20058
rect 36084 19994 36136 20000
rect 36544 20052 36596 20058
rect 36544 19994 36596 20000
rect 36636 20052 36688 20058
rect 36636 19994 36688 20000
rect 35164 19984 35216 19990
rect 35164 19926 35216 19932
rect 35072 19848 35124 19854
rect 35072 19790 35124 19796
rect 35084 19514 35112 19790
rect 35176 19514 35204 19926
rect 35256 19916 35308 19922
rect 35256 19858 35308 19864
rect 35268 19514 35296 19858
rect 35072 19508 35124 19514
rect 35072 19450 35124 19456
rect 35164 19508 35216 19514
rect 35164 19450 35216 19456
rect 35256 19508 35308 19514
rect 35256 19450 35308 19456
rect 33876 19372 33928 19378
rect 34428 19372 34480 19378
rect 33876 19314 33928 19320
rect 34348 19332 34428 19360
rect 33508 18896 33560 18902
rect 33508 18838 33560 18844
rect 33784 18896 33836 18902
rect 33784 18838 33836 18844
rect 33520 18766 33548 18838
rect 33692 18828 33744 18834
rect 33692 18770 33744 18776
rect 33416 18760 33468 18766
rect 33416 18702 33468 18708
rect 33508 18760 33560 18766
rect 33508 18702 33560 18708
rect 33232 18692 33284 18698
rect 33232 18634 33284 18640
rect 33244 18426 33272 18634
rect 33232 18420 33284 18426
rect 33232 18362 33284 18368
rect 32220 18284 32272 18290
rect 32220 18226 32272 18232
rect 32312 18284 32364 18290
rect 33152 18278 33364 18306
rect 32312 18226 32364 18232
rect 31024 18216 31076 18222
rect 31024 18158 31076 18164
rect 30840 17740 30892 17746
rect 30840 17682 30892 17688
rect 30748 16788 30800 16794
rect 30748 16730 30800 16736
rect 30852 16538 30880 17682
rect 30932 16992 30984 16998
rect 30932 16934 30984 16940
rect 30944 16794 30972 16934
rect 30932 16788 30984 16794
rect 30932 16730 30984 16736
rect 30852 16510 30972 16538
rect 30746 16280 30802 16289
rect 30746 16215 30802 16224
rect 30564 16040 30616 16046
rect 30564 15982 30616 15988
rect 30656 16040 30708 16046
rect 30656 15982 30708 15988
rect 30576 15706 30604 15982
rect 30564 15700 30616 15706
rect 30564 15642 30616 15648
rect 30564 15496 30616 15502
rect 30564 15438 30616 15444
rect 30576 15162 30604 15438
rect 30564 15156 30616 15162
rect 30564 15098 30616 15104
rect 30472 15020 30524 15026
rect 30472 14962 30524 14968
rect 30196 14544 30248 14550
rect 30196 14486 30248 14492
rect 30288 14408 30340 14414
rect 30668 14362 30696 15982
rect 30288 14350 30340 14356
rect 30300 13462 30328 14350
rect 30576 14334 30696 14362
rect 30380 13796 30432 13802
rect 30380 13738 30432 13744
rect 30288 13456 30340 13462
rect 30392 13433 30420 13738
rect 30288 13398 30340 13404
rect 30378 13424 30434 13433
rect 30378 13359 30434 13368
rect 30472 13388 30524 13394
rect 30472 13330 30524 13336
rect 30104 13320 30156 13326
rect 30104 13262 30156 13268
rect 30288 13320 30340 13326
rect 30288 13262 30340 13268
rect 30116 12850 30144 13262
rect 30300 12986 30328 13262
rect 30288 12980 30340 12986
rect 30288 12922 30340 12928
rect 30104 12844 30156 12850
rect 30104 12786 30156 12792
rect 30288 12640 30340 12646
rect 30288 12582 30340 12588
rect 30300 12434 30328 12582
rect 30208 12406 30328 12434
rect 30012 11892 30064 11898
rect 30012 11834 30064 11840
rect 29828 11756 29880 11762
rect 29828 11698 29880 11704
rect 29920 11756 29972 11762
rect 29920 11698 29972 11704
rect 30208 11694 30236 12406
rect 30288 12164 30340 12170
rect 30288 12106 30340 12112
rect 30300 11898 30328 12106
rect 30288 11892 30340 11898
rect 30288 11834 30340 11840
rect 30288 11756 30340 11762
rect 30288 11698 30340 11704
rect 30196 11688 30248 11694
rect 30196 11630 30248 11636
rect 29736 11144 29788 11150
rect 29736 11086 29788 11092
rect 29828 11144 29880 11150
rect 29828 11086 29880 11092
rect 29552 10668 29604 10674
rect 29552 10610 29604 10616
rect 29644 10668 29696 10674
rect 29644 10610 29696 10616
rect 29460 10532 29512 10538
rect 29460 10474 29512 10480
rect 29368 9648 29420 9654
rect 29368 9590 29420 9596
rect 29472 9586 29500 10474
rect 29564 10198 29592 10610
rect 29552 10192 29604 10198
rect 29552 10134 29604 10140
rect 29564 9926 29592 10134
rect 29552 9920 29604 9926
rect 29552 9862 29604 9868
rect 29460 9580 29512 9586
rect 29460 9522 29512 9528
rect 29550 9480 29606 9489
rect 29550 9415 29606 9424
rect 29564 8974 29592 9415
rect 29552 8968 29604 8974
rect 29552 8910 29604 8916
rect 29366 8120 29422 8129
rect 29366 8055 29422 8064
rect 29184 6792 29236 6798
rect 29184 6734 29236 6740
rect 29092 4752 29144 4758
rect 29092 4694 29144 4700
rect 28540 4480 28592 4486
rect 28540 4422 28592 4428
rect 27712 3528 27764 3534
rect 27712 3470 27764 3476
rect 28264 3528 28316 3534
rect 28264 3470 28316 3476
rect 27344 3188 27396 3194
rect 27344 3130 27396 3136
rect 28552 3126 28580 4422
rect 29104 3942 29132 4694
rect 29092 3936 29144 3942
rect 29092 3878 29144 3884
rect 29380 3738 29408 8055
rect 29656 7886 29684 10610
rect 29748 10266 29776 11086
rect 29840 10810 29868 11086
rect 29828 10804 29880 10810
rect 29828 10746 29880 10752
rect 30012 10668 30064 10674
rect 30012 10610 30064 10616
rect 29736 10260 29788 10266
rect 29736 10202 29788 10208
rect 29736 10124 29788 10130
rect 29736 10066 29788 10072
rect 29748 8090 29776 10066
rect 29920 9580 29972 9586
rect 29920 9522 29972 9528
rect 29932 9450 29960 9522
rect 29920 9444 29972 9450
rect 29920 9386 29972 9392
rect 29826 9344 29882 9353
rect 29932 9330 29960 9386
rect 29882 9302 29960 9330
rect 29826 9279 29882 9288
rect 29920 8968 29972 8974
rect 29920 8910 29972 8916
rect 29932 8634 29960 8910
rect 29920 8628 29972 8634
rect 29920 8570 29972 8576
rect 29736 8084 29788 8090
rect 29736 8026 29788 8032
rect 30024 7970 30052 10610
rect 30104 9648 30156 9654
rect 30104 9590 30156 9596
rect 30116 9178 30144 9590
rect 30300 9586 30328 11698
rect 30484 11642 30512 13330
rect 30576 13326 30604 14334
rect 30656 14272 30708 14278
rect 30656 14214 30708 14220
rect 30668 13462 30696 14214
rect 30656 13456 30708 13462
rect 30656 13398 30708 13404
rect 30564 13320 30616 13326
rect 30564 13262 30616 13268
rect 30392 11626 30512 11642
rect 30380 11620 30512 11626
rect 30432 11614 30512 11620
rect 30380 11562 30432 11568
rect 30392 11218 30420 11562
rect 30576 11286 30604 13262
rect 30564 11280 30616 11286
rect 30564 11222 30616 11228
rect 30380 11212 30432 11218
rect 30380 11154 30432 11160
rect 30668 10130 30696 13398
rect 30760 13376 30788 16215
rect 30840 15496 30892 15502
rect 30840 15438 30892 15444
rect 30852 15162 30880 15438
rect 30840 15156 30892 15162
rect 30840 15098 30892 15104
rect 30760 13348 30880 13376
rect 30748 13252 30800 13258
rect 30748 13194 30800 13200
rect 30760 11218 30788 13194
rect 30852 12306 30880 13348
rect 30840 12300 30892 12306
rect 30840 12242 30892 12248
rect 30748 11212 30800 11218
rect 30748 11154 30800 11160
rect 30840 11144 30892 11150
rect 30840 11086 30892 11092
rect 30380 10124 30432 10130
rect 30380 10066 30432 10072
rect 30656 10124 30708 10130
rect 30656 10066 30708 10072
rect 30288 9580 30340 9586
rect 30288 9522 30340 9528
rect 30300 9217 30328 9522
rect 30286 9208 30342 9217
rect 30104 9172 30156 9178
rect 30286 9143 30342 9152
rect 30104 9114 30156 9120
rect 30196 8968 30248 8974
rect 30196 8910 30248 8916
rect 30208 8634 30236 8910
rect 30196 8628 30248 8634
rect 30196 8570 30248 8576
rect 29932 7942 30052 7970
rect 29644 7880 29696 7886
rect 29644 7822 29696 7828
rect 29552 7404 29604 7410
rect 29552 7346 29604 7352
rect 29564 6662 29592 7346
rect 29656 7342 29684 7822
rect 29736 7744 29788 7750
rect 29736 7686 29788 7692
rect 29644 7336 29696 7342
rect 29644 7278 29696 7284
rect 29552 6656 29604 6662
rect 29552 6598 29604 6604
rect 29644 5704 29696 5710
rect 29644 5646 29696 5652
rect 29656 5370 29684 5646
rect 29644 5364 29696 5370
rect 29644 5306 29696 5312
rect 29460 4480 29512 4486
rect 29460 4422 29512 4428
rect 29472 4214 29500 4422
rect 29748 4282 29776 7686
rect 29932 7478 29960 7942
rect 30012 7880 30064 7886
rect 30012 7822 30064 7828
rect 30024 7546 30052 7822
rect 30012 7540 30064 7546
rect 30012 7482 30064 7488
rect 29920 7472 29972 7478
rect 29920 7414 29972 7420
rect 29828 7404 29880 7410
rect 29828 7346 29880 7352
rect 30104 7404 30156 7410
rect 30104 7346 30156 7352
rect 29840 7274 29868 7346
rect 29828 7268 29880 7274
rect 29828 7210 29880 7216
rect 29840 6934 29868 7210
rect 30116 7206 30144 7346
rect 30104 7200 30156 7206
rect 30104 7142 30156 7148
rect 29828 6928 29880 6934
rect 29828 6870 29880 6876
rect 29828 6656 29880 6662
rect 29828 6598 29880 6604
rect 29840 6458 29868 6598
rect 29828 6452 29880 6458
rect 29828 6394 29880 6400
rect 30196 6316 30248 6322
rect 30196 6258 30248 6264
rect 30012 6112 30064 6118
rect 30012 6054 30064 6060
rect 30024 5778 30052 6054
rect 30012 5772 30064 5778
rect 30012 5714 30064 5720
rect 30208 5370 30236 6258
rect 30196 5364 30248 5370
rect 30196 5306 30248 5312
rect 30392 5250 30420 10066
rect 30472 9376 30524 9382
rect 30472 9318 30524 9324
rect 30484 9042 30512 9318
rect 30852 9178 30880 11086
rect 30840 9172 30892 9178
rect 30840 9114 30892 9120
rect 30472 9036 30524 9042
rect 30472 8978 30524 8984
rect 30564 8900 30616 8906
rect 30564 8842 30616 8848
rect 30576 8090 30604 8842
rect 30564 8084 30616 8090
rect 30564 8026 30616 8032
rect 30852 7954 30880 9114
rect 30944 8566 30972 16510
rect 31036 12170 31064 18158
rect 31208 17672 31260 17678
rect 31208 17614 31260 17620
rect 31116 16448 31168 16454
rect 31116 16390 31168 16396
rect 31128 15026 31156 16390
rect 31116 15020 31168 15026
rect 31116 14962 31168 14968
rect 31116 14816 31168 14822
rect 31116 14758 31168 14764
rect 31128 13190 31156 14758
rect 31116 13184 31168 13190
rect 31116 13126 31168 13132
rect 31024 12164 31076 12170
rect 31024 12106 31076 12112
rect 31036 10810 31064 12106
rect 31128 11150 31156 13126
rect 31116 11144 31168 11150
rect 31116 11086 31168 11092
rect 31024 10804 31076 10810
rect 31024 10746 31076 10752
rect 30932 8560 30984 8566
rect 30932 8502 30984 8508
rect 30944 8090 30972 8502
rect 30932 8084 30984 8090
rect 30932 8026 30984 8032
rect 30840 7948 30892 7954
rect 30840 7890 30892 7896
rect 30472 7880 30524 7886
rect 30472 7822 30524 7828
rect 30484 7546 30512 7822
rect 30472 7540 30524 7546
rect 30472 7482 30524 7488
rect 30472 6724 30524 6730
rect 30472 6666 30524 6672
rect 30484 5370 30512 6666
rect 31024 5704 31076 5710
rect 31024 5646 31076 5652
rect 30472 5364 30524 5370
rect 30472 5306 30524 5312
rect 30300 5234 30420 5250
rect 30288 5228 30420 5234
rect 30340 5222 30420 5228
rect 30288 5170 30340 5176
rect 29736 4276 29788 4282
rect 29736 4218 29788 4224
rect 31036 4214 31064 5646
rect 29460 4208 29512 4214
rect 29460 4150 29512 4156
rect 31024 4208 31076 4214
rect 31024 4150 31076 4156
rect 29368 3732 29420 3738
rect 29368 3674 29420 3680
rect 31220 3602 31248 17614
rect 31300 17604 31352 17610
rect 31300 17546 31352 17552
rect 31312 13954 31340 17546
rect 32232 17134 32260 18226
rect 32220 17128 32272 17134
rect 32220 17070 32272 17076
rect 32232 16794 32260 17070
rect 32220 16788 32272 16794
rect 32220 16730 32272 16736
rect 32324 16538 32352 18226
rect 33140 18148 33192 18154
rect 33140 18090 33192 18096
rect 33152 17202 33180 18090
rect 33140 17196 33192 17202
rect 33140 17138 33192 17144
rect 33232 17196 33284 17202
rect 33232 17138 33284 17144
rect 33048 16992 33100 16998
rect 33048 16934 33100 16940
rect 33060 16658 33088 16934
rect 33048 16652 33100 16658
rect 33048 16594 33100 16600
rect 32140 16510 32352 16538
rect 32680 16584 32732 16590
rect 32680 16526 32732 16532
rect 32034 16280 32090 16289
rect 32034 16215 32090 16224
rect 32048 16114 32076 16215
rect 32036 16108 32088 16114
rect 32036 16050 32088 16056
rect 31668 15020 31720 15026
rect 31668 14962 31720 14968
rect 31392 14340 31444 14346
rect 31392 14282 31444 14288
rect 31404 14074 31432 14282
rect 31392 14068 31444 14074
rect 31392 14010 31444 14016
rect 31312 13926 31432 13954
rect 31300 13796 31352 13802
rect 31300 13738 31352 13744
rect 31312 12782 31340 13738
rect 31300 12776 31352 12782
rect 31300 12718 31352 12724
rect 31404 12730 31432 13926
rect 31484 13320 31536 13326
rect 31484 13262 31536 13268
rect 31496 12918 31524 13262
rect 31484 12912 31536 12918
rect 31484 12854 31536 12860
rect 31404 12702 31524 12730
rect 31392 12640 31444 12646
rect 31392 12582 31444 12588
rect 31300 12436 31352 12442
rect 31300 12378 31352 12384
rect 31312 11762 31340 12378
rect 31404 12374 31432 12582
rect 31392 12368 31444 12374
rect 31392 12310 31444 12316
rect 31300 11756 31352 11762
rect 31300 11698 31352 11704
rect 31496 11234 31524 12702
rect 31680 12170 31708 14962
rect 31944 13320 31996 13326
rect 31944 13262 31996 13268
rect 31956 12986 31984 13262
rect 32036 13184 32088 13190
rect 32036 13126 32088 13132
rect 32048 12986 32076 13126
rect 31944 12980 31996 12986
rect 31944 12922 31996 12928
rect 32036 12980 32088 12986
rect 32036 12922 32088 12928
rect 31668 12164 31720 12170
rect 31668 12106 31720 12112
rect 31404 11206 31524 11234
rect 31300 10464 31352 10470
rect 31300 10406 31352 10412
rect 31312 10130 31340 10406
rect 31300 10124 31352 10130
rect 31300 10066 31352 10072
rect 31300 9988 31352 9994
rect 31300 9930 31352 9936
rect 31312 9518 31340 9930
rect 31300 9512 31352 9518
rect 31300 9454 31352 9460
rect 31404 7546 31432 11206
rect 31576 10804 31628 10810
rect 31576 10746 31628 10752
rect 31588 9994 31616 10746
rect 31680 10441 31708 12106
rect 31666 10432 31722 10441
rect 31666 10367 31722 10376
rect 31576 9988 31628 9994
rect 31576 9930 31628 9936
rect 31588 9110 31616 9930
rect 31576 9104 31628 9110
rect 31576 9046 31628 9052
rect 31588 7698 31616 9046
rect 31680 8634 31708 10367
rect 31852 10124 31904 10130
rect 31852 10066 31904 10072
rect 31668 8628 31720 8634
rect 31668 8570 31720 8576
rect 31864 8498 31892 10066
rect 31944 9512 31996 9518
rect 31944 9454 31996 9460
rect 31956 9178 31984 9454
rect 31944 9172 31996 9178
rect 31944 9114 31996 9120
rect 31852 8492 31904 8498
rect 31852 8434 31904 8440
rect 31668 8288 31720 8294
rect 31668 8230 31720 8236
rect 31680 7818 31708 8230
rect 31864 7886 31892 8434
rect 31852 7880 31904 7886
rect 31852 7822 31904 7828
rect 31668 7812 31720 7818
rect 31668 7754 31720 7760
rect 31496 7670 31616 7698
rect 31392 7540 31444 7546
rect 31392 7482 31444 7488
rect 31496 5914 31524 7670
rect 31576 7540 31628 7546
rect 31576 7482 31628 7488
rect 31484 5908 31536 5914
rect 31484 5850 31536 5856
rect 31484 5704 31536 5710
rect 31484 5646 31536 5652
rect 31392 5568 31444 5574
rect 31392 5510 31444 5516
rect 31404 5370 31432 5510
rect 31496 5370 31524 5646
rect 31392 5364 31444 5370
rect 31392 5306 31444 5312
rect 31484 5364 31536 5370
rect 31484 5306 31536 5312
rect 31588 5030 31616 7482
rect 31680 7410 31708 7754
rect 32036 7472 32088 7478
rect 32036 7414 32088 7420
rect 31668 7404 31720 7410
rect 31668 7346 31720 7352
rect 31944 7200 31996 7206
rect 31944 7142 31996 7148
rect 31956 6798 31984 7142
rect 31944 6792 31996 6798
rect 31944 6734 31996 6740
rect 32048 5642 32076 7414
rect 31760 5636 31812 5642
rect 31760 5578 31812 5584
rect 32036 5636 32088 5642
rect 32036 5578 32088 5584
rect 31772 5098 31800 5578
rect 32048 5370 32076 5578
rect 32036 5364 32088 5370
rect 32036 5306 32088 5312
rect 31760 5092 31812 5098
rect 31760 5034 31812 5040
rect 31576 5024 31628 5030
rect 31576 4966 31628 4972
rect 31208 3596 31260 3602
rect 31208 3538 31260 3544
rect 27160 3120 27212 3126
rect 27160 3062 27212 3068
rect 28540 3120 28592 3126
rect 28540 3062 28592 3068
rect 26700 3052 26752 3058
rect 26700 2994 26752 3000
rect 31024 3052 31076 3058
rect 31024 2994 31076 3000
rect 26332 2916 26384 2922
rect 26332 2858 26384 2864
rect 26516 2916 26568 2922
rect 26516 2858 26568 2864
rect 26424 2848 26476 2854
rect 26476 2796 26740 2802
rect 26424 2790 26740 2796
rect 26436 2774 26740 2790
rect 25240 2746 25360 2774
rect 24674 2615 24730 2624
rect 25136 2644 25188 2650
rect 19800 2586 19852 2592
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 16212 2508 16264 2514
rect 16212 2450 16264 2456
rect 19708 2508 19760 2514
rect 19708 2450 19760 2456
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 2044 2372 2096 2378
rect 2044 2314 2096 2320
rect 3976 2372 4028 2378
rect 3976 2314 4028 2320
rect 6552 2372 6604 2378
rect 6552 2314 6604 2320
rect 1490 2136 1546 2145
rect 1490 2071 1546 2080
rect 2056 1170 2084 2314
rect 3988 1170 4016 2314
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 6564 1170 6592 2314
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 11164 1442 11192 2246
rect 1964 1142 2084 1170
rect 3896 1142 4016 1170
rect 6472 1142 6592 1170
rect 10980 1414 11192 1442
rect 1964 800 1992 1142
rect 3896 800 3924 1142
rect 6472 800 6500 1142
rect 10980 800 11008 1414
rect 13004 1306 13032 2382
rect 14384 2378 14412 2450
rect 24688 2446 24716 2615
rect 25136 2586 25188 2592
rect 25240 2514 25268 2746
rect 25228 2508 25280 2514
rect 25228 2450 25280 2456
rect 26712 2446 26740 2774
rect 31036 2582 31064 2994
rect 31220 2774 31248 3538
rect 32140 3058 32168 16510
rect 32692 16250 32720 16526
rect 33244 16250 33272 17138
rect 33336 16250 33364 18278
rect 33428 18154 33456 18702
rect 33520 18290 33548 18702
rect 33508 18284 33560 18290
rect 33508 18226 33560 18232
rect 33704 18222 33732 18770
rect 33888 18426 33916 19314
rect 34348 18970 34376 19332
rect 34428 19314 34480 19320
rect 34612 19372 34664 19378
rect 34612 19314 34664 19320
rect 34336 18964 34388 18970
rect 34336 18906 34388 18912
rect 34060 18896 34112 18902
rect 34060 18838 34112 18844
rect 34072 18766 34100 18838
rect 34060 18760 34112 18766
rect 34060 18702 34112 18708
rect 33876 18420 33928 18426
rect 33876 18362 33928 18368
rect 34348 18222 34376 18906
rect 34624 18902 34652 19314
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35360 18970 35388 19994
rect 35992 19848 36044 19854
rect 35992 19790 36044 19796
rect 35440 19712 35492 19718
rect 35440 19654 35492 19660
rect 35452 19378 35480 19654
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 35440 19372 35492 19378
rect 35440 19314 35492 19320
rect 36004 19310 36032 19790
rect 35992 19304 36044 19310
rect 35992 19246 36044 19252
rect 35348 18964 35400 18970
rect 35348 18906 35400 18912
rect 34612 18896 34664 18902
rect 34612 18838 34664 18844
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 37292 18222 37320 22066
rect 37372 18760 37424 18766
rect 37372 18702 37424 18708
rect 33692 18216 33744 18222
rect 33692 18158 33744 18164
rect 34336 18216 34388 18222
rect 34336 18158 34388 18164
rect 37280 18216 37332 18222
rect 37280 18158 37332 18164
rect 33416 18148 33468 18154
rect 33416 18090 33468 18096
rect 32680 16244 32732 16250
rect 32680 16186 32732 16192
rect 33232 16244 33284 16250
rect 33232 16186 33284 16192
rect 33324 16244 33376 16250
rect 33324 16186 33376 16192
rect 33140 16108 33192 16114
rect 33140 16050 33192 16056
rect 32404 15496 32456 15502
rect 32404 15438 32456 15444
rect 32416 15026 32444 15438
rect 32588 15360 32640 15366
rect 32588 15302 32640 15308
rect 32404 15020 32456 15026
rect 32404 14962 32456 14968
rect 32600 14958 32628 15302
rect 33048 15020 33100 15026
rect 33048 14962 33100 14968
rect 32588 14952 32640 14958
rect 32588 14894 32640 14900
rect 33060 14618 33088 14962
rect 32496 14612 32548 14618
rect 32496 14554 32548 14560
rect 33048 14612 33100 14618
rect 33048 14554 33100 14560
rect 32508 14074 32536 14554
rect 33152 14482 33180 16050
rect 33508 15564 33560 15570
rect 33508 15506 33560 15512
rect 33324 15360 33376 15366
rect 33324 15302 33376 15308
rect 33336 14958 33364 15302
rect 33324 14952 33376 14958
rect 33324 14894 33376 14900
rect 33520 14804 33548 15506
rect 33600 14816 33652 14822
rect 33520 14776 33600 14804
rect 33140 14476 33192 14482
rect 33140 14418 33192 14424
rect 33324 14476 33376 14482
rect 33324 14418 33376 14424
rect 32496 14068 32548 14074
rect 32496 14010 32548 14016
rect 32680 13728 32732 13734
rect 32680 13670 32732 13676
rect 32312 13184 32364 13190
rect 32312 13126 32364 13132
rect 32324 12986 32352 13126
rect 32312 12980 32364 12986
rect 32312 12922 32364 12928
rect 32496 11008 32548 11014
rect 32496 10950 32548 10956
rect 32508 10674 32536 10950
rect 32588 10736 32640 10742
rect 32588 10678 32640 10684
rect 32496 10668 32548 10674
rect 32496 10610 32548 10616
rect 32508 10266 32536 10610
rect 32600 10606 32628 10678
rect 32692 10606 32720 13670
rect 32588 10600 32640 10606
rect 32588 10542 32640 10548
rect 32680 10600 32732 10606
rect 32680 10542 32732 10548
rect 32496 10260 32548 10266
rect 32496 10202 32548 10208
rect 32600 9450 32628 10542
rect 33152 10062 33180 14418
rect 33232 13252 33284 13258
rect 33232 13194 33284 13200
rect 33244 10606 33272 13194
rect 33336 12434 33364 14418
rect 33520 14346 33548 14776
rect 33600 14758 33652 14764
rect 33508 14340 33560 14346
rect 33508 14282 33560 14288
rect 33704 14226 33732 18158
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 37384 17882 37412 18702
rect 37568 18306 37596 30330
rect 37648 21548 37700 21554
rect 37648 21490 37700 21496
rect 37660 18970 37688 21490
rect 37832 21344 37884 21350
rect 37832 21286 37884 21292
rect 37844 21185 37872 21286
rect 37830 21176 37886 21185
rect 37830 21111 37886 21120
rect 38292 19372 38344 19378
rect 38292 19314 38344 19320
rect 37740 19168 37792 19174
rect 38304 19145 38332 19314
rect 37740 19110 37792 19116
rect 38290 19136 38346 19145
rect 37648 18964 37700 18970
rect 37648 18906 37700 18912
rect 37568 18278 37688 18306
rect 37372 17876 37424 17882
rect 37372 17818 37424 17824
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 33968 17128 34020 17134
rect 33968 17070 34020 17076
rect 33980 16522 34008 17070
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 33968 16516 34020 16522
rect 33968 16458 34020 16464
rect 33784 16244 33836 16250
rect 33784 16186 33836 16192
rect 33796 14278 33824 16186
rect 33876 16040 33928 16046
rect 33876 15982 33928 15988
rect 33520 14198 33732 14226
rect 33784 14272 33836 14278
rect 33784 14214 33836 14220
rect 33336 12406 33456 12434
rect 33428 12306 33456 12406
rect 33416 12300 33468 12306
rect 33416 12242 33468 12248
rect 33232 10600 33284 10606
rect 33232 10542 33284 10548
rect 33324 10600 33376 10606
rect 33324 10542 33376 10548
rect 33140 10056 33192 10062
rect 33140 9998 33192 10004
rect 32772 9920 32824 9926
rect 32772 9862 32824 9868
rect 32784 9586 32812 9862
rect 32772 9580 32824 9586
rect 32772 9522 32824 9528
rect 32588 9444 32640 9450
rect 32588 9386 32640 9392
rect 32404 9376 32456 9382
rect 32404 9318 32456 9324
rect 32772 9376 32824 9382
rect 32772 9318 32824 9324
rect 32416 9178 32444 9318
rect 32404 9172 32456 9178
rect 32404 9114 32456 9120
rect 32680 8968 32732 8974
rect 32680 8910 32732 8916
rect 32692 8634 32720 8910
rect 32680 8628 32732 8634
rect 32680 8570 32732 8576
rect 32784 8514 32812 9318
rect 32692 8486 32812 8514
rect 32312 7744 32364 7750
rect 32312 7686 32364 7692
rect 32324 7546 32352 7686
rect 32312 7540 32364 7546
rect 32312 7482 32364 7488
rect 32404 7336 32456 7342
rect 32404 7278 32456 7284
rect 32416 7002 32444 7278
rect 32404 6996 32456 7002
rect 32404 6938 32456 6944
rect 32692 5166 32720 8486
rect 33244 7818 33272 10542
rect 33336 9722 33364 10542
rect 33324 9716 33376 9722
rect 33324 9658 33376 9664
rect 33324 9512 33376 9518
rect 33428 9500 33456 12242
rect 33520 9654 33548 14198
rect 33796 14074 33824 14214
rect 33784 14068 33836 14074
rect 33784 14010 33836 14016
rect 33600 13864 33652 13870
rect 33600 13806 33652 13812
rect 33612 13394 33640 13806
rect 33888 13394 33916 15982
rect 33980 15434 34008 16458
rect 34428 16448 34480 16454
rect 34428 16390 34480 16396
rect 34440 16250 34468 16390
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 34428 16244 34480 16250
rect 34428 16186 34480 16192
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 33968 15428 34020 15434
rect 33968 15370 34020 15376
rect 33980 15162 34008 15370
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 33968 15156 34020 15162
rect 33968 15098 34020 15104
rect 33980 14482 34008 15098
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 33968 14476 34020 14482
rect 33968 14418 34020 14424
rect 33980 13938 34008 14418
rect 37660 14414 37688 18278
rect 37752 17270 37780 19110
rect 38290 19071 38346 19080
rect 37740 17264 37792 17270
rect 37740 17206 37792 17212
rect 38292 14544 38344 14550
rect 38292 14486 38344 14492
rect 37648 14408 37700 14414
rect 38304 14385 38332 14486
rect 37648 14350 37700 14356
rect 38290 14376 38346 14385
rect 38290 14311 38346 14320
rect 35440 14272 35492 14278
rect 35440 14214 35492 14220
rect 35452 14074 35480 14214
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 35440 14068 35492 14074
rect 35440 14010 35492 14016
rect 33968 13932 34020 13938
rect 33968 13874 34020 13880
rect 33600 13388 33652 13394
rect 33600 13330 33652 13336
rect 33876 13388 33928 13394
rect 33876 13330 33928 13336
rect 33692 13184 33744 13190
rect 33692 13126 33744 13132
rect 33598 12744 33654 12753
rect 33598 12679 33654 12688
rect 33612 12170 33640 12679
rect 33704 12374 33732 13126
rect 33980 12850 34008 13874
rect 34060 13728 34112 13734
rect 34060 13670 34112 13676
rect 34072 13530 34100 13670
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34060 13524 34112 13530
rect 34060 13466 34112 13472
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 33968 12844 34020 12850
rect 33968 12786 34020 12792
rect 33980 12434 34008 12786
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 33980 12406 34100 12434
rect 33692 12368 33744 12374
rect 33692 12310 33744 12316
rect 33600 12164 33652 12170
rect 33600 12106 33652 12112
rect 33612 11694 33640 12106
rect 34072 11830 34100 12406
rect 37646 12336 37702 12345
rect 37646 12271 37702 12280
rect 34152 12096 34204 12102
rect 34152 12038 34204 12044
rect 34520 12096 34572 12102
rect 34520 12038 34572 12044
rect 34164 11898 34192 12038
rect 34152 11892 34204 11898
rect 34152 11834 34204 11840
rect 34532 11830 34560 12038
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 34060 11824 34112 11830
rect 34060 11766 34112 11772
rect 34520 11824 34572 11830
rect 34520 11766 34572 11772
rect 37660 11762 37688 12271
rect 37648 11756 37700 11762
rect 37648 11698 37700 11704
rect 33600 11688 33652 11694
rect 33600 11630 33652 11636
rect 37830 11656 37886 11665
rect 37830 11591 37832 11600
rect 37884 11591 37886 11600
rect 37832 11562 37884 11568
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 34520 10464 34572 10470
rect 34520 10406 34572 10412
rect 34532 9654 34560 10406
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35072 9920 35124 9926
rect 35072 9862 35124 9868
rect 33508 9648 33560 9654
rect 33508 9590 33560 9596
rect 34520 9648 34572 9654
rect 34520 9590 34572 9596
rect 33692 9580 33744 9586
rect 33692 9522 33744 9528
rect 33376 9472 33456 9500
rect 33324 9454 33376 9460
rect 33704 9042 33732 9522
rect 35084 9518 35112 9862
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 34428 9512 34480 9518
rect 34428 9454 34480 9460
rect 35072 9512 35124 9518
rect 35072 9454 35124 9460
rect 34440 9178 34468 9454
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34428 9172 34480 9178
rect 34428 9114 34480 9120
rect 33692 9036 33744 9042
rect 33692 8978 33744 8984
rect 33704 8906 33732 8978
rect 33692 8900 33744 8906
rect 33692 8842 33744 8848
rect 33232 7812 33284 7818
rect 33232 7754 33284 7760
rect 33704 7478 33732 8842
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 33692 7472 33744 7478
rect 33692 7414 33744 7420
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 32680 5160 32732 5166
rect 32680 5102 32732 5108
rect 32692 4758 32720 5102
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 32680 4752 32732 4758
rect 32680 4694 32732 4700
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 37464 3528 37516 3534
rect 37464 3470 37516 3476
rect 36912 3392 36964 3398
rect 36912 3334 36964 3340
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 36924 3058 36952 3334
rect 32128 3052 32180 3058
rect 32128 2994 32180 3000
rect 36912 3052 36964 3058
rect 36912 2994 36964 3000
rect 37280 2848 37332 2854
rect 37280 2790 37332 2796
rect 31128 2746 31248 2774
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 31024 2576 31076 2582
rect 31024 2518 31076 2524
rect 31128 2514 31156 2746
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 31116 2508 31168 2514
rect 31116 2450 31168 2456
rect 37292 2446 37320 2790
rect 24676 2440 24728 2446
rect 24676 2382 24728 2388
rect 26700 2440 26752 2446
rect 26700 2382 26752 2388
rect 31024 2440 31076 2446
rect 35532 2440 35584 2446
rect 31024 2382 31076 2388
rect 35452 2388 35532 2394
rect 37280 2440 37332 2446
rect 35452 2382 35584 2388
rect 35714 2408 35770 2417
rect 14372 2372 14424 2378
rect 15568 2372 15620 2378
rect 14372 2314 14424 2320
rect 15488 2332 15568 2360
rect 12912 1278 13032 1306
rect 12912 800 12940 1278
rect 15488 800 15516 2332
rect 15568 2314 15620 2320
rect 20260 2304 20312 2310
rect 24584 2304 24636 2310
rect 20260 2246 20312 2252
rect 24504 2264 24584 2292
rect 19996 870 20116 898
rect 19996 800 20024 870
rect 18 0 74 800
rect 1950 0 2006 800
rect 3882 0 3938 800
rect 6458 0 6514 800
rect 8390 0 8446 800
rect 10966 0 11022 800
rect 12898 0 12954 800
rect 15474 0 15530 800
rect 17406 0 17462 800
rect 19982 0 20038 800
rect 20088 762 20116 870
rect 20272 762 20300 2246
rect 24504 800 24532 2264
rect 24584 2246 24636 2252
rect 26424 2304 26476 2310
rect 26424 2246 26476 2252
rect 26436 800 26464 2246
rect 31036 1306 31064 2382
rect 30944 1278 31064 1306
rect 35452 2366 35572 2382
rect 30944 800 30972 1278
rect 35452 800 35480 2366
rect 37280 2382 37332 2388
rect 35714 2343 35770 2352
rect 35728 2310 35756 2343
rect 35716 2304 35768 2310
rect 35716 2246 35768 2252
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 37476 1850 37504 3470
rect 37832 2848 37884 2854
rect 37884 2796 37964 2802
rect 37832 2790 37964 2796
rect 37844 2774 37964 2790
rect 37740 2304 37792 2310
rect 37740 2246 37792 2252
rect 37752 2145 37780 2246
rect 37738 2136 37794 2145
rect 37738 2071 37794 2080
rect 37384 1822 37504 1850
rect 37384 800 37412 1822
rect 20088 734 20300 762
rect 21914 0 21970 800
rect 24490 0 24546 800
rect 26422 0 26478 800
rect 28998 0 29054 800
rect 30930 0 30986 800
rect 32862 0 32918 800
rect 35438 0 35494 800
rect 37370 0 37426 800
rect 37936 105 37964 2774
rect 37922 96 37978 105
rect 37922 31 37978 40
<< via2 >>
rect 1122 39480 1178 39536
rect 938 37440 994 37496
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 35600 39194 35656 39196
rect 35680 39194 35736 39196
rect 35760 39194 35816 39196
rect 35840 39194 35896 39196
rect 35600 39142 35646 39194
rect 35646 39142 35656 39194
rect 35680 39142 35710 39194
rect 35710 39142 35722 39194
rect 35722 39142 35736 39194
rect 35760 39142 35774 39194
rect 35774 39142 35786 39194
rect 35786 39142 35816 39194
rect 35840 39142 35850 39194
rect 35850 39142 35896 39194
rect 35600 39140 35656 39142
rect 35680 39140 35736 39142
rect 35760 39140 35816 39142
rect 35840 39140 35896 39142
rect 37186 40160 37242 40216
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 938 34720 994 34776
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 938 25900 994 25936
rect 938 25880 940 25900
rect 940 25880 992 25900
rect 992 25880 994 25900
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4618 29144 4674 29200
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 5078 29144 5134 29200
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 938 21120 994 21176
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 938 18400 994 18456
rect 938 16360 994 16416
rect 3146 20848 3202 20904
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 3146 19388 3148 19408
rect 3148 19388 3200 19408
rect 3200 19388 3202 19408
rect 3146 19352 3202 19388
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 6642 24792 6698 24848
rect 11610 35264 11666 35320
rect 6090 21548 6146 21584
rect 6090 21528 6092 21548
rect 6092 21528 6144 21548
rect 6144 21528 6146 21548
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 1490 13640 1546 13696
rect 938 11600 994 11656
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4066 11600 4122 11656
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 938 4120 994 4176
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 6918 23704 6974 23760
rect 11978 34720 12034 34776
rect 7470 24520 7526 24576
rect 7930 20476 7932 20496
rect 7932 20476 7984 20496
rect 7984 20476 7986 20496
rect 7930 20440 7986 20476
rect 8298 19780 8354 19816
rect 8298 19760 8300 19780
rect 8300 19760 8352 19780
rect 8352 19760 8354 19780
rect 8206 12416 8262 12472
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 8850 21956 8906 21992
rect 8850 21936 8852 21956
rect 8852 21936 8904 21956
rect 8904 21936 8906 21956
rect 12438 35808 12494 35864
rect 12990 35572 12992 35592
rect 12992 35572 13044 35592
rect 13044 35572 13046 35592
rect 12990 35536 13046 35572
rect 10414 21936 10470 21992
rect 10506 21392 10562 21448
rect 10414 17720 10470 17776
rect 10506 17312 10562 17368
rect 10966 19216 11022 19272
rect 10874 18944 10930 19000
rect 11150 17992 11206 18048
rect 11058 17212 11060 17232
rect 11060 17212 11112 17232
rect 11112 17212 11114 17232
rect 11058 17176 11114 17212
rect 11058 15000 11114 15056
rect 10874 13640 10930 13696
rect 10782 13232 10838 13288
rect 9126 4528 9182 4584
rect 10874 12416 10930 12472
rect 10138 8200 10194 8256
rect 11150 10684 11152 10704
rect 11152 10684 11204 10704
rect 11204 10684 11206 10704
rect 11150 10648 11206 10684
rect 11150 9560 11206 9616
rect 11242 9424 11298 9480
rect 11702 21392 11758 21448
rect 11610 19624 11666 19680
rect 11702 19080 11758 19136
rect 11518 14728 11574 14784
rect 11702 15136 11758 15192
rect 12162 29008 12218 29064
rect 12530 30368 12586 30424
rect 13726 31456 13782 31512
rect 13818 31048 13874 31104
rect 11978 21956 12034 21992
rect 11978 21936 11980 21956
rect 11980 21936 12032 21956
rect 12032 21936 12034 21956
rect 12346 20712 12402 20768
rect 12438 19216 12494 19272
rect 13174 25744 13230 25800
rect 12898 25356 12954 25392
rect 12898 25336 12900 25356
rect 12900 25336 12952 25356
rect 12952 25336 12954 25356
rect 13910 24520 13966 24576
rect 12070 15444 12072 15464
rect 12072 15444 12124 15464
rect 12124 15444 12126 15464
rect 12070 15408 12126 15444
rect 11426 9424 11482 9480
rect 11886 13368 11942 13424
rect 11978 12844 12034 12880
rect 11978 12824 11980 12844
rect 11980 12824 12032 12844
rect 12032 12824 12034 12844
rect 11794 10512 11850 10568
rect 11978 9424 12034 9480
rect 12070 9152 12126 9208
rect 12438 9288 12494 9344
rect 10966 3440 11022 3496
rect 11610 3848 11666 3904
rect 12622 10240 12678 10296
rect 12806 17332 12862 17368
rect 12806 17312 12808 17332
rect 12808 17312 12860 17332
rect 12860 17312 12862 17332
rect 13174 18264 13230 18320
rect 13082 10104 13138 10160
rect 13542 17060 13598 17096
rect 13542 17040 13544 17060
rect 13544 17040 13596 17060
rect 13596 17040 13598 17060
rect 14830 31204 14886 31240
rect 14830 31184 14832 31204
rect 14832 31184 14884 31204
rect 14884 31184 14886 31204
rect 15198 31084 15200 31104
rect 15200 31084 15252 31104
rect 15252 31084 15254 31104
rect 15198 31048 15254 31084
rect 14922 26288 14978 26344
rect 14554 25880 14610 25936
rect 15106 24656 15162 24712
rect 14554 23432 14610 23488
rect 14370 19624 14426 19680
rect 14278 19080 14334 19136
rect 14094 17992 14150 18048
rect 14554 21392 14610 21448
rect 14830 21392 14886 21448
rect 14646 19660 14648 19680
rect 14648 19660 14700 19680
rect 14700 19660 14702 19680
rect 14646 19624 14702 19660
rect 14370 16904 14426 16960
rect 15106 24520 15162 24576
rect 15382 24148 15384 24168
rect 15384 24148 15436 24168
rect 15436 24148 15438 24168
rect 15382 24112 15438 24148
rect 15566 31476 15622 31512
rect 15566 31456 15568 31476
rect 15568 31456 15620 31476
rect 15620 31456 15622 31476
rect 15566 30368 15622 30424
rect 16118 35536 16174 35592
rect 19338 35944 19394 36000
rect 16670 31184 16726 31240
rect 16854 26460 16856 26480
rect 16856 26460 16908 26480
rect 16908 26460 16910 26480
rect 16854 26424 16910 26460
rect 16394 25916 16396 25936
rect 16396 25916 16448 25936
rect 16448 25916 16450 25936
rect 16394 25880 16450 25916
rect 16118 23024 16174 23080
rect 13634 11736 13690 11792
rect 13358 10648 13414 10704
rect 12622 3848 12678 3904
rect 13818 11212 13874 11248
rect 13818 11192 13820 11212
rect 13820 11192 13872 11212
rect 13872 11192 13874 11212
rect 14186 12960 14242 13016
rect 13542 9288 13598 9344
rect 13726 9424 13782 9480
rect 13910 9596 13912 9616
rect 13912 9596 13964 9616
rect 13964 9596 13966 9616
rect 13910 9560 13966 9596
rect 14002 7248 14058 7304
rect 14554 13096 14610 13152
rect 14462 10920 14518 10976
rect 14554 10784 14610 10840
rect 14278 9832 14334 9888
rect 14002 6196 14004 6216
rect 14004 6196 14056 6216
rect 14056 6196 14058 6216
rect 14002 6160 14058 6196
rect 14370 4120 14426 4176
rect 14278 3984 14334 4040
rect 15014 11464 15070 11520
rect 14922 11192 14978 11248
rect 14922 9152 14978 9208
rect 15198 10512 15254 10568
rect 15658 19624 15714 19680
rect 15382 12436 15438 12472
rect 15382 12416 15384 12436
rect 15384 12416 15436 12436
rect 15436 12416 15438 12436
rect 15382 12280 15438 12336
rect 16762 24148 16764 24168
rect 16764 24148 16816 24168
rect 16816 24148 16818 24168
rect 16762 24112 16818 24148
rect 16302 18944 16358 19000
rect 15658 11600 15714 11656
rect 15566 11092 15568 11112
rect 15568 11092 15620 11112
rect 15620 11092 15622 11112
rect 15566 11056 15622 11092
rect 15474 10648 15530 10704
rect 17038 22092 17094 22128
rect 17038 22072 17040 22092
rect 17040 22072 17092 22092
rect 17092 22072 17094 22092
rect 17038 21800 17094 21856
rect 17498 30776 17554 30832
rect 17498 25236 17500 25256
rect 17500 25236 17552 25256
rect 17552 25236 17554 25256
rect 17498 25200 17554 25236
rect 16486 19796 16488 19816
rect 16488 19796 16540 19816
rect 16540 19796 16542 19816
rect 16486 19760 16542 19796
rect 16946 19624 17002 19680
rect 16394 18264 16450 18320
rect 16302 18128 16358 18184
rect 15842 12164 15898 12200
rect 15842 12144 15844 12164
rect 15844 12144 15896 12164
rect 15896 12144 15898 12164
rect 16118 13388 16174 13424
rect 16118 13368 16120 13388
rect 16120 13368 16172 13388
rect 16172 13368 16174 13388
rect 16670 17992 16726 18048
rect 16486 17040 16542 17096
rect 16302 11328 16358 11384
rect 16302 11056 16358 11112
rect 16118 10784 16174 10840
rect 16854 17196 16910 17232
rect 16854 17176 16856 17196
rect 16856 17176 16908 17196
rect 16908 17176 16910 17196
rect 17958 25744 18014 25800
rect 18602 30368 18658 30424
rect 18326 26444 18382 26480
rect 18326 26424 18328 26444
rect 18328 26424 18380 26444
rect 18380 26424 18382 26444
rect 17866 24928 17922 24984
rect 17774 22072 17830 22128
rect 17682 21800 17738 21856
rect 17498 21392 17554 21448
rect 16946 14864 17002 14920
rect 16946 12824 17002 12880
rect 16854 12280 16910 12336
rect 16854 10648 16910 10704
rect 17498 15136 17554 15192
rect 17774 15408 17830 15464
rect 17774 15136 17830 15192
rect 18970 34720 19026 34776
rect 18602 23060 18604 23080
rect 18604 23060 18656 23080
rect 18656 23060 18658 23080
rect 18602 23024 18658 23060
rect 18418 19624 18474 19680
rect 18050 17620 18052 17640
rect 18052 17620 18104 17640
rect 18104 17620 18106 17640
rect 18050 17584 18106 17620
rect 17774 13796 17830 13832
rect 17774 13776 17776 13796
rect 17776 13776 17828 13796
rect 17828 13776 17830 13796
rect 16486 9444 16542 9480
rect 16486 9424 16488 9444
rect 16488 9424 16540 9444
rect 16540 9424 16542 9444
rect 16946 10512 17002 10568
rect 16946 9832 17002 9888
rect 17038 9696 17094 9752
rect 16762 7656 16818 7712
rect 17038 8336 17094 8392
rect 17130 7828 17132 7848
rect 17132 7828 17184 7848
rect 17184 7828 17186 7848
rect 17130 7792 17186 7828
rect 17406 10004 17408 10024
rect 17408 10004 17460 10024
rect 17460 10004 17462 10024
rect 17406 9968 17462 10004
rect 17314 9052 17316 9072
rect 17316 9052 17368 9072
rect 17368 9052 17370 9072
rect 17314 9016 17370 9052
rect 17406 7520 17462 7576
rect 17222 7404 17278 7440
rect 17222 7384 17224 7404
rect 17224 7384 17276 7404
rect 17276 7384 17278 7404
rect 18418 16360 18474 16416
rect 18418 15580 18420 15600
rect 18420 15580 18472 15600
rect 18472 15580 18474 15600
rect 18418 15544 18474 15580
rect 18418 15444 18420 15464
rect 18420 15444 18472 15464
rect 18472 15444 18474 15464
rect 18418 15408 18474 15444
rect 18326 12416 18382 12472
rect 18234 11600 18290 11656
rect 19062 25372 19064 25392
rect 19064 25372 19116 25392
rect 19116 25372 19118 25392
rect 19062 25336 19118 25372
rect 20534 36080 20590 36136
rect 19798 26424 19854 26480
rect 19798 26288 19854 26344
rect 19890 25236 19892 25256
rect 19892 25236 19944 25256
rect 19944 25236 19946 25256
rect 19890 25200 19946 25236
rect 19522 25064 19578 25120
rect 19430 21548 19486 21584
rect 19430 21528 19432 21548
rect 19432 21528 19484 21548
rect 19484 21528 19486 21548
rect 19430 20748 19432 20768
rect 19432 20748 19484 20768
rect 19484 20748 19486 20768
rect 19430 20712 19486 20748
rect 20074 23296 20130 23352
rect 20350 32680 20406 32736
rect 20534 32408 20590 32464
rect 20718 25744 20774 25800
rect 20718 24792 20774 24848
rect 20534 23840 20590 23896
rect 19890 21800 19946 21856
rect 19246 19216 19302 19272
rect 19614 19352 19670 19408
rect 21362 23060 21364 23080
rect 21364 23060 21416 23080
rect 21416 23060 21418 23080
rect 21362 23024 21418 23060
rect 21270 22616 21326 22672
rect 20350 20848 20406 20904
rect 19246 18264 19302 18320
rect 19154 18128 19210 18184
rect 19154 16904 19210 16960
rect 19338 16632 19394 16688
rect 19246 15680 19302 15736
rect 19062 15580 19064 15600
rect 19064 15580 19116 15600
rect 19116 15580 19118 15600
rect 19062 15544 19118 15580
rect 19154 14456 19210 14512
rect 18418 11772 18420 11792
rect 18420 11772 18472 11792
rect 18472 11772 18474 11792
rect 18418 11736 18474 11772
rect 17866 7248 17922 7304
rect 18602 11328 18658 11384
rect 18510 9560 18566 9616
rect 18234 9016 18290 9072
rect 18970 10784 19026 10840
rect 19798 16496 19854 16552
rect 20902 21020 20904 21040
rect 20904 21020 20956 21040
rect 20956 21020 20958 21040
rect 20902 20984 20958 21020
rect 21822 32680 21878 32736
rect 22006 32680 22062 32736
rect 22282 31456 22338 31512
rect 22650 32444 22652 32464
rect 22652 32444 22704 32464
rect 22704 32444 22706 32464
rect 22650 32408 22706 32444
rect 22006 29144 22062 29200
rect 21178 19780 21234 19816
rect 21178 19760 21180 19780
rect 21180 19760 21232 19780
rect 21232 19760 21234 19780
rect 21546 19352 21602 19408
rect 20902 18264 20958 18320
rect 20810 17992 20866 18048
rect 19706 14728 19762 14784
rect 18694 8200 18750 8256
rect 18510 6160 18566 6216
rect 15842 3596 15898 3632
rect 15842 3576 15844 3596
rect 15844 3576 15896 3596
rect 15896 3576 15898 3596
rect 17590 3984 17646 4040
rect 18878 10548 18880 10568
rect 18880 10548 18932 10568
rect 18932 10548 18934 10568
rect 18878 10512 18934 10548
rect 18878 9968 18934 10024
rect 19246 9016 19302 9072
rect 19062 8336 19118 8392
rect 18970 7792 19026 7848
rect 19154 7656 19210 7712
rect 19062 7248 19118 7304
rect 19614 10104 19670 10160
rect 19430 6432 19486 6488
rect 18878 3576 18934 3632
rect 18786 3440 18842 3496
rect 19614 9152 19670 9208
rect 19614 8916 19616 8936
rect 19616 8916 19668 8936
rect 19668 8916 19670 8936
rect 19614 8880 19670 8916
rect 19614 8492 19670 8528
rect 19614 8472 19616 8492
rect 19616 8472 19668 8492
rect 19668 8472 19670 8492
rect 19982 14356 19984 14376
rect 19984 14356 20036 14376
rect 20036 14356 20038 14376
rect 19982 14320 20038 14356
rect 20258 14592 20314 14648
rect 20166 13388 20222 13424
rect 20166 13368 20168 13388
rect 20168 13368 20220 13388
rect 20220 13368 20222 13388
rect 20258 13096 20314 13152
rect 20166 12960 20222 13016
rect 20074 11736 20130 11792
rect 19890 10920 19946 10976
rect 22006 25100 22008 25120
rect 22008 25100 22060 25120
rect 22060 25100 22062 25120
rect 22006 25064 22062 25100
rect 22282 23568 22338 23624
rect 22466 23432 22522 23488
rect 22190 21972 22192 21992
rect 22192 21972 22244 21992
rect 22244 21972 22246 21992
rect 22190 21936 22246 21972
rect 22558 19352 22614 19408
rect 23662 30368 23718 30424
rect 22742 22752 22798 22808
rect 21822 18400 21878 18456
rect 20626 15156 20682 15192
rect 20626 15136 20628 15156
rect 20628 15136 20680 15156
rect 20680 15136 20682 15156
rect 21546 15680 21602 15736
rect 20626 14728 20682 14784
rect 20534 9052 20536 9072
rect 20536 9052 20588 9072
rect 20588 9052 20590 9072
rect 20534 9016 20590 9052
rect 20442 8608 20498 8664
rect 20810 8900 20866 8936
rect 20810 8880 20812 8900
rect 20812 8880 20864 8900
rect 20864 8880 20866 8900
rect 20994 9172 21050 9208
rect 20994 9152 20996 9172
rect 20996 9152 21048 9172
rect 21048 9152 21050 9172
rect 20902 8492 20958 8528
rect 20902 8472 20904 8492
rect 20904 8472 20956 8492
rect 20956 8472 20958 8492
rect 20718 7520 20774 7576
rect 22926 17856 22982 17912
rect 24950 36080 25006 36136
rect 23386 23704 23442 23760
rect 24398 32000 24454 32056
rect 24214 26308 24270 26344
rect 24214 26288 24216 26308
rect 24216 26288 24268 26308
rect 24268 26288 24270 26308
rect 24122 24928 24178 24984
rect 23938 23840 23994 23896
rect 24122 24656 24178 24712
rect 23662 23568 23718 23624
rect 23754 23432 23810 23488
rect 24122 23840 24178 23896
rect 21914 14864 21970 14920
rect 22282 12552 22338 12608
rect 22926 17604 22982 17640
rect 22926 17584 22928 17604
rect 22928 17584 22980 17604
rect 22980 17584 22982 17604
rect 22558 15564 22614 15600
rect 22558 15544 22560 15564
rect 22560 15544 22612 15564
rect 22612 15544 22614 15564
rect 22098 11872 22154 11928
rect 22374 12180 22376 12200
rect 22376 12180 22428 12200
rect 22428 12180 22430 12200
rect 22374 12144 22430 12180
rect 22558 12824 22614 12880
rect 21914 11600 21970 11656
rect 21454 11056 21510 11112
rect 21270 10784 21326 10840
rect 21270 9696 21326 9752
rect 21178 9016 21234 9072
rect 21270 8880 21326 8936
rect 21822 11228 21824 11248
rect 21824 11228 21876 11248
rect 21876 11228 21878 11248
rect 21822 11192 21878 11228
rect 21546 9968 21602 10024
rect 21730 9832 21786 9888
rect 21454 8492 21510 8528
rect 21454 8472 21456 8492
rect 21456 8472 21508 8492
rect 21508 8472 21510 8492
rect 21454 8200 21510 8256
rect 22098 11056 22154 11112
rect 22098 10920 22154 10976
rect 22558 10648 22614 10704
rect 22834 15544 22890 15600
rect 23386 16768 23442 16824
rect 23570 15408 23626 15464
rect 23478 13640 23534 13696
rect 22742 10240 22798 10296
rect 22650 9560 22706 9616
rect 22926 10140 22928 10160
rect 22928 10140 22980 10160
rect 22980 10140 22982 10160
rect 22926 10104 22982 10140
rect 23018 8608 23074 8664
rect 24030 17584 24086 17640
rect 25594 35944 25650 36000
rect 25594 34584 25650 34640
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 35600 38106 35656 38108
rect 35680 38106 35736 38108
rect 35760 38106 35816 38108
rect 35840 38106 35896 38108
rect 35600 38054 35646 38106
rect 35646 38054 35656 38106
rect 35680 38054 35710 38106
rect 35710 38054 35722 38106
rect 35722 38054 35736 38106
rect 35760 38054 35774 38106
rect 35774 38054 35786 38106
rect 35786 38054 35816 38106
rect 35840 38054 35850 38106
rect 35850 38054 35896 38106
rect 35600 38052 35656 38054
rect 35680 38052 35736 38054
rect 35760 38052 35816 38054
rect 35840 38052 35896 38054
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 37830 37440 37886 37496
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 24766 22616 24822 22672
rect 25318 23704 25374 23760
rect 25594 23296 25650 23352
rect 24766 20440 24822 20496
rect 25410 21528 25466 21584
rect 23478 11464 23534 11520
rect 23478 10784 23534 10840
rect 23662 10512 23718 10568
rect 23938 14592 23994 14648
rect 24122 11772 24124 11792
rect 24124 11772 24176 11792
rect 24176 11772 24178 11792
rect 24122 11736 24178 11772
rect 24490 16496 24546 16552
rect 24306 16088 24362 16144
rect 24306 13796 24362 13832
rect 24306 13776 24308 13796
rect 24308 13776 24360 13796
rect 24360 13776 24362 13796
rect 24306 12724 24308 12744
rect 24308 12724 24360 12744
rect 24360 12724 24362 12744
rect 24306 12688 24362 12724
rect 26330 29552 26386 29608
rect 25962 24792 26018 24848
rect 26698 26288 26754 26344
rect 26330 22772 26386 22808
rect 26330 22752 26332 22772
rect 26332 22752 26384 22772
rect 26384 22752 26386 22772
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 37830 35436 37832 35456
rect 37832 35436 37884 35456
rect 37884 35436 37886 35456
rect 37830 35400 37886 35436
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 28630 32680 28686 32736
rect 28078 29280 28134 29336
rect 28078 29008 28134 29064
rect 26422 21800 26478 21856
rect 26330 21428 26332 21448
rect 26332 21428 26384 21448
rect 26384 21428 26386 21448
rect 26330 21392 26386 21428
rect 27250 23860 27306 23896
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 28722 29588 28724 29608
rect 28724 29588 28776 29608
rect 28776 29588 28778 29608
rect 28722 29552 28778 29588
rect 27250 23840 27252 23860
rect 27252 23840 27304 23860
rect 27304 23840 27306 23860
rect 27894 21392 27950 21448
rect 26790 20748 26792 20768
rect 26792 20748 26844 20768
rect 26844 20748 26846 20768
rect 26790 20712 26846 20748
rect 27526 20712 27582 20768
rect 28998 29280 29054 29336
rect 25226 16088 25282 16144
rect 24858 13096 24914 13152
rect 24398 11600 24454 11656
rect 23846 10260 23902 10296
rect 23846 10240 23848 10260
rect 23848 10240 23900 10260
rect 23900 10240 23902 10260
rect 21914 7404 21970 7440
rect 21914 7384 21916 7404
rect 21916 7384 21968 7404
rect 21968 7384 21970 7404
rect 21638 6704 21694 6760
rect 21914 6316 21970 6352
rect 21914 6296 21916 6316
rect 21916 6296 21968 6316
rect 21968 6296 21970 6316
rect 22558 6296 22614 6352
rect 22926 6432 22982 6488
rect 23294 6976 23350 7032
rect 23478 6840 23534 6896
rect 23754 8880 23810 8936
rect 23294 5480 23350 5536
rect 23846 7520 23902 7576
rect 24766 10920 24822 10976
rect 24674 9596 24676 9616
rect 24676 9596 24728 9616
rect 24728 9596 24730 9616
rect 24674 9560 24730 9596
rect 24398 9152 24454 9208
rect 24306 8472 24362 8528
rect 24582 3440 24638 3496
rect 25502 15308 25504 15328
rect 25504 15308 25556 15328
rect 25556 15308 25558 15328
rect 25502 15272 25558 15308
rect 25410 14320 25466 14376
rect 25778 16108 25834 16144
rect 25778 16088 25780 16108
rect 25780 16088 25832 16108
rect 25832 16088 25834 16108
rect 25778 15428 25834 15464
rect 25778 15408 25780 15428
rect 25780 15408 25832 15428
rect 25832 15408 25834 15428
rect 25778 15272 25834 15328
rect 25134 13096 25190 13152
rect 25042 12844 25098 12880
rect 25042 12824 25044 12844
rect 25044 12824 25096 12844
rect 25096 12824 25098 12844
rect 25042 11872 25098 11928
rect 25318 12980 25374 13016
rect 25318 12960 25320 12980
rect 25320 12960 25372 12980
rect 25372 12960 25374 12980
rect 25778 13232 25834 13288
rect 25962 15680 26018 15736
rect 25410 12552 25466 12608
rect 25502 12416 25558 12472
rect 25502 11636 25504 11656
rect 25504 11636 25556 11656
rect 25556 11636 25558 11656
rect 25502 11600 25558 11636
rect 25502 11092 25504 11112
rect 25504 11092 25556 11112
rect 25556 11092 25558 11112
rect 25502 11056 25558 11092
rect 25502 10784 25558 10840
rect 24858 9968 24914 10024
rect 25134 9560 25190 9616
rect 25410 10376 25466 10432
rect 25594 10104 25650 10160
rect 25686 9696 25742 9752
rect 26146 15408 26202 15464
rect 25962 10784 26018 10840
rect 26330 16532 26332 16552
rect 26332 16532 26384 16552
rect 26384 16532 26386 16552
rect 26330 16496 26386 16532
rect 26330 15544 26386 15600
rect 26882 16496 26938 16552
rect 26790 15680 26846 15736
rect 26882 15544 26938 15600
rect 26422 12960 26478 13016
rect 26422 12824 26478 12880
rect 26974 12980 27030 13016
rect 26974 12960 26976 12980
rect 26976 12960 27028 12980
rect 27028 12960 27030 12980
rect 26514 12280 26570 12336
rect 26330 11056 26386 11112
rect 26054 9832 26110 9888
rect 26146 9580 26202 9616
rect 26146 9560 26148 9580
rect 26148 9560 26200 9580
rect 26200 9560 26202 9580
rect 26790 9560 26846 9616
rect 25226 7384 25282 7440
rect 25410 7112 25466 7168
rect 25502 6724 25558 6760
rect 25870 7112 25926 7168
rect 25502 6704 25504 6724
rect 25504 6704 25556 6724
rect 25556 6704 25558 6724
rect 25870 6432 25926 6488
rect 25594 6316 25650 6352
rect 25594 6296 25596 6316
rect 25596 6296 25648 6316
rect 25648 6296 25650 6316
rect 26514 6976 26570 7032
rect 25226 3848 25282 3904
rect 24674 2624 24730 2680
rect 28722 18264 28778 18320
rect 27526 17604 27582 17640
rect 27526 17584 27528 17604
rect 27528 17584 27580 17604
rect 27580 17584 27582 17604
rect 27526 16632 27582 16688
rect 27066 10920 27122 10976
rect 27342 10240 27398 10296
rect 28078 16088 28134 16144
rect 28722 16632 28778 16688
rect 27894 14864 27950 14920
rect 28262 13912 28318 13968
rect 28170 12144 28226 12200
rect 26790 4936 26846 4992
rect 27894 10104 27950 10160
rect 27710 9016 27766 9072
rect 27710 7928 27766 7984
rect 28630 12144 28686 12200
rect 28998 12708 29054 12744
rect 28998 12688 29000 12708
rect 29000 12688 29052 12708
rect 29052 12688 29054 12708
rect 28814 10784 28870 10840
rect 28538 10260 28594 10296
rect 28538 10240 28540 10260
rect 28540 10240 28592 10260
rect 28592 10240 28594 10260
rect 28446 9968 28502 10024
rect 28630 10104 28686 10160
rect 28906 10512 28962 10568
rect 28998 9560 29054 9616
rect 29550 25880 29606 25936
rect 29366 11872 29422 11928
rect 30286 20304 30342 20360
rect 29826 16244 29882 16280
rect 29826 16224 29828 16244
rect 29828 16224 29880 16244
rect 29880 16224 29882 16244
rect 29826 12688 29882 12744
rect 31482 29280 31538 29336
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 32218 25900 32274 25936
rect 32218 25880 32220 25900
rect 32220 25880 32272 25900
rect 32272 25880 32274 25900
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 31206 20324 31262 20360
rect 31206 20304 31208 20324
rect 31208 20304 31260 20324
rect 31260 20304 31262 20324
rect 33782 26288 33838 26344
rect 32402 20440 32458 20496
rect 30102 15000 30158 15056
rect 30562 16768 30618 16824
rect 34150 29008 34206 29064
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 35162 29280 35218 29336
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 36450 28464 36506 28520
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 33874 23024 33930 23080
rect 34426 23840 34482 23896
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 36818 29144 36874 29200
rect 37278 28464 37334 28520
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34886 22516 34888 22536
rect 34888 22516 34940 22536
rect 34940 22516 34942 22536
rect 34886 22480 34942 22516
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34242 19760 34298 19816
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 36266 22636 36322 22672
rect 36266 22616 36268 22636
rect 36268 22616 36320 22636
rect 36320 22616 36322 22636
rect 36266 22500 36322 22536
rect 36266 22480 36268 22500
rect 36268 22480 36320 22500
rect 36320 22480 36322 22500
rect 38290 32680 38346 32736
rect 30746 16224 30802 16280
rect 30378 13368 30434 13424
rect 29550 9424 29606 9480
rect 29366 8064 29422 8120
rect 29826 9288 29882 9344
rect 30286 9152 30342 9208
rect 32034 16224 32090 16280
rect 31666 10376 31722 10432
rect 1490 2080 1546 2136
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 37830 21120 37886 21176
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 38290 19080 38346 19136
rect 38290 14320 38346 14376
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 33598 12688 33654 12744
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 37646 12280 37702 12336
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 37830 11620 37886 11656
rect 37830 11600 37832 11620
rect 37832 11600 37884 11620
rect 37884 11600 37886 11620
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35714 2352 35770 2408
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
rect 37738 2080 37794 2136
rect 37922 40 37978 96
<< metal3 >>
rect 37181 40218 37247 40221
rect 38621 40218 39421 40248
rect 37181 40216 39421 40218
rect 37181 40160 37186 40216
rect 37242 40160 39421 40216
rect 37181 40158 39421 40160
rect 37181 40155 37247 40158
rect 38621 40128 39421 40158
rect 0 39538 800 39568
rect 1117 39538 1183 39541
rect 0 39536 1183 39538
rect 0 39480 1122 39536
rect 1178 39480 1183 39536
rect 0 39478 1183 39480
rect 0 39448 800 39478
rect 1117 39475 1183 39478
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 35590 39200 35906 39201
rect 35590 39136 35596 39200
rect 35660 39136 35676 39200
rect 35740 39136 35756 39200
rect 35820 39136 35836 39200
rect 35900 39136 35906 39200
rect 35590 39135 35906 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 35590 38112 35906 38113
rect 35590 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35906 38112
rect 35590 38047 35906 38048
rect 4210 37568 4526 37569
rect 0 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 933 37498 999 37501
rect 0 37496 999 37498
rect 0 37440 938 37496
rect 994 37440 999 37496
rect 0 37438 999 37440
rect 0 37408 800 37438
rect 933 37435 999 37438
rect 37825 37498 37891 37501
rect 38621 37498 39421 37528
rect 37825 37496 39421 37498
rect 37825 37440 37830 37496
rect 37886 37440 39421 37496
rect 37825 37438 39421 37440
rect 37825 37435 37891 37438
rect 38621 37408 39421 37438
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 20529 36138 20595 36141
rect 24945 36138 25011 36141
rect 20529 36136 25011 36138
rect 20529 36080 20534 36136
rect 20590 36080 24950 36136
rect 25006 36080 25011 36136
rect 20529 36078 25011 36080
rect 20529 36075 20595 36078
rect 24945 36075 25011 36078
rect 19333 36002 19399 36005
rect 25589 36002 25655 36005
rect 19333 36000 25655 36002
rect 19333 35944 19338 36000
rect 19394 35944 25594 36000
rect 25650 35944 25655 36000
rect 19333 35942 25655 35944
rect 19333 35939 19399 35942
rect 25589 35939 25655 35942
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 12433 35868 12499 35869
rect 12382 35866 12388 35868
rect 12342 35806 12388 35866
rect 12452 35864 12499 35868
rect 12494 35808 12499 35864
rect 12382 35804 12388 35806
rect 12452 35804 12499 35808
rect 12433 35803 12499 35804
rect 12985 35594 13051 35597
rect 16113 35594 16179 35597
rect 12985 35592 16179 35594
rect 12985 35536 12990 35592
rect 13046 35536 16118 35592
rect 16174 35536 16179 35592
rect 12985 35534 16179 35536
rect 12985 35531 13051 35534
rect 16113 35531 16179 35534
rect 37825 35458 37891 35461
rect 38621 35458 39421 35488
rect 37825 35456 39421 35458
rect 37825 35400 37830 35456
rect 37886 35400 39421 35456
rect 37825 35398 39421 35400
rect 37825 35395 37891 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 38621 35368 39421 35398
rect 34930 35327 35246 35328
rect 11605 35324 11671 35325
rect 11605 35322 11652 35324
rect 11560 35320 11652 35322
rect 11560 35264 11610 35320
rect 11560 35262 11652 35264
rect 11605 35260 11652 35262
rect 11716 35260 11722 35324
rect 11605 35259 11671 35260
rect 4870 34848 5186 34849
rect 0 34778 800 34808
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 933 34778 999 34781
rect 0 34776 999 34778
rect 0 34720 938 34776
rect 994 34720 999 34776
rect 0 34718 999 34720
rect 0 34688 800 34718
rect 933 34715 999 34718
rect 11973 34778 12039 34781
rect 18965 34778 19031 34781
rect 11973 34776 19031 34778
rect 11973 34720 11978 34776
rect 12034 34720 18970 34776
rect 19026 34720 19031 34776
rect 11973 34718 19031 34720
rect 11973 34715 12039 34718
rect 18965 34715 19031 34718
rect 25589 34642 25655 34645
rect 25998 34642 26004 34644
rect 25589 34640 26004 34642
rect 25589 34584 25594 34640
rect 25650 34584 26004 34640
rect 25589 34582 26004 34584
rect 25589 34579 25655 34582
rect 25998 34580 26004 34582
rect 26068 34580 26074 34644
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 0 32648 800 32768
rect 20345 32738 20411 32741
rect 21817 32738 21883 32741
rect 20345 32736 21883 32738
rect 20345 32680 20350 32736
rect 20406 32680 21822 32736
rect 21878 32680 21883 32736
rect 20345 32678 21883 32680
rect 20345 32675 20411 32678
rect 21817 32675 21883 32678
rect 22001 32738 22067 32741
rect 28625 32738 28691 32741
rect 29126 32738 29132 32740
rect 22001 32736 29132 32738
rect 22001 32680 22006 32736
rect 22062 32680 28630 32736
rect 28686 32680 29132 32736
rect 22001 32678 29132 32680
rect 22001 32675 22067 32678
rect 28625 32675 28691 32678
rect 29126 32676 29132 32678
rect 29196 32676 29202 32740
rect 38285 32738 38351 32741
rect 38621 32738 39421 32768
rect 38285 32736 39421 32738
rect 38285 32680 38290 32736
rect 38346 32680 39421 32736
rect 38285 32678 39421 32680
rect 38285 32675 38351 32678
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 38621 32648 39421 32678
rect 35590 32607 35906 32608
rect 20529 32466 20595 32469
rect 22645 32466 22711 32469
rect 20529 32464 22711 32466
rect 20529 32408 20534 32464
rect 20590 32408 22650 32464
rect 22706 32408 22711 32464
rect 20529 32406 22711 32408
rect 20529 32403 20595 32406
rect 22645 32403 22711 32406
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 24393 32058 24459 32061
rect 26734 32058 26740 32060
rect 24393 32056 26740 32058
rect 24393 32000 24398 32056
rect 24454 32000 26740 32056
rect 24393 31998 26740 32000
rect 24393 31995 24459 31998
rect 26734 31996 26740 31998
rect 26804 31996 26810 32060
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 13721 31514 13787 31517
rect 15561 31514 15627 31517
rect 22277 31516 22343 31517
rect 22277 31514 22324 31516
rect 13721 31512 15627 31514
rect 13721 31456 13726 31512
rect 13782 31456 15566 31512
rect 15622 31456 15627 31512
rect 13721 31454 15627 31456
rect 22232 31512 22324 31514
rect 22232 31456 22282 31512
rect 22232 31454 22324 31456
rect 13721 31451 13787 31454
rect 15561 31451 15627 31454
rect 22277 31452 22324 31454
rect 22388 31452 22394 31516
rect 22277 31451 22343 31452
rect 14825 31242 14891 31245
rect 16665 31242 16731 31245
rect 14825 31240 16731 31242
rect 14825 31184 14830 31240
rect 14886 31184 16670 31240
rect 16726 31184 16731 31240
rect 14825 31182 16731 31184
rect 14825 31179 14891 31182
rect 16665 31179 16731 31182
rect 13813 31106 13879 31109
rect 15193 31106 15259 31109
rect 13813 31104 15259 31106
rect 13813 31048 13818 31104
rect 13874 31048 15198 31104
rect 15254 31048 15259 31104
rect 13813 31046 15259 31048
rect 13813 31043 13879 31046
rect 15193 31043 15259 31046
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 17493 30834 17559 30837
rect 20110 30834 20116 30836
rect 17493 30832 20116 30834
rect 17493 30776 17498 30832
rect 17554 30776 20116 30832
rect 17493 30774 20116 30776
rect 17493 30771 17559 30774
rect 20110 30772 20116 30774
rect 20180 30772 20186 30836
rect 0 30608 800 30728
rect 38621 30608 39421 30728
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 12198 30364 12204 30428
rect 12268 30426 12274 30428
rect 12525 30426 12591 30429
rect 12268 30424 12591 30426
rect 12268 30368 12530 30424
rect 12586 30368 12591 30424
rect 12268 30366 12591 30368
rect 12268 30364 12274 30366
rect 12525 30363 12591 30366
rect 15561 30426 15627 30429
rect 18597 30428 18663 30429
rect 17534 30426 17540 30428
rect 15561 30424 17540 30426
rect 15561 30368 15566 30424
rect 15622 30368 17540 30424
rect 15561 30366 17540 30368
rect 15561 30363 15627 30366
rect 17534 30364 17540 30366
rect 17604 30364 17610 30428
rect 18597 30426 18644 30428
rect 18552 30424 18644 30426
rect 18552 30368 18602 30424
rect 18552 30366 18644 30368
rect 18597 30364 18644 30366
rect 18708 30364 18714 30428
rect 23657 30426 23723 30429
rect 25446 30426 25452 30428
rect 23657 30424 25452 30426
rect 23657 30368 23662 30424
rect 23718 30368 25452 30424
rect 23657 30366 25452 30368
rect 18597 30363 18663 30364
rect 23657 30363 23723 30366
rect 25446 30364 25452 30366
rect 25516 30364 25522 30428
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 26325 29610 26391 29613
rect 28717 29610 28783 29613
rect 26325 29608 28783 29610
rect 26325 29552 26330 29608
rect 26386 29552 28722 29608
rect 28778 29552 28783 29608
rect 26325 29550 28783 29552
rect 26325 29547 26391 29550
rect 28717 29547 28783 29550
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 28073 29338 28139 29341
rect 28993 29338 29059 29341
rect 28073 29336 29059 29338
rect 28073 29280 28078 29336
rect 28134 29280 28998 29336
rect 29054 29280 29059 29336
rect 28073 29278 29059 29280
rect 28073 29275 28139 29278
rect 28993 29275 29059 29278
rect 31477 29338 31543 29341
rect 35157 29338 35223 29341
rect 31477 29336 35223 29338
rect 31477 29280 31482 29336
rect 31538 29280 35162 29336
rect 35218 29280 35223 29336
rect 31477 29278 35223 29280
rect 31477 29275 31543 29278
rect 35157 29275 35223 29278
rect 4613 29202 4679 29205
rect 5073 29202 5139 29205
rect 4613 29200 5139 29202
rect 4613 29144 4618 29200
rect 4674 29144 5078 29200
rect 5134 29144 5139 29200
rect 4613 29142 5139 29144
rect 4613 29139 4679 29142
rect 5073 29139 5139 29142
rect 22001 29202 22067 29205
rect 36813 29202 36879 29205
rect 22001 29200 36879 29202
rect 22001 29144 22006 29200
rect 22062 29144 36818 29200
rect 36874 29144 36879 29200
rect 22001 29142 36879 29144
rect 22001 29139 22067 29142
rect 36813 29139 36879 29142
rect 12157 29066 12223 29069
rect 12382 29066 12388 29068
rect 12157 29064 12388 29066
rect 12157 29008 12162 29064
rect 12218 29008 12388 29064
rect 12157 29006 12388 29008
rect 12157 29003 12223 29006
rect 12382 29004 12388 29006
rect 12452 29004 12458 29068
rect 28073 29066 28139 29069
rect 34145 29066 34211 29069
rect 28073 29064 34211 29066
rect 28073 29008 28078 29064
rect 28134 29008 34150 29064
rect 34206 29008 34211 29064
rect 28073 29006 34211 29008
rect 28073 29003 28139 29006
rect 34145 29003 34211 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 36445 28522 36511 28525
rect 37273 28522 37339 28525
rect 36445 28520 37339 28522
rect 36445 28464 36450 28520
rect 36506 28464 37278 28520
rect 37334 28464 37339 28520
rect 36445 28462 37339 28464
rect 36445 28459 36511 28462
rect 37273 28459 37339 28462
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 0 27888 800 28008
rect 38621 27888 39421 28008
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 35590 27167 35906 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 16849 26482 16915 26485
rect 18321 26482 18387 26485
rect 16849 26480 18387 26482
rect 16849 26424 16854 26480
rect 16910 26424 18326 26480
rect 18382 26424 18387 26480
rect 16849 26422 18387 26424
rect 16849 26419 16915 26422
rect 18321 26419 18387 26422
rect 19793 26482 19859 26485
rect 21030 26482 21036 26484
rect 19793 26480 21036 26482
rect 19793 26424 19798 26480
rect 19854 26424 21036 26480
rect 19793 26422 21036 26424
rect 19793 26419 19859 26422
rect 21030 26420 21036 26422
rect 21100 26420 21106 26484
rect 14406 26284 14412 26348
rect 14476 26346 14482 26348
rect 14917 26346 14983 26349
rect 19793 26348 19859 26349
rect 14476 26344 14983 26346
rect 14476 26288 14922 26344
rect 14978 26288 14983 26344
rect 14476 26286 14983 26288
rect 14476 26284 14482 26286
rect 14917 26283 14983 26286
rect 19742 26284 19748 26348
rect 19812 26346 19859 26348
rect 24209 26346 24275 26349
rect 24710 26346 24716 26348
rect 19812 26344 19904 26346
rect 19854 26288 19904 26344
rect 19812 26286 19904 26288
rect 24209 26344 24716 26346
rect 24209 26288 24214 26344
rect 24270 26288 24716 26344
rect 24209 26286 24716 26288
rect 19812 26284 19859 26286
rect 19793 26283 19859 26284
rect 24209 26283 24275 26286
rect 24710 26284 24716 26286
rect 24780 26284 24786 26348
rect 26693 26346 26759 26349
rect 33777 26346 33843 26349
rect 26693 26344 33843 26346
rect 26693 26288 26698 26344
rect 26754 26288 33782 26344
rect 33838 26288 33843 26344
rect 26693 26286 33843 26288
rect 26693 26283 26759 26286
rect 33777 26283 33843 26286
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 0 25938 800 25968
rect 933 25938 999 25941
rect 14549 25940 14615 25941
rect 14549 25938 14596 25940
rect 0 25936 999 25938
rect 0 25880 938 25936
rect 994 25880 999 25936
rect 0 25878 999 25880
rect 14508 25936 14596 25938
rect 14660 25938 14666 25940
rect 16389 25938 16455 25941
rect 14660 25936 16455 25938
rect 14508 25880 14554 25936
rect 14660 25880 16394 25936
rect 16450 25880 16455 25936
rect 14508 25878 14596 25880
rect 0 25848 800 25878
rect 933 25875 999 25878
rect 14549 25876 14596 25878
rect 14660 25878 16455 25880
rect 14660 25876 14666 25878
rect 14549 25875 14615 25876
rect 16389 25875 16455 25878
rect 29545 25938 29611 25941
rect 32213 25938 32279 25941
rect 29545 25936 32279 25938
rect 29545 25880 29550 25936
rect 29606 25880 32218 25936
rect 32274 25880 32279 25936
rect 29545 25878 32279 25880
rect 29545 25875 29611 25878
rect 32213 25875 32279 25878
rect 38621 25848 39421 25968
rect 13169 25802 13235 25805
rect 17953 25802 18019 25805
rect 20713 25802 20779 25805
rect 13169 25800 20779 25802
rect 13169 25744 13174 25800
rect 13230 25744 17958 25800
rect 18014 25744 20718 25800
rect 20774 25744 20779 25800
rect 13169 25742 20779 25744
rect 13169 25739 13235 25742
rect 17953 25739 18019 25742
rect 20713 25739 20779 25742
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 12893 25394 12959 25397
rect 19057 25394 19123 25397
rect 12893 25392 19123 25394
rect 12893 25336 12898 25392
rect 12954 25336 19062 25392
rect 19118 25336 19123 25392
rect 12893 25334 19123 25336
rect 12893 25331 12959 25334
rect 19057 25331 19123 25334
rect 17493 25258 17559 25261
rect 19885 25258 19951 25261
rect 17493 25256 19951 25258
rect 17493 25200 17498 25256
rect 17554 25200 19890 25256
rect 19946 25200 19951 25256
rect 17493 25198 19951 25200
rect 17493 25195 17559 25198
rect 19885 25195 19951 25198
rect 19517 25122 19583 25125
rect 22001 25122 22067 25125
rect 19517 25120 22067 25122
rect 19517 25064 19522 25120
rect 19578 25064 22006 25120
rect 22062 25064 22067 25120
rect 19517 25062 22067 25064
rect 19517 25059 19583 25062
rect 22001 25059 22067 25062
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 17718 24924 17724 24988
rect 17788 24986 17794 24988
rect 17861 24986 17927 24989
rect 17788 24984 17927 24986
rect 17788 24928 17866 24984
rect 17922 24928 17927 24984
rect 17788 24926 17927 24928
rect 17788 24924 17794 24926
rect 17861 24923 17927 24926
rect 24117 24986 24183 24989
rect 30966 24986 30972 24988
rect 24117 24984 30972 24986
rect 24117 24928 24122 24984
rect 24178 24928 30972 24984
rect 24117 24926 30972 24928
rect 24117 24923 24183 24926
rect 30966 24924 30972 24926
rect 31036 24924 31042 24988
rect 6637 24850 6703 24853
rect 20713 24850 20779 24853
rect 25957 24852 26023 24853
rect 25957 24850 26004 24852
rect 6637 24848 20779 24850
rect 6637 24792 6642 24848
rect 6698 24792 20718 24848
rect 20774 24792 20779 24848
rect 6637 24790 20779 24792
rect 25912 24848 26004 24850
rect 25912 24792 25962 24848
rect 25912 24790 26004 24792
rect 6637 24787 6703 24790
rect 20713 24787 20779 24790
rect 25957 24788 26004 24790
rect 26068 24788 26074 24852
rect 25957 24787 26023 24788
rect 15101 24714 15167 24717
rect 24117 24714 24183 24717
rect 15101 24712 24183 24714
rect 15101 24656 15106 24712
rect 15162 24656 24122 24712
rect 24178 24656 24183 24712
rect 15101 24654 24183 24656
rect 15101 24651 15167 24654
rect 24117 24651 24183 24654
rect 7465 24578 7531 24581
rect 13905 24578 13971 24581
rect 15101 24578 15167 24581
rect 7465 24576 15167 24578
rect 7465 24520 7470 24576
rect 7526 24520 13910 24576
rect 13966 24520 15106 24576
rect 15162 24520 15167 24576
rect 7465 24518 15167 24520
rect 7465 24515 7531 24518
rect 13905 24515 13971 24518
rect 15101 24515 15167 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 15377 24170 15443 24173
rect 16757 24170 16823 24173
rect 15377 24168 16823 24170
rect 15377 24112 15382 24168
rect 15438 24112 16762 24168
rect 16818 24112 16823 24168
rect 15377 24110 16823 24112
rect 15377 24107 15443 24110
rect 16757 24107 16823 24110
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 20529 23898 20595 23901
rect 23933 23898 23999 23901
rect 24117 23900 24183 23901
rect 24117 23898 24164 23900
rect 20529 23896 23999 23898
rect 20529 23840 20534 23896
rect 20590 23840 23938 23896
rect 23994 23840 23999 23896
rect 20529 23838 23999 23840
rect 24072 23896 24164 23898
rect 24072 23840 24122 23896
rect 24072 23838 24164 23840
rect 20529 23835 20595 23838
rect 23933 23835 23999 23838
rect 24117 23836 24164 23838
rect 24228 23836 24234 23900
rect 27245 23898 27311 23901
rect 34421 23898 34487 23901
rect 27245 23896 34487 23898
rect 27245 23840 27250 23896
rect 27306 23840 34426 23896
rect 34482 23840 34487 23896
rect 27245 23838 34487 23840
rect 24117 23835 24183 23836
rect 27245 23835 27311 23838
rect 34421 23835 34487 23838
rect 38621 23808 39421 23928
rect 6913 23762 6979 23765
rect 23381 23762 23447 23765
rect 23606 23762 23612 23764
rect 6913 23760 23306 23762
rect 6913 23704 6918 23760
rect 6974 23704 23306 23760
rect 6913 23702 23306 23704
rect 6913 23699 6979 23702
rect 22277 23626 22343 23629
rect 22686 23626 22692 23628
rect 22277 23624 22692 23626
rect 22277 23568 22282 23624
rect 22338 23568 22692 23624
rect 22277 23566 22692 23568
rect 22277 23563 22343 23566
rect 22686 23564 22692 23566
rect 22756 23564 22762 23628
rect 13118 23428 13124 23492
rect 13188 23490 13194 23492
rect 14549 23490 14615 23493
rect 13188 23488 14615 23490
rect 13188 23432 14554 23488
rect 14610 23432 14615 23488
rect 13188 23430 14615 23432
rect 13188 23428 13194 23430
rect 14549 23427 14615 23430
rect 22461 23492 22527 23493
rect 22461 23488 22508 23492
rect 22572 23490 22578 23492
rect 23246 23490 23306 23702
rect 23381 23760 23612 23762
rect 23381 23704 23386 23760
rect 23442 23704 23612 23760
rect 23381 23702 23612 23704
rect 23381 23699 23447 23702
rect 23606 23700 23612 23702
rect 23676 23762 23682 23764
rect 25313 23762 25379 23765
rect 23676 23760 25379 23762
rect 23676 23704 25318 23760
rect 25374 23704 25379 23760
rect 23676 23702 25379 23704
rect 23676 23700 23682 23702
rect 25313 23699 25379 23702
rect 23657 23626 23723 23629
rect 26918 23626 26924 23628
rect 23657 23624 26924 23626
rect 23657 23568 23662 23624
rect 23718 23568 26924 23624
rect 23657 23566 26924 23568
rect 23657 23563 23723 23566
rect 26918 23564 26924 23566
rect 26988 23564 26994 23628
rect 23749 23492 23815 23493
rect 23749 23490 23796 23492
rect 22461 23432 22466 23488
rect 22461 23428 22508 23432
rect 22572 23430 22618 23490
rect 23246 23488 23796 23490
rect 23246 23432 23754 23488
rect 23246 23430 23796 23432
rect 22572 23428 22578 23430
rect 23749 23428 23796 23430
rect 23860 23428 23866 23492
rect 22461 23427 22527 23428
rect 23749 23427 23815 23428
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 20069 23354 20135 23357
rect 25589 23354 25655 23357
rect 20069 23352 25655 23354
rect 20069 23296 20074 23352
rect 20130 23296 25594 23352
rect 25650 23296 25655 23352
rect 20069 23294 25655 23296
rect 20069 23291 20135 23294
rect 25589 23291 25655 23294
rect 0 23128 800 23248
rect 16113 23082 16179 23085
rect 18597 23082 18663 23085
rect 16113 23080 18663 23082
rect 16113 23024 16118 23080
rect 16174 23024 18602 23080
rect 18658 23024 18663 23080
rect 16113 23022 18663 23024
rect 16113 23019 16179 23022
rect 18597 23019 18663 23022
rect 21357 23082 21423 23085
rect 33869 23082 33935 23085
rect 21357 23080 33935 23082
rect 21357 23024 21362 23080
rect 21418 23024 33874 23080
rect 33930 23024 33935 23080
rect 21357 23022 33935 23024
rect 21357 23019 21423 23022
rect 33869 23019 33935 23022
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 22737 22810 22803 22813
rect 26325 22810 26391 22813
rect 22737 22808 26391 22810
rect 22737 22752 22742 22808
rect 22798 22752 26330 22808
rect 26386 22752 26391 22808
rect 22737 22750 26391 22752
rect 22737 22747 22803 22750
rect 26325 22747 26391 22750
rect 21265 22674 21331 22677
rect 24761 22674 24827 22677
rect 36261 22674 36327 22677
rect 21265 22672 36327 22674
rect 21265 22616 21270 22672
rect 21326 22616 24766 22672
rect 24822 22616 36266 22672
rect 36322 22616 36327 22672
rect 21265 22614 36327 22616
rect 21265 22611 21331 22614
rect 24761 22611 24827 22614
rect 36261 22611 36327 22614
rect 34881 22538 34947 22541
rect 36261 22538 36327 22541
rect 34881 22536 36327 22538
rect 34881 22480 34886 22536
rect 34942 22480 36266 22536
rect 36322 22480 36327 22536
rect 34881 22478 36327 22480
rect 34881 22475 34947 22478
rect 36261 22475 36327 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 17033 22130 17099 22133
rect 17769 22130 17835 22133
rect 17033 22128 17835 22130
rect 17033 22072 17038 22128
rect 17094 22072 17774 22128
rect 17830 22072 17835 22128
rect 17033 22070 17835 22072
rect 17033 22067 17099 22070
rect 17769 22067 17835 22070
rect 8845 21994 8911 21997
rect 10409 21994 10475 21997
rect 8845 21992 10475 21994
rect 8845 21936 8850 21992
rect 8906 21936 10414 21992
rect 10470 21936 10475 21992
rect 8845 21934 10475 21936
rect 8845 21931 8911 21934
rect 10409 21931 10475 21934
rect 11973 21994 12039 21997
rect 22185 21994 22251 21997
rect 11973 21992 22251 21994
rect 11973 21936 11978 21992
rect 12034 21936 22190 21992
rect 22246 21936 22251 21992
rect 11973 21934 22251 21936
rect 11973 21931 12039 21934
rect 22185 21931 22251 21934
rect 17033 21858 17099 21861
rect 17677 21858 17743 21861
rect 17033 21856 17743 21858
rect 17033 21800 17038 21856
rect 17094 21800 17682 21856
rect 17738 21800 17743 21856
rect 17033 21798 17743 21800
rect 17033 21795 17099 21798
rect 17677 21795 17743 21798
rect 19885 21858 19951 21861
rect 26417 21858 26483 21861
rect 19885 21856 26483 21858
rect 19885 21800 19890 21856
rect 19946 21800 26422 21856
rect 26478 21800 26483 21856
rect 19885 21798 26483 21800
rect 19885 21795 19951 21798
rect 26417 21795 26483 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 35590 21727 35906 21728
rect 6085 21586 6151 21589
rect 19425 21586 19491 21589
rect 6085 21584 19491 21586
rect 6085 21528 6090 21584
rect 6146 21528 19430 21584
rect 19486 21528 19491 21584
rect 6085 21526 19491 21528
rect 6085 21523 6151 21526
rect 19425 21523 19491 21526
rect 25405 21588 25471 21589
rect 25405 21584 25452 21588
rect 25516 21586 25522 21588
rect 25405 21528 25410 21584
rect 25405 21524 25452 21528
rect 25516 21526 25562 21586
rect 25516 21524 25522 21526
rect 25405 21523 25471 21524
rect 10501 21450 10567 21453
rect 11697 21450 11763 21453
rect 14549 21450 14615 21453
rect 10501 21448 14615 21450
rect 10501 21392 10506 21448
rect 10562 21392 11702 21448
rect 11758 21392 14554 21448
rect 14610 21392 14615 21448
rect 10501 21390 14615 21392
rect 10501 21387 10567 21390
rect 11697 21387 11763 21390
rect 14549 21387 14615 21390
rect 14825 21450 14891 21453
rect 17493 21450 17559 21453
rect 14825 21448 17559 21450
rect 14825 21392 14830 21448
rect 14886 21392 17498 21448
rect 17554 21392 17559 21448
rect 14825 21390 17559 21392
rect 14825 21387 14891 21390
rect 17493 21387 17559 21390
rect 26325 21450 26391 21453
rect 27889 21450 27955 21453
rect 26325 21448 27955 21450
rect 26325 21392 26330 21448
rect 26386 21392 27894 21448
rect 27950 21392 27955 21448
rect 26325 21390 27955 21392
rect 26325 21387 26391 21390
rect 27889 21387 27955 21390
rect 4210 21248 4526 21249
rect 0 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 933 21178 999 21181
rect 0 21176 999 21178
rect 0 21120 938 21176
rect 994 21120 999 21176
rect 0 21118 999 21120
rect 0 21088 800 21118
rect 933 21115 999 21118
rect 37825 21178 37891 21181
rect 38621 21178 39421 21208
rect 37825 21176 39421 21178
rect 37825 21120 37830 21176
rect 37886 21120 39421 21176
rect 37825 21118 39421 21120
rect 37825 21115 37891 21118
rect 38621 21088 39421 21118
rect 18822 20980 18828 21044
rect 18892 21042 18898 21044
rect 20897 21042 20963 21045
rect 18892 21040 20963 21042
rect 18892 20984 20902 21040
rect 20958 20984 20963 21040
rect 18892 20982 20963 20984
rect 18892 20980 18898 20982
rect 20897 20979 20963 20982
rect 3141 20906 3207 20909
rect 20345 20906 20411 20909
rect 3141 20904 20411 20906
rect 3141 20848 3146 20904
rect 3202 20848 20350 20904
rect 20406 20848 20411 20904
rect 3141 20846 20411 20848
rect 3141 20843 3207 20846
rect 20345 20843 20411 20846
rect 12341 20770 12407 20773
rect 19425 20770 19491 20773
rect 12341 20768 19491 20770
rect 12341 20712 12346 20768
rect 12402 20712 19430 20768
rect 19486 20712 19491 20768
rect 12341 20710 19491 20712
rect 12341 20707 12407 20710
rect 19425 20707 19491 20710
rect 26785 20770 26851 20773
rect 27102 20770 27108 20772
rect 26785 20768 27108 20770
rect 26785 20712 26790 20768
rect 26846 20712 27108 20768
rect 26785 20710 27108 20712
rect 26785 20707 26851 20710
rect 27102 20708 27108 20710
rect 27172 20770 27178 20772
rect 27521 20770 27587 20773
rect 27172 20768 27587 20770
rect 27172 20712 27526 20768
rect 27582 20712 27587 20768
rect 27172 20710 27587 20712
rect 27172 20708 27178 20710
rect 27521 20707 27587 20710
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 7925 20498 7991 20501
rect 24761 20498 24827 20501
rect 32397 20498 32463 20501
rect 7925 20496 32463 20498
rect 7925 20440 7930 20496
rect 7986 20440 24766 20496
rect 24822 20440 32402 20496
rect 32458 20440 32463 20496
rect 7925 20438 32463 20440
rect 7925 20435 7991 20438
rect 24761 20435 24827 20438
rect 32397 20435 32463 20438
rect 30281 20362 30347 20365
rect 31201 20362 31267 20365
rect 30281 20360 31267 20362
rect 30281 20304 30286 20360
rect 30342 20304 31206 20360
rect 31262 20304 31267 20360
rect 30281 20302 31267 20304
rect 30281 20299 30347 20302
rect 31201 20299 31267 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 8293 19818 8359 19821
rect 16481 19818 16547 19821
rect 8293 19816 16547 19818
rect 8293 19760 8298 19816
rect 8354 19760 16486 19816
rect 16542 19760 16547 19816
rect 8293 19758 16547 19760
rect 8293 19755 8359 19758
rect 16481 19755 16547 19758
rect 21173 19818 21239 19821
rect 34237 19818 34303 19821
rect 21173 19816 34303 19818
rect 21173 19760 21178 19816
rect 21234 19760 34242 19816
rect 34298 19760 34303 19816
rect 21173 19758 34303 19760
rect 21173 19755 21239 19758
rect 34237 19755 34303 19758
rect 11605 19682 11671 19685
rect 14365 19682 14431 19685
rect 11605 19680 14431 19682
rect 11605 19624 11610 19680
rect 11666 19624 14370 19680
rect 14426 19624 14431 19680
rect 11605 19622 14431 19624
rect 11605 19619 11671 19622
rect 14365 19619 14431 19622
rect 14641 19682 14707 19685
rect 15653 19682 15719 19685
rect 14641 19680 15719 19682
rect 14641 19624 14646 19680
rect 14702 19624 15658 19680
rect 15714 19624 15719 19680
rect 14641 19622 15719 19624
rect 14641 19619 14707 19622
rect 15653 19619 15719 19622
rect 16941 19682 17007 19685
rect 18413 19682 18479 19685
rect 16941 19680 18479 19682
rect 16941 19624 16946 19680
rect 17002 19624 18418 19680
rect 18474 19624 18479 19680
rect 16941 19622 18479 19624
rect 16941 19619 17007 19622
rect 18413 19619 18479 19622
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 3141 19410 3207 19413
rect 19609 19410 19675 19413
rect 21541 19410 21607 19413
rect 3141 19408 21607 19410
rect 3141 19352 3146 19408
rect 3202 19352 19614 19408
rect 19670 19352 21546 19408
rect 21602 19352 21607 19408
rect 3141 19350 21607 19352
rect 3141 19347 3207 19350
rect 19609 19347 19675 19350
rect 21541 19347 21607 19350
rect 22553 19410 22619 19413
rect 23238 19410 23244 19412
rect 22553 19408 23244 19410
rect 22553 19352 22558 19408
rect 22614 19352 23244 19408
rect 22553 19350 23244 19352
rect 22553 19347 22619 19350
rect 23238 19348 23244 19350
rect 23308 19348 23314 19412
rect 10961 19274 11027 19277
rect 12433 19274 12499 19277
rect 10961 19272 12499 19274
rect 10961 19216 10966 19272
rect 11022 19216 12438 19272
rect 12494 19216 12499 19272
rect 10961 19214 12499 19216
rect 10961 19211 11027 19214
rect 12433 19211 12499 19214
rect 16430 19212 16436 19276
rect 16500 19274 16506 19276
rect 19241 19274 19307 19277
rect 16500 19272 19307 19274
rect 16500 19216 19246 19272
rect 19302 19216 19307 19272
rect 16500 19214 19307 19216
rect 16500 19212 16506 19214
rect 19241 19211 19307 19214
rect 11697 19138 11763 19141
rect 14273 19138 14339 19141
rect 11697 19136 14339 19138
rect 11697 19080 11702 19136
rect 11758 19080 14278 19136
rect 14334 19080 14339 19136
rect 11697 19078 14339 19080
rect 11697 19075 11763 19078
rect 14273 19075 14339 19078
rect 38285 19138 38351 19141
rect 38621 19138 39421 19168
rect 38285 19136 39421 19138
rect 38285 19080 38290 19136
rect 38346 19080 39421 19136
rect 38285 19078 39421 19080
rect 38285 19075 38351 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 38621 19048 39421 19078
rect 34930 19007 35246 19008
rect 10869 19002 10935 19005
rect 16297 19002 16363 19005
rect 10869 19000 16363 19002
rect 10869 18944 10874 19000
rect 10930 18944 16302 19000
rect 16358 18944 16363 19000
rect 10869 18942 16363 18944
rect 10869 18939 10935 18942
rect 16297 18939 16363 18942
rect 4870 18528 5186 18529
rect 0 18458 800 18488
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 933 18458 999 18461
rect 0 18456 999 18458
rect 0 18400 938 18456
rect 994 18400 999 18456
rect 0 18398 999 18400
rect 0 18368 800 18398
rect 933 18395 999 18398
rect 21817 18458 21883 18461
rect 28206 18458 28212 18460
rect 21817 18456 28212 18458
rect 21817 18400 21822 18456
rect 21878 18400 28212 18456
rect 21817 18398 28212 18400
rect 21817 18395 21883 18398
rect 28206 18396 28212 18398
rect 28276 18396 28282 18460
rect 13169 18322 13235 18325
rect 16389 18322 16455 18325
rect 19241 18324 19307 18325
rect 19190 18322 19196 18324
rect 13169 18320 16455 18322
rect 13169 18264 13174 18320
rect 13230 18264 16394 18320
rect 16450 18264 16455 18320
rect 13169 18262 16455 18264
rect 19150 18262 19196 18322
rect 19260 18320 19307 18324
rect 19302 18264 19307 18320
rect 13169 18259 13235 18262
rect 16389 18259 16455 18262
rect 19190 18260 19196 18262
rect 19260 18260 19307 18264
rect 19241 18259 19307 18260
rect 20897 18322 20963 18325
rect 28717 18322 28783 18325
rect 20897 18320 28783 18322
rect 20897 18264 20902 18320
rect 20958 18264 28722 18320
rect 28778 18264 28783 18320
rect 20897 18262 28783 18264
rect 20897 18259 20963 18262
rect 28717 18259 28783 18262
rect 16297 18186 16363 18189
rect 19149 18186 19215 18189
rect 16297 18184 19215 18186
rect 16297 18128 16302 18184
rect 16358 18128 19154 18184
rect 19210 18128 19215 18184
rect 16297 18126 19215 18128
rect 16297 18123 16363 18126
rect 19149 18123 19215 18126
rect 11145 18050 11211 18053
rect 14089 18050 14155 18053
rect 11145 18048 14155 18050
rect 11145 17992 11150 18048
rect 11206 17992 14094 18048
rect 14150 17992 14155 18048
rect 11145 17990 14155 17992
rect 11145 17987 11211 17990
rect 14089 17987 14155 17990
rect 16665 18050 16731 18053
rect 20805 18050 20871 18053
rect 16665 18048 20871 18050
rect 16665 17992 16670 18048
rect 16726 17992 20810 18048
rect 20866 17992 20871 18048
rect 16665 17990 20871 17992
rect 16665 17987 16731 17990
rect 20805 17987 20871 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 22921 17914 22987 17917
rect 22050 17912 22987 17914
rect 22050 17856 22926 17912
rect 22982 17856 22987 17912
rect 22050 17854 22987 17856
rect 10409 17778 10475 17781
rect 22050 17778 22110 17854
rect 22921 17851 22987 17854
rect 10409 17776 22110 17778
rect 10409 17720 10414 17776
rect 10470 17720 22110 17776
rect 10409 17718 22110 17720
rect 10409 17715 10475 17718
rect 18045 17642 18111 17645
rect 22921 17642 22987 17645
rect 18045 17640 22987 17642
rect 18045 17584 18050 17640
rect 18106 17584 22926 17640
rect 22982 17584 22987 17640
rect 18045 17582 22987 17584
rect 18045 17579 18111 17582
rect 22921 17579 22987 17582
rect 24025 17642 24091 17645
rect 27521 17642 27587 17645
rect 24025 17640 27587 17642
rect 24025 17584 24030 17640
rect 24086 17584 27526 17640
rect 27582 17584 27587 17640
rect 24025 17582 27587 17584
rect 24025 17579 24091 17582
rect 27521 17579 27587 17582
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 10501 17370 10567 17373
rect 12801 17370 12867 17373
rect 10501 17368 12867 17370
rect 10501 17312 10506 17368
rect 10562 17312 12806 17368
rect 12862 17312 12867 17368
rect 10501 17310 12867 17312
rect 10501 17307 10567 17310
rect 12801 17307 12867 17310
rect 11053 17234 11119 17237
rect 16849 17234 16915 17237
rect 11053 17232 16915 17234
rect 11053 17176 11058 17232
rect 11114 17176 16854 17232
rect 16910 17176 16915 17232
rect 11053 17174 16915 17176
rect 11053 17171 11119 17174
rect 16849 17171 16915 17174
rect 13537 17098 13603 17101
rect 16481 17098 16547 17101
rect 13537 17096 16547 17098
rect 13537 17040 13542 17096
rect 13598 17040 16486 17096
rect 16542 17040 16547 17096
rect 13537 17038 16547 17040
rect 13537 17035 13603 17038
rect 16481 17035 16547 17038
rect 14365 16962 14431 16965
rect 19149 16962 19215 16965
rect 14365 16960 19215 16962
rect 14365 16904 14370 16960
rect 14426 16904 19154 16960
rect 19210 16904 19215 16960
rect 14365 16902 19215 16904
rect 14365 16899 14431 16902
rect 19149 16899 19215 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 23381 16826 23447 16829
rect 30557 16826 30623 16829
rect 23381 16824 30623 16826
rect 23381 16768 23386 16824
rect 23442 16768 30562 16824
rect 30618 16768 30623 16824
rect 23381 16766 30623 16768
rect 23381 16763 23447 16766
rect 30557 16763 30623 16766
rect 19333 16690 19399 16693
rect 27521 16690 27587 16693
rect 28717 16692 28783 16693
rect 28717 16690 28764 16692
rect 19333 16688 27587 16690
rect 19333 16632 19338 16688
rect 19394 16632 27526 16688
rect 27582 16632 27587 16688
rect 19333 16630 27587 16632
rect 28672 16688 28764 16690
rect 28672 16632 28722 16688
rect 28672 16630 28764 16632
rect 19333 16627 19399 16630
rect 27521 16627 27587 16630
rect 28717 16628 28764 16630
rect 28828 16628 28834 16692
rect 28717 16627 28783 16628
rect 19793 16554 19859 16557
rect 24485 16554 24551 16557
rect 26325 16554 26391 16557
rect 19793 16552 26391 16554
rect 19793 16496 19798 16552
rect 19854 16496 24490 16552
rect 24546 16496 26330 16552
rect 26386 16496 26391 16552
rect 19793 16494 26391 16496
rect 19793 16491 19859 16494
rect 24485 16491 24551 16494
rect 26325 16491 26391 16494
rect 26734 16492 26740 16556
rect 26804 16554 26810 16556
rect 26877 16554 26943 16557
rect 26804 16552 26943 16554
rect 26804 16496 26882 16552
rect 26938 16496 26943 16552
rect 26804 16494 26943 16496
rect 26804 16492 26810 16494
rect 26877 16491 26943 16494
rect 0 16418 800 16448
rect 933 16418 999 16421
rect 0 16416 999 16418
rect 0 16360 938 16416
rect 994 16360 999 16416
rect 0 16358 999 16360
rect 0 16328 800 16358
rect 933 16355 999 16358
rect 13670 16356 13676 16420
rect 13740 16418 13746 16420
rect 18413 16418 18479 16421
rect 13740 16416 18479 16418
rect 13740 16360 18418 16416
rect 18474 16360 18479 16416
rect 13740 16358 18479 16360
rect 13740 16356 13746 16358
rect 18413 16355 18479 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 38621 16328 39421 16448
rect 35590 16287 35906 16288
rect 29821 16282 29887 16285
rect 30741 16282 30807 16285
rect 32029 16282 32095 16285
rect 29821 16280 32095 16282
rect 29821 16224 29826 16280
rect 29882 16224 30746 16280
rect 30802 16224 32034 16280
rect 32090 16224 32095 16280
rect 29821 16222 32095 16224
rect 29821 16219 29887 16222
rect 30741 16219 30807 16222
rect 32029 16219 32095 16222
rect 24301 16146 24367 16149
rect 25221 16146 25287 16149
rect 24301 16144 25287 16146
rect 24301 16088 24306 16144
rect 24362 16088 25226 16144
rect 25282 16088 25287 16144
rect 24301 16086 25287 16088
rect 24301 16083 24367 16086
rect 25221 16083 25287 16086
rect 25773 16146 25839 16149
rect 28073 16146 28139 16149
rect 25773 16144 28139 16146
rect 25773 16088 25778 16144
rect 25834 16088 28078 16144
rect 28134 16088 28139 16144
rect 25773 16086 28139 16088
rect 25773 16083 25839 16086
rect 28073 16083 28139 16086
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19241 15738 19307 15741
rect 21541 15738 21607 15741
rect 19241 15736 21607 15738
rect 19241 15680 19246 15736
rect 19302 15680 21546 15736
rect 21602 15680 21607 15736
rect 19241 15678 21607 15680
rect 19241 15675 19307 15678
rect 21541 15675 21607 15678
rect 25957 15738 26023 15741
rect 26785 15738 26851 15741
rect 25957 15736 26851 15738
rect 25957 15680 25962 15736
rect 26018 15680 26790 15736
rect 26846 15680 26851 15736
rect 25957 15678 26851 15680
rect 25957 15675 26023 15678
rect 26785 15675 26851 15678
rect 18413 15602 18479 15605
rect 19057 15602 19123 15605
rect 22553 15602 22619 15605
rect 18413 15600 19123 15602
rect 18413 15544 18418 15600
rect 18474 15544 19062 15600
rect 19118 15544 19123 15600
rect 18413 15542 19123 15544
rect 18413 15539 18479 15542
rect 19057 15539 19123 15542
rect 19290 15600 22619 15602
rect 19290 15544 22558 15600
rect 22614 15544 22619 15600
rect 19290 15542 22619 15544
rect 12065 15466 12131 15469
rect 17769 15466 17835 15469
rect 18413 15466 18479 15469
rect 19290 15466 19350 15542
rect 22553 15539 22619 15542
rect 22829 15602 22895 15605
rect 26325 15602 26391 15605
rect 22829 15600 26391 15602
rect 22829 15544 22834 15600
rect 22890 15544 26330 15600
rect 26386 15544 26391 15600
rect 22829 15542 26391 15544
rect 22829 15539 22895 15542
rect 26325 15539 26391 15542
rect 26877 15602 26943 15605
rect 27286 15602 27292 15604
rect 26877 15600 27292 15602
rect 26877 15544 26882 15600
rect 26938 15544 27292 15600
rect 26877 15542 27292 15544
rect 26877 15539 26943 15542
rect 27286 15540 27292 15542
rect 27356 15540 27362 15604
rect 12065 15464 19350 15466
rect 12065 15408 12070 15464
rect 12126 15408 17774 15464
rect 17830 15408 18418 15464
rect 18474 15408 19350 15464
rect 12065 15406 19350 15408
rect 23565 15466 23631 15469
rect 25773 15466 25839 15469
rect 26141 15466 26207 15469
rect 23565 15464 25839 15466
rect 23565 15408 23570 15464
rect 23626 15408 25778 15464
rect 25834 15408 25839 15464
rect 23565 15406 25839 15408
rect 12065 15403 12131 15406
rect 17769 15403 17835 15406
rect 18413 15403 18479 15406
rect 23565 15403 23631 15406
rect 25773 15403 25839 15406
rect 26006 15464 26207 15466
rect 26006 15408 26146 15464
rect 26202 15408 26207 15464
rect 26006 15406 26207 15408
rect 25262 15268 25268 15332
rect 25332 15330 25338 15332
rect 25497 15330 25563 15333
rect 25332 15328 25563 15330
rect 25332 15272 25502 15328
rect 25558 15272 25563 15328
rect 25332 15270 25563 15272
rect 25332 15268 25338 15270
rect 25497 15267 25563 15270
rect 25773 15330 25839 15333
rect 26006 15330 26066 15406
rect 26141 15403 26207 15406
rect 25773 15328 26066 15330
rect 25773 15272 25778 15328
rect 25834 15272 26066 15328
rect 25773 15270 26066 15272
rect 25773 15267 25839 15270
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 11462 15132 11468 15196
rect 11532 15194 11538 15196
rect 11697 15194 11763 15197
rect 17493 15196 17559 15197
rect 17493 15194 17540 15196
rect 11532 15192 11763 15194
rect 11532 15136 11702 15192
rect 11758 15136 11763 15192
rect 11532 15134 11763 15136
rect 17448 15192 17540 15194
rect 17448 15136 17498 15192
rect 17448 15134 17540 15136
rect 11532 15132 11538 15134
rect 11697 15131 11763 15134
rect 17493 15132 17540 15134
rect 17604 15132 17610 15196
rect 17769 15194 17835 15197
rect 20621 15194 20687 15197
rect 17769 15192 20687 15194
rect 17769 15136 17774 15192
rect 17830 15136 20626 15192
rect 20682 15136 20687 15192
rect 17769 15134 20687 15136
rect 17493 15131 17559 15132
rect 17769 15131 17835 15134
rect 20621 15131 20687 15134
rect 11053 15058 11119 15061
rect 30097 15058 30163 15061
rect 11053 15056 30163 15058
rect 11053 15000 11058 15056
rect 11114 15000 30102 15056
rect 30158 15000 30163 15056
rect 11053 14998 30163 15000
rect 11053 14995 11119 14998
rect 30097 14995 30163 14998
rect 16941 14922 17007 14925
rect 21909 14922 21975 14925
rect 27889 14922 27955 14925
rect 16941 14920 27955 14922
rect 16941 14864 16946 14920
rect 17002 14864 21914 14920
rect 21970 14864 27894 14920
rect 27950 14864 27955 14920
rect 16941 14862 27955 14864
rect 16941 14859 17007 14862
rect 21909 14859 21975 14862
rect 27889 14859 27955 14862
rect 11513 14786 11579 14789
rect 11646 14786 11652 14788
rect 11513 14784 11652 14786
rect 11513 14728 11518 14784
rect 11574 14728 11652 14784
rect 11513 14726 11652 14728
rect 11513 14723 11579 14726
rect 11646 14724 11652 14726
rect 11716 14724 11722 14788
rect 19701 14786 19767 14789
rect 20621 14786 20687 14789
rect 19701 14784 20687 14786
rect 19701 14728 19706 14784
rect 19762 14728 20626 14784
rect 20682 14728 20687 14784
rect 19701 14726 20687 14728
rect 19701 14723 19767 14726
rect 20621 14723 20687 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 20253 14650 20319 14653
rect 23933 14650 23999 14653
rect 20253 14648 23999 14650
rect 20253 14592 20258 14648
rect 20314 14592 23938 14648
rect 23994 14592 23999 14648
rect 20253 14590 23999 14592
rect 20253 14587 20319 14590
rect 23933 14587 23999 14590
rect 19149 14516 19215 14517
rect 19149 14514 19196 14516
rect 19104 14512 19196 14514
rect 19104 14456 19154 14512
rect 19104 14454 19196 14456
rect 19149 14452 19196 14454
rect 19260 14452 19266 14516
rect 19149 14451 19215 14452
rect 19977 14378 20043 14381
rect 25405 14378 25471 14381
rect 19977 14376 25471 14378
rect 19977 14320 19982 14376
rect 20038 14320 25410 14376
rect 25466 14320 25471 14376
rect 19977 14318 25471 14320
rect 19977 14315 20043 14318
rect 25405 14315 25471 14318
rect 38285 14378 38351 14381
rect 38621 14378 39421 14408
rect 38285 14376 39421 14378
rect 38285 14320 38290 14376
rect 38346 14320 39421 14376
rect 38285 14318 39421 14320
rect 38285 14315 38351 14318
rect 38621 14288 39421 14318
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 28257 13970 28323 13973
rect 28390 13970 28396 13972
rect 28257 13968 28396 13970
rect 28257 13912 28262 13968
rect 28318 13912 28396 13968
rect 28257 13910 28396 13912
rect 28257 13907 28323 13910
rect 28390 13908 28396 13910
rect 28460 13908 28466 13972
rect 17769 13834 17835 13837
rect 24301 13834 24367 13837
rect 17769 13832 24367 13834
rect 17769 13776 17774 13832
rect 17830 13776 24306 13832
rect 24362 13776 24367 13832
rect 17769 13774 24367 13776
rect 17769 13771 17835 13774
rect 24301 13771 24367 13774
rect 0 13698 800 13728
rect 1485 13698 1551 13701
rect 0 13696 1551 13698
rect 0 13640 1490 13696
rect 1546 13640 1551 13696
rect 0 13638 1551 13640
rect 0 13608 800 13638
rect 1485 13635 1551 13638
rect 10869 13698 10935 13701
rect 23473 13698 23539 13701
rect 10869 13696 23539 13698
rect 10869 13640 10874 13696
rect 10930 13640 23478 13696
rect 23534 13640 23539 13696
rect 10869 13638 23539 13640
rect 10869 13635 10935 13638
rect 23473 13635 23539 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 11881 13426 11947 13429
rect 12014 13426 12020 13428
rect 11881 13424 12020 13426
rect 11881 13368 11886 13424
rect 11942 13368 12020 13424
rect 11881 13366 12020 13368
rect 11881 13363 11947 13366
rect 12014 13364 12020 13366
rect 12084 13426 12090 13428
rect 16113 13426 16179 13429
rect 12084 13424 16179 13426
rect 12084 13368 16118 13424
rect 16174 13368 16179 13424
rect 12084 13366 16179 13368
rect 12084 13364 12090 13366
rect 16113 13363 16179 13366
rect 20161 13426 20227 13429
rect 30373 13426 30439 13429
rect 20161 13424 30439 13426
rect 20161 13368 20166 13424
rect 20222 13368 30378 13424
rect 30434 13368 30439 13424
rect 20161 13366 30439 13368
rect 20161 13363 20227 13366
rect 30373 13363 30439 13366
rect 10777 13290 10843 13293
rect 25773 13290 25839 13293
rect 10777 13288 25839 13290
rect 10777 13232 10782 13288
rect 10838 13232 25778 13288
rect 25834 13232 25839 13288
rect 10777 13230 25839 13232
rect 10777 13227 10843 13230
rect 25773 13227 25839 13230
rect 14549 13154 14615 13157
rect 14774 13154 14780 13156
rect 14549 13152 14780 13154
rect 14549 13096 14554 13152
rect 14610 13096 14780 13152
rect 14549 13094 14780 13096
rect 14549 13091 14615 13094
rect 14774 13092 14780 13094
rect 14844 13092 14850 13156
rect 20253 13154 20319 13157
rect 24853 13154 24919 13157
rect 25129 13154 25195 13157
rect 20253 13152 22110 13154
rect 20253 13096 20258 13152
rect 20314 13096 22110 13152
rect 20253 13094 22110 13096
rect 20253 13091 20319 13094
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 14181 13018 14247 13021
rect 20161 13018 20227 13021
rect 14181 13016 20227 13018
rect 14181 12960 14186 13016
rect 14242 12960 20166 13016
rect 20222 12960 20227 13016
rect 14181 12958 20227 12960
rect 14181 12955 14247 12958
rect 20161 12955 20227 12958
rect 11973 12882 12039 12885
rect 16941 12882 17007 12885
rect 11973 12880 17007 12882
rect 11973 12824 11978 12880
rect 12034 12824 16946 12880
rect 17002 12824 17007 12880
rect 11973 12822 17007 12824
rect 11973 12819 12039 12822
rect 16941 12819 17007 12822
rect 22050 12746 22110 13094
rect 24853 13152 25195 13154
rect 24853 13096 24858 13152
rect 24914 13096 25134 13152
rect 25190 13096 25195 13152
rect 24853 13094 25195 13096
rect 24853 13091 24919 13094
rect 25129 13091 25195 13094
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 25313 13018 25379 13021
rect 26417 13018 26483 13021
rect 26969 13018 27035 13021
rect 25313 13016 26066 13018
rect 25313 12960 25318 13016
rect 25374 12960 26066 13016
rect 25313 12958 26066 12960
rect 25313 12955 25379 12958
rect 22553 12882 22619 12885
rect 25037 12882 25103 12885
rect 26006 12882 26066 12958
rect 26417 13016 27035 13018
rect 26417 12960 26422 13016
rect 26478 12960 26974 13016
rect 27030 12960 27035 13016
rect 26417 12958 27035 12960
rect 26417 12955 26483 12958
rect 26969 12955 27035 12958
rect 26417 12882 26483 12885
rect 22553 12880 25882 12882
rect 22553 12824 22558 12880
rect 22614 12824 25042 12880
rect 25098 12824 25882 12880
rect 22553 12822 25882 12824
rect 26006 12880 26483 12882
rect 26006 12824 26422 12880
rect 26478 12824 26483 12880
rect 26006 12822 26483 12824
rect 22553 12819 22619 12822
rect 25037 12819 25103 12822
rect 24301 12746 24367 12749
rect 25630 12746 25636 12748
rect 22050 12744 25636 12746
rect 22050 12688 24306 12744
rect 24362 12688 25636 12744
rect 22050 12686 25636 12688
rect 24301 12683 24367 12686
rect 25630 12684 25636 12686
rect 25700 12684 25706 12748
rect 22277 12612 22343 12613
rect 22277 12608 22324 12612
rect 22388 12610 22394 12612
rect 22277 12552 22282 12608
rect 22277 12548 22324 12552
rect 22388 12550 22434 12610
rect 22388 12548 22394 12550
rect 25262 12548 25268 12612
rect 25332 12610 25338 12612
rect 25405 12610 25471 12613
rect 25332 12608 25471 12610
rect 25332 12552 25410 12608
rect 25466 12552 25471 12608
rect 25332 12550 25471 12552
rect 25332 12548 25338 12550
rect 22277 12547 22343 12548
rect 25405 12547 25471 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 8201 12474 8267 12477
rect 10869 12474 10935 12477
rect 8201 12472 10935 12474
rect 8201 12416 8206 12472
rect 8262 12416 10874 12472
rect 10930 12416 10935 12472
rect 8201 12414 10935 12416
rect 8201 12411 8267 12414
rect 10869 12411 10935 12414
rect 15377 12474 15443 12477
rect 18321 12474 18387 12477
rect 15377 12472 18387 12474
rect 15377 12416 15382 12472
rect 15438 12416 18326 12472
rect 18382 12416 18387 12472
rect 15377 12414 18387 12416
rect 15377 12411 15443 12414
rect 18321 12411 18387 12414
rect 25497 12474 25563 12477
rect 25822 12474 25882 12822
rect 26417 12819 26483 12822
rect 28993 12746 29059 12749
rect 29821 12746 29887 12749
rect 33593 12746 33659 12749
rect 28993 12744 33659 12746
rect 28993 12688 28998 12744
rect 29054 12688 29826 12744
rect 29882 12688 33598 12744
rect 33654 12688 33659 12744
rect 28993 12686 33659 12688
rect 28993 12683 29059 12686
rect 29821 12683 29887 12686
rect 33593 12683 33659 12686
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 25497 12472 25882 12474
rect 25497 12416 25502 12472
rect 25558 12416 25882 12472
rect 25497 12414 25882 12416
rect 25497 12411 25563 12414
rect 15377 12338 15443 12341
rect 16849 12338 16915 12341
rect 15377 12336 16915 12338
rect 15377 12280 15382 12336
rect 15438 12280 16854 12336
rect 16910 12280 16915 12336
rect 15377 12278 16915 12280
rect 15377 12275 15443 12278
rect 16849 12275 16915 12278
rect 25814 12276 25820 12340
rect 25884 12338 25890 12340
rect 26509 12338 26575 12341
rect 25884 12336 26575 12338
rect 25884 12280 26514 12336
rect 26570 12280 26575 12336
rect 25884 12278 26575 12280
rect 25884 12276 25890 12278
rect 26509 12275 26575 12278
rect 30966 12276 30972 12340
rect 31036 12338 31042 12340
rect 37641 12338 37707 12341
rect 31036 12336 37707 12338
rect 31036 12280 37646 12336
rect 37702 12280 37707 12336
rect 31036 12278 37707 12280
rect 31036 12276 31042 12278
rect 37641 12275 37707 12278
rect 15837 12202 15903 12205
rect 16430 12202 16436 12204
rect 15837 12200 16436 12202
rect 15837 12144 15842 12200
rect 15898 12144 16436 12200
rect 15837 12142 16436 12144
rect 15837 12139 15903 12142
rect 16430 12140 16436 12142
rect 16500 12140 16506 12204
rect 22369 12202 22435 12205
rect 28165 12202 28231 12205
rect 28625 12202 28691 12205
rect 22369 12200 28691 12202
rect 22369 12144 22374 12200
rect 22430 12144 28170 12200
rect 28226 12144 28630 12200
rect 28686 12144 28691 12200
rect 22369 12142 28691 12144
rect 22369 12139 22435 12142
rect 28165 12139 28231 12142
rect 28625 12139 28691 12142
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 22093 11930 22159 11933
rect 25037 11930 25103 11933
rect 22093 11928 25103 11930
rect 22093 11872 22098 11928
rect 22154 11872 25042 11928
rect 25098 11872 25103 11928
rect 22093 11870 25103 11872
rect 22093 11867 22159 11870
rect 25037 11867 25103 11870
rect 28758 11868 28764 11932
rect 28828 11930 28834 11932
rect 29361 11930 29427 11933
rect 28828 11928 29427 11930
rect 28828 11872 29366 11928
rect 29422 11872 29427 11928
rect 28828 11870 29427 11872
rect 28828 11868 28834 11870
rect 29361 11867 29427 11870
rect 13629 11794 13695 11797
rect 18413 11794 18479 11797
rect 13629 11792 18479 11794
rect 13629 11736 13634 11792
rect 13690 11736 18418 11792
rect 18474 11736 18479 11792
rect 13629 11734 18479 11736
rect 13629 11731 13695 11734
rect 18413 11731 18479 11734
rect 20069 11796 20135 11797
rect 20069 11792 20116 11796
rect 20180 11794 20186 11796
rect 24117 11794 24183 11797
rect 28390 11794 28396 11796
rect 20069 11736 20074 11792
rect 20069 11732 20116 11736
rect 20180 11734 20226 11794
rect 24117 11792 28396 11794
rect 24117 11736 24122 11792
rect 24178 11736 28396 11792
rect 24117 11734 28396 11736
rect 20180 11732 20186 11734
rect 20069 11731 20135 11732
rect 24117 11731 24183 11734
rect 28390 11732 28396 11734
rect 28460 11732 28466 11796
rect 0 11658 800 11688
rect 933 11658 999 11661
rect 0 11656 999 11658
rect 0 11600 938 11656
rect 994 11600 999 11656
rect 0 11598 999 11600
rect 0 11568 800 11598
rect 933 11595 999 11598
rect 4061 11658 4127 11661
rect 13118 11658 13124 11660
rect 4061 11656 13124 11658
rect 4061 11600 4066 11656
rect 4122 11600 13124 11656
rect 4061 11598 13124 11600
rect 4061 11595 4127 11598
rect 13118 11596 13124 11598
rect 13188 11596 13194 11660
rect 15653 11658 15719 11661
rect 18229 11658 18295 11661
rect 15653 11656 18295 11658
rect 15653 11600 15658 11656
rect 15714 11600 18234 11656
rect 18290 11600 18295 11656
rect 15653 11598 18295 11600
rect 15653 11595 15719 11598
rect 18229 11595 18295 11598
rect 21909 11658 21975 11661
rect 24393 11658 24459 11661
rect 25497 11658 25563 11661
rect 21909 11656 25563 11658
rect 21909 11600 21914 11656
rect 21970 11600 24398 11656
rect 24454 11600 25502 11656
rect 25558 11600 25563 11656
rect 21909 11598 25563 11600
rect 21909 11595 21975 11598
rect 24393 11595 24459 11598
rect 25497 11595 25563 11598
rect 37825 11658 37891 11661
rect 38621 11658 39421 11688
rect 37825 11656 39421 11658
rect 37825 11600 37830 11656
rect 37886 11600 39421 11656
rect 37825 11598 39421 11600
rect 37825 11595 37891 11598
rect 38621 11568 39421 11598
rect 15009 11522 15075 11525
rect 23473 11522 23539 11525
rect 15009 11520 23539 11522
rect 15009 11464 15014 11520
rect 15070 11464 23478 11520
rect 23534 11464 23539 11520
rect 15009 11462 23539 11464
rect 15009 11459 15075 11462
rect 23473 11459 23539 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 16297 11386 16363 11389
rect 18597 11386 18663 11389
rect 16297 11384 18663 11386
rect 16297 11328 16302 11384
rect 16358 11328 18602 11384
rect 18658 11328 18663 11384
rect 16297 11326 18663 11328
rect 16297 11323 16363 11326
rect 18597 11323 18663 11326
rect 13813 11250 13879 11253
rect 14917 11250 14983 11253
rect 21817 11250 21883 11253
rect 13813 11248 13922 11250
rect 13813 11192 13818 11248
rect 13874 11192 13922 11248
rect 13813 11187 13922 11192
rect 14917 11248 21883 11250
rect 14917 11192 14922 11248
rect 14978 11192 21822 11248
rect 21878 11192 21883 11248
rect 14917 11190 21883 11192
rect 14917 11187 14983 11190
rect 21817 11187 21883 11190
rect 13862 11116 13922 11187
rect 13854 11052 13860 11116
rect 13924 11052 13930 11116
rect 15561 11114 15627 11117
rect 16297 11114 16363 11117
rect 21449 11114 21515 11117
rect 22093 11116 22159 11117
rect 22093 11114 22140 11116
rect 15561 11112 21515 11114
rect 15561 11056 15566 11112
rect 15622 11056 16302 11112
rect 16358 11056 21454 11112
rect 21510 11056 21515 11112
rect 15561 11054 21515 11056
rect 22012 11112 22140 11114
rect 22204 11114 22210 11116
rect 25497 11114 25563 11117
rect 26325 11114 26391 11117
rect 22204 11112 26391 11114
rect 22012 11056 22098 11112
rect 22204 11056 25502 11112
rect 25558 11056 26330 11112
rect 26386 11056 26391 11112
rect 22012 11054 22140 11056
rect 15561 11051 15627 11054
rect 16297 11051 16363 11054
rect 21449 11051 21515 11054
rect 22093 11052 22140 11054
rect 22204 11054 26391 11056
rect 22204 11052 22210 11054
rect 22093 11051 22159 11052
rect 25497 11051 25563 11054
rect 26325 11051 26391 11054
rect 14457 10978 14523 10981
rect 19885 10978 19951 10981
rect 14457 10976 19951 10978
rect 14457 10920 14462 10976
rect 14518 10920 19890 10976
rect 19946 10920 19951 10976
rect 14457 10918 19951 10920
rect 14457 10915 14523 10918
rect 19885 10915 19951 10918
rect 22093 10978 22159 10981
rect 22502 10978 22508 10980
rect 22093 10976 22508 10978
rect 22093 10920 22098 10976
rect 22154 10920 22508 10976
rect 22093 10918 22508 10920
rect 22093 10915 22159 10918
rect 22502 10916 22508 10918
rect 22572 10916 22578 10980
rect 24761 10978 24827 10981
rect 27061 10978 27127 10981
rect 24761 10976 27127 10978
rect 24761 10920 24766 10976
rect 24822 10920 27066 10976
rect 27122 10920 27127 10976
rect 24761 10918 27127 10920
rect 24761 10915 24827 10918
rect 27061 10915 27127 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 35590 10847 35906 10848
rect 14549 10842 14615 10845
rect 16113 10842 16179 10845
rect 18965 10842 19031 10845
rect 14549 10840 16179 10842
rect 14549 10784 14554 10840
rect 14610 10784 16118 10840
rect 16174 10784 16179 10840
rect 14549 10782 16179 10784
rect 14549 10779 14615 10782
rect 16113 10779 16179 10782
rect 16254 10840 19031 10842
rect 16254 10784 18970 10840
rect 19026 10784 19031 10840
rect 16254 10782 19031 10784
rect 11145 10706 11211 10709
rect 13353 10706 13419 10709
rect 11145 10704 13419 10706
rect 11145 10648 11150 10704
rect 11206 10648 13358 10704
rect 13414 10648 13419 10704
rect 11145 10646 13419 10648
rect 11145 10643 11211 10646
rect 13353 10643 13419 10646
rect 15469 10706 15535 10709
rect 16254 10706 16314 10782
rect 18965 10779 19031 10782
rect 21265 10842 21331 10845
rect 23473 10842 23539 10845
rect 21265 10840 23539 10842
rect 21265 10784 21270 10840
rect 21326 10784 23478 10840
rect 23534 10784 23539 10840
rect 21265 10782 23539 10784
rect 21265 10779 21331 10782
rect 23473 10779 23539 10782
rect 25497 10842 25563 10845
rect 25957 10842 26023 10845
rect 28809 10842 28875 10845
rect 25497 10840 26023 10842
rect 25497 10784 25502 10840
rect 25558 10784 25962 10840
rect 26018 10784 26023 10840
rect 25497 10782 26023 10784
rect 25497 10779 25563 10782
rect 25957 10779 26023 10782
rect 28766 10840 28875 10842
rect 28766 10784 28814 10840
rect 28870 10784 28875 10840
rect 28766 10779 28875 10784
rect 16849 10706 16915 10709
rect 22553 10708 22619 10709
rect 22502 10706 22508 10708
rect 15469 10704 16314 10706
rect 15469 10648 15474 10704
rect 15530 10648 16314 10704
rect 15469 10646 16314 10648
rect 16392 10704 16915 10706
rect 16392 10648 16854 10704
rect 16910 10648 16915 10704
rect 16392 10646 16915 10648
rect 22462 10646 22508 10706
rect 22572 10704 22619 10708
rect 22614 10648 22619 10704
rect 15469 10643 15535 10646
rect 11789 10570 11855 10573
rect 12198 10570 12204 10572
rect 11789 10568 12204 10570
rect 11789 10512 11794 10568
rect 11850 10512 12204 10568
rect 11789 10510 12204 10512
rect 11789 10507 11855 10510
rect 12198 10508 12204 10510
rect 12268 10508 12274 10572
rect 15193 10570 15259 10573
rect 16392 10570 16452 10646
rect 16849 10643 16915 10646
rect 22502 10644 22508 10646
rect 22572 10644 22619 10648
rect 22553 10643 22619 10644
rect 15193 10568 16452 10570
rect 15193 10512 15198 10568
rect 15254 10512 16452 10568
rect 15193 10510 16452 10512
rect 16941 10570 17007 10573
rect 18873 10570 18939 10573
rect 16941 10568 18939 10570
rect 16941 10512 16946 10568
rect 17002 10512 18878 10568
rect 18934 10512 18939 10568
rect 16941 10510 18939 10512
rect 15193 10507 15259 10510
rect 16941 10507 17007 10510
rect 18873 10507 18939 10510
rect 23657 10570 23723 10573
rect 28766 10570 28826 10779
rect 28901 10570 28967 10573
rect 23657 10568 28967 10570
rect 23657 10512 23662 10568
rect 23718 10512 28906 10568
rect 28962 10512 28967 10568
rect 23657 10510 28967 10512
rect 23657 10507 23723 10510
rect 28901 10507 28967 10510
rect 25405 10434 25471 10437
rect 31661 10434 31727 10437
rect 25405 10432 31727 10434
rect 25405 10376 25410 10432
rect 25466 10376 31666 10432
rect 31722 10376 31727 10432
rect 25405 10374 31727 10376
rect 25405 10371 25471 10374
rect 31661 10371 31727 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 12617 10298 12683 10301
rect 22737 10298 22803 10301
rect 23841 10298 23907 10301
rect 11884 10296 23907 10298
rect 11884 10240 12622 10296
rect 12678 10240 22742 10296
rect 22798 10240 23846 10296
rect 23902 10240 23907 10296
rect 11884 10238 23907 10240
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 11884 9754 11944 10238
rect 12617 10235 12683 10238
rect 22737 10235 22803 10238
rect 23841 10235 23907 10238
rect 27337 10298 27403 10301
rect 28533 10298 28599 10301
rect 27337 10296 28599 10298
rect 27337 10240 27342 10296
rect 27398 10240 28538 10296
rect 28594 10240 28599 10296
rect 27337 10238 28599 10240
rect 27337 10235 27403 10238
rect 28533 10235 28599 10238
rect 13077 10162 13143 10165
rect 19609 10162 19675 10165
rect 22921 10162 22987 10165
rect 25589 10164 25655 10165
rect 25589 10162 25636 10164
rect 13077 10160 22987 10162
rect 13077 10104 13082 10160
rect 13138 10104 19614 10160
rect 19670 10104 22926 10160
rect 22982 10104 22987 10160
rect 13077 10102 22987 10104
rect 25544 10160 25636 10162
rect 25544 10104 25594 10160
rect 25544 10102 25636 10104
rect 13077 10099 13143 10102
rect 19609 10099 19675 10102
rect 22921 10099 22987 10102
rect 25589 10100 25636 10102
rect 25700 10100 25706 10164
rect 27889 10162 27955 10165
rect 28625 10162 28691 10165
rect 27889 10160 28691 10162
rect 27889 10104 27894 10160
rect 27950 10104 28630 10160
rect 28686 10104 28691 10160
rect 27889 10102 28691 10104
rect 25589 10099 25655 10100
rect 27889 10099 27955 10102
rect 28625 10099 28691 10102
rect 17401 10026 17467 10029
rect 18873 10026 18939 10029
rect 17401 10024 18939 10026
rect 17401 9968 17406 10024
rect 17462 9968 18878 10024
rect 18934 9968 18939 10024
rect 17401 9966 18939 9968
rect 17401 9963 17467 9966
rect 18873 9963 18939 9966
rect 21541 10026 21607 10029
rect 24853 10026 24919 10029
rect 28441 10028 28507 10029
rect 21541 10024 24919 10026
rect 21541 9968 21546 10024
rect 21602 9968 24858 10024
rect 24914 9968 24919 10024
rect 21541 9966 24919 9968
rect 21541 9963 21607 9966
rect 24853 9963 24919 9966
rect 28390 9964 28396 10028
rect 28460 10026 28507 10028
rect 28460 10024 28552 10026
rect 28502 9968 28552 10024
rect 28460 9966 28552 9968
rect 28460 9964 28507 9966
rect 28441 9963 28507 9964
rect 14273 9890 14339 9893
rect 16941 9890 17007 9893
rect 14273 9888 17007 9890
rect 14273 9832 14278 9888
rect 14334 9832 16946 9888
rect 17002 9832 17007 9888
rect 14273 9830 17007 9832
rect 14273 9827 14339 9830
rect 16941 9827 17007 9830
rect 21725 9890 21791 9893
rect 26049 9890 26115 9893
rect 21725 9888 26115 9890
rect 21725 9832 21730 9888
rect 21786 9832 26054 9888
rect 26110 9832 26115 9888
rect 21725 9830 26115 9832
rect 21725 9827 21791 9830
rect 26049 9827 26115 9830
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 11838 9694 11944 9754
rect 17033 9754 17099 9757
rect 21265 9754 21331 9757
rect 17033 9752 21331 9754
rect 17033 9696 17038 9752
rect 17094 9696 21270 9752
rect 21326 9696 21331 9752
rect 17033 9694 21331 9696
rect 11145 9618 11211 9621
rect 11462 9618 11468 9620
rect 11145 9616 11468 9618
rect 11145 9560 11150 9616
rect 11206 9560 11468 9616
rect 11145 9558 11468 9560
rect 11145 9555 11211 9558
rect 11462 9556 11468 9558
rect 11532 9556 11538 9620
rect 11237 9482 11303 9485
rect 11421 9482 11487 9485
rect 11237 9480 11487 9482
rect 11237 9424 11242 9480
rect 11298 9424 11426 9480
rect 11482 9424 11487 9480
rect 11237 9422 11487 9424
rect 11838 9482 11898 9694
rect 17033 9691 17099 9694
rect 21265 9691 21331 9694
rect 25681 9754 25747 9757
rect 25998 9754 26004 9756
rect 25681 9752 26004 9754
rect 25681 9696 25686 9752
rect 25742 9696 26004 9752
rect 25681 9694 26004 9696
rect 25681 9691 25747 9694
rect 25998 9692 26004 9694
rect 26068 9692 26074 9756
rect 13118 9556 13124 9620
rect 13188 9618 13194 9620
rect 13905 9618 13971 9621
rect 13188 9616 13971 9618
rect 13188 9560 13910 9616
rect 13966 9560 13971 9616
rect 13188 9558 13971 9560
rect 13188 9556 13194 9558
rect 13905 9555 13971 9558
rect 18505 9618 18571 9621
rect 22645 9620 22711 9621
rect 18638 9618 18644 9620
rect 18505 9616 18644 9618
rect 18505 9560 18510 9616
rect 18566 9560 18644 9616
rect 18505 9558 18644 9560
rect 18505 9555 18571 9558
rect 18638 9556 18644 9558
rect 18708 9556 18714 9620
rect 22645 9618 22692 9620
rect 22600 9616 22692 9618
rect 22600 9560 22650 9616
rect 22600 9558 22692 9560
rect 22645 9556 22692 9558
rect 22756 9556 22762 9620
rect 24669 9618 24735 9621
rect 25129 9618 25195 9621
rect 24669 9616 25195 9618
rect 24669 9560 24674 9616
rect 24730 9560 25134 9616
rect 25190 9560 25195 9616
rect 24669 9558 25195 9560
rect 22645 9555 22711 9556
rect 24669 9555 24735 9558
rect 25129 9555 25195 9558
rect 25814 9556 25820 9620
rect 25884 9618 25890 9620
rect 26141 9618 26207 9621
rect 25884 9616 26207 9618
rect 25884 9560 26146 9616
rect 26202 9560 26207 9616
rect 25884 9558 26207 9560
rect 25884 9556 25890 9558
rect 26141 9555 26207 9558
rect 26785 9618 26851 9621
rect 27102 9618 27108 9620
rect 26785 9616 27108 9618
rect 26785 9560 26790 9616
rect 26846 9560 27108 9616
rect 26785 9558 27108 9560
rect 26785 9555 26851 9558
rect 27102 9556 27108 9558
rect 27172 9556 27178 9620
rect 28993 9618 29059 9621
rect 29126 9618 29132 9620
rect 28993 9616 29132 9618
rect 28993 9560 28998 9616
rect 29054 9560 29132 9616
rect 28993 9558 29132 9560
rect 28993 9555 29059 9558
rect 29126 9556 29132 9558
rect 29196 9556 29202 9620
rect 38621 9528 39421 9648
rect 11973 9482 12039 9485
rect 13721 9484 13787 9485
rect 11838 9480 12039 9482
rect 11838 9424 11978 9480
rect 12034 9424 12039 9480
rect 11838 9422 12039 9424
rect 11237 9419 11303 9422
rect 11421 9419 11487 9422
rect 11973 9419 12039 9422
rect 13670 9420 13676 9484
rect 13740 9482 13787 9484
rect 16481 9482 16547 9485
rect 29545 9482 29611 9485
rect 13740 9480 13832 9482
rect 13782 9424 13832 9480
rect 13740 9422 13832 9424
rect 16481 9480 29611 9482
rect 16481 9424 16486 9480
rect 16542 9424 29550 9480
rect 29606 9424 29611 9480
rect 16481 9422 29611 9424
rect 13740 9420 13787 9422
rect 13721 9419 13787 9420
rect 16481 9419 16547 9422
rect 29545 9419 29611 9422
rect 12433 9346 12499 9349
rect 13537 9346 13603 9349
rect 12433 9344 28090 9346
rect 12433 9288 12438 9344
rect 12494 9288 13542 9344
rect 13598 9288 28090 9344
rect 12433 9286 28090 9288
rect 12433 9283 12499 9286
rect 13537 9283 13603 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 12065 9212 12131 9213
rect 12014 9148 12020 9212
rect 12084 9210 12131 9212
rect 12084 9208 12176 9210
rect 12126 9152 12176 9208
rect 12084 9150 12176 9152
rect 12084 9148 12131 9150
rect 14774 9148 14780 9212
rect 14844 9210 14850 9212
rect 14917 9210 14983 9213
rect 14844 9208 14983 9210
rect 14844 9152 14922 9208
rect 14978 9152 14983 9208
rect 14844 9150 14983 9152
rect 14844 9148 14850 9150
rect 12065 9147 12131 9148
rect 14917 9147 14983 9150
rect 19609 9210 19675 9213
rect 20989 9212 21055 9213
rect 19742 9210 19748 9212
rect 19609 9208 19748 9210
rect 19609 9152 19614 9208
rect 19670 9152 19748 9208
rect 19609 9150 19748 9152
rect 19609 9147 19675 9150
rect 19742 9148 19748 9150
rect 19812 9148 19818 9212
rect 20989 9210 21036 9212
rect 20944 9208 21036 9210
rect 20944 9152 20994 9208
rect 20944 9150 21036 9152
rect 20989 9148 21036 9150
rect 21100 9148 21106 9212
rect 21950 9148 21956 9212
rect 22020 9210 22026 9212
rect 24393 9210 24459 9213
rect 22020 9208 24459 9210
rect 22020 9152 24398 9208
rect 24454 9152 24459 9208
rect 22020 9150 24459 9152
rect 28030 9210 28090 9286
rect 28206 9284 28212 9348
rect 28276 9346 28282 9348
rect 29821 9346 29887 9349
rect 28276 9344 29887 9346
rect 28276 9288 29826 9344
rect 29882 9288 29887 9344
rect 28276 9286 29887 9288
rect 28276 9284 28282 9286
rect 29821 9283 29887 9286
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 30281 9210 30347 9213
rect 28030 9208 30347 9210
rect 28030 9152 30286 9208
rect 30342 9152 30347 9208
rect 28030 9150 30347 9152
rect 22020 9148 22026 9150
rect 20989 9147 21055 9148
rect 24393 9147 24459 9150
rect 30281 9147 30347 9150
rect 17309 9074 17375 9077
rect 18229 9074 18295 9077
rect 17309 9072 18295 9074
rect 17309 9016 17314 9072
rect 17370 9016 18234 9072
rect 18290 9016 18295 9072
rect 17309 9014 18295 9016
rect 17309 9011 17375 9014
rect 18229 9011 18295 9014
rect 19241 9074 19307 9077
rect 20529 9074 20595 9077
rect 19241 9072 20595 9074
rect 19241 9016 19246 9072
rect 19302 9016 20534 9072
rect 20590 9016 20595 9072
rect 19241 9014 20595 9016
rect 19241 9011 19307 9014
rect 20529 9011 20595 9014
rect 21173 9074 21239 9077
rect 27705 9074 27771 9077
rect 21173 9072 27771 9074
rect 21173 9016 21178 9072
rect 21234 9016 27710 9072
rect 27766 9016 27771 9072
rect 21173 9014 27771 9016
rect 21173 9011 21239 9014
rect 27705 9011 27771 9014
rect 0 8848 800 8968
rect 19609 8938 19675 8941
rect 20805 8938 20871 8941
rect 19609 8936 20871 8938
rect 19609 8880 19614 8936
rect 19670 8880 20810 8936
rect 20866 8880 20871 8936
rect 19609 8878 20871 8880
rect 19609 8875 19675 8878
rect 20805 8875 20871 8878
rect 21265 8938 21331 8941
rect 23749 8938 23815 8941
rect 21265 8936 23815 8938
rect 21265 8880 21270 8936
rect 21326 8880 23754 8936
rect 23810 8880 23815 8936
rect 21265 8878 23815 8880
rect 21265 8875 21331 8878
rect 23749 8875 23815 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 20437 8666 20503 8669
rect 23013 8666 23079 8669
rect 20437 8664 23079 8666
rect 20437 8608 20442 8664
rect 20498 8608 23018 8664
rect 23074 8608 23079 8664
rect 20437 8606 23079 8608
rect 20437 8603 20503 8606
rect 23013 8603 23079 8606
rect 19609 8530 19675 8533
rect 20897 8530 20963 8533
rect 19609 8528 20963 8530
rect 19609 8472 19614 8528
rect 19670 8472 20902 8528
rect 20958 8472 20963 8528
rect 19609 8470 20963 8472
rect 19609 8467 19675 8470
rect 20897 8467 20963 8470
rect 21449 8530 21515 8533
rect 24301 8530 24367 8533
rect 21449 8528 24367 8530
rect 21449 8472 21454 8528
rect 21510 8472 24306 8528
rect 24362 8472 24367 8528
rect 21449 8470 24367 8472
rect 21449 8467 21515 8470
rect 24301 8467 24367 8470
rect 17033 8394 17099 8397
rect 19057 8394 19123 8397
rect 17033 8392 19123 8394
rect 17033 8336 17038 8392
rect 17094 8336 19062 8392
rect 19118 8336 19123 8392
rect 17033 8334 19123 8336
rect 17033 8331 17099 8334
rect 19057 8331 19123 8334
rect 10133 8258 10199 8261
rect 12934 8258 12940 8260
rect 10133 8256 12940 8258
rect 10133 8200 10138 8256
rect 10194 8200 12940 8256
rect 10133 8198 12940 8200
rect 10133 8195 10199 8198
rect 12934 8196 12940 8198
rect 13004 8196 13010 8260
rect 18689 8258 18755 8261
rect 18822 8258 18828 8260
rect 18689 8256 18828 8258
rect 18689 8200 18694 8256
rect 18750 8200 18828 8256
rect 18689 8198 18828 8200
rect 18689 8195 18755 8198
rect 18822 8196 18828 8198
rect 18892 8196 18898 8260
rect 21449 8258 21515 8261
rect 22502 8258 22508 8260
rect 21449 8256 22508 8258
rect 21449 8200 21454 8256
rect 21510 8200 22508 8256
rect 21449 8198 22508 8200
rect 21449 8195 21515 8198
rect 22502 8196 22508 8198
rect 22572 8196 22578 8260
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 23790 8060 23796 8124
rect 23860 8122 23866 8124
rect 29361 8122 29427 8125
rect 23860 8120 29427 8122
rect 23860 8064 29366 8120
rect 29422 8064 29427 8120
rect 23860 8062 29427 8064
rect 23860 8060 23866 8062
rect 29361 8059 29427 8062
rect 27286 7924 27292 7988
rect 27356 7986 27362 7988
rect 27705 7986 27771 7989
rect 27356 7984 27771 7986
rect 27356 7928 27710 7984
rect 27766 7928 27771 7984
rect 27356 7926 27771 7928
rect 27356 7924 27362 7926
rect 27705 7923 27771 7926
rect 17125 7850 17191 7853
rect 18965 7850 19031 7853
rect 17125 7848 19031 7850
rect 17125 7792 17130 7848
rect 17186 7792 18970 7848
rect 19026 7792 19031 7848
rect 17125 7790 19031 7792
rect 17125 7787 17191 7790
rect 18965 7787 19031 7790
rect 16757 7714 16823 7717
rect 19149 7714 19215 7717
rect 16757 7712 19215 7714
rect 16757 7656 16762 7712
rect 16818 7656 19154 7712
rect 19210 7656 19215 7712
rect 16757 7654 19215 7656
rect 16757 7651 16823 7654
rect 19149 7651 19215 7654
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 17401 7578 17467 7581
rect 20713 7578 20779 7581
rect 23841 7578 23907 7581
rect 17401 7576 23907 7578
rect 17401 7520 17406 7576
rect 17462 7520 20718 7576
rect 20774 7520 23846 7576
rect 23902 7520 23907 7576
rect 17401 7518 23907 7520
rect 17401 7515 17467 7518
rect 20713 7515 20779 7518
rect 23841 7515 23907 7518
rect 17217 7442 17283 7445
rect 21909 7442 21975 7445
rect 25221 7442 25287 7445
rect 25814 7442 25820 7444
rect 17217 7440 25820 7442
rect 17217 7384 17222 7440
rect 17278 7384 21914 7440
rect 21970 7384 25226 7440
rect 25282 7384 25820 7440
rect 17217 7382 25820 7384
rect 17217 7379 17283 7382
rect 21909 7379 21975 7382
rect 25221 7379 25287 7382
rect 25814 7380 25820 7382
rect 25884 7380 25890 7444
rect 13854 7244 13860 7308
rect 13924 7306 13930 7308
rect 13997 7306 14063 7309
rect 13924 7304 14063 7306
rect 13924 7248 14002 7304
rect 14058 7248 14063 7304
rect 13924 7246 14063 7248
rect 13924 7244 13930 7246
rect 13997 7243 14063 7246
rect 17861 7306 17927 7309
rect 19057 7306 19123 7309
rect 17861 7304 19123 7306
rect 17861 7248 17866 7304
rect 17922 7248 19062 7304
rect 19118 7248 19123 7304
rect 17861 7246 19123 7248
rect 17861 7243 17927 7246
rect 19057 7243 19123 7246
rect 25405 7170 25471 7173
rect 25865 7170 25931 7173
rect 25405 7168 25931 7170
rect 25405 7112 25410 7168
rect 25466 7112 25870 7168
rect 25926 7112 25931 7168
rect 25405 7110 25931 7112
rect 25405 7107 25471 7110
rect 25865 7107 25931 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 23289 7034 23355 7037
rect 26509 7034 26575 7037
rect 23289 7032 26575 7034
rect 23289 6976 23294 7032
rect 23350 6976 26514 7032
rect 26570 6976 26575 7032
rect 23289 6974 26575 6976
rect 23289 6971 23355 6974
rect 26509 6971 26575 6974
rect 0 6808 800 6928
rect 23473 6898 23539 6901
rect 23606 6898 23612 6900
rect 23473 6896 23612 6898
rect 23473 6840 23478 6896
rect 23534 6840 23612 6896
rect 23473 6838 23612 6840
rect 23473 6835 23539 6838
rect 23606 6836 23612 6838
rect 23676 6836 23682 6900
rect 38621 6808 39421 6928
rect 21633 6762 21699 6765
rect 25497 6762 25563 6765
rect 21633 6760 25563 6762
rect 21633 6704 21638 6760
rect 21694 6704 25502 6760
rect 25558 6704 25563 6760
rect 21633 6702 25563 6704
rect 21633 6699 21699 6702
rect 25497 6699 25563 6702
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 19425 6490 19491 6493
rect 22921 6490 22987 6493
rect 25865 6490 25931 6493
rect 25998 6490 26004 6492
rect 19425 6488 26004 6490
rect 19425 6432 19430 6488
rect 19486 6432 22926 6488
rect 22982 6432 25870 6488
rect 25926 6432 26004 6488
rect 19425 6430 26004 6432
rect 19425 6427 19491 6430
rect 22921 6427 22987 6430
rect 25865 6427 25931 6430
rect 25998 6428 26004 6430
rect 26068 6428 26074 6492
rect 21909 6354 21975 6357
rect 22134 6354 22140 6356
rect 21909 6352 22140 6354
rect 21909 6296 21914 6352
rect 21970 6296 22140 6352
rect 21909 6294 22140 6296
rect 21909 6291 21975 6294
rect 22134 6292 22140 6294
rect 22204 6292 22210 6356
rect 22553 6354 22619 6357
rect 25589 6356 25655 6357
rect 25589 6354 25636 6356
rect 22553 6352 25636 6354
rect 22553 6296 22558 6352
rect 22614 6296 25594 6352
rect 22553 6294 25636 6296
rect 22553 6291 22619 6294
rect 25589 6292 25636 6294
rect 25700 6292 25706 6356
rect 25589 6291 25655 6292
rect 13997 6218 14063 6221
rect 18505 6218 18571 6221
rect 13997 6216 18571 6218
rect 13997 6160 14002 6216
rect 14058 6160 18510 6216
rect 18566 6160 18571 6216
rect 13997 6158 18571 6160
rect 13997 6155 14063 6158
rect 18505 6155 18571 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 23289 5540 23355 5541
rect 23238 5476 23244 5540
rect 23308 5538 23355 5540
rect 23308 5536 23400 5538
rect 23350 5480 23400 5536
rect 23308 5478 23400 5480
rect 23308 5476 23355 5478
rect 23289 5475 23355 5476
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 26785 4994 26851 4997
rect 26918 4994 26924 4996
rect 26785 4992 26924 4994
rect 26785 4936 26790 4992
rect 26846 4936 26924 4992
rect 26785 4934 26924 4936
rect 26785 4931 26851 4934
rect 26918 4932 26924 4934
rect 26988 4932 26994 4996
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 38621 4768 39421 4888
rect 9121 4586 9187 4589
rect 22318 4586 22324 4588
rect 9121 4584 22324 4586
rect 9121 4528 9126 4584
rect 9182 4528 22324 4584
rect 9121 4526 22324 4528
rect 9121 4523 9187 4526
rect 22318 4524 22324 4526
rect 22388 4524 22394 4588
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 0 4178 800 4208
rect 933 4178 999 4181
rect 0 4176 999 4178
rect 0 4120 938 4176
rect 994 4120 999 4176
rect 0 4118 999 4120
rect 0 4088 800 4118
rect 933 4115 999 4118
rect 14365 4178 14431 4181
rect 14590 4178 14596 4180
rect 14365 4176 14596 4178
rect 14365 4120 14370 4176
rect 14426 4120 14596 4176
rect 14365 4118 14596 4120
rect 14365 4115 14431 4118
rect 14590 4116 14596 4118
rect 14660 4116 14666 4180
rect 14273 4042 14339 4045
rect 14406 4042 14412 4044
rect 14273 4040 14412 4042
rect 14273 3984 14278 4040
rect 14334 3984 14412 4040
rect 14273 3982 14412 3984
rect 14273 3979 14339 3982
rect 14406 3980 14412 3982
rect 14476 3980 14482 4044
rect 17585 4042 17651 4045
rect 17718 4042 17724 4044
rect 17585 4040 17724 4042
rect 17585 3984 17590 4040
rect 17646 3984 17724 4040
rect 17585 3982 17724 3984
rect 17585 3979 17651 3982
rect 17718 3980 17724 3982
rect 17788 3980 17794 4044
rect 11605 3908 11671 3909
rect 11605 3906 11652 3908
rect 11524 3904 11652 3906
rect 11716 3906 11722 3908
rect 12617 3906 12683 3909
rect 25221 3906 25287 3909
rect 11716 3904 25287 3906
rect 11524 3848 11610 3904
rect 11716 3848 12622 3904
rect 12678 3848 25226 3904
rect 25282 3848 25287 3904
rect 11524 3846 11652 3848
rect 11605 3844 11652 3846
rect 11716 3846 25287 3848
rect 11716 3844 11722 3846
rect 11605 3843 11671 3844
rect 12617 3843 12683 3846
rect 25221 3843 25287 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 15837 3634 15903 3637
rect 18873 3634 18939 3637
rect 15837 3632 18939 3634
rect 15837 3576 15842 3632
rect 15898 3576 18878 3632
rect 18934 3576 18939 3632
rect 15837 3574 18939 3576
rect 15837 3571 15903 3574
rect 18873 3571 18939 3574
rect 10961 3498 11027 3501
rect 18781 3498 18847 3501
rect 24577 3498 24643 3501
rect 10961 3496 24643 3498
rect 10961 3440 10966 3496
rect 11022 3440 18786 3496
rect 18842 3440 24582 3496
rect 24638 3440 24643 3496
rect 10961 3438 24643 3440
rect 10961 3435 11027 3438
rect 18781 3435 18847 3438
rect 24577 3435 24643 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 24669 2684 24735 2685
rect 24669 2680 24716 2684
rect 24780 2682 24786 2684
rect 24669 2624 24674 2680
rect 24669 2620 24716 2624
rect 24780 2622 24826 2682
rect 24780 2620 24786 2622
rect 24669 2619 24735 2620
rect 24158 2348 24164 2412
rect 24228 2410 24234 2412
rect 35709 2410 35775 2413
rect 24228 2408 35775 2410
rect 24228 2352 35714 2408
rect 35770 2352 35775 2408
rect 24228 2350 35775 2352
rect 24228 2348 24234 2350
rect 35709 2347 35775 2350
rect 4870 2208 5186 2209
rect 0 2138 800 2168
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
rect 1485 2138 1551 2141
rect 0 2136 1551 2138
rect 0 2080 1490 2136
rect 1546 2080 1551 2136
rect 0 2078 1551 2080
rect 0 2048 800 2078
rect 1485 2075 1551 2078
rect 37733 2138 37799 2141
rect 38621 2138 39421 2168
rect 37733 2136 39421 2138
rect 37733 2080 37738 2136
rect 37794 2080 39421 2136
rect 37733 2078 39421 2080
rect 37733 2075 37799 2078
rect 38621 2048 39421 2078
rect 37917 98 37983 101
rect 38621 98 39421 128
rect 37917 96 39421 98
rect 37917 40 37922 96
rect 37978 40 39421 96
rect 37917 38 39421 40
rect 37917 35 37983 38
rect 38621 8 39421 38
<< via3 >>
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 35596 39196 35660 39200
rect 35596 39140 35600 39196
rect 35600 39140 35656 39196
rect 35656 39140 35660 39196
rect 35596 39136 35660 39140
rect 35676 39196 35740 39200
rect 35676 39140 35680 39196
rect 35680 39140 35736 39196
rect 35736 39140 35740 39196
rect 35676 39136 35740 39140
rect 35756 39196 35820 39200
rect 35756 39140 35760 39196
rect 35760 39140 35816 39196
rect 35816 39140 35820 39196
rect 35756 39136 35820 39140
rect 35836 39196 35900 39200
rect 35836 39140 35840 39196
rect 35840 39140 35896 39196
rect 35896 39140 35900 39196
rect 35836 39136 35900 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 35596 38108 35660 38112
rect 35596 38052 35600 38108
rect 35600 38052 35656 38108
rect 35656 38052 35660 38108
rect 35596 38048 35660 38052
rect 35676 38108 35740 38112
rect 35676 38052 35680 38108
rect 35680 38052 35736 38108
rect 35736 38052 35740 38108
rect 35676 38048 35740 38052
rect 35756 38108 35820 38112
rect 35756 38052 35760 38108
rect 35760 38052 35816 38108
rect 35816 38052 35820 38108
rect 35756 38048 35820 38052
rect 35836 38108 35900 38112
rect 35836 38052 35840 38108
rect 35840 38052 35896 38108
rect 35896 38052 35900 38108
rect 35836 38048 35900 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 12388 35864 12452 35868
rect 12388 35808 12438 35864
rect 12438 35808 12452 35864
rect 12388 35804 12452 35808
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 11652 35320 11716 35324
rect 11652 35264 11666 35320
rect 11666 35264 11716 35320
rect 11652 35260 11716 35264
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 26004 34580 26068 34644
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 29132 32676 29196 32740
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 26740 31996 26804 32060
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 22324 31512 22388 31516
rect 22324 31456 22338 31512
rect 22338 31456 22388 31512
rect 22324 31452 22388 31456
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 20116 30772 20180 30836
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 12204 30364 12268 30428
rect 17540 30364 17604 30428
rect 18644 30424 18708 30428
rect 18644 30368 18658 30424
rect 18658 30368 18708 30424
rect 18644 30364 18708 30368
rect 25452 30364 25516 30428
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 12388 29004 12452 29068
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 21036 26420 21100 26484
rect 14412 26284 14476 26348
rect 19748 26344 19812 26348
rect 19748 26288 19798 26344
rect 19798 26288 19812 26344
rect 19748 26284 19812 26288
rect 24716 26284 24780 26348
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 14596 25936 14660 25940
rect 14596 25880 14610 25936
rect 14610 25880 14660 25936
rect 14596 25876 14660 25880
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 17724 24924 17788 24988
rect 30972 24924 31036 24988
rect 26004 24848 26068 24852
rect 26004 24792 26018 24848
rect 26018 24792 26068 24848
rect 26004 24788 26068 24792
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 24164 23896 24228 23900
rect 24164 23840 24178 23896
rect 24178 23840 24228 23896
rect 24164 23836 24228 23840
rect 22692 23564 22756 23628
rect 13124 23428 13188 23492
rect 22508 23488 22572 23492
rect 23612 23700 23676 23764
rect 26924 23564 26988 23628
rect 22508 23432 22522 23488
rect 22522 23432 22572 23488
rect 22508 23428 22572 23432
rect 23796 23488 23860 23492
rect 23796 23432 23810 23488
rect 23810 23432 23860 23488
rect 23796 23428 23860 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 25452 21584 25516 21588
rect 25452 21528 25466 21584
rect 25466 21528 25516 21584
rect 25452 21524 25516 21528
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 18828 20980 18892 21044
rect 27108 20708 27172 20772
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 23244 19348 23308 19412
rect 16436 19212 16500 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 28212 18396 28276 18460
rect 19196 18320 19260 18324
rect 19196 18264 19246 18320
rect 19246 18264 19260 18320
rect 19196 18260 19260 18264
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 28764 16688 28828 16692
rect 28764 16632 28778 16688
rect 28778 16632 28828 16688
rect 28764 16628 28828 16632
rect 26740 16492 26804 16556
rect 13676 16356 13740 16420
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 27292 15540 27356 15604
rect 25268 15268 25332 15332
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 11468 15132 11532 15196
rect 17540 15192 17604 15196
rect 17540 15136 17554 15192
rect 17554 15136 17604 15192
rect 17540 15132 17604 15136
rect 11652 14724 11716 14788
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19196 14512 19260 14516
rect 19196 14456 19210 14512
rect 19210 14456 19260 14512
rect 19196 14452 19260 14456
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 28396 13908 28460 13972
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 12020 13364 12084 13428
rect 14780 13092 14844 13156
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 25636 12684 25700 12748
rect 22324 12608 22388 12612
rect 22324 12552 22338 12608
rect 22338 12552 22388 12608
rect 22324 12548 22388 12552
rect 25268 12548 25332 12612
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 25820 12276 25884 12340
rect 30972 12276 31036 12340
rect 16436 12140 16500 12204
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 28764 11868 28828 11932
rect 20116 11792 20180 11796
rect 20116 11736 20130 11792
rect 20130 11736 20180 11792
rect 20116 11732 20180 11736
rect 28396 11732 28460 11796
rect 13124 11596 13188 11660
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 13860 11052 13924 11116
rect 22140 11112 22204 11116
rect 22140 11056 22154 11112
rect 22154 11056 22204 11112
rect 22140 11052 22204 11056
rect 22508 10916 22572 10980
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 22508 10704 22572 10708
rect 22508 10648 22558 10704
rect 22558 10648 22572 10704
rect 12204 10508 12268 10572
rect 22508 10644 22572 10648
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 25636 10160 25700 10164
rect 25636 10104 25650 10160
rect 25650 10104 25700 10160
rect 25636 10100 25700 10104
rect 28396 10024 28460 10028
rect 28396 9968 28446 10024
rect 28446 9968 28460 10024
rect 28396 9964 28460 9968
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 11468 9556 11532 9620
rect 26004 9692 26068 9756
rect 13124 9556 13188 9620
rect 18644 9556 18708 9620
rect 22692 9616 22756 9620
rect 22692 9560 22706 9616
rect 22706 9560 22756 9616
rect 22692 9556 22756 9560
rect 25820 9556 25884 9620
rect 27108 9556 27172 9620
rect 29132 9556 29196 9620
rect 13676 9480 13740 9484
rect 13676 9424 13726 9480
rect 13726 9424 13740 9480
rect 13676 9420 13740 9424
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 12020 9208 12084 9212
rect 12020 9152 12070 9208
rect 12070 9152 12084 9208
rect 12020 9148 12084 9152
rect 14780 9148 14844 9212
rect 19748 9148 19812 9212
rect 21036 9208 21100 9212
rect 21036 9152 21050 9208
rect 21050 9152 21100 9208
rect 21036 9148 21100 9152
rect 21956 9148 22020 9212
rect 28212 9284 28276 9348
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 12940 8196 13004 8260
rect 18828 8196 18892 8260
rect 22508 8196 22572 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 23796 8060 23860 8124
rect 27292 7924 27356 7988
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 25820 7380 25884 7444
rect 13860 7244 13924 7308
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 23612 6836 23676 6900
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 26004 6428 26068 6492
rect 22140 6292 22204 6356
rect 25636 6352 25700 6356
rect 25636 6296 25650 6352
rect 25650 6296 25700 6352
rect 25636 6292 25700 6296
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 23244 5536 23308 5540
rect 23244 5480 23294 5536
rect 23294 5480 23308 5536
rect 23244 5476 23308 5480
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 26924 4932 26988 4996
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 22324 4524 22388 4588
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 14596 4116 14660 4180
rect 14412 3980 14476 4044
rect 17724 3980 17788 4044
rect 11652 3904 11716 3908
rect 11652 3848 11666 3904
rect 11666 3848 11716 3904
rect 11652 3844 11716 3848
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 24716 2680 24780 2684
rect 24716 2624 24730 2680
rect 24730 2624 24780 2680
rect 24716 2620 24780 2624
rect 24164 2348 24228 2412
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 38656 4528 39216
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36260 4528 36416
rect 4208 36024 4250 36260
rect 4486 36024 4528 36260
rect 4208 35392 4528 36024
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 39200 5188 39216
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 36920 5188 36960
rect 4868 36684 4910 36920
rect 5146 36684 5188 36920
rect 4868 35936 5188 36684
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 34928 38656 35248 39216
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36260 35248 36416
rect 34928 36024 34970 36260
rect 35206 36024 35248 36260
rect 12387 35868 12453 35869
rect 12387 35804 12388 35868
rect 12452 35804 12453 35868
rect 12387 35803 12453 35804
rect 11651 35324 11717 35325
rect 11651 35260 11652 35324
rect 11716 35260 11717 35324
rect 11651 35259 11717 35260
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 11467 15196 11533 15197
rect 11467 15132 11468 15196
rect 11532 15132 11533 15196
rect 11467 15131 11533 15132
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 11470 9621 11530 15131
rect 11654 14789 11714 35259
rect 12203 30428 12269 30429
rect 12203 30364 12204 30428
rect 12268 30364 12269 30428
rect 12203 30363 12269 30364
rect 11651 14788 11717 14789
rect 11651 14724 11652 14788
rect 11716 14724 11717 14788
rect 11651 14723 11717 14724
rect 11467 9620 11533 9621
rect 11467 9556 11468 9620
rect 11532 9556 11533 9620
rect 11467 9555 11533 9556
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 6284 5188 6496
rect 4868 6048 4910 6284
rect 5146 6048 5188 6284
rect 4868 5472 5188 6048
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 11654 3909 11714 14723
rect 12019 13428 12085 13429
rect 12019 13364 12020 13428
rect 12084 13364 12085 13428
rect 12019 13363 12085 13364
rect 12022 9213 12082 13363
rect 12206 10573 12266 30363
rect 12390 29069 12450 35803
rect 34928 35392 35248 36024
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 26003 34644 26069 34645
rect 26003 34580 26004 34644
rect 26068 34580 26069 34644
rect 26003 34579 26069 34580
rect 22323 31516 22389 31517
rect 22323 31452 22324 31516
rect 22388 31452 22389 31516
rect 22323 31451 22389 31452
rect 20115 30836 20181 30837
rect 20115 30772 20116 30836
rect 20180 30772 20181 30836
rect 20115 30771 20181 30772
rect 17539 30428 17605 30429
rect 17539 30364 17540 30428
rect 17604 30364 17605 30428
rect 17539 30363 17605 30364
rect 18643 30428 18709 30429
rect 18643 30364 18644 30428
rect 18708 30364 18709 30428
rect 18643 30363 18709 30364
rect 12387 29068 12453 29069
rect 12387 29004 12388 29068
rect 12452 29004 12453 29068
rect 12387 29003 12453 29004
rect 14411 26348 14477 26349
rect 14411 26284 14412 26348
rect 14476 26284 14477 26348
rect 14411 26283 14477 26284
rect 13123 23492 13189 23493
rect 13123 23428 13124 23492
rect 13188 23428 13189 23492
rect 13123 23427 13189 23428
rect 13126 12450 13186 23427
rect 13675 16420 13741 16421
rect 13675 16356 13676 16420
rect 13740 16356 13741 16420
rect 13675 16355 13741 16356
rect 12942 12390 13186 12450
rect 12203 10572 12269 10573
rect 12203 10508 12204 10572
rect 12268 10508 12269 10572
rect 12203 10507 12269 10508
rect 12019 9212 12085 9213
rect 12019 9148 12020 9212
rect 12084 9148 12085 9212
rect 12019 9147 12085 9148
rect 12942 8261 13002 12390
rect 13123 11660 13189 11661
rect 13123 11596 13124 11660
rect 13188 11596 13189 11660
rect 13123 11595 13189 11596
rect 13126 9621 13186 11595
rect 13123 9620 13189 9621
rect 13123 9556 13124 9620
rect 13188 9556 13189 9620
rect 13123 9555 13189 9556
rect 13678 9485 13738 16355
rect 13859 11116 13925 11117
rect 13859 11052 13860 11116
rect 13924 11052 13925 11116
rect 13859 11051 13925 11052
rect 13675 9484 13741 9485
rect 13675 9420 13676 9484
rect 13740 9420 13741 9484
rect 13675 9419 13741 9420
rect 12939 8260 13005 8261
rect 12939 8196 12940 8260
rect 13004 8196 13005 8260
rect 12939 8195 13005 8196
rect 13862 7309 13922 11051
rect 13859 7308 13925 7309
rect 13859 7244 13860 7308
rect 13924 7244 13925 7308
rect 13859 7243 13925 7244
rect 14414 4045 14474 26283
rect 14595 25940 14661 25941
rect 14595 25876 14596 25940
rect 14660 25876 14661 25940
rect 14595 25875 14661 25876
rect 14598 4181 14658 25875
rect 16435 19276 16501 19277
rect 16435 19212 16436 19276
rect 16500 19212 16501 19276
rect 16435 19211 16501 19212
rect 14779 13156 14845 13157
rect 14779 13092 14780 13156
rect 14844 13092 14845 13156
rect 14779 13091 14845 13092
rect 14782 9213 14842 13091
rect 16438 12205 16498 19211
rect 17542 15197 17602 30363
rect 17723 24988 17789 24989
rect 17723 24924 17724 24988
rect 17788 24924 17789 24988
rect 17723 24923 17789 24924
rect 17539 15196 17605 15197
rect 17539 15132 17540 15196
rect 17604 15132 17605 15196
rect 17539 15131 17605 15132
rect 16435 12204 16501 12205
rect 16435 12140 16436 12204
rect 16500 12140 16501 12204
rect 16435 12139 16501 12140
rect 14779 9212 14845 9213
rect 14779 9148 14780 9212
rect 14844 9148 14845 9212
rect 14779 9147 14845 9148
rect 14595 4180 14661 4181
rect 14595 4116 14596 4180
rect 14660 4116 14661 4180
rect 14595 4115 14661 4116
rect 17726 4045 17786 24923
rect 18646 9621 18706 30363
rect 19747 26348 19813 26349
rect 19747 26284 19748 26348
rect 19812 26284 19813 26348
rect 19747 26283 19813 26284
rect 18827 21044 18893 21045
rect 18827 20980 18828 21044
rect 18892 20980 18893 21044
rect 18827 20979 18893 20980
rect 18643 9620 18709 9621
rect 18643 9556 18644 9620
rect 18708 9556 18709 9620
rect 18643 9555 18709 9556
rect 18830 8261 18890 20979
rect 19195 18324 19261 18325
rect 19195 18260 19196 18324
rect 19260 18260 19261 18324
rect 19195 18259 19261 18260
rect 19198 14517 19258 18259
rect 19195 14516 19261 14517
rect 19195 14452 19196 14516
rect 19260 14452 19261 14516
rect 19195 14451 19261 14452
rect 19750 9213 19810 26283
rect 20118 11797 20178 30771
rect 21035 26484 21101 26485
rect 21035 26420 21036 26484
rect 21100 26420 21101 26484
rect 21035 26419 21101 26420
rect 20115 11796 20181 11797
rect 20115 11732 20116 11796
rect 20180 11732 20181 11796
rect 20115 11731 20181 11732
rect 21038 9213 21098 26419
rect 22326 18730 22386 31451
rect 25451 30428 25517 30429
rect 25451 30364 25452 30428
rect 25516 30364 25517 30428
rect 25451 30363 25517 30364
rect 24715 26348 24781 26349
rect 24715 26284 24716 26348
rect 24780 26284 24781 26348
rect 24715 26283 24781 26284
rect 24163 23900 24229 23901
rect 24163 23836 24164 23900
rect 24228 23836 24229 23900
rect 24163 23835 24229 23836
rect 23611 23764 23677 23765
rect 23611 23700 23612 23764
rect 23676 23700 23677 23764
rect 23611 23699 23677 23700
rect 22691 23628 22757 23629
rect 22691 23564 22692 23628
rect 22756 23564 22757 23628
rect 22691 23563 22757 23564
rect 22507 23492 22573 23493
rect 22507 23428 22508 23492
rect 22572 23428 22573 23492
rect 22507 23427 22573 23428
rect 21958 18670 22386 18730
rect 21958 9213 22018 18670
rect 22323 12612 22389 12613
rect 22323 12548 22324 12612
rect 22388 12548 22389 12612
rect 22323 12547 22389 12548
rect 22139 11116 22205 11117
rect 22139 11052 22140 11116
rect 22204 11052 22205 11116
rect 22139 11051 22205 11052
rect 19747 9212 19813 9213
rect 19747 9148 19748 9212
rect 19812 9148 19813 9212
rect 19747 9147 19813 9148
rect 21035 9212 21101 9213
rect 21035 9148 21036 9212
rect 21100 9148 21101 9212
rect 21035 9147 21101 9148
rect 21955 9212 22021 9213
rect 21955 9148 21956 9212
rect 22020 9148 22021 9212
rect 21955 9147 22021 9148
rect 18827 8260 18893 8261
rect 18827 8196 18828 8260
rect 18892 8196 18893 8260
rect 18827 8195 18893 8196
rect 22142 6357 22202 11051
rect 22139 6356 22205 6357
rect 22139 6292 22140 6356
rect 22204 6292 22205 6356
rect 22139 6291 22205 6292
rect 22326 4589 22386 12547
rect 22510 10981 22570 23427
rect 22507 10980 22573 10981
rect 22507 10916 22508 10980
rect 22572 10916 22573 10980
rect 22507 10915 22573 10916
rect 22507 10708 22573 10709
rect 22507 10644 22508 10708
rect 22572 10644 22573 10708
rect 22507 10643 22573 10644
rect 22510 8261 22570 10643
rect 22694 9621 22754 23563
rect 23243 19412 23309 19413
rect 23243 19348 23244 19412
rect 23308 19348 23309 19412
rect 23243 19347 23309 19348
rect 22691 9620 22757 9621
rect 22691 9556 22692 9620
rect 22756 9556 22757 9620
rect 22691 9555 22757 9556
rect 22507 8260 22573 8261
rect 22507 8196 22508 8260
rect 22572 8196 22573 8260
rect 22507 8195 22573 8196
rect 23246 5541 23306 19347
rect 23614 6901 23674 23699
rect 23795 23492 23861 23493
rect 23795 23428 23796 23492
rect 23860 23428 23861 23492
rect 23795 23427 23861 23428
rect 23798 8125 23858 23427
rect 23795 8124 23861 8125
rect 23795 8060 23796 8124
rect 23860 8060 23861 8124
rect 23795 8059 23861 8060
rect 23611 6900 23677 6901
rect 23611 6836 23612 6900
rect 23676 6836 23677 6900
rect 23611 6835 23677 6836
rect 23243 5540 23309 5541
rect 23243 5476 23244 5540
rect 23308 5476 23309 5540
rect 23243 5475 23309 5476
rect 22323 4588 22389 4589
rect 22323 4524 22324 4588
rect 22388 4524 22389 4588
rect 22323 4523 22389 4524
rect 14411 4044 14477 4045
rect 14411 3980 14412 4044
rect 14476 3980 14477 4044
rect 14411 3979 14477 3980
rect 17723 4044 17789 4045
rect 17723 3980 17724 4044
rect 17788 3980 17789 4044
rect 17723 3979 17789 3980
rect 11651 3908 11717 3909
rect 11651 3844 11652 3908
rect 11716 3844 11717 3908
rect 11651 3843 11717 3844
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 24166 2413 24226 23835
rect 24718 2685 24778 26283
rect 25454 21589 25514 30363
rect 26006 24853 26066 34579
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 29131 32740 29197 32741
rect 29131 32676 29132 32740
rect 29196 32676 29197 32740
rect 29131 32675 29197 32676
rect 26739 32060 26805 32061
rect 26739 31996 26740 32060
rect 26804 31996 26805 32060
rect 26739 31995 26805 31996
rect 26003 24852 26069 24853
rect 26003 24788 26004 24852
rect 26068 24788 26069 24852
rect 26003 24787 26069 24788
rect 25451 21588 25517 21589
rect 25451 21524 25452 21588
rect 25516 21524 25517 21588
rect 25451 21523 25517 21524
rect 26742 16557 26802 31995
rect 26923 23628 26989 23629
rect 26923 23564 26924 23628
rect 26988 23564 26989 23628
rect 26923 23563 26989 23564
rect 26739 16556 26805 16557
rect 26739 16492 26740 16556
rect 26804 16492 26805 16556
rect 26739 16491 26805 16492
rect 25267 15332 25333 15333
rect 25267 15268 25268 15332
rect 25332 15268 25333 15332
rect 25267 15267 25333 15268
rect 25270 12613 25330 15267
rect 25635 12748 25701 12749
rect 25635 12684 25636 12748
rect 25700 12684 25701 12748
rect 25635 12683 25701 12684
rect 25267 12612 25333 12613
rect 25267 12548 25268 12612
rect 25332 12548 25333 12612
rect 25267 12547 25333 12548
rect 25638 10165 25698 12683
rect 25819 12340 25885 12341
rect 25819 12276 25820 12340
rect 25884 12276 25885 12340
rect 25819 12275 25885 12276
rect 25635 10164 25701 10165
rect 25635 10100 25636 10164
rect 25700 10100 25701 10164
rect 25635 10099 25701 10100
rect 25638 6357 25698 10099
rect 25822 9621 25882 12275
rect 26003 9756 26069 9757
rect 26003 9692 26004 9756
rect 26068 9692 26069 9756
rect 26003 9691 26069 9692
rect 25819 9620 25885 9621
rect 25819 9556 25820 9620
rect 25884 9556 25885 9620
rect 25819 9555 25885 9556
rect 25822 7445 25882 9555
rect 25819 7444 25885 7445
rect 25819 7380 25820 7444
rect 25884 7380 25885 7444
rect 25819 7379 25885 7380
rect 26006 6493 26066 9691
rect 26003 6492 26069 6493
rect 26003 6428 26004 6492
rect 26068 6428 26069 6492
rect 26003 6427 26069 6428
rect 25635 6356 25701 6357
rect 25635 6292 25636 6356
rect 25700 6292 25701 6356
rect 25635 6291 25701 6292
rect 26926 4997 26986 23563
rect 27107 20772 27173 20773
rect 27107 20708 27108 20772
rect 27172 20708 27173 20772
rect 27107 20707 27173 20708
rect 27110 9621 27170 20707
rect 28211 18460 28277 18461
rect 28211 18396 28212 18460
rect 28276 18396 28277 18460
rect 28211 18395 28277 18396
rect 27291 15604 27357 15605
rect 27291 15540 27292 15604
rect 27356 15540 27357 15604
rect 27291 15539 27357 15540
rect 27107 9620 27173 9621
rect 27107 9556 27108 9620
rect 27172 9556 27173 9620
rect 27107 9555 27173 9556
rect 27294 7989 27354 15539
rect 28214 9349 28274 18395
rect 28763 16692 28829 16693
rect 28763 16628 28764 16692
rect 28828 16628 28829 16692
rect 28763 16627 28829 16628
rect 28395 13972 28461 13973
rect 28395 13908 28396 13972
rect 28460 13908 28461 13972
rect 28395 13907 28461 13908
rect 28398 11797 28458 13907
rect 28766 11933 28826 16627
rect 28763 11932 28829 11933
rect 28763 11868 28764 11932
rect 28828 11868 28829 11932
rect 28763 11867 28829 11868
rect 28395 11796 28461 11797
rect 28395 11732 28396 11796
rect 28460 11732 28461 11796
rect 28395 11731 28461 11732
rect 28398 10029 28458 11731
rect 28395 10028 28461 10029
rect 28395 9964 28396 10028
rect 28460 9964 28461 10028
rect 28395 9963 28461 9964
rect 29134 9621 29194 32675
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 30971 24988 31037 24989
rect 30971 24924 30972 24988
rect 31036 24924 31037 24988
rect 30971 24923 31037 24924
rect 30974 12341 31034 24923
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 30971 12340 31037 12341
rect 30971 12276 30972 12340
rect 31036 12276 31037 12340
rect 30971 12275 31037 12276
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 29131 9620 29197 9621
rect 29131 9556 29132 9620
rect 29196 9556 29197 9620
rect 29131 9555 29197 9556
rect 28211 9348 28277 9349
rect 28211 9284 28212 9348
rect 28276 9284 28277 9348
rect 28211 9283 28277 9284
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 27291 7988 27357 7989
rect 27291 7924 27292 7988
rect 27356 7924 27357 7988
rect 27291 7923 27357 7924
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5624 35248 5952
rect 34928 5388 34970 5624
rect 35206 5388 35248 5624
rect 26923 4996 26989 4997
rect 26923 4932 26924 4996
rect 26988 4932 26989 4996
rect 26923 4931 26989 4932
rect 34928 4928 35248 5388
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 24715 2684 24781 2685
rect 24715 2620 24716 2684
rect 24780 2620 24781 2684
rect 24715 2619 24781 2620
rect 24163 2412 24229 2413
rect 24163 2348 24164 2412
rect 24228 2348 24229 2412
rect 24163 2347 24229 2348
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 2128 35248 2688
rect 35588 39200 35908 39216
rect 35588 39136 35596 39200
rect 35660 39136 35676 39200
rect 35740 39136 35756 39200
rect 35820 39136 35836 39200
rect 35900 39136 35908 39200
rect 35588 38112 35908 39136
rect 35588 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35908 38112
rect 35588 37024 35908 38048
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 36920 35908 36960
rect 35588 36684 35630 36920
rect 35866 36684 35908 36920
rect 35588 35936 35908 36684
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35588 29408 35908 30432
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35588 25056 35908 26080
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35588 18528 35908 19552
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 6284 35908 6496
rect 35588 6048 35630 6284
rect 35866 6048 35908 6284
rect 35588 5472 35908 6048
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
<< via4 >>
rect 4250 36024 4486 36260
rect 4250 5388 4486 5624
rect 4910 36684 5146 36920
rect 34970 36024 35206 36260
rect 4910 6048 5146 6284
rect 34970 5388 35206 5624
rect 35630 36684 35866 36920
rect 35630 6048 35866 6284
<< metal5 >>
rect 1056 36920 38320 36962
rect 1056 36684 4910 36920
rect 5146 36684 35630 36920
rect 35866 36684 38320 36920
rect 1056 36642 38320 36684
rect 1056 36260 38320 36302
rect 1056 36024 4250 36260
rect 4486 36024 34970 36260
rect 35206 36024 38320 36260
rect 1056 35982 38320 36024
rect 1056 6284 38320 6326
rect 1056 6048 4910 6284
rect 5146 6048 35630 6284
rect 35866 6048 38320 6284
rect 1056 6006 38320 6048
rect 1056 5624 38320 5666
rect 1056 5388 4250 5624
rect 4486 5388 34970 5624
rect 35206 5388 38320 5624
rect 1056 5346 38320 5388
use sky130_fd_sc_hd__inv_2  _1276_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9292 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _1277_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _1278_
timestamp 1688980957
transform 1 0 8372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1279_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13800 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _1280_
timestamp 1688980957
transform 1 0 7176 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_2  _1281_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14904 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _1282_
timestamp 1688980957
transform 1 0 4140 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__or2_1  _1283_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13064 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1284_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11040 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1285_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4968 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _1286_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_8  _1287_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15364 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  _1288_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28152 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_2  _1289_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13800 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_4  _1290_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12052 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__a21boi_1  _1291_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1292_
timestamp 1688980957
transform 1 0 12236 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _1293_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7176 0 -1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__nand3b_2  _1294_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15180 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1295_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _1296_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14720 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__and2b_1  _1297_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7820 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1298_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15824 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1299_
timestamp 1688980957
transform 1 0 7912 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_4  _1300_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8464 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__or4bb_1  _1301_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o221ai_4  _1302_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7912 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_8  _1303_
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__a221oi_2  _1304_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17296 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1305_
timestamp 1688980957
transform 1 0 12788 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1306_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12052 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1307_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13524 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1308_
timestamp 1688980957
transform 1 0 18492 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1309_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20424 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1310_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20792 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1311_
timestamp 1688980957
transform 1 0 15456 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _1312_
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_16  _1313_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23000 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__nand2_1  _1314_
timestamp 1688980957
transform -1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1315_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1316_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4324 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1317_
timestamp 1688980957
transform 1 0 4600 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1318_
timestamp 1688980957
transform 1 0 8372 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1319_
timestamp 1688980957
transform 1 0 8096 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1320_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9016 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1321_
timestamp 1688980957
transform 1 0 9752 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_4  _1322_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12512 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__o211a_1  _1323_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10948 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1324_
timestamp 1688980957
transform 1 0 12052 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _1325_
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _1326_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10120 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1327_
timestamp 1688980957
transform -1 0 13156 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _1328_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20516 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1329_
timestamp 1688980957
transform 1 0 10672 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _1330_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 2062 592
use sky130_fd_sc_hd__o211a_1  _1331_
timestamp 1688980957
transform -1 0 12880 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _1332_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13064 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_8  _1333_
timestamp 1688980957
transform 1 0 19688 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_4  _1334_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23736 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _1335_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1336_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14536 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _1337_
timestamp 1688980957
transform 1 0 15732 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1338_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18308 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_4  _1339_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17940 0 -1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_1  _1340_
timestamp 1688980957
transform 1 0 19780 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1341_
timestamp 1688980957
transform 1 0 20056 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_2  _1342_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15916 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1343_
timestamp 1688980957
transform -1 0 18216 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _1344_
timestamp 1688980957
transform 1 0 16928 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1345_
timestamp 1688980957
transform 1 0 18216 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1346_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1347_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18400 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1348_
timestamp 1688980957
transform 1 0 17572 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1349_
timestamp 1688980957
transform 1 0 16008 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _1350_
timestamp 1688980957
transform -1 0 13708 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_8  _1351_
timestamp 1688980957
transform 1 0 19136 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_1  _1352_
timestamp 1688980957
transform 1 0 13524 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1353_
timestamp 1688980957
transform -1 0 14812 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _1354_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12144 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1355_
timestamp 1688980957
transform 1 0 14260 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_4  _1356_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16008 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_4  _1357_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1358_
timestamp 1688980957
transform 1 0 9016 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1359_
timestamp 1688980957
transform 1 0 12328 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1360_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13432 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_4  _1361_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13892 0 -1 16320
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_8  _1362_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21620 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_8  _1363_
timestamp 1688980957
transform 1 0 22448 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__o22ai_1  _1364_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13156 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_8  _1365_
timestamp 1688980957
transform 1 0 20056 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__a21oi_2  _1366_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _1367_
timestamp 1688980957
transform 1 0 27692 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1368_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11960 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_8  _1369_
timestamp 1688980957
transform 1 0 22172 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__a211o_1  _1370_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11960 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1371_
timestamp 1688980957
transform -1 0 12420 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1372_
timestamp 1688980957
transform 1 0 12420 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1373_
timestamp 1688980957
transform -1 0 16560 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1374_
timestamp 1688980957
transform 1 0 15548 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1375_
timestamp 1688980957
transform 1 0 15272 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1376_
timestamp 1688980957
transform 1 0 15640 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1377_
timestamp 1688980957
transform 1 0 17296 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1378_
timestamp 1688980957
transform 1 0 17664 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _1379_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17848 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1380_
timestamp 1688980957
transform 1 0 11592 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1381_
timestamp 1688980957
transform 1 0 11500 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1382_
timestamp 1688980957
transform -1 0 11500 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1383_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12236 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1384_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18492 0 -1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__a221o_1  _1385_
timestamp 1688980957
transform 1 0 17296 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1386_
timestamp 1688980957
transform 1 0 18584 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _1387_
timestamp 1688980957
transform -1 0 18768 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1388_
timestamp 1688980957
transform -1 0 12880 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1389_
timestamp 1688980957
transform 1 0 11684 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1390_
timestamp 1688980957
transform -1 0 12236 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1391_
timestamp 1688980957
transform 1 0 12420 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1392_
timestamp 1688980957
transform 1 0 18492 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1393_
timestamp 1688980957
transform 1 0 19136 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1394_
timestamp 1688980957
transform 1 0 19596 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1395_
timestamp 1688980957
transform 1 0 20608 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1396_
timestamp 1688980957
transform -1 0 26036 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1397_
timestamp 1688980957
transform 1 0 24748 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_4  _1398_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25944 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _1399_
timestamp 1688980957
transform -1 0 28060 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1400_
timestamp 1688980957
transform 1 0 28796 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1401_
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_2  _1402_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28428 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1403_
timestamp 1688980957
transform -1 0 22172 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1404_
timestamp 1688980957
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1405_
timestamp 1688980957
transform 1 0 24012 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1406_
timestamp 1688980957
transform -1 0 25300 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1407_
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1408_
timestamp 1688980957
transform 1 0 24840 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1409_
timestamp 1688980957
transform -1 0 26588 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1410_
timestamp 1688980957
transform -1 0 26956 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1411_
timestamp 1688980957
transform -1 0 24472 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1412_
timestamp 1688980957
transform 1 0 24104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1413_
timestamp 1688980957
transform 1 0 24472 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1414_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24288 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1415_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14260 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1416_
timestamp 1688980957
transform -1 0 13248 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1417_
timestamp 1688980957
transform -1 0 12696 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _1418_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19136 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _1419_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17388 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a31oi_4  _1420_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__o211a_2  _1421_
timestamp 1688980957
transform -1 0 23276 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1422_
timestamp 1688980957
transform 1 0 24656 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _1423_
timestamp 1688980957
transform -1 0 22908 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1424_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19228 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _1425_
timestamp 1688980957
transform -1 0 22540 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1426_
timestamp 1688980957
transform -1 0 25668 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1427_
timestamp 1688980957
transform 1 0 24564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1428_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_4  _1429_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23552 0 -1 17408
box -38 -48 1326 592
use sky130_fd_sc_hd__nor4_1  _1430_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 21344 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1431_
timestamp 1688980957
transform -1 0 26864 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1432_
timestamp 1688980957
transform 1 0 20792 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_2  _1433_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26128 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1434_
timestamp 1688980957
transform 1 0 25576 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1435_
timestamp 1688980957
transform 1 0 26312 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1436_
timestamp 1688980957
transform 1 0 26956 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1437_
timestamp 1688980957
transform 1 0 21160 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _1438_
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__o211ai_4  _1439_
timestamp 1688980957
transform -1 0 28888 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _1440_
timestamp 1688980957
transform 1 0 25024 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1441_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14996 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1442_
timestamp 1688980957
transform 1 0 15180 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _1443_
timestamp 1688980957
transform 1 0 13708 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1444_
timestamp 1688980957
transform 1 0 23644 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1445_
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _1446_
timestamp 1688980957
transform 1 0 16192 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1447_
timestamp 1688980957
transform 1 0 15364 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1448_
timestamp 1688980957
transform 1 0 27968 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1449_
timestamp 1688980957
transform -1 0 28980 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1450_
timestamp 1688980957
transform 1 0 14720 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1451_
timestamp 1688980957
transform 1 0 24196 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _1452_
timestamp 1688980957
transform 1 0 24748 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1453_
timestamp 1688980957
transform -1 0 27692 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1454_
timestamp 1688980957
transform 1 0 27232 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1455_
timestamp 1688980957
transform 1 0 27508 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1456_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28336 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1457_
timestamp 1688980957
transform -1 0 30176 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1458_
timestamp 1688980957
transform 1 0 31096 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1459_
timestamp 1688980957
transform -1 0 29992 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _1460_
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _1461_
timestamp 1688980957
transform -1 0 29440 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1462_
timestamp 1688980957
transform -1 0 29808 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1463_
timestamp 1688980957
transform -1 0 31004 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1464_
timestamp 1688980957
transform 1 0 29716 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1465_
timestamp 1688980957
transform 1 0 17480 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1466_
timestamp 1688980957
transform 1 0 17020 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1467_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18492 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1468_
timestamp 1688980957
transform -1 0 19872 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1469_
timestamp 1688980957
transform 1 0 17664 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1470_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1471_
timestamp 1688980957
transform 1 0 17848 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1472_
timestamp 1688980957
transform 1 0 17020 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _1473_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19044 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_8  _1474_
timestamp 1688980957
transform 1 0 27784 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__and3_2  _1475_
timestamp 1688980957
transform 1 0 21896 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1476_
timestamp 1688980957
transform -1 0 15824 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1477_
timestamp 1688980957
transform 1 0 15272 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1478_
timestamp 1688980957
transform -1 0 17112 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1479_
timestamp 1688980957
transform 1 0 15088 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1480_
timestamp 1688980957
transform 1 0 15732 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1481_
timestamp 1688980957
transform 1 0 16560 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1482_
timestamp 1688980957
transform -1 0 17112 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1483_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14444 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1484_
timestamp 1688980957
transform 1 0 14168 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1485_
timestamp 1688980957
transform -1 0 15916 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1486_
timestamp 1688980957
transform -1 0 19964 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _1487_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16652 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1488_
timestamp 1688980957
transform 1 0 19412 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_4  _1489_
timestamp 1688980957
transform -1 0 21252 0 1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_1  _1490_
timestamp 1688980957
transform 1 0 36800 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1491_
timestamp 1688980957
transform 1 0 14812 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1492_
timestamp 1688980957
transform 1 0 15364 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1493_
timestamp 1688980957
transform -1 0 16560 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1494_
timestamp 1688980957
transform 1 0 15088 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1495_
timestamp 1688980957
transform 1 0 15732 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1496_
timestamp 1688980957
transform 1 0 16376 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1497_
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1498_
timestamp 1688980957
transform -1 0 14628 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1499_
timestamp 1688980957
transform 1 0 14628 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1500_
timestamp 1688980957
transform -1 0 16284 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1501_
timestamp 1688980957
transform -1 0 16560 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_2  _1502_
timestamp 1688980957
transform 1 0 20608 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1503_
timestamp 1688980957
transform 1 0 17204 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1504_
timestamp 1688980957
transform 1 0 16836 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1505_
timestamp 1688980957
transform -1 0 18308 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1506_
timestamp 1688980957
transform 1 0 17020 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1507_
timestamp 1688980957
transform 1 0 18400 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1508_
timestamp 1688980957
transform 1 0 18124 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1509_
timestamp 1688980957
transform 1 0 17664 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1510_
timestamp 1688980957
transform 1 0 16836 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1511_
timestamp 1688980957
transform -1 0 18768 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1512_
timestamp 1688980957
transform 1 0 28520 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1513_
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1514_
timestamp 1688980957
transform 1 0 35420 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1515_
timestamp 1688980957
transform -1 0 24840 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1516_
timestamp 1688980957
transform -1 0 25392 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1517_
timestamp 1688980957
transform 1 0 24840 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1518_
timestamp 1688980957
transform -1 0 25760 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1519_
timestamp 1688980957
transform -1 0 26312 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1520_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25116 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1521_
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1522_
timestamp 1688980957
transform -1 0 26588 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1523_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26036 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1524_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25944 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_4  _1525_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25208 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__or2_1  _1526_
timestamp 1688980957
transform 1 0 34408 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1527_
timestamp 1688980957
transform -1 0 32660 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1528_
timestamp 1688980957
transform 1 0 27784 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _1529_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1530_
timestamp 1688980957
transform 1 0 27508 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1531_
timestamp 1688980957
transform 1 0 26956 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1532_
timestamp 1688980957
transform -1 0 28336 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a2111oi_1  _1533_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28336 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1534_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1535_
timestamp 1688980957
transform -1 0 29992 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1536_
timestamp 1688980957
transform 1 0 29716 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _1537_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30176 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1538_
timestamp 1688980957
transform -1 0 30176 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1539_
timestamp 1688980957
transform 1 0 34316 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1540_
timestamp 1688980957
transform 1 0 36156 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1541_
timestamp 1688980957
transform -1 0 34316 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _1542_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33304 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1543_
timestamp 1688980957
transform 1 0 19412 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _1544_
timestamp 1688980957
transform 1 0 24196 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1545_
timestamp 1688980957
transform 1 0 27140 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1546_
timestamp 1688980957
transform 1 0 27784 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1547_
timestamp 1688980957
transform 1 0 28704 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1548_
timestamp 1688980957
transform 1 0 28060 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1549_
timestamp 1688980957
transform 1 0 27876 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1550_
timestamp 1688980957
transform -1 0 29164 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1551_
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1552_
timestamp 1688980957
transform 1 0 29808 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1553_
timestamp 1688980957
transform -1 0 31096 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1554_
timestamp 1688980957
transform 1 0 28612 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_1  _1555_
timestamp 1688980957
transform -1 0 25484 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1556_
timestamp 1688980957
transform 1 0 25484 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_1  _1557_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26036 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o2111a_1  _1558_
timestamp 1688980957
transform -1 0 24656 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o2111a_1  _1559_
timestamp 1688980957
transform -1 0 25208 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _1560_
timestamp 1688980957
transform 1 0 24656 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _1561_
timestamp 1688980957
transform -1 0 26128 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1562_
timestamp 1688980957
transform 1 0 25760 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1563_
timestamp 1688980957
transform 1 0 25944 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1564_
timestamp 1688980957
transform 1 0 26588 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1565_
timestamp 1688980957
transform -1 0 27416 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1566_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27140 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1567_
timestamp 1688980957
transform -1 0 32108 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1568_
timestamp 1688980957
transform 1 0 33212 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1569_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 36156 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1570_
timestamp 1688980957
transform -1 0 37444 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1571_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35604 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1572_
timestamp 1688980957
transform 1 0 24748 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1573_
timestamp 1688980957
transform -1 0 25116 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1574_
timestamp 1688980957
transform 1 0 24932 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1575_
timestamp 1688980957
transform -1 0 26404 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _1576_
timestamp 1688980957
transform -1 0 26220 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1577_
timestamp 1688980957
transform 1 0 25576 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1578_
timestamp 1688980957
transform -1 0 27600 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _1579_
timestamp 1688980957
transform -1 0 26956 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1580_
timestamp 1688980957
transform 1 0 30176 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1581_
timestamp 1688980957
transform 1 0 28336 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1582_
timestamp 1688980957
transform 1 0 23644 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1583_
timestamp 1688980957
transform 1 0 27876 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1584_
timestamp 1688980957
transform 1 0 27232 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1585_
timestamp 1688980957
transform -1 0 29164 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1586_
timestamp 1688980957
transform 1 0 27692 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1587_
timestamp 1688980957
transform -1 0 28336 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1588_
timestamp 1688980957
transform 1 0 28612 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1589_
timestamp 1688980957
transform 1 0 29256 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1590_
timestamp 1688980957
transform 1 0 30176 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1591_
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1592_
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1593_
timestamp 1688980957
transform -1 0 31004 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1594_
timestamp 1688980957
transform 1 0 31096 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1595_
timestamp 1688980957
transform 1 0 31740 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _1596_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35696 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1597_
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1598_
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1599_
timestamp 1688980957
transform 1 0 22264 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1600_
timestamp 1688980957
transform 1 0 21528 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _1601_
timestamp 1688980957
transform -1 0 22632 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1602_
timestamp 1688980957
transform -1 0 23736 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1603_
timestamp 1688980957
transform 1 0 22724 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _1604_
timestamp 1688980957
transform -1 0 23644 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1605_
timestamp 1688980957
transform 1 0 25300 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1606_
timestamp 1688980957
transform 1 0 22080 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1607_
timestamp 1688980957
transform 1 0 22540 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1608_
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1609_
timestamp 1688980957
transform 1 0 21068 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1610_
timestamp 1688980957
transform 1 0 21528 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1611_
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1612_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22448 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1613_
timestamp 1688980957
transform 1 0 22080 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1614_
timestamp 1688980957
transform 1 0 22724 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1615_
timestamp 1688980957
transform -1 0 23920 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1616_
timestamp 1688980957
transform 1 0 22540 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _1617_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23092 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_4  _1618_
timestamp 1688980957
transform 1 0 24840 0 -1 25024
box -38 -48 2062 592
use sky130_fd_sc_hd__a22oi_1  _1619_
timestamp 1688980957
transform -1 0 20516 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1620_
timestamp 1688980957
transform 1 0 17572 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _1621_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18400 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _1622_
timestamp 1688980957
transform 1 0 20516 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1623_
timestamp 1688980957
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1624_
timestamp 1688980957
transform -1 0 20332 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1625_
timestamp 1688980957
transform -1 0 20976 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1626_
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_2  _1627_
timestamp 1688980957
transform 1 0 19412 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1628_
timestamp 1688980957
transform 1 0 24472 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1629_
timestamp 1688980957
transform -1 0 22724 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1630_
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1631_
timestamp 1688980957
transform 1 0 18860 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1632_
timestamp 1688980957
transform 1 0 21068 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1633_
timestamp 1688980957
transform -1 0 22448 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1634_
timestamp 1688980957
transform 1 0 20976 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1635_
timestamp 1688980957
transform 1 0 21712 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1636_
timestamp 1688980957
transform -1 0 22632 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1637_
timestamp 1688980957
transform 1 0 19872 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1638_
timestamp 1688980957
transform 1 0 20884 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1639_
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_4  _1640_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23092 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__xnor2_4  _1641_
timestamp 1688980957
transform 1 0 25668 0 1 30464
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _1642_
timestamp 1688980957
transform -1 0 28796 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1643_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29808 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1644_
timestamp 1688980957
transform 1 0 25300 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1645_
timestamp 1688980957
transform 1 0 25760 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1646_
timestamp 1688980957
transform -1 0 26128 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1647_
timestamp 1688980957
transform 1 0 28980 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1648_
timestamp 1688980957
transform 1 0 29716 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1649_
timestamp 1688980957
transform -1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1650_
timestamp 1688980957
transform 1 0 24932 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1651_
timestamp 1688980957
transform 1 0 23552 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1652_
timestamp 1688980957
transform 1 0 22632 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1653_
timestamp 1688980957
transform 1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1654_
timestamp 1688980957
transform -1 0 19504 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1655_
timestamp 1688980957
transform 1 0 19596 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1656_
timestamp 1688980957
transform 1 0 18768 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1657_
timestamp 1688980957
transform 1 0 18492 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1658_
timestamp 1688980957
transform 1 0 17204 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1659_
timestamp 1688980957
transform 1 0 17204 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1660_
timestamp 1688980957
transform 1 0 17940 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _1661_
timestamp 1688980957
transform -1 0 18216 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1662_
timestamp 1688980957
transform 1 0 12144 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1663_
timestamp 1688980957
transform 1 0 12788 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1664_
timestamp 1688980957
transform 1 0 11868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1665_
timestamp 1688980957
transform 1 0 12328 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1666_
timestamp 1688980957
transform 1 0 13432 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1667_
timestamp 1688980957
transform -1 0 14352 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1668_
timestamp 1688980957
transform -1 0 14260 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1669_
timestamp 1688980957
transform -1 0 13984 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1670_
timestamp 1688980957
transform 1 0 19964 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1671_
timestamp 1688980957
transform 1 0 20884 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_4  _1672_
timestamp 1688980957
transform -1 0 21620 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _1673_
timestamp 1688980957
transform -1 0 24196 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1674_
timestamp 1688980957
transform -1 0 23368 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _1675_
timestamp 1688980957
transform 1 0 23092 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1676_
timestamp 1688980957
transform 1 0 13156 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1677_
timestamp 1688980957
transform 1 0 14904 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1678_
timestamp 1688980957
transform -1 0 14904 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1679_
timestamp 1688980957
transform 1 0 14812 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1680_
timestamp 1688980957
transform 1 0 15364 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1681_
timestamp 1688980957
transform -1 0 15548 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1682_
timestamp 1688980957
transform -1 0 14904 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1683_
timestamp 1688980957
transform -1 0 17296 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1684_
timestamp 1688980957
transform -1 0 16652 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1685_
timestamp 1688980957
transform 1 0 19780 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1686_
timestamp 1688980957
transform 1 0 20516 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1687_
timestamp 1688980957
transform 1 0 19596 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1688_
timestamp 1688980957
transform -1 0 21068 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1689_
timestamp 1688980957
transform -1 0 20424 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1690_
timestamp 1688980957
transform -1 0 21068 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1691_
timestamp 1688980957
transform -1 0 19872 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1692_
timestamp 1688980957
transform -1 0 20516 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1693_
timestamp 1688980957
transform 1 0 19964 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1694_
timestamp 1688980957
transform 1 0 19780 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1695_
timestamp 1688980957
transform 1 0 19872 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1696_
timestamp 1688980957
transform -1 0 18400 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1697_
timestamp 1688980957
transform 1 0 13524 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1698_
timestamp 1688980957
transform -1 0 14812 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1699_
timestamp 1688980957
transform -1 0 14352 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1700_
timestamp 1688980957
transform 1 0 14352 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _1701_
timestamp 1688980957
transform 1 0 15272 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__and3b_4  _1702_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12696 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_2  _1703_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16192 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1704_
timestamp 1688980957
transform 1 0 22724 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _1705_
timestamp 1688980957
transform 1 0 22448 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__o211ai_4  _1706_
timestamp 1688980957
transform 1 0 21896 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_8  _1707_
timestamp 1688980957
transform -1 0 25392 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_2  _1708_
timestamp 1688980957
transform 1 0 20976 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_2  _1709_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17664 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1710_
timestamp 1688980957
transform 1 0 18124 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1711_
timestamp 1688980957
transform 1 0 22172 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1712_
timestamp 1688980957
transform -1 0 22632 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1713_
timestamp 1688980957
transform 1 0 23552 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1714_
timestamp 1688980957
transform 1 0 32844 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _1715_
timestamp 1688980957
transform -1 0 37996 0 1 23936
box -38 -48 2062 592
use sky130_fd_sc_hd__o211a_1  _1716_
timestamp 1688980957
transform -1 0 33856 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_2  _1717_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30912 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1718_
timestamp 1688980957
transform -1 0 33948 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1719_
timestamp 1688980957
transform 1 0 32936 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1720_
timestamp 1688980957
transform 1 0 33580 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1721_
timestamp 1688980957
transform 1 0 33028 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1722_
timestamp 1688980957
transform 1 0 33028 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1723_
timestamp 1688980957
transform -1 0 31556 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1724_
timestamp 1688980957
transform 1 0 25024 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1725_
timestamp 1688980957
transform 1 0 26128 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1726_
timestamp 1688980957
transform 1 0 26128 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1727_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26588 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1728_
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1729_
timestamp 1688980957
transform -1 0 30084 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_2  _1730_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29256 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1731_
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1732_
timestamp 1688980957
transform 1 0 30084 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1733_
timestamp 1688980957
transform -1 0 26220 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1734_
timestamp 1688980957
transform -1 0 26864 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1735_
timestamp 1688980957
transform -1 0 27692 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1736_
timestamp 1688980957
transform -1 0 27508 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _1737_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27784 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1738_
timestamp 1688980957
transform -1 0 25116 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1739_
timestamp 1688980957
transform -1 0 22356 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1740_
timestamp 1688980957
transform 1 0 21436 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1741_
timestamp 1688980957
transform 1 0 17940 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1742_
timestamp 1688980957
transform -1 0 19136 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1743_
timestamp 1688980957
transform 1 0 17940 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1744_
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1745_
timestamp 1688980957
transform -1 0 15272 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1746_
timestamp 1688980957
transform 1 0 15916 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1747_
timestamp 1688980957
transform -1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1748_
timestamp 1688980957
transform 1 0 17020 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1749_
timestamp 1688980957
transform 1 0 24104 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _1750_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24472 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1751_
timestamp 1688980957
transform 1 0 24196 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__o22ai_4  _1752_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19136 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _1753_
timestamp 1688980957
transform 1 0 25668 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1754_
timestamp 1688980957
transform -1 0 26864 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1755_
timestamp 1688980957
transform 1 0 26128 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1756_
timestamp 1688980957
transform -1 0 26772 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1757_
timestamp 1688980957
transform 1 0 25208 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1758_
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1759_
timestamp 1688980957
transform -1 0 29900 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1760_
timestamp 1688980957
transform 1 0 29164 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1761_
timestamp 1688980957
transform -1 0 30176 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1762_
timestamp 1688980957
transform 1 0 35144 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1763_
timestamp 1688980957
transform -1 0 36340 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1764_
timestamp 1688980957
transform -1 0 37352 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1765_
timestamp 1688980957
transform -1 0 36892 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1766_
timestamp 1688980957
transform -1 0 31924 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1767_
timestamp 1688980957
transform 1 0 30452 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1768_
timestamp 1688980957
transform -1 0 31556 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1769_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 36156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1770_
timestamp 1688980957
transform -1 0 36800 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1771_
timestamp 1688980957
transform 1 0 35972 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1772_
timestamp 1688980957
transform 1 0 36156 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1773_
timestamp 1688980957
transform 1 0 35696 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1774_
timestamp 1688980957
transform 1 0 36340 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1775_
timestamp 1688980957
transform 1 0 32384 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1776_
timestamp 1688980957
transform 1 0 34132 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _1777_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 32016 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1778_
timestamp 1688980957
transform -1 0 30268 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1779_
timestamp 1688980957
transform -1 0 27600 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _1780_
timestamp 1688980957
transform 1 0 21988 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1781_
timestamp 1688980957
transform -1 0 26128 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1782_
timestamp 1688980957
transform -1 0 31464 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1783_
timestamp 1688980957
transform -1 0 26680 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1784_
timestamp 1688980957
transform 1 0 26680 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1785_
timestamp 1688980957
transform -1 0 33028 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1786_
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1787_
timestamp 1688980957
transform -1 0 28060 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1788_
timestamp 1688980957
transform 1 0 27508 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1789_
timestamp 1688980957
transform 1 0 28244 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1790_
timestamp 1688980957
transform -1 0 32476 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1791_
timestamp 1688980957
transform -1 0 31832 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1792_
timestamp 1688980957
transform 1 0 31004 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_1  _1793_
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1794_
timestamp 1688980957
transform 1 0 32844 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1795_
timestamp 1688980957
transform 1 0 33396 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1796_
timestamp 1688980957
transform 1 0 33764 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1797_
timestamp 1688980957
transform 1 0 34868 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _1798_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 30728 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1799_
timestamp 1688980957
transform 1 0 30176 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1800_
timestamp 1688980957
transform -1 0 35236 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1801_
timestamp 1688980957
transform -1 0 35972 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1802_
timestamp 1688980957
transform -1 0 34500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1803_
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1804_
timestamp 1688980957
transform 1 0 35604 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _1805_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33672 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1806_
timestamp 1688980957
transform -1 0 29440 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1807_
timestamp 1688980957
transform -1 0 28980 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1808_
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  _1809_
timestamp 1688980957
transform -1 0 16560 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__a2111oi_1  _1810_
timestamp 1688980957
transform 1 0 27692 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1811_
timestamp 1688980957
transform -1 0 27048 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1812_
timestamp 1688980957
transform -1 0 31096 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1813_
timestamp 1688980957
transform 1 0 30176 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1814_
timestamp 1688980957
transform 1 0 28060 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1815_
timestamp 1688980957
transform 1 0 26220 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1816_
timestamp 1688980957
transform 1 0 25760 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1817_
timestamp 1688980957
transform 1 0 23460 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1818_
timestamp 1688980957
transform 1 0 26496 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1819_
timestamp 1688980957
transform 1 0 27324 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1820_
timestamp 1688980957
transform -1 0 28060 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _1821_
timestamp 1688980957
transform -1 0 23000 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1822_
timestamp 1688980957
transform 1 0 26496 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1823_
timestamp 1688980957
transform 1 0 26128 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1824_
timestamp 1688980957
transform -1 0 32200 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1825_
timestamp 1688980957
transform 1 0 27600 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_4  _1826_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26864 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1827_
timestamp 1688980957
transform -1 0 27508 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1828_
timestamp 1688980957
transform 1 0 27048 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1829_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1830_
timestamp 1688980957
transform -1 0 27324 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1831_
timestamp 1688980957
transform 1 0 23460 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1832_
timestamp 1688980957
transform -1 0 29256 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1833_
timestamp 1688980957
transform 1 0 28796 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1834_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28152 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1835_
timestamp 1688980957
transform 1 0 27600 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1836_
timestamp 1688980957
transform 1 0 27692 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1837_
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1838_
timestamp 1688980957
transform -1 0 27232 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1839_
timestamp 1688980957
transform -1 0 28704 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _1840_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1841_
timestamp 1688980957
transform 1 0 16928 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1842_
timestamp 1688980957
transform 1 0 17204 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1843_
timestamp 1688980957
transform 1 0 10764 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1844_
timestamp 1688980957
transform -1 0 10672 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1845_
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _1846_
timestamp 1688980957
transform -1 0 11132 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1847_
timestamp 1688980957
transform 1 0 10212 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1848_
timestamp 1688980957
transform 1 0 10028 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1849_
timestamp 1688980957
transform -1 0 10120 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1850_
timestamp 1688980957
transform -1 0 11684 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _1851_
timestamp 1688980957
transform 1 0 9476 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1852_
timestamp 1688980957
transform -1 0 9200 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1853_
timestamp 1688980957
transform -1 0 10304 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1854_
timestamp 1688980957
transform -1 0 9568 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1855_
timestamp 1688980957
transform -1 0 9844 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1856_
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1857_
timestamp 1688980957
transform 1 0 9476 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1858_
timestamp 1688980957
transform -1 0 10764 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1859_
timestamp 1688980957
transform -1 0 10120 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_4  _1860_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9844 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__nor2_8  _1861_
timestamp 1688980957
transform 1 0 9384 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _1862_
timestamp 1688980957
transform 1 0 18216 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1863_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1864_
timestamp 1688980957
transform 1 0 30268 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1865_
timestamp 1688980957
transform 1 0 29624 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1866_
timestamp 1688980957
transform -1 0 31740 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1867_
timestamp 1688980957
transform -1 0 30636 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1868_
timestamp 1688980957
transform 1 0 29624 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1869_
timestamp 1688980957
transform 1 0 28244 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1870_
timestamp 1688980957
transform -1 0 28152 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1871_
timestamp 1688980957
transform 1 0 27600 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _1872_
timestamp 1688980957
transform 1 0 27876 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _1873_
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1874_
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1875_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27048 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1876_
timestamp 1688980957
transform 1 0 28060 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1877_
timestamp 1688980957
transform -1 0 28428 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1878_
timestamp 1688980957
transform 1 0 28336 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _1879_
timestamp 1688980957
transform -1 0 30176 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1880_
timestamp 1688980957
transform -1 0 29348 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1881_
timestamp 1688980957
transform 1 0 15548 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1882_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14904 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1883_
timestamp 1688980957
transform -1 0 16192 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1884_
timestamp 1688980957
transform -1 0 14720 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1885_
timestamp 1688980957
transform 1 0 6348 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1886_
timestamp 1688980957
transform 1 0 5244 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1887_
timestamp 1688980957
transform -1 0 35144 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1888_
timestamp 1688980957
transform -1 0 35144 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1889_
timestamp 1688980957
transform 1 0 30912 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1890_
timestamp 1688980957
transform -1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1891_
timestamp 1688980957
transform 1 0 29348 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1892_
timestamp 1688980957
transform -1 0 30176 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1893_
timestamp 1688980957
transform -1 0 30912 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1894_
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1895_
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1896_
timestamp 1688980957
transform 1 0 32200 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1897_
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1898_
timestamp 1688980957
transform -1 0 33672 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _1899_
timestamp 1688980957
transform -1 0 34408 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1900_
timestamp 1688980957
transform 1 0 14812 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1901_
timestamp 1688980957
transform -1 0 16468 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1902_
timestamp 1688980957
transform 1 0 15088 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1903_
timestamp 1688980957
transform -1 0 16008 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1904_
timestamp 1688980957
transform 1 0 15548 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1905_
timestamp 1688980957
transform 1 0 15916 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1906_
timestamp 1688980957
transform 1 0 16560 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _1907_
timestamp 1688980957
transform -1 0 13616 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1908_
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1909_
timestamp 1688980957
transform 1 0 4140 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1910_
timestamp 1688980957
transform 1 0 33672 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1911_
timestamp 1688980957
transform 1 0 36432 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1912_
timestamp 1688980957
transform -1 0 36432 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1913_
timestamp 1688980957
transform -1 0 35420 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1914_
timestamp 1688980957
transform 1 0 31740 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1915_
timestamp 1688980957
transform 1 0 29348 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1916_
timestamp 1688980957
transform 1 0 25576 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1917_
timestamp 1688980957
transform 1 0 30912 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1918_
timestamp 1688980957
transform 1 0 29716 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1919_
timestamp 1688980957
transform 1 0 30728 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1920_
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1921_
timestamp 1688980957
transform 1 0 30452 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1922_
timestamp 1688980957
transform -1 0 31832 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1923_
timestamp 1688980957
transform -1 0 32844 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o221ai_1  _1924_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33764 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1925_
timestamp 1688980957
transform 1 0 35144 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _1926_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34224 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1927_
timestamp 1688980957
transform 1 0 16008 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1928_
timestamp 1688980957
transform 1 0 15364 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1929_
timestamp 1688980957
transform 1 0 15640 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1930_
timestamp 1688980957
transform -1 0 16284 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1931_
timestamp 1688980957
transform 1 0 10396 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1932_
timestamp 1688980957
transform 1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1933_
timestamp 1688980957
transform 1 0 36892 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1934_
timestamp 1688980957
transform -1 0 36984 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1935_
timestamp 1688980957
transform 1 0 36064 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1936_
timestamp 1688980957
transform 1 0 35052 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1937_
timestamp 1688980957
transform -1 0 36708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1938_
timestamp 1688980957
transform -1 0 37904 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__o22a_1  _1939_
timestamp 1688980957
transform -1 0 31096 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1940_
timestamp 1688980957
transform -1 0 31924 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1941_
timestamp 1688980957
transform 1 0 32200 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1942_
timestamp 1688980957
transform -1 0 33304 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1943_
timestamp 1688980957
transform 1 0 33672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1944_
timestamp 1688980957
transform -1 0 34960 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1945_
timestamp 1688980957
transform -1 0 34592 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _1946_
timestamp 1688980957
transform 1 0 34408 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _1947_
timestamp 1688980957
transform -1 0 19228 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1948_
timestamp 1688980957
transform 1 0 18308 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1949_
timestamp 1688980957
transform -1 0 18032 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_2  _1950_
timestamp 1688980957
transform 1 0 17572 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1951_
timestamp 1688980957
transform -1 0 15180 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1952_
timestamp 1688980957
transform 1 0 5336 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1953_
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1954_
timestamp 1688980957
transform -1 0 35696 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1955_
timestamp 1688980957
transform -1 0 34960 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1956_
timestamp 1688980957
transform -1 0 36984 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1957_
timestamp 1688980957
transform -1 0 36892 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1958_
timestamp 1688980957
transform 1 0 36708 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1959_
timestamp 1688980957
transform -1 0 37168 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1960_
timestamp 1688980957
transform 1 0 33212 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1961_
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1962_
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1963_
timestamp 1688980957
transform -1 0 33212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1964_
timestamp 1688980957
transform -1 0 32476 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1965_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32844 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1966_
timestamp 1688980957
transform 1 0 36432 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1967_
timestamp 1688980957
transform -1 0 36616 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_2  _1968_
timestamp 1688980957
transform 1 0 34960 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1969_
timestamp 1688980957
transform 1 0 20332 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1970_
timestamp 1688980957
transform 1 0 20056 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1971_
timestamp 1688980957
transform 1 0 19780 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1972_
timestamp 1688980957
transform 1 0 19320 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1973_
timestamp 1688980957
transform -1 0 16468 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1974_
timestamp 1688980957
transform -1 0 16376 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1975_
timestamp 1688980957
transform 1 0 5244 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1976_
timestamp 1688980957
transform 1 0 4876 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1977_
timestamp 1688980957
transform 1 0 33856 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1978_
timestamp 1688980957
transform 1 0 35512 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1979_
timestamp 1688980957
transform -1 0 35696 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1980_
timestamp 1688980957
transform -1 0 35420 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1981_
timestamp 1688980957
transform 1 0 32844 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1982_
timestamp 1688980957
transform 1 0 33764 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1983_
timestamp 1688980957
transform 1 0 33948 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1984_
timestamp 1688980957
transform -1 0 32384 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1985_
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1986_
timestamp 1688980957
transform -1 0 33396 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _1987_
timestamp 1688980957
transform 1 0 33396 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1988_
timestamp 1688980957
transform 1 0 34776 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1989_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34960 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1990_
timestamp 1688980957
transform 1 0 23092 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1991_
timestamp 1688980957
transform 1 0 22172 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1992_
timestamp 1688980957
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _1993_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 22448 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1994_
timestamp 1688980957
transform -1 0 21160 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1995_
timestamp 1688980957
transform 1 0 23092 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1996_
timestamp 1688980957
transform -1 0 25300 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1997_
timestamp 1688980957
transform 1 0 25116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1998_
timestamp 1688980957
transform 1 0 30084 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1999_
timestamp 1688980957
transform -1 0 32016 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2000_
timestamp 1688980957
transform -1 0 30912 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2001_
timestamp 1688980957
transform 1 0 31464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _2002_
timestamp 1688980957
transform 1 0 30728 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _2003_
timestamp 1688980957
transform -1 0 30544 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _2004_
timestamp 1688980957
transform 1 0 31280 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2005_
timestamp 1688980957
transform -1 0 30084 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2006_
timestamp 1688980957
transform -1 0 28980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2007_
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2008_
timestamp 1688980957
transform 1 0 30084 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_2  _2009_
timestamp 1688980957
transform -1 0 31280 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2010_
timestamp 1688980957
transform -1 0 24656 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2011_
timestamp 1688980957
transform 1 0 23092 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2012_
timestamp 1688980957
transform -1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2013_
timestamp 1688980957
transform -1 0 24196 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _2014_
timestamp 1688980957
transform 1 0 24196 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2015_
timestamp 1688980957
transform 1 0 22816 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2016_
timestamp 1688980957
transform -1 0 30636 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2017_
timestamp 1688980957
transform -1 0 30912 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2018_
timestamp 1688980957
transform 1 0 9752 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _2019_
timestamp 1688980957
transform 1 0 10212 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2020_
timestamp 1688980957
transform 1 0 19320 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2021_
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2022_
timestamp 1688980957
transform 1 0 6532 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2023_
timestamp 1688980957
transform 1 0 5152 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2024_
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2025_
timestamp 1688980957
transform 1 0 5612 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2026_
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2027_
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2028_
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2029_
timestamp 1688980957
transform 1 0 5888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2030_
timestamp 1688980957
transform 1 0 7544 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2031_
timestamp 1688980957
transform 1 0 7176 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2032_
timestamp 1688980957
transform -1 0 27232 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2033_
timestamp 1688980957
transform -1 0 27508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2034_
timestamp 1688980957
transform -1 0 30820 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2035_
timestamp 1688980957
transform -1 0 30820 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _2036_
timestamp 1688980957
transform -1 0 13800 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _2037_
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and4_2  _2038_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12880 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2039_
timestamp 1688980957
transform -1 0 24104 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2040_
timestamp 1688980957
transform -1 0 10120 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2041_
timestamp 1688980957
transform -1 0 9016 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2042_
timestamp 1688980957
transform -1 0 9292 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _2043_
timestamp 1688980957
transform 1 0 9568 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _2044_
timestamp 1688980957
transform 1 0 10120 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_4  _2045_
timestamp 1688980957
transform -1 0 11960 0 1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _2046_
timestamp 1688980957
transform 1 0 21896 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2047_
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2048_
timestamp 1688980957
transform -1 0 15180 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2049_
timestamp 1688980957
transform 1 0 15548 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2050_
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _2051_
timestamp 1688980957
transform 1 0 24104 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2052_
timestamp 1688980957
transform -1 0 34040 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2053_
timestamp 1688980957
transform -1 0 34592 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _2054_
timestamp 1688980957
transform 1 0 21252 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2055_
timestamp 1688980957
transform 1 0 32384 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2056_
timestamp 1688980957
transform -1 0 32660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _2057_
timestamp 1688980957
transform 1 0 13800 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2058_
timestamp 1688980957
transform 1 0 14904 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2059_
timestamp 1688980957
transform 1 0 14996 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2060_
timestamp 1688980957
transform -1 0 17296 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2061_
timestamp 1688980957
transform 1 0 11500 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2062_
timestamp 1688980957
transform 1 0 10488 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _2063_
timestamp 1688980957
transform 1 0 23644 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2064_
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2065_
timestamp 1688980957
transform -1 0 31556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2066_
timestamp 1688980957
transform 1 0 20608 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2067_
timestamp 1688980957
transform 1 0 33212 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2068_
timestamp 1688980957
transform -1 0 33304 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2069_
timestamp 1688980957
transform 1 0 8464 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2070_
timestamp 1688980957
transform 1 0 8832 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _2071_
timestamp 1688980957
transform 1 0 9936 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _2072_
timestamp 1688980957
transform 1 0 10120 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2073_
timestamp 1688980957
transform 1 0 17112 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2074_
timestamp 1688980957
transform -1 0 16560 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2075_
timestamp 1688980957
transform 1 0 7544 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2076_
timestamp 1688980957
transform 1 0 7268 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2077_
timestamp 1688980957
transform 1 0 7636 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2078_
timestamp 1688980957
transform 1 0 7268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2079_
timestamp 1688980957
transform -1 0 12696 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2080_
timestamp 1688980957
transform 1 0 12328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2081_
timestamp 1688980957
transform 1 0 8004 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2082_
timestamp 1688980957
transform 1 0 7636 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2083_
timestamp 1688980957
transform 1 0 7268 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2084_
timestamp 1688980957
transform 1 0 6808 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2085_
timestamp 1688980957
transform -1 0 26772 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2086_
timestamp 1688980957
transform -1 0 26680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2087_
timestamp 1688980957
transform 1 0 23368 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2088_
timestamp 1688980957
transform 1 0 23184 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _2089_
timestamp 1688980957
transform -1 0 11408 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _2090_
timestamp 1688980957
transform 1 0 22908 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2091_
timestamp 1688980957
transform 1 0 22172 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2092_
timestamp 1688980957
transform 1 0 19596 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2093_
timestamp 1688980957
transform -1 0 19596 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2094_
timestamp 1688980957
transform -1 0 32016 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2095_
timestamp 1688980957
transform -1 0 32016 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2096_
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2097_
timestamp 1688980957
transform 1 0 31188 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2098_
timestamp 1688980957
transform 1 0 13432 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2099_
timestamp 1688980957
transform 1 0 12328 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2100_
timestamp 1688980957
transform 1 0 13156 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2101_
timestamp 1688980957
transform 1 0 12788 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2102_
timestamp 1688980957
transform 1 0 29992 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2103_
timestamp 1688980957
transform 1 0 29992 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2104_
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2105_
timestamp 1688980957
transform 1 0 31372 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _2106_
timestamp 1688980957
transform 1 0 9292 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _2107_
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2108_
timestamp 1688980957
transform -1 0 20516 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2109_
timestamp 1688980957
transform 1 0 20516 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2110_
timestamp 1688980957
transform 1 0 9108 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2111_
timestamp 1688980957
transform 1 0 7728 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2112_
timestamp 1688980957
transform 1 0 9292 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2113_
timestamp 1688980957
transform 1 0 9016 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2114_
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2115_
timestamp 1688980957
transform 1 0 14904 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2116_
timestamp 1688980957
transform 1 0 9752 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2117_
timestamp 1688980957
transform 1 0 9476 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2118_
timestamp 1688980957
transform 1 0 8924 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2119_
timestamp 1688980957
transform -1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2120_
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2121_
timestamp 1688980957
transform -1 0 27232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2122_
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2123_
timestamp 1688980957
transform -1 0 27232 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _2124_
timestamp 1688980957
transform -1 0 12788 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2125_
timestamp 1688980957
transform -1 0 24288 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2126_
timestamp 1688980957
transform -1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2127_
timestamp 1688980957
transform 1 0 13892 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2128_
timestamp 1688980957
transform 1 0 13524 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2129_
timestamp 1688980957
transform 1 0 33304 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2130_
timestamp 1688980957
transform -1 0 33304 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2131_
timestamp 1688980957
transform -1 0 33948 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2132_
timestamp 1688980957
transform -1 0 34224 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2133_
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2134_
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2135_
timestamp 1688980957
transform 1 0 14444 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2136_
timestamp 1688980957
transform 1 0 13064 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2137_
timestamp 1688980957
transform -1 0 32016 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2138_
timestamp 1688980957
transform -1 0 31832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2139_
timestamp 1688980957
transform 1 0 33212 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2140_
timestamp 1688980957
transform 1 0 33212 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2141_
timestamp 1688980957
transform -1 0 17756 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2142_
timestamp 1688980957
transform -1 0 17480 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2143_
timestamp 1688980957
transform 1 0 22172 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2144_
timestamp 1688980957
transform 1 0 10028 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2145_
timestamp 1688980957
transform 1 0 9292 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2146_
timestamp 1688980957
transform 1 0 9568 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2147_
timestamp 1688980957
transform 1 0 9476 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _2148_
timestamp 1688980957
transform -1 0 10120 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_2  _2149_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10212 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_2  _2150_
timestamp 1688980957
transform -1 0 10764 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2151_
timestamp 1688980957
transform 1 0 21988 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2152_
timestamp 1688980957
transform -1 0 22080 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2153_
timestamp 1688980957
transform -1 0 28796 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2154_
timestamp 1688980957
transform 1 0 15824 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2155_
timestamp 1688980957
transform 1 0 17940 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2156_
timestamp 1688980957
transform 1 0 18308 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2157_
timestamp 1688980957
transform -1 0 20240 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2158_
timestamp 1688980957
transform -1 0 18308 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2159_
timestamp 1688980957
transform -1 0 17756 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2160_
timestamp 1688980957
transform 1 0 18492 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2161_
timestamp 1688980957
transform -1 0 19136 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2162_
timestamp 1688980957
transform 1 0 19136 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2163_
timestamp 1688980957
transform 1 0 29532 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2164_
timestamp 1688980957
transform 1 0 29624 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2165_
timestamp 1688980957
transform -1 0 13984 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2166_
timestamp 1688980957
transform 1 0 17020 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _2167_
timestamp 1688980957
transform -1 0 25024 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2168_
timestamp 1688980957
transform -1 0 33580 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2169_
timestamp 1688980957
transform 1 0 33948 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2170_
timestamp 1688980957
transform 1 0 35604 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2171_
timestamp 1688980957
transform 1 0 36524 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2172_
timestamp 1688980957
transform 1 0 33672 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2173_
timestamp 1688980957
transform 1 0 34132 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2174_
timestamp 1688980957
transform -1 0 37904 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2175_
timestamp 1688980957
transform 1 0 36156 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2176_
timestamp 1688980957
transform 1 0 32936 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2177_
timestamp 1688980957
transform -1 0 32568 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2178_
timestamp 1688980957
transform -1 0 32292 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _2179_
timestamp 1688980957
transform 1 0 32476 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _2180_
timestamp 1688980957
transform -1 0 37996 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _2181_
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2182_
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2183_
timestamp 1688980957
transform -1 0 20792 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2184_
timestamp 1688980957
transform 1 0 19964 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2185_
timestamp 1688980957
transform 1 0 20424 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2186_
timestamp 1688980957
transform -1 0 20424 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2187_
timestamp 1688980957
transform -1 0 27784 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2188_
timestamp 1688980957
transform 1 0 28060 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2189_
timestamp 1688980957
transform -1 0 29164 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2190_
timestamp 1688980957
transform 1 0 23736 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2191_
timestamp 1688980957
transform -1 0 25024 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2192_
timestamp 1688980957
transform 1 0 20608 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2193_
timestamp 1688980957
transform -1 0 21528 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2194_
timestamp 1688980957
transform 1 0 21252 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2195_
timestamp 1688980957
transform 1 0 22080 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2196_
timestamp 1688980957
transform 1 0 22540 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_4  _2197_
timestamp 1688980957
transform -1 0 35420 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__a21oi_1  _2198_
timestamp 1688980957
transform -1 0 23184 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2199_
timestamp 1688980957
transform 1 0 22356 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2200_
timestamp 1688980957
transform 1 0 18400 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2201_
timestamp 1688980957
transform 1 0 19320 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2202_
timestamp 1688980957
transform 1 0 19688 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2203_
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2204_
timestamp 1688980957
transform 1 0 20516 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2205_
timestamp 1688980957
transform 1 0 21160 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2206_
timestamp 1688980957
transform 1 0 22080 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2207_
timestamp 1688980957
transform 1 0 22908 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_2  _2208_
timestamp 1688980957
transform 1 0 22172 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _2209_
timestamp 1688980957
transform -1 0 17572 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2210_
timestamp 1688980957
transform -1 0 17664 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2211_
timestamp 1688980957
transform 1 0 17664 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2212_
timestamp 1688980957
transform -1 0 29440 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2213_
timestamp 1688980957
transform 1 0 28704 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2214_
timestamp 1688980957
transform 1 0 25668 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2215_
timestamp 1688980957
transform -1 0 25760 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2216_
timestamp 1688980957
transform -1 0 28060 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2217_
timestamp 1688980957
transform 1 0 24748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2218_
timestamp 1688980957
transform -1 0 26036 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2219_
timestamp 1688980957
transform -1 0 28704 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _2220_
timestamp 1688980957
transform 1 0 27232 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _2221_
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2222_
timestamp 1688980957
transform -1 0 19964 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2223_
timestamp 1688980957
transform 1 0 19412 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2224_
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _2225_
timestamp 1688980957
transform -1 0 19780 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2226_
timestamp 1688980957
transform 1 0 23920 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2227_
timestamp 1688980957
transform -1 0 24472 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2228_
timestamp 1688980957
transform -1 0 25208 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2229_
timestamp 1688980957
transform -1 0 25116 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2230_
timestamp 1688980957
transform -1 0 3680 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _2231_
timestamp 1688980957
transform 1 0 3956 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _2232_
timestamp 1688980957
transform -1 0 5428 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _2233_
timestamp 1688980957
transform -1 0 5060 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2234_
timestamp 1688980957
transform 1 0 3312 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2235_
timestamp 1688980957
transform -1 0 4968 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _2236_
timestamp 1688980957
transform -1 0 10028 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_2  _2237_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5244 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _2238_
timestamp 1688980957
transform -1 0 4508 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _2239_
timestamp 1688980957
transform -1 0 3588 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2240_
timestamp 1688980957
transform -1 0 4600 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2241_
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2242_
timestamp 1688980957
transform -1 0 4968 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _2243_
timestamp 1688980957
transform -1 0 12420 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _2244_
timestamp 1688980957
transform -1 0 12328 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2245_
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _2246_
timestamp 1688980957
transform 1 0 7084 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2247_
timestamp 1688980957
transform -1 0 7360 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2248_
timestamp 1688980957
transform 1 0 6624 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _2249_
timestamp 1688980957
transform 1 0 7084 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2250_
timestamp 1688980957
transform -1 0 8280 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2251_
timestamp 1688980957
transform 1 0 6348 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2252_
timestamp 1688980957
transform -1 0 5980 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _2253_
timestamp 1688980957
transform -1 0 7084 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2254_
timestamp 1688980957
transform -1 0 7728 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2255_
timestamp 1688980957
transform -1 0 7544 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2256_
timestamp 1688980957
transform 1 0 5612 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2257_
timestamp 1688980957
transform -1 0 5060 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _2258_
timestamp 1688980957
transform -1 0 5704 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _2259_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7268 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _2260_
timestamp 1688980957
transform -1 0 6072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2261_
timestamp 1688980957
transform -1 0 6900 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2262_
timestamp 1688980957
transform -1 0 6992 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _2263_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6072 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2264_
timestamp 1688980957
transform 1 0 6808 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2265_
timestamp 1688980957
transform 1 0 5060 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2266_
timestamp 1688980957
transform 1 0 4600 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2267_
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2268_
timestamp 1688980957
transform -1 0 4416 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2269_
timestamp 1688980957
transform -1 0 4048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2270_
timestamp 1688980957
transform 1 0 2208 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__buf_8  _2271_
timestamp 1688980957
transform -1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _2272_
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2273_
timestamp 1688980957
transform -1 0 37628 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2274_
timestamp 1688980957
transform 1 0 30820 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2275_
timestamp 1688980957
transform -1 0 31924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2276_
timestamp 1688980957
transform -1 0 5152 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2277_
timestamp 1688980957
transform 1 0 1932 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2278_
timestamp 1688980957
transform -1 0 5612 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2279_
timestamp 1688980957
transform 1 0 1748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2280_
timestamp 1688980957
transform -1 0 12512 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2281_
timestamp 1688980957
transform -1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2282_
timestamp 1688980957
transform -1 0 4600 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2283_
timestamp 1688980957
transform 1 0 1748 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2284_
timestamp 1688980957
transform 1 0 30544 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2285_
timestamp 1688980957
transform -1 0 37628 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2286_
timestamp 1688980957
transform 1 0 19320 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2287_
timestamp 1688980957
transform -1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_2  _2288_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14444 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _2289_
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_8  _2290_
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _2291_
timestamp 1688980957
transform 1 0 16100 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2292_
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2293_
timestamp 1688980957
transform 1 0 12788 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _2294_
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2295_
timestamp 1688980957
transform -1 0 19780 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2296_
timestamp 1688980957
transform 1 0 18860 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2297_
timestamp 1688980957
transform 1 0 18952 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2298_
timestamp 1688980957
transform -1 0 21160 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2299_
timestamp 1688980957
transform 1 0 19964 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2300_
timestamp 1688980957
transform 1 0 22724 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2301_
timestamp 1688980957
transform -1 0 24196 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2302_
timestamp 1688980957
transform 1 0 22908 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2303_
timestamp 1688980957
transform -1 0 24288 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2304_
timestamp 1688980957
transform -1 0 25484 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2305_
timestamp 1688980957
transform -1 0 25668 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2306_
timestamp 1688980957
transform 1 0 25024 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2307_
timestamp 1688980957
transform 1 0 25208 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2308_
timestamp 1688980957
transform 1 0 25484 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2309_
timestamp 1688980957
transform -1 0 26680 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2310_
timestamp 1688980957
transform 1 0 16008 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2311_
timestamp 1688980957
transform 1 0 15824 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2312_
timestamp 1688980957
transform 1 0 14904 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2313_
timestamp 1688980957
transform -1 0 14536 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2314_
timestamp 1688980957
transform 1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2315_
timestamp 1688980957
transform -1 0 13524 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2316_
timestamp 1688980957
transform -1 0 13524 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2317_
timestamp 1688980957
transform 1 0 1748 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2318_
timestamp 1688980957
transform 1 0 19872 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2319_
timestamp 1688980957
transform -1 0 20792 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2320_
timestamp 1688980957
transform 1 0 13524 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2321_
timestamp 1688980957
transform -1 0 14904 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2322_
timestamp 1688980957
transform 1 0 12512 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2323_
timestamp 1688980957
transform -1 0 14812 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2324_
timestamp 1688980957
transform 1 0 13064 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2325_
timestamp 1688980957
transform 1 0 12972 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2326_
timestamp 1688980957
transform 1 0 12788 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2327_
timestamp 1688980957
transform 1 0 13248 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _2328_
timestamp 1688980957
transform 1 0 13248 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2329_
timestamp 1688980957
transform -1 0 13248 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2330_
timestamp 1688980957
transform -1 0 2024 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _2331_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2332_
timestamp 1688980957
transform 1 0 12512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2333_
timestamp 1688980957
transform 1 0 28152 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2334_
timestamp 1688980957
transform -1 0 37168 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2335_
timestamp 1688980957
transform 1 0 28612 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2336_
timestamp 1688980957
transform -1 0 37628 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2337_
timestamp 1688980957
transform -1 0 11868 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2338_
timestamp 1688980957
transform 1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2339_
timestamp 1688980957
transform -1 0 11684 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2340_
timestamp 1688980957
transform 1 0 1932 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2341_
timestamp 1688980957
transform 1 0 28060 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2342_
timestamp 1688980957
transform -1 0 33672 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2343_
timestamp 1688980957
transform -1 0 12052 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2344_
timestamp 1688980957
transform 1 0 11408 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2345_
timestamp 1688980957
transform -1 0 12512 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2346_
timestamp 1688980957
transform 1 0 10212 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2347_
timestamp 1688980957
transform 1 0 25300 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2348_
timestamp 1688980957
transform -1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2349_
timestamp 1688980957
transform 1 0 2300 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2350_
timestamp 1688980957
transform 1 0 1748 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2351_
timestamp 1688980957
transform -1 0 5060 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2352_
timestamp 1688980957
transform 1 0 3128 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2353_
timestamp 1688980957
transform 1 0 3220 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2354_
timestamp 1688980957
transform 1 0 1840 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2355_
timestamp 1688980957
transform 1 0 5796 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2356_
timestamp 1688980957
transform 1 0 5888 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2357_
timestamp 1688980957
transform 1 0 6808 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2358_
timestamp 1688980957
transform -1 0 6992 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2359_
timestamp 1688980957
transform 1 0 6624 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2360_
timestamp 1688980957
transform -1 0 6624 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2361_
timestamp 1688980957
transform -1 0 5612 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2362_
timestamp 1688980957
transform 1 0 4692 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2363_
timestamp 1688980957
transform 1 0 4416 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2364_
timestamp 1688980957
transform -1 0 8464 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2365_
timestamp 1688980957
transform 1 0 8464 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2366_
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2367_
timestamp 1688980957
transform 1 0 8096 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2368_
timestamp 1688980957
transform -1 0 8004 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2369_
timestamp 1688980957
transform 1 0 8004 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2370_
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2371_
timestamp 1688980957
transform 1 0 8280 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2372_
timestamp 1688980957
transform -1 0 5152 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2373_
timestamp 1688980957
transform 1 0 4508 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2374_
timestamp 1688980957
transform 1 0 5060 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2375_
timestamp 1688980957
transform 1 0 4600 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2376_
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2377_
timestamp 1688980957
transform 1 0 5612 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2378_
timestamp 1688980957
transform 1 0 3680 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2379_
timestamp 1688980957
transform 1 0 2944 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2380_
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2381_
timestamp 1688980957
transform 1 0 3312 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2382_
timestamp 1688980957
transform 1 0 6440 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2383_
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2384_
timestamp 1688980957
transform 1 0 8004 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2385_
timestamp 1688980957
transform -1 0 8004 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2386_
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2387_
timestamp 1688980957
transform 1 0 2300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2388_
timestamp 1688980957
transform -1 0 9752 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2389_
timestamp 1688980957
transform -1 0 9476 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2390_
timestamp 1688980957
transform 1 0 5152 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2391_
timestamp 1688980957
transform 1 0 4784 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2392_
timestamp 1688980957
transform 1 0 6716 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2393_
timestamp 1688980957
transform 1 0 6440 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2394_
timestamp 1688980957
transform 1 0 4324 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2395_
timestamp 1688980957
transform 1 0 4048 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2396_
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2397_
timestamp 1688980957
transform 1 0 1932 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2398_
timestamp 1688980957
transform 1 0 7268 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2399_
timestamp 1688980957
transform 1 0 6992 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2400_
timestamp 1688980957
transform 1 0 9016 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2401_
timestamp 1688980957
transform -1 0 8924 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2402_
timestamp 1688980957
transform 1 0 2576 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2403_
timestamp 1688980957
transform 1 0 1932 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2404_
timestamp 1688980957
transform -1 0 11132 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2405_
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2406_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2407_
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2408__8
timestamp 1688980957
transform -1 0 25576 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2409__9
timestamp 1688980957
transform -1 0 29072 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2410__10
timestamp 1688980957
transform -1 0 17848 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2411__11
timestamp 1688980957
transform -1 0 12512 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2412__12
timestamp 1688980957
transform -1 0 30544 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2413__13
timestamp 1688980957
transform 1 0 29716 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2414__14
timestamp 1688980957
transform 1 0 19412 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2415__15
timestamp 1688980957
transform 1 0 21528 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2416__16
timestamp 1688980957
transform -1 0 33028 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2417__17
timestamp 1688980957
transform -1 0 32476 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2418__18
timestamp 1688980957
transform -1 0 12972 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2419__19
timestamp 1688980957
transform -1 0 13156 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2420__20
timestamp 1688980957
transform 1 0 33396 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2421__21
timestamp 1688980957
transform 1 0 35328 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2422__22
timestamp 1688980957
transform -1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2423__23
timestamp 1688980957
transform -1 0 24288 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2424__24
timestamp 1688980957
transform 1 0 26496 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2425__25
timestamp 1688980957
transform -1 0 27784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2426__26
timestamp 1688980957
transform -1 0 8832 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2427_
timestamp 1688980957
transform 1 0 6900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2428__27
timestamp 1688980957
transform -1 0 9476 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2429__28
timestamp 1688980957
transform 1 0 14628 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2430__29
timestamp 1688980957
transform -1 0 9016 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2431__30
timestamp 1688980957
transform -1 0 7544 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2432__31
timestamp 1688980957
transform -1 0 21068 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2433__32
timestamp 1688980957
transform 1 0 30820 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2434__33
timestamp 1688980957
transform -1 0 29992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2435__34
timestamp 1688980957
transform -1 0 12604 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2436__35
timestamp 1688980957
transform -1 0 11960 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2437__36
timestamp 1688980957
transform 1 0 30728 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2438__37
timestamp 1688980957
transform 1 0 32200 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2439__38
timestamp 1688980957
transform -1 0 20700 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2440__39
timestamp 1688980957
transform -1 0 22172 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2441__40
timestamp 1688980957
transform -1 0 22816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2442__41
timestamp 1688980957
transform -1 0 27324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2443__42
timestamp 1688980957
transform -1 0 6716 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2444__43
timestamp 1688980957
transform 1 0 6716 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2445__44
timestamp 1688980957
transform -1 0 12328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2446__45
timestamp 1688980957
transform -1 0 6716 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2447_
timestamp 1688980957
transform 1 0 5336 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2448__46
timestamp 1688980957
transform 1 0 6440 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2449__47
timestamp 1688980957
transform -1 0 17020 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2450__48
timestamp 1688980957
transform -1 0 33672 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2451__49
timestamp 1688980957
transform -1 0 31832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2452__50
timestamp 1688980957
transform -1 0 10028 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2453__51
timestamp 1688980957
transform -1 0 15088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2454__52
timestamp 1688980957
transform -1 0 33028 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2455__53
timestamp 1688980957
transform 1 0 34040 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2456__54
timestamp 1688980957
transform -1 0 15088 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2457__55
timestamp 1688980957
transform -1 0 21068 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2458__56
timestamp 1688980957
transform -1 0 31188 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2459__57
timestamp 1688980957
transform -1 0 28152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2460__58
timestamp 1688980957
transform 1 0 6440 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2461__59
timestamp 1688980957
transform 1 0 5152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2462__60
timestamp 1688980957
transform -1 0 10580 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2463__61
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2464__62
timestamp 1688980957
transform -1 0 4968 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2465__63
timestamp 1688980957
transform 1 0 19504 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2466__64
timestamp 1688980957
transform 1 0 30360 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2467__1
timestamp 1688980957
transform 1 0 23920 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2468__2
timestamp 1688980957
transform 1 0 4048 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2469__3
timestamp 1688980957
transform -1 0 4692 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2470__4
timestamp 1688980957
transform 1 0 9016 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2471__5
timestamp 1688980957
transform -1 0 4048 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2472__6
timestamp 1688980957
transform 1 0 4416 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2473__7
timestamp 1688980957
transform 1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2474_
timestamp 1688980957
transform 1 0 12420 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2475_
timestamp 1688980957
transform 1 0 13524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2476_
timestamp 1688980957
transform -1 0 20332 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2477_
timestamp 1688980957
transform -1 0 26128 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2478_
timestamp 1688980957
transform 1 0 19504 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2479_
timestamp 1688980957
transform -1 0 16928 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2480_
timestamp 1688980957
transform 1 0 18124 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2481_
timestamp 1688980957
transform 1 0 18492 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2482_
timestamp 1688980957
transform 1 0 17204 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2483_
timestamp 1688980957
transform 1 0 17480 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2484_
timestamp 1688980957
transform 1 0 18400 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2485_
timestamp 1688980957
transform 1 0 17664 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2486_
timestamp 1688980957
transform -1 0 18676 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2487_
timestamp 1688980957
transform -1 0 18124 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _2488_
timestamp 1688980957
transform -1 0 18676 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o41a_1  _2489_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _2490_
timestamp 1688980957
transform 1 0 16284 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2491_
timestamp 1688980957
transform 1 0 16928 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _2492_
timestamp 1688980957
transform 1 0 15364 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2493_
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _2494_
timestamp 1688980957
transform -1 0 14628 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _2495_
timestamp 1688980957
transform 1 0 15640 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _2496_
timestamp 1688980957
transform -1 0 17020 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _2497_
timestamp 1688980957
transform -1 0 20056 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_8  _2498_
timestamp 1688980957
transform -1 0 5796 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _2499_
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2500_
timestamp 1688980957
transform 1 0 18492 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2501_
timestamp 1688980957
transform -1 0 24840 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2502_
timestamp 1688980957
transform 1 0 25392 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _2503_
timestamp 1688980957
transform 1 0 22540 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2504_
timestamp 1688980957
transform 1 0 23276 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2505_
timestamp 1688980957
transform 1 0 22540 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2506_
timestamp 1688980957
transform 1 0 22264 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2507_
timestamp 1688980957
transform -1 0 21436 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2508_
timestamp 1688980957
transform -1 0 21528 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2509_
timestamp 1688980957
transform -1 0 22448 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2510_
timestamp 1688980957
transform -1 0 21804 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2511_
timestamp 1688980957
transform 1 0 20700 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2512_
timestamp 1688980957
transform 1 0 20332 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2513_
timestamp 1688980957
transform 1 0 20056 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2514_
timestamp 1688980957
transform -1 0 21160 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2515_
timestamp 1688980957
transform 1 0 22448 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2516_
timestamp 1688980957
transform 1 0 22724 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2517_
timestamp 1688980957
transform 1 0 22448 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2518_
timestamp 1688980957
transform -1 0 22448 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2519_
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2520_
timestamp 1688980957
transform 1 0 20976 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2521_
timestamp 1688980957
transform -1 0 26036 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _2522_
timestamp 1688980957
transform 1 0 24932 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2523_
timestamp 1688980957
transform 1 0 25208 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2524_
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2525_
timestamp 1688980957
transform 1 0 23736 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2526_
timestamp 1688980957
transform 1 0 25944 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2527_
timestamp 1688980957
transform 1 0 24932 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _2528_
timestamp 1688980957
transform -1 0 26036 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2529_
timestamp 1688980957
transform -1 0 26036 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2530_
timestamp 1688980957
transform -1 0 25392 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2531_
timestamp 1688980957
transform 1 0 24840 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2532_
timestamp 1688980957
transform 1 0 24380 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2533_
timestamp 1688980957
transform -1 0 24288 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2534_
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2535_
timestamp 1688980957
transform -1 0 17756 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2536_
timestamp 1688980957
transform 1 0 17940 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2537_
timestamp 1688980957
transform -1 0 18124 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2538_
timestamp 1688980957
transform 1 0 18124 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2539_
timestamp 1688980957
transform 1 0 17572 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2540_
timestamp 1688980957
transform 1 0 17572 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2541_
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _2542_
timestamp 1688980957
transform 1 0 16100 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2543_
timestamp 1688980957
transform 1 0 16744 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2544_
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2545_
timestamp 1688980957
transform 1 0 15548 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2546_
timestamp 1688980957
transform -1 0 16560 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2547_
timestamp 1688980957
transform 1 0 16100 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2548_
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _2549_
timestamp 1688980957
transform -1 0 15824 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _2550_
timestamp 1688980957
transform 1 0 16376 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2551_
timestamp 1688980957
transform 1 0 14904 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2552_
timestamp 1688980957
transform 1 0 14628 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2553_
timestamp 1688980957
transform 1 0 12512 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2554_
timestamp 1688980957
transform -1 0 12052 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2555_
timestamp 1688980957
transform -1 0 12512 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2556_
timestamp 1688980957
transform 1 0 11316 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2557_
timestamp 1688980957
transform 1 0 10580 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2558_
timestamp 1688980957
transform 1 0 10028 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2559_
timestamp 1688980957
transform -1 0 13340 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2560_
timestamp 1688980957
transform 1 0 13432 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2561_
timestamp 1688980957
transform -1 0 13432 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2562_
timestamp 1688980957
transform -1 0 12788 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2563_
timestamp 1688980957
transform -1 0 12972 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2564_
timestamp 1688980957
transform -1 0 13248 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2565_
timestamp 1688980957
transform -1 0 11408 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2566_
timestamp 1688980957
transform 1 0 12052 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2567_
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2568_
timestamp 1688980957
transform 1 0 9384 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2569_
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2570_
timestamp 1688980957
transform 1 0 11684 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2571_
timestamp 1688980957
transform -1 0 12696 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2572_
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2573_
timestamp 1688980957
transform 1 0 10396 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2574_
timestamp 1688980957
transform 1 0 9752 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2575_
timestamp 1688980957
transform -1 0 11868 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2576_
timestamp 1688980957
transform 1 0 11132 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2577_
timestamp 1688980957
transform 1 0 11592 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _2578_
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2579_
timestamp 1688980957
transform 1 0 10304 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2580_
timestamp 1688980957
transform 1 0 9752 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2581_
timestamp 1688980957
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2582_
timestamp 1688980957
transform 1 0 11408 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2583_
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2584_
timestamp 1688980957
transform 1 0 10120 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2585_
timestamp 1688980957
transform 1 0 9660 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2586_
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2587_
timestamp 1688980957
transform -1 0 12788 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2588_
timestamp 1688980957
transform 1 0 11316 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2589_
timestamp 1688980957
transform -1 0 11316 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _2590_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2591_
timestamp 1688980957
transform 1 0 1840 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2592_
timestamp 1688980957
transform -1 0 3404 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2593_
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2594_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5152 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2595_
timestamp 1688980957
transform 1 0 6992 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2596_
timestamp 1688980957
transform 1 0 6348 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2597_
timestamp 1688980957
transform 1 0 4048 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2598_
timestamp 1688980957
transform 1 0 7636 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2599_
timestamp 1688980957
transform 1 0 6992 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2600_
timestamp 1688980957
transform 1 0 6992 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2601_
timestamp 1688980957
transform 1 0 8004 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2602_
timestamp 1688980957
transform 1 0 4048 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2603_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5060 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2604_
timestamp 1688980957
transform 1 0 1840 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2605_
timestamp 1688980957
transform 1 0 2760 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2606_
timestamp 1688980957
transform 1 0 5704 0 1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2607_
timestamp 1688980957
transform 1 0 8004 0 -1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2608_
timestamp 1688980957
transform 1 0 1564 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2609_
timestamp 1688980957
transform 1 0 9476 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2610_
timestamp 1688980957
transform 1 0 4324 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2611_
timestamp 1688980957
transform 1 0 6164 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2612_
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2613_
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2614_
timestamp 1688980957
transform 1 0 6624 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2615_
timestamp 1688980957
transform 1 0 8924 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2616_
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2617_
timestamp 1688980957
transform 1 0 11132 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2618_
timestamp 1688980957
transform 1 0 25208 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2619_
timestamp 1688980957
transform 1 0 28704 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2620_
timestamp 1688980957
transform 1 0 17020 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2621_
timestamp 1688980957
transform 1 0 12144 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2622_
timestamp 1688980957
transform 1 0 30176 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2623_
timestamp 1688980957
transform 1 0 29992 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2624_
timestamp 1688980957
transform 1 0 19688 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2625_
timestamp 1688980957
transform 1 0 22080 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2626_
timestamp 1688980957
transform 1 0 32660 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2627_
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2628_
timestamp 1688980957
transform 1 0 11960 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2629_
timestamp 1688980957
transform 1 0 12788 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2630_
timestamp 1688980957
transform -1 0 35144 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2631_
timestamp 1688980957
transform -1 0 35420 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2632_
timestamp 1688980957
transform 1 0 12972 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2633_
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2634_
timestamp 1688980957
transform 1 0 26772 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2635_
timestamp 1688980957
transform 1 0 27416 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2636_
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2637_
timestamp 1688980957
transform 1 0 9108 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2638_
timestamp 1688980957
transform 1 0 14536 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2639_
timestamp 1688980957
transform 1 0 8648 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2640_
timestamp 1688980957
transform 1 0 7176 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2641_
timestamp 1688980957
transform 1 0 19780 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2642_
timestamp 1688980957
transform 1 0 31096 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2643_
timestamp 1688980957
transform 1 0 29624 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2644_
timestamp 1688980957
transform 1 0 12236 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2645_
timestamp 1688980957
transform 1 0 11592 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2646_
timestamp 1688980957
transform 1 0 31004 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2647_
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2648_
timestamp 1688980957
transform 1 0 19596 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2649_
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2650_
timestamp 1688980957
transform 1 0 22448 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2651_
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2652_
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2653_
timestamp 1688980957
transform 1 0 6992 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2654_
timestamp 1688980957
transform 1 0 11868 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2655_
timestamp 1688980957
transform 1 0 6716 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2656_
timestamp 1688980957
transform 1 0 6716 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2657_
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2658_
timestamp 1688980957
transform 1 0 33304 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2659_
timestamp 1688980957
transform 1 0 31464 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2660_
timestamp 1688980957
transform 1 0 9568 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2661_
timestamp 1688980957
transform 1 0 14720 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2662_
timestamp 1688980957
transform 1 0 32660 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2663_
timestamp 1688980957
transform -1 0 35144 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2664_
timestamp 1688980957
transform 1 0 14720 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2665_
timestamp 1688980957
transform 1 0 21068 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2666_
timestamp 1688980957
transform 1 0 30820 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2667_
timestamp 1688980957
transform 1 0 27784 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2668_
timestamp 1688980957
transform 1 0 6716 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2669_
timestamp 1688980957
transform 1 0 5428 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2670_
timestamp 1688980957
transform 1 0 10212 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2671_
timestamp 1688980957
transform 1 0 5152 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2672_
timestamp 1688980957
transform 1 0 4600 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2673_
timestamp 1688980957
transform 1 0 18952 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2674_
timestamp 1688980957
transform 1 0 30636 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2675_
timestamp 1688980957
transform 1 0 23828 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2676_
timestamp 1688980957
transform 1 0 4324 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2677_
timestamp 1688980957
transform 1 0 4140 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2678_
timestamp 1688980957
transform 1 0 9292 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2679_
timestamp 1688980957
transform 1 0 3496 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2680_
timestamp 1688980957
transform 1 0 4692 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2681_
timestamp 1688980957
transform 1 0 17296 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2682_
timestamp 1688980957
transform 1 0 18124 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2683_
timestamp 1688980957
transform 1 0 21804 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2684_
timestamp 1688980957
transform 1 0 19688 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2685_
timestamp 1688980957
transform 1 0 20700 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2686_
timestamp 1688980957
transform 1 0 23276 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2687_
timestamp 1688980957
transform 1 0 24380 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2688_
timestamp 1688980957
transform 1 0 17296 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2689_
timestamp 1688980957
transform 1 0 14996 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2690_
timestamp 1688980957
transform 1 0 14168 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2691_
timestamp 1688980957
transform 1 0 9476 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2692_
timestamp 1688980957
transform 1 0 12788 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2693_
timestamp 1688980957
transform 1 0 8188 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2694_
timestamp 1688980957
transform 1 0 9200 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2695_
timestamp 1688980957
transform 1 0 9292 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2696_
timestamp 1688980957
transform 1 0 9108 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2697_
timestamp 1688980957
transform 1 0 11500 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2698_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5520 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2699_
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2700_
timestamp 1688980957
transform -1 0 5612 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2701_
timestamp 1688980957
transform -1 0 6900 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2702_
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2703_
timestamp 1688980957
transform 1 0 2116 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0514_
timestamp 1688980957
transform 1 0 13892 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0515_
timestamp 1688980957
transform 1 0 22264 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0516_
timestamp 1688980957
transform 1 0 19320 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0517_
timestamp 1688980957
transform 1 0 19044 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1688980957
transform 1 0 12972 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0514_
timestamp 1688980957
transform -1 0 9660 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0515_
timestamp 1688980957
transform -1 0 17480 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0516_
timestamp 1688980957
transform -1 0 14812 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0517_
timestamp 1688980957
transform -1 0 14812 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0514_
timestamp 1688980957
transform -1 0 14536 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0515_
timestamp 1688980957
transform 1 0 26036 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0516_
timestamp 1688980957
transform 1 0 23368 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0517_
timestamp 1688980957
transform 1 0 23368 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1688980957
transform -1 0 8096 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1688980957
transform -1 0 7084 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1688980957
transform 1 0 12972 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  fanout58
timestamp 1688980957
transform 1 0 14076 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout59
timestamp 1688980957
transform -1 0 19136 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout60
timestamp 1688980957
transform 1 0 30636 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  fanout61
timestamp 1688980957
transform 1 0 33672 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout62
timestamp 1688980957
transform -1 0 13800 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  fanout63
timestamp 1688980957
transform 1 0 15364 0 1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout64
timestamp 1688980957
transform -1 0 35236 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_16 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_37
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1688980957
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_77
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_97 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_105
timestamp 1688980957
transform 1 0 10764 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_127
timestamp 1688980957
transform 1 0 12788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_153 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_172
timestamp 1688980957
transform 1 0 16928 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_184
timestamp 1688980957
transform 1 0 18032 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_212
timestamp 1688980957
transform 1 0 20608 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_264
timestamp 1688980957
transform 1 0 25392 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_276
timestamp 1688980957
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_287
timestamp 1688980957
transform 1 0 27508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_299
timestamp 1688980957
transform 1 0 28612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 1688980957
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_331
timestamp 1688980957
transform 1 0 31556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_335
timestamp 1688980957
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1688980957
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_373
timestamp 1688980957
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_378
timestamp 1688980957
transform 1 0 35880 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_390
timestamp 1688980957
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_399
timestamp 1688980957
transform 1 0 37812 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_12
timestamp 1688980957
transform 1 0 2208 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_24
timestamp 1688980957
transform 1 0 3312 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_36
timestamp 1688980957
transform 1 0 4416 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_48
timestamp 1688980957
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_61
timestamp 1688980957
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_65
timestamp 1688980957
transform 1 0 7084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_77
timestamp 1688980957
transform 1 0 8188 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_89
timestamp 1688980957
transform 1 0 9292 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_98
timestamp 1688980957
transform 1 0 10120 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_110
timestamp 1688980957
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_175
timestamp 1688980957
transform 1 0 17204 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_197
timestamp 1688980957
transform 1 0 19228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_246
timestamp 1688980957
transform 1 0 23736 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_278
timestamp 1688980957
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_301
timestamp 1688980957
transform 1 0 28796 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_313
timestamp 1688980957
transform 1 0 29900 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_321
timestamp 1688980957
transform 1 0 30636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_328
timestamp 1688980957
transform 1 0 31280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_61
timestamp 1688980957
transform 1 0 6716 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_66
timestamp 1688980957
transform 1 0 7176 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_78
timestamp 1688980957
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_146
timestamp 1688980957
transform 1 0 14536 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_162
timestamp 1688980957
transform 1 0 16008 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_170
timestamp 1688980957
transform 1 0 16744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_201
timestamp 1688980957
transform 1 0 19596 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_217
timestamp 1688980957
transform 1 0 21068 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_225
timestamp 1688980957
transform 1 0 21804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_232
timestamp 1688980957
transform 1 0 22448 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_244
timestamp 1688980957
transform 1 0 23552 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_268
timestamp 1688980957
transform 1 0 25760 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_279
timestamp 1688980957
transform 1 0 26772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_285
timestamp 1688980957
transform 1 0 27324 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_293
timestamp 1688980957
transform 1 0 28060 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_299
timestamp 1688980957
transform 1 0 28612 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_399
timestamp 1688980957
transform 1 0 37812 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_190
timestamp 1688980957
transform 1 0 18584 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_202
timestamp 1688980957
transform 1 0 19688 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_214
timestamp 1688980957
transform 1 0 20792 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_222
timestamp 1688980957
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_228
timestamp 1688980957
transform 1 0 22080 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_240
timestamp 1688980957
transform 1 0 23184 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_252
timestamp 1688980957
transform 1 0 24288 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_264
timestamp 1688980957
transform 1 0 25392 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_276
timestamp 1688980957
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_311
timestamp 1688980957
transform 1 0 29716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_323
timestamp 1688980957
transform 1 0 30820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_7
timestamp 1688980957
transform 1 0 1748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_19
timestamp 1688980957
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_88
timestamp 1688980957
transform 1 0 9200 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_100
timestamp 1688980957
transform 1 0 10304 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_112
timestamp 1688980957
transform 1 0 11408 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_124
timestamp 1688980957
transform 1 0 12512 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_132
timestamp 1688980957
transform 1 0 13248 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_136
timestamp 1688980957
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_149
timestamp 1688980957
transform 1 0 14812 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_154
timestamp 1688980957
transform 1 0 15272 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_166
timestamp 1688980957
transform 1 0 16376 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_173
timestamp 1688980957
transform 1 0 17020 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_185
timestamp 1688980957
transform 1 0 18124 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 1688980957
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_207
timestamp 1688980957
transform 1 0 20148 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_213
timestamp 1688980957
transform 1 0 20700 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_274
timestamp 1688980957
transform 1 0 26312 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_284
timestamp 1688980957
transform 1 0 27232 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_10
timestamp 1688980957
transform 1 0 2024 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_22
timestamp 1688980957
transform 1 0 3128 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_34
timestamp 1688980957
transform 1 0 4232 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_49
timestamp 1688980957
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_65
timestamp 1688980957
transform 1 0 7084 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_70
timestamp 1688980957
transform 1 0 7544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_80
timestamp 1688980957
transform 1 0 8464 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_108
timestamp 1688980957
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_122
timestamp 1688980957
transform 1 0 12328 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_126
timestamp 1688980957
transform 1 0 12696 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_147
timestamp 1688980957
transform 1 0 14628 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_215
timestamp 1688980957
transform 1 0 20884 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_235
timestamp 1688980957
transform 1 0 22724 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_252
timestamp 1688980957
transform 1 0 24288 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_264
timestamp 1688980957
transform 1 0 25392 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_276
timestamp 1688980957
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_290
timestamp 1688980957
transform 1 0 27784 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_294
timestamp 1688980957
transform 1 0 28152 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_306
timestamp 1688980957
transform 1 0 29256 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_310
timestamp 1688980957
transform 1 0 29624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_323
timestamp 1688980957
transform 1 0 30820 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_327
timestamp 1688980957
transform 1 0 31188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_334
timestamp 1688980957
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_346
timestamp 1688980957
transform 1 0 32936 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_358
timestamp 1688980957
transform 1 0 34040 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_370
timestamp 1688980957
transform 1 0 35144 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_382
timestamp 1688980957
transform 1 0 36248 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_390
timestamp 1688980957
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_49
timestamp 1688980957
transform 1 0 5612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_57
timestamp 1688980957
transform 1 0 6348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_98
timestamp 1688980957
transform 1 0 10120 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_125
timestamp 1688980957
transform 1 0 12604 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_131
timestamp 1688980957
transform 1 0 13156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_159
timestamp 1688980957
transform 1 0 15732 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_171
timestamp 1688980957
transform 1 0 16836 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_182
timestamp 1688980957
transform 1 0 17848 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_194
timestamp 1688980957
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_203
timestamp 1688980957
transform 1 0 19780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_215
timestamp 1688980957
transform 1 0 20884 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_227
timestamp 1688980957
transform 1 0 21988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_239
timestamp 1688980957
transform 1 0 23092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_264
timestamp 1688980957
transform 1 0 25392 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_276
timestamp 1688980957
transform 1 0 26496 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_288
timestamp 1688980957
transform 1 0 27600 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_300
timestamp 1688980957
transform 1 0 28704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_351
timestamp 1688980957
transform 1 0 33396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_86
timestamp 1688980957
transform 1 0 9016 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_98
timestamp 1688980957
transform 1 0 10120 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_103
timestamp 1688980957
transform 1 0 10580 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_143
timestamp 1688980957
transform 1 0 14260 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_152
timestamp 1688980957
transform 1 0 15088 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_164
timestamp 1688980957
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_187
timestamp 1688980957
transform 1 0 18308 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_199
timestamp 1688980957
transform 1 0 19412 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_208
timestamp 1688980957
transform 1 0 20240 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_216
timestamp 1688980957
transform 1 0 20976 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_234
timestamp 1688980957
transform 1 0 22632 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_245
timestamp 1688980957
transform 1 0 23644 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_274
timestamp 1688980957
transform 1 0 26312 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_294
timestamp 1688980957
transform 1 0 28152 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_306
timestamp 1688980957
transform 1 0 29256 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_68
timestamp 1688980957
transform 1 0 7360 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_80
timestamp 1688980957
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_118
timestamp 1688980957
transform 1 0 11960 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_130
timestamp 1688980957
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_138
timestamp 1688980957
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_155
timestamp 1688980957
transform 1 0 15364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_167
timestamp 1688980957
transform 1 0 16468 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_178
timestamp 1688980957
transform 1 0 17480 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_184
timestamp 1688980957
transform 1 0 18032 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_193
timestamp 1688980957
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_205
timestamp 1688980957
transform 1 0 19964 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_212
timestamp 1688980957
transform 1 0 20608 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_220
timestamp 1688980957
transform 1 0 21344 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_246
timestamp 1688980957
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_268
timestamp 1688980957
transform 1 0 25760 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_304
timestamp 1688980957
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_314
timestamp 1688980957
transform 1 0 29992 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_326
timestamp 1688980957
transform 1 0 31096 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_330
timestamp 1688980957
transform 1 0 31464 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_334
timestamp 1688980957
transform 1 0 31832 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_346
timestamp 1688980957
transform 1 0 32936 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_358
timestamp 1688980957
transform 1 0 34040 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_66
timestamp 1688980957
transform 1 0 7176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_70
timestamp 1688980957
transform 1 0 7544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_74
timestamp 1688980957
transform 1 0 7912 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_84
timestamp 1688980957
transform 1 0 8832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_108
timestamp 1688980957
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_124
timestamp 1688980957
transform 1 0 12512 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_128
timestamp 1688980957
transform 1 0 12880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_195
timestamp 1688980957
transform 1 0 19044 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_203
timestamp 1688980957
transform 1 0 19780 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_222
timestamp 1688980957
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_232
timestamp 1688980957
transform 1 0 22448 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_262
timestamp 1688980957
transform 1 0 25208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_275
timestamp 1688980957
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_308
timestamp 1688980957
transform 1 0 29440 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_319
timestamp 1688980957
transform 1 0 30452 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_358
timestamp 1688980957
transform 1 0 34040 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_370
timestamp 1688980957
transform 1 0 35144 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_382
timestamp 1688980957
transform 1 0 36248 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_390
timestamp 1688980957
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_44
timestamp 1688980957
transform 1 0 5152 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_55
timestamp 1688980957
transform 1 0 6164 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_103
timestamp 1688980957
transform 1 0 10580 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_111
timestamp 1688980957
transform 1 0 11316 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_149
timestamp 1688980957
transform 1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_171
timestamp 1688980957
transform 1 0 16836 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_175
timestamp 1688980957
transform 1 0 17204 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_184
timestamp 1688980957
transform 1 0 18032 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_192
timestamp 1688980957
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_217
timestamp 1688980957
transform 1 0 21068 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_229
timestamp 1688980957
transform 1 0 22172 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_240
timestamp 1688980957
transform 1 0 23184 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_263
timestamp 1688980957
transform 1 0 25300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_275
timestamp 1688980957
transform 1 0 26404 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_287
timestamp 1688980957
transform 1 0 27508 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_293
timestamp 1688980957
transform 1 0 28060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_305
timestamp 1688980957
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_322
timestamp 1688980957
transform 1 0 30728 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_334
timestamp 1688980957
transform 1 0 31832 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_341
timestamp 1688980957
transform 1 0 32476 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_353
timestamp 1688980957
transform 1 0 33580 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_361
timestamp 1688980957
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_156
timestamp 1688980957
transform 1 0 15456 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_177
timestamp 1688980957
transform 1 0 17388 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_186
timestamp 1688980957
transform 1 0 18216 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_198
timestamp 1688980957
transform 1 0 19320 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_202
timestamp 1688980957
transform 1 0 19688 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_232
timestamp 1688980957
transform 1 0 22448 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_248
timestamp 1688980957
transform 1 0 23920 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_260
timestamp 1688980957
transform 1 0 25024 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_284
timestamp 1688980957
transform 1 0 27232 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_288
timestamp 1688980957
transform 1 0 27600 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_303
timestamp 1688980957
transform 1 0 28980 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_315
timestamp 1688980957
transform 1 0 30084 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_320
timestamp 1688980957
transform 1 0 30544 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_332
timestamp 1688980957
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_343
timestamp 1688980957
transform 1 0 32660 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_347
timestamp 1688980957
transform 1 0 33028 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_359
timestamp 1688980957
transform 1 0 34132 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_371
timestamp 1688980957
transform 1 0 35236 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_383
timestamp 1688980957
transform 1 0 36340 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_35
timestamp 1688980957
transform 1 0 4324 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_39
timestamp 1688980957
transform 1 0 4692 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_51
timestamp 1688980957
transform 1 0 5796 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_63
timestamp 1688980957
transform 1 0 6900 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_75
timestamp 1688980957
transform 1 0 8004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_101
timestamp 1688980957
transform 1 0 10396 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_122
timestamp 1688980957
transform 1 0 12328 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_154
timestamp 1688980957
transform 1 0 15272 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_181
timestamp 1688980957
transform 1 0 17756 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_190
timestamp 1688980957
transform 1 0 18584 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_229
timestamp 1688980957
transform 1 0 22172 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_238
timestamp 1688980957
transform 1 0 23000 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_250
timestamp 1688980957
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_274
timestamp 1688980957
transform 1 0 26312 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_286
timestamp 1688980957
transform 1 0 27416 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_293
timestamp 1688980957
transform 1 0 28060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_305
timestamp 1688980957
transform 1 0 29164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_336
timestamp 1688980957
transform 1 0 32016 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_78
timestamp 1688980957
transform 1 0 8280 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_90
timestamp 1688980957
transform 1 0 9384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_117
timestamp 1688980957
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_159
timestamp 1688980957
transform 1 0 15732 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_189
timestamp 1688980957
transform 1 0 18492 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_197
timestamp 1688980957
transform 1 0 19228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_218
timestamp 1688980957
transform 1 0 21160 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_238
timestamp 1688980957
transform 1 0 23000 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_244
timestamp 1688980957
transform 1 0 23552 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_252
timestamp 1688980957
transform 1 0 24288 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_261
timestamp 1688980957
transform 1 0 25116 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_275
timestamp 1688980957
transform 1 0 26404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1688980957
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_288
timestamp 1688980957
transform 1 0 27600 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_300
timestamp 1688980957
transform 1 0 28704 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_308
timestamp 1688980957
transform 1 0 29440 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_317
timestamp 1688980957
transform 1 0 30268 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_331
timestamp 1688980957
transform 1 0 31556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1688980957
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_370
timestamp 1688980957
transform 1 0 35144 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_382
timestamp 1688980957
transform 1 0 36248 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_390
timestamp 1688980957
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_61
timestamp 1688980957
transform 1 0 6716 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_76
timestamp 1688980957
transform 1 0 8096 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_106
timestamp 1688980957
transform 1 0 10856 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_118
timestamp 1688980957
transform 1 0 11960 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_129
timestamp 1688980957
transform 1 0 12972 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_137
timestamp 1688980957
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_185
timestamp 1688980957
transform 1 0 18124 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_193
timestamp 1688980957
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_213
timestamp 1688980957
transform 1 0 20700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_225
timestamp 1688980957
transform 1 0 21804 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_234
timestamp 1688980957
transform 1 0 22632 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_242
timestamp 1688980957
transform 1 0 23368 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1688980957
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_267
timestamp 1688980957
transform 1 0 25668 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_298
timestamp 1688980957
transform 1 0 28520 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_304
timestamp 1688980957
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_321
timestamp 1688980957
transform 1 0 30636 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_346
timestamp 1688980957
transform 1 0 32936 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_350
timestamp 1688980957
transform 1 0 33304 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_354
timestamp 1688980957
transform 1 0 33672 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_362
timestamp 1688980957
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_365
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_377
timestamp 1688980957
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_389
timestamp 1688980957
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_39
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_44
timestamp 1688980957
transform 1 0 5152 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1688980957
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_79
timestamp 1688980957
transform 1 0 8372 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_97
timestamp 1688980957
transform 1 0 10028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp 1688980957
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_128
timestamp 1688980957
transform 1 0 12880 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_136
timestamp 1688980957
transform 1 0 13616 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_145
timestamp 1688980957
transform 1 0 14444 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_151
timestamp 1688980957
transform 1 0 14996 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_166
timestamp 1688980957
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_221
timestamp 1688980957
transform 1 0 21436 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_231
timestamp 1688980957
transform 1 0 22356 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_262
timestamp 1688980957
transform 1 0 25208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_274
timestamp 1688980957
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_305
timestamp 1688980957
transform 1 0 29164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_313
timestamp 1688980957
transform 1 0 29900 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_325
timestamp 1688980957
transform 1 0 31004 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_330
timestamp 1688980957
transform 1 0 31464 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_346
timestamp 1688980957
transform 1 0 32936 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_360
timestamp 1688980957
transform 1 0 34224 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_372
timestamp 1688980957
transform 1 0 35328 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_384
timestamp 1688980957
transform 1 0 36432 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_393
timestamp 1688980957
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_37
timestamp 1688980957
transform 1 0 4508 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_44
timestamp 1688980957
transform 1 0 5152 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_56
timestamp 1688980957
transform 1 0 6256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1688980957
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_107
timestamp 1688980957
transform 1 0 10948 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_122
timestamp 1688980957
transform 1 0 12328 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_126
timestamp 1688980957
transform 1 0 12696 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_130
timestamp 1688980957
transform 1 0 13064 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_150
timestamp 1688980957
transform 1 0 14904 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_173
timestamp 1688980957
transform 1 0 17020 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_184
timestamp 1688980957
transform 1 0 18032 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_204
timestamp 1688980957
transform 1 0 19872 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_247
timestamp 1688980957
transform 1 0 23828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1688980957
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_264
timestamp 1688980957
transform 1 0 25392 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_281
timestamp 1688980957
transform 1 0 26956 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_289
timestamp 1688980957
transform 1 0 27692 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1688980957
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1688980957
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_323
timestamp 1688980957
transform 1 0 30820 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_335
timestamp 1688980957
transform 1 0 31924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_347
timestamp 1688980957
transform 1 0 33028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_359
timestamp 1688980957
transform 1 0 34132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 1688980957
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_365
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_377
timestamp 1688980957
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_389
timestamp 1688980957
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_12
timestamp 1688980957
transform 1 0 2208 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_24
timestamp 1688980957
transform 1 0 3312 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_36
timestamp 1688980957
transform 1 0 4416 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_48
timestamp 1688980957
transform 1 0 5520 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_52
timestamp 1688980957
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_117
timestamp 1688980957
transform 1 0 11868 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1688980957
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_174
timestamp 1688980957
transform 1 0 17112 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_196
timestamp 1688980957
transform 1 0 19136 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_208
timestamp 1688980957
transform 1 0 20240 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_219
timestamp 1688980957
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1688980957
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_263
timestamp 1688980957
transform 1 0 25300 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_275
timestamp 1688980957
transform 1 0 26404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1688980957
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1688980957
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_305
timestamp 1688980957
transform 1 0 29164 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_316
timestamp 1688980957
transform 1 0 30176 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_330
timestamp 1688980957
transform 1 0 31464 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_370
timestamp 1688980957
transform 1 0 35144 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_382
timestamp 1688980957
transform 1 0 36248 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_390
timestamp 1688980957
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_393
timestamp 1688980957
transform 1 0 37260 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_36
timestamp 1688980957
transform 1 0 4416 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_40
timestamp 1688980957
transform 1 0 4784 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_67
timestamp 1688980957
transform 1 0 7268 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_79
timestamp 1688980957
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_89
timestamp 1688980957
transform 1 0 9292 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_115
timestamp 1688980957
transform 1 0 11684 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_121
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_125
timestamp 1688980957
transform 1 0 12604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_137
timestamp 1688980957
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_174
timestamp 1688980957
transform 1 0 17112 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_182
timestamp 1688980957
transform 1 0 17848 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_192
timestamp 1688980957
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 1688980957
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_221
timestamp 1688980957
transform 1 0 21436 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_225
timestamp 1688980957
transform 1 0 21804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_248
timestamp 1688980957
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_267
timestamp 1688980957
transform 1 0 25668 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_279
timestamp 1688980957
transform 1 0 26772 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1688980957
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 1688980957
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1688980957
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_309
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_335
timestamp 1688980957
transform 1 0 31924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_347
timestamp 1688980957
transform 1 0 33028 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 1688980957
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 1688980957
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_23
timestamp 1688980957
transform 1 0 3220 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_49
timestamp 1688980957
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_77
timestamp 1688980957
transform 1 0 8188 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 1688980957
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_119
timestamp 1688980957
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_127
timestamp 1688980957
transform 1 0 12788 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_150
timestamp 1688980957
transform 1 0 14904 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_162
timestamp 1688980957
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1688980957
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_193
timestamp 1688980957
transform 1 0 18860 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_197
timestamp 1688980957
transform 1 0 19228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_221
timestamp 1688980957
transform 1 0 21436 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_229
timestamp 1688980957
transform 1 0 22172 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_250
timestamp 1688980957
transform 1 0 24104 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_254
timestamp 1688980957
transform 1 0 24472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_297
timestamp 1688980957
transform 1 0 28428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_305
timestamp 1688980957
transform 1 0 29164 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_314
timestamp 1688980957
transform 1 0 29992 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_326
timestamp 1688980957
transform 1 0 31096 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_357
timestamp 1688980957
transform 1 0 33948 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_369
timestamp 1688980957
transform 1 0 35052 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_381
timestamp 1688980957
transform 1 0 36156 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_389
timestamp 1688980957
transform 1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_393
timestamp 1688980957
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_32
timestamp 1688980957
transform 1 0 4048 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_40
timestamp 1688980957
transform 1 0 4784 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_50
timestamp 1688980957
transform 1 0 5704 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1688980957
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_91
timestamp 1688980957
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 1688980957
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_156
timestamp 1688980957
transform 1 0 15456 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_166
timestamp 1688980957
transform 1 0 16376 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_174
timestamp 1688980957
transform 1 0 17112 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 1688980957
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_213
timestamp 1688980957
transform 1 0 20700 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_225
timestamp 1688980957
transform 1 0 21804 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_237
timestamp 1688980957
transform 1 0 22908 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_249
timestamp 1688980957
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_263
timestamp 1688980957
transform 1 0 25300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_286
timestamp 1688980957
transform 1 0 27416 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_303
timestamp 1688980957
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1688980957
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_336
timestamp 1688980957
transform 1 0 32016 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_341
timestamp 1688980957
transform 1 0 32476 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_359
timestamp 1688980957
transform 1 0 34132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 1688980957
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_377
timestamp 1688980957
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_389
timestamp 1688980957
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_9
timestamp 1688980957
transform 1 0 1932 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_21
timestamp 1688980957
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_33
timestamp 1688980957
transform 1 0 4140 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_42
timestamp 1688980957
transform 1 0 4968 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_47
timestamp 1688980957
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_65
timestamp 1688980957
transform 1 0 7084 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_70
timestamp 1688980957
transform 1 0 7544 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_82
timestamp 1688980957
transform 1 0 8648 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_94
timestamp 1688980957
transform 1 0 9752 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_105
timestamp 1688980957
transform 1 0 10764 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_133
timestamp 1688980957
transform 1 0 13340 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_138
timestamp 1688980957
transform 1 0 13800 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_177
timestamp 1688980957
transform 1 0 17388 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_186
timestamp 1688980957
transform 1 0 18216 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_192
timestamp 1688980957
transform 1 0 18768 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_200
timestamp 1688980957
transform 1 0 19504 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_212
timestamp 1688980957
transform 1 0 20608 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_216
timestamp 1688980957
transform 1 0 20976 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_222
timestamp 1688980957
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_232
timestamp 1688980957
transform 1 0 22448 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_236
timestamp 1688980957
transform 1 0 22816 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_251
timestamp 1688980957
transform 1 0 24196 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_263
timestamp 1688980957
transform 1 0 25300 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_275
timestamp 1688980957
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1688980957
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_292
timestamp 1688980957
transform 1 0 27968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_304
timestamp 1688980957
transform 1 0 29072 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_308
timestamp 1688980957
transform 1 0 29440 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_316
timestamp 1688980957
transform 1 0 30176 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_328
timestamp 1688980957
transform 1 0 31280 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_332
timestamp 1688980957
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_346
timestamp 1688980957
transform 1 0 32936 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_373
timestamp 1688980957
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_385
timestamp 1688980957
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 1688980957
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_393
timestamp 1688980957
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_68
timestamp 1688980957
transform 1 0 7360 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_79
timestamp 1688980957
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_93
timestamp 1688980957
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_110
timestamp 1688980957
transform 1 0 11224 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_125
timestamp 1688980957
transform 1 0 12604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_137
timestamp 1688980957
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_152
timestamp 1688980957
transform 1 0 15088 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_164
timestamp 1688980957
transform 1 0 16192 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_176
timestamp 1688980957
transform 1 0 17296 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_186
timestamp 1688980957
transform 1 0 18216 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1688980957
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_211
timestamp 1688980957
transform 1 0 20516 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_215
timestamp 1688980957
transform 1 0 20884 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_223
timestamp 1688980957
transform 1 0 21620 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_230
timestamp 1688980957
transform 1 0 22264 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1688980957
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1688980957
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_298
timestamp 1688980957
transform 1 0 28520 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_306
timestamp 1688980957
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_321
timestamp 1688980957
transform 1 0 30636 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_347
timestamp 1688980957
transform 1 0 33028 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_358
timestamp 1688980957
transform 1 0 34040 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_365
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_371
timestamp 1688980957
transform 1 0 35236 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_375
timestamp 1688980957
transform 1 0 35604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_387
timestamp 1688980957
transform 1 0 36708 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_395
timestamp 1688980957
transform 1 0 37444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_10
timestamp 1688980957
transform 1 0 2024 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_22
timestamp 1688980957
transform 1 0 3128 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_34
timestamp 1688980957
transform 1 0 4232 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_46
timestamp 1688980957
transform 1 0 5336 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 1688980957
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_65
timestamp 1688980957
transform 1 0 7084 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_96
timestamp 1688980957
transform 1 0 9936 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1688980957
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_117
timestamp 1688980957
transform 1 0 11868 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1688980957
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_137
timestamp 1688980957
transform 1 0 13708 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_145
timestamp 1688980957
transform 1 0 14444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_162
timestamp 1688980957
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_173
timestamp 1688980957
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_195
timestamp 1688980957
transform 1 0 19044 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_209
timestamp 1688980957
transform 1 0 20332 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_218
timestamp 1688980957
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_230
timestamp 1688980957
transform 1 0 22264 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_238
timestamp 1688980957
transform 1 0 23000 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_243
timestamp 1688980957
transform 1 0 23460 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_265
timestamp 1688980957
transform 1 0 25484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_269
timestamp 1688980957
transform 1 0 25852 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_277
timestamp 1688980957
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_305
timestamp 1688980957
transform 1 0 29164 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_313
timestamp 1688980957
transform 1 0 29900 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_323
timestamp 1688980957
transform 1 0 30820 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_327
timestamp 1688980957
transform 1 0 31188 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 1688980957
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_345
timestamp 1688980957
transform 1 0 32844 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_370
timestamp 1688980957
transform 1 0 35144 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_382
timestamp 1688980957
transform 1 0 36248 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_390
timestamp 1688980957
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_393
timestamp 1688980957
transform 1 0 37260 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_35
timestamp 1688980957
transform 1 0 4324 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_62
timestamp 1688980957
transform 1 0 6808 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_66
timestamp 1688980957
transform 1 0 7176 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_70
timestamp 1688980957
transform 1 0 7544 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_75
timestamp 1688980957
transform 1 0 8004 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_93
timestamp 1688980957
transform 1 0 9660 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_100
timestamp 1688980957
transform 1 0 10304 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_108
timestamp 1688980957
transform 1 0 11040 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_123
timestamp 1688980957
transform 1 0 12420 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_131
timestamp 1688980957
transform 1 0 13156 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_153
timestamp 1688980957
transform 1 0 15180 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_192
timestamp 1688980957
transform 1 0 18768 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_223
timestamp 1688980957
transform 1 0 21620 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_229
timestamp 1688980957
transform 1 0 22172 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_235
timestamp 1688980957
transform 1 0 22724 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_247
timestamp 1688980957
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_257
timestamp 1688980957
transform 1 0 24748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_281
timestamp 1688980957
transform 1 0 26956 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_305
timestamp 1688980957
transform 1 0 29164 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_316
timestamp 1688980957
transform 1 0 30176 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_344
timestamp 1688980957
transform 1 0 32752 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_350
timestamp 1688980957
transform 1 0 33304 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_354
timestamp 1688980957
transform 1 0 33672 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_362
timestamp 1688980957
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_365
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_377
timestamp 1688980957
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_389
timestamp 1688980957
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_12
timestamp 1688980957
transform 1 0 2208 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_24
timestamp 1688980957
transform 1 0 3312 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_33
timestamp 1688980957
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_48
timestamp 1688980957
transform 1 0 5520 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_82
timestamp 1688980957
transform 1 0 8648 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_88
timestamp 1688980957
transform 1 0 9200 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_104
timestamp 1688980957
transform 1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_121
timestamp 1688980957
transform 1 0 12236 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_139
timestamp 1688980957
transform 1 0 13892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_155
timestamp 1688980957
transform 1 0 15364 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_173
timestamp 1688980957
transform 1 0 17020 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_193
timestamp 1688980957
transform 1 0 18860 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_216
timestamp 1688980957
transform 1 0 20976 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_234
timestamp 1688980957
transform 1 0 22632 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_246
timestamp 1688980957
transform 1 0 23736 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_263
timestamp 1688980957
transform 1 0 25300 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_267
timestamp 1688980957
transform 1 0 25668 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_276
timestamp 1688980957
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_289
timestamp 1688980957
transform 1 0 27692 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_296
timestamp 1688980957
transform 1 0 28336 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_326
timestamp 1688980957
transform 1 0 31096 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_334
timestamp 1688980957
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_337
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_343
timestamp 1688980957
transform 1 0 32660 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_347
timestamp 1688980957
transform 1 0 33028 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_358
timestamp 1688980957
transform 1 0 34040 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_370
timestamp 1688980957
transform 1 0 35144 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_382
timestamp 1688980957
transform 1 0 36248 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_390
timestamp 1688980957
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_393
timestamp 1688980957
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_7
timestamp 1688980957
transform 1 0 1748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_44
timestamp 1688980957
transform 1 0 5152 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_56
timestamp 1688980957
transform 1 0 6256 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_66
timestamp 1688980957
transform 1 0 7176 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_80
timestamp 1688980957
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_88
timestamp 1688980957
transform 1 0 9200 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_124
timestamp 1688980957
transform 1 0 12512 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_132
timestamp 1688980957
transform 1 0 13248 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_151
timestamp 1688980957
transform 1 0 14996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_163
timestamp 1688980957
transform 1 0 16100 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_171
timestamp 1688980957
transform 1 0 16836 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_192
timestamp 1688980957
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1688980957
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_221
timestamp 1688980957
transform 1 0 21436 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_241
timestamp 1688980957
transform 1 0 23276 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_249
timestamp 1688980957
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_265
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_269
timestamp 1688980957
transform 1 0 25852 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_282
timestamp 1688980957
transform 1 0 27048 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_294
timestamp 1688980957
transform 1 0 28152 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_306
timestamp 1688980957
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_317
timestamp 1688980957
transform 1 0 30268 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_342
timestamp 1688980957
transform 1 0 32568 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_365
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_377
timestamp 1688980957
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_389
timestamp 1688980957
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_19
timestamp 1688980957
transform 1 0 2852 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_23
timestamp 1688980957
transform 1 0 3220 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_31
timestamp 1688980957
transform 1 0 3956 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_52
timestamp 1688980957
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_68
timestamp 1688980957
transform 1 0 7360 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_95
timestamp 1688980957
transform 1 0 9844 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_108
timestamp 1688980957
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_132
timestamp 1688980957
transform 1 0 13248 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_136
timestamp 1688980957
transform 1 0 13616 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_145
timestamp 1688980957
transform 1 0 14444 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_151
timestamp 1688980957
transform 1 0 14996 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1688980957
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1688980957
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_178
timestamp 1688980957
transform 1 0 17480 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_197
timestamp 1688980957
transform 1 0 19228 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_209
timestamp 1688980957
transform 1 0 20332 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_220
timestamp 1688980957
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_229
timestamp 1688980957
transform 1 0 22172 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_244
timestamp 1688980957
transform 1 0 23552 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_265
timestamp 1688980957
transform 1 0 25484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_277
timestamp 1688980957
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_290
timestamp 1688980957
transform 1 0 27784 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_302
timestamp 1688980957
transform 1 0 28888 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_310
timestamp 1688980957
transform 1 0 29624 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_324
timestamp 1688980957
transform 1 0 30912 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_352
timestamp 1688980957
transform 1 0 33488 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_371
timestamp 1688980957
transform 1 0 35236 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_383
timestamp 1688980957
transform 1 0 36340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 1688980957
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_393
timestamp 1688980957
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_37
timestamp 1688980957
transform 1 0 4508 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1688980957
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_97
timestamp 1688980957
transform 1 0 10028 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_107
timestamp 1688980957
transform 1 0 10948 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_119
timestamp 1688980957
transform 1 0 12052 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_126
timestamp 1688980957
transform 1 0 12696 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_138
timestamp 1688980957
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_147
timestamp 1688980957
transform 1 0 14628 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_176
timestamp 1688980957
transform 1 0 17296 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_227
timestamp 1688980957
transform 1 0 21988 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_246
timestamp 1688980957
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_271
timestamp 1688980957
transform 1 0 26036 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_275
timestamp 1688980957
transform 1 0 26404 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1688980957
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_319
timestamp 1688980957
transform 1 0 30452 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_325
timestamp 1688980957
transform 1 0 31004 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_337
timestamp 1688980957
transform 1 0 32108 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_349
timestamp 1688980957
transform 1 0 33212 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_361
timestamp 1688980957
transform 1 0 34316 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_377
timestamp 1688980957
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_389
timestamp 1688980957
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_37
timestamp 1688980957
transform 1 0 4508 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_52
timestamp 1688980957
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_65
timestamp 1688980957
transform 1 0 7084 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_88
timestamp 1688980957
transform 1 0 9200 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_96
timestamp 1688980957
transform 1 0 9936 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_102
timestamp 1688980957
transform 1 0 10488 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_110
timestamp 1688980957
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1688980957
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_137
timestamp 1688980957
transform 1 0 13708 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_149
timestamp 1688980957
transform 1 0 14812 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_157
timestamp 1688980957
transform 1 0 15548 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_183
timestamp 1688980957
transform 1 0 17940 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_195
timestamp 1688980957
transform 1 0 19044 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_203
timestamp 1688980957
transform 1 0 19780 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1688980957
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_230
timestamp 1688980957
transform 1 0 22264 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_258
timestamp 1688980957
transform 1 0 24840 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_262
timestamp 1688980957
transform 1 0 25208 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_272
timestamp 1688980957
transform 1 0 26128 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_284
timestamp 1688980957
transform 1 0 27232 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_296
timestamp 1688980957
transform 1 0 28336 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_333
timestamp 1688980957
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_342
timestamp 1688980957
transform 1 0 32568 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_356
timestamp 1688980957
transform 1 0 33856 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_368
timestamp 1688980957
transform 1 0 34960 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_380
timestamp 1688980957
transform 1 0 36064 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_393
timestamp 1688980957
transform 1 0 37260 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_16
timestamp 1688980957
transform 1 0 2576 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_38
timestamp 1688980957
transform 1 0 4600 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_46
timestamp 1688980957
transform 1 0 5336 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_52
timestamp 1688980957
transform 1 0 5888 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_64
timestamp 1688980957
transform 1 0 6992 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_72
timestamp 1688980957
transform 1 0 7728 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_82
timestamp 1688980957
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_103
timestamp 1688980957
transform 1 0 10580 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_115
timestamp 1688980957
transform 1 0 11684 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_119
timestamp 1688980957
transform 1 0 12052 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_134
timestamp 1688980957
transform 1 0 13432 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_162
timestamp 1688980957
transform 1 0 16008 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_176
timestamp 1688980957
transform 1 0 17296 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_188
timestamp 1688980957
transform 1 0 18400 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_239
timestamp 1688980957
transform 1 0 23092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_261
timestamp 1688980957
transform 1 0 25116 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_273
timestamp 1688980957
transform 1 0 26220 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_285
timestamp 1688980957
transform 1 0 27324 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_297
timestamp 1688980957
transform 1 0 28428 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_304
timestamp 1688980957
transform 1 0 29072 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_321
timestamp 1688980957
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_333
timestamp 1688980957
transform 1 0 31740 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_339
timestamp 1688980957
transform 1 0 32292 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_343
timestamp 1688980957
transform 1 0 32660 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_347
timestamp 1688980957
transform 1 0 33028 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_365
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_377
timestamp 1688980957
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_389
timestamp 1688980957
transform 1 0 36892 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_393
timestamp 1688980957
transform 1 0 37260 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_397
timestamp 1688980957
transform 1 0 37628 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_24
timestamp 1688980957
transform 1 0 3312 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_44
timestamp 1688980957
transform 1 0 5152 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_66
timestamp 1688980957
transform 1 0 7176 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_78
timestamp 1688980957
transform 1 0 8280 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_90
timestamp 1688980957
transform 1 0 9384 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_101
timestamp 1688980957
transform 1 0 10396 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_109
timestamp 1688980957
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_122
timestamp 1688980957
transform 1 0 12328 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_131
timestamp 1688980957
transform 1 0 13156 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_141
timestamp 1688980957
transform 1 0 14076 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_145
timestamp 1688980957
transform 1 0 14444 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_149
timestamp 1688980957
transform 1 0 14812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_162
timestamp 1688980957
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_194
timestamp 1688980957
transform 1 0 18952 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_206
timestamp 1688980957
transform 1 0 20056 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_218
timestamp 1688980957
transform 1 0 21160 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_236
timestamp 1688980957
transform 1 0 22816 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_248
timestamp 1688980957
transform 1 0 23920 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_256
timestamp 1688980957
transform 1 0 24656 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_261
timestamp 1688980957
transform 1 0 25116 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_266
timestamp 1688980957
transform 1 0 25576 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_276
timestamp 1688980957
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_286
timestamp 1688980957
transform 1 0 27416 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_306
timestamp 1688980957
transform 1 0 29256 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_318
timestamp 1688980957
transform 1 0 30360 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_322
timestamp 1688980957
transform 1 0 30728 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_328
timestamp 1688980957
transform 1 0 31280 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_335
timestamp 1688980957
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_349
timestamp 1688980957
transform 1 0 33212 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_360
timestamp 1688980957
transform 1 0 34224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_371
timestamp 1688980957
transform 1 0 35236 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_376
timestamp 1688980957
transform 1 0 35696 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_388
timestamp 1688980957
transform 1 0 36800 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_393
timestamp 1688980957
transform 1 0 37260 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_397
timestamp 1688980957
transform 1 0 37628 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_12
timestamp 1688980957
transform 1 0 2208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_25
timestamp 1688980957
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_50
timestamp 1688980957
transform 1 0 5704 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_54
timestamp 1688980957
transform 1 0 6072 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_76
timestamp 1688980957
transform 1 0 8096 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_89
timestamp 1688980957
transform 1 0 9292 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_105
timestamp 1688980957
transform 1 0 10764 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_117
timestamp 1688980957
transform 1 0 11868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_128
timestamp 1688980957
transform 1 0 12880 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_137
timestamp 1688980957
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_149
timestamp 1688980957
transform 1 0 14812 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_183
timestamp 1688980957
transform 1 0 17940 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_219
timestamp 1688980957
transform 1 0 21252 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_249
timestamp 1688980957
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_302
timestamp 1688980957
transform 1 0 28888 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_331
timestamp 1688980957
transform 1 0 31556 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_337
timestamp 1688980957
transform 1 0 32108 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_358
timestamp 1688980957
transform 1 0 34040 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_365
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_389
timestamp 1688980957
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1688980957
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_70
timestamp 1688980957
transform 1 0 7544 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_83
timestamp 1688980957
transform 1 0 8740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_95
timestamp 1688980957
transform 1 0 9844 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_103
timestamp 1688980957
transform 1 0 10580 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1688980957
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_125
timestamp 1688980957
transform 1 0 12604 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_129
timestamp 1688980957
transform 1 0 12972 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_143
timestamp 1688980957
transform 1 0 14260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_155
timestamp 1688980957
transform 1 0 15364 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 1688980957
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_182
timestamp 1688980957
transform 1 0 17848 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_188
timestamp 1688980957
transform 1 0 18400 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_192
timestamp 1688980957
transform 1 0 18768 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 1688980957
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_238
timestamp 1688980957
transform 1 0 23000 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_244
timestamp 1688980957
transform 1 0 23552 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_254
timestamp 1688980957
transform 1 0 24472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_258
timestamp 1688980957
transform 1 0 24840 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_266
timestamp 1688980957
transform 1 0 25576 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_272
timestamp 1688980957
transform 1 0 26128 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_287
timestamp 1688980957
transform 1 0 27508 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_322
timestamp 1688980957
transform 1 0 30728 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_349
timestamp 1688980957
transform 1 0 33212 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_360
timestamp 1688980957
transform 1 0 34224 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_372
timestamp 1688980957
transform 1 0 35328 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_384
timestamp 1688980957
transform 1 0 36432 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_393
timestamp 1688980957
transform 1 0 37260 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_23
timestamp 1688980957
transform 1 0 3220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_76
timestamp 1688980957
transform 1 0 8096 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_91
timestamp 1688980957
transform 1 0 9476 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_98
timestamp 1688980957
transform 1 0 10120 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_106
timestamp 1688980957
transform 1 0 10856 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_124
timestamp 1688980957
transform 1 0 12512 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_132
timestamp 1688980957
transform 1 0 13248 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_149
timestamp 1688980957
transform 1 0 14812 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_168
timestamp 1688980957
transform 1 0 16560 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_180
timestamp 1688980957
transform 1 0 17664 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_192
timestamp 1688980957
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_223
timestamp 1688980957
transform 1 0 21620 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_235
timestamp 1688980957
transform 1 0 22724 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_247
timestamp 1688980957
transform 1 0 23828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1688980957
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_268
timestamp 1688980957
transform 1 0 25760 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_280
timestamp 1688980957
transform 1 0 26864 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_285
timestamp 1688980957
transform 1 0 27324 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_297
timestamp 1688980957
transform 1 0 28428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_305
timestamp 1688980957
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_320
timestamp 1688980957
transform 1 0 30544 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_334
timestamp 1688980957
transform 1 0 31832 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_342
timestamp 1688980957
transform 1 0 32568 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_352
timestamp 1688980957
transform 1 0 33488 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_363
timestamp 1688980957
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_368
timestamp 1688980957
transform 1 0 34960 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_380
timestamp 1688980957
transform 1 0 36064 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_395
timestamp 1688980957
transform 1 0 37444 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_12
timestamp 1688980957
transform 1 0 2208 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_41
timestamp 1688980957
transform 1 0 4876 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_53
timestamp 1688980957
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_60
timestamp 1688980957
transform 1 0 6624 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_72
timestamp 1688980957
transform 1 0 7728 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_80
timestamp 1688980957
transform 1 0 8464 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_88
timestamp 1688980957
transform 1 0 9200 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_105
timestamp 1688980957
transform 1 0 10764 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_135
timestamp 1688980957
transform 1 0 13524 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_152
timestamp 1688980957
transform 1 0 15088 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_178
timestamp 1688980957
transform 1 0 17480 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_188
timestamp 1688980957
transform 1 0 18400 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_196
timestamp 1688980957
transform 1 0 19136 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_220
timestamp 1688980957
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_231
timestamp 1688980957
transform 1 0 22356 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_245
timestamp 1688980957
transform 1 0 23644 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_249
timestamp 1688980957
transform 1 0 24012 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_255
timestamp 1688980957
transform 1 0 24564 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_263
timestamp 1688980957
transform 1 0 25300 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_293
timestamp 1688980957
transform 1 0 28060 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_297
timestamp 1688980957
transform 1 0 28428 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_303
timestamp 1688980957
transform 1 0 28980 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_315
timestamp 1688980957
transform 1 0 30084 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_327
timestamp 1688980957
transform 1 0 31188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_335
timestamp 1688980957
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_349
timestamp 1688980957
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_361
timestamp 1688980957
transform 1 0 34316 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_367
timestamp 1688980957
transform 1 0 34868 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_371
timestamp 1688980957
transform 1 0 35236 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_383
timestamp 1688980957
transform 1 0 36340 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_393
timestamp 1688980957
transform 1 0 37260 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_38
timestamp 1688980957
transform 1 0 4600 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_43
timestamp 1688980957
transform 1 0 5060 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_49
timestamp 1688980957
transform 1 0 5612 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_73
timestamp 1688980957
transform 1 0 7820 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_92
timestamp 1688980957
transform 1 0 9568 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_100
timestamp 1688980957
transform 1 0 10304 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_112
timestamp 1688980957
transform 1 0 11408 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_126
timestamp 1688980957
transform 1 0 12696 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_130
timestamp 1688980957
transform 1 0 13064 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_138
timestamp 1688980957
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_146
timestamp 1688980957
transform 1 0 14536 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_154
timestamp 1688980957
transform 1 0 15272 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_164
timestamp 1688980957
transform 1 0 16192 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_172
timestamp 1688980957
transform 1 0 16928 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_191
timestamp 1688980957
transform 1 0 18676 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_218
timestamp 1688980957
transform 1 0 21160 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_248
timestamp 1688980957
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_272
timestamp 1688980957
transform 1 0 26128 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_282
timestamp 1688980957
transform 1 0 27048 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_304
timestamp 1688980957
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_316
timestamp 1688980957
transform 1 0 30176 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_328
timestamp 1688980957
transform 1 0 31280 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_340
timestamp 1688980957
transform 1 0 32384 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 1688980957
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 1688980957
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_365
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_379
timestamp 1688980957
transform 1 0 35972 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_391
timestamp 1688980957
transform 1 0 37076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_399
timestamp 1688980957
transform 1 0 37812 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1688980957
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_67
timestamp 1688980957
transform 1 0 7268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_79
timestamp 1688980957
transform 1 0 8372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_85
timestamp 1688980957
transform 1 0 8924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_93
timestamp 1688980957
transform 1 0 9660 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_97
timestamp 1688980957
transform 1 0 10028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_109
timestamp 1688980957
transform 1 0 11132 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_122
timestamp 1688980957
transform 1 0 12328 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_134
timestamp 1688980957
transform 1 0 13432 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_138
timestamp 1688980957
transform 1 0 13800 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_147
timestamp 1688980957
transform 1 0 14628 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_162
timestamp 1688980957
transform 1 0 16008 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_172
timestamp 1688980957
transform 1 0 16928 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_181
timestamp 1688980957
transform 1 0 17756 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_191
timestamp 1688980957
transform 1 0 18676 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_199
timestamp 1688980957
transform 1 0 19412 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_206
timestamp 1688980957
transform 1 0 20056 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_210
timestamp 1688980957
transform 1 0 20424 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_218
timestamp 1688980957
transform 1 0 21160 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_271
timestamp 1688980957
transform 1 0 26036 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_277
timestamp 1688980957
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_286
timestamp 1688980957
transform 1 0 27416 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_294
timestamp 1688980957
transform 1 0 28152 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_300
timestamp 1688980957
transform 1 0 28704 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_345
timestamp 1688980957
transform 1 0 32844 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_353
timestamp 1688980957
transform 1 0 33580 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_357
timestamp 1688980957
transform 1 0 33948 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_382
timestamp 1688980957
transform 1 0 36248 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_389
timestamp 1688980957
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_400
timestamp 1688980957
transform 1 0 37904 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_23
timestamp 1688980957
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_32
timestamp 1688980957
transform 1 0 4048 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_36
timestamp 1688980957
transform 1 0 4416 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_48
timestamp 1688980957
transform 1 0 5520 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_60
timestamp 1688980957
transform 1 0 6624 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_76
timestamp 1688980957
transform 1 0 8096 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_97
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_101
timestamp 1688980957
transform 1 0 10396 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_130
timestamp 1688980957
transform 1 0 13064 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_138
timestamp 1688980957
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_145
timestamp 1688980957
transform 1 0 14444 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_155
timestamp 1688980957
transform 1 0 15364 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_164
timestamp 1688980957
transform 1 0 16192 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_192
timestamp 1688980957
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_209
timestamp 1688980957
transform 1 0 20332 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_221
timestamp 1688980957
transform 1 0 21436 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_229
timestamp 1688980957
transform 1 0 22172 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_238
timestamp 1688980957
transform 1 0 23000 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_250
timestamp 1688980957
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_261
timestamp 1688980957
transform 1 0 25116 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_273
timestamp 1688980957
transform 1 0 26220 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_281
timestamp 1688980957
transform 1 0 26956 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_287
timestamp 1688980957
transform 1 0 27508 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_295
timestamp 1688980957
transform 1 0 28244 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_306
timestamp 1688980957
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_320
timestamp 1688980957
transform 1 0 30544 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_328
timestamp 1688980957
transform 1 0 31280 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_339
timestamp 1688980957
transform 1 0 32292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_351
timestamp 1688980957
transform 1 0 33396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 1688980957
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_365
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_377
timestamp 1688980957
transform 1 0 35788 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_383
timestamp 1688980957
transform 1 0 36340 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_392
timestamp 1688980957
transform 1 0 37168 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_400
timestamp 1688980957
transform 1 0 37904 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_10
timestamp 1688980957
transform 1 0 2024 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_48
timestamp 1688980957
transform 1 0 5520 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_92
timestamp 1688980957
transform 1 0 9568 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_104
timestamp 1688980957
transform 1 0 10672 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_136
timestamp 1688980957
transform 1 0 13616 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_146
timestamp 1688980957
transform 1 0 14536 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_158
timestamp 1688980957
transform 1 0 15640 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_166
timestamp 1688980957
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_178
timestamp 1688980957
transform 1 0 17480 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_186
timestamp 1688980957
transform 1 0 18216 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_191
timestamp 1688980957
transform 1 0 18676 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_203
timestamp 1688980957
transform 1 0 19780 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_211
timestamp 1688980957
transform 1 0 20516 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_219
timestamp 1688980957
transform 1 0 21252 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1688980957
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_237
timestamp 1688980957
transform 1 0 22908 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_253
timestamp 1688980957
transform 1 0 24380 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_261
timestamp 1688980957
transform 1 0 25116 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_271
timestamp 1688980957
transform 1 0 26036 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1688980957
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 1688980957
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_305
timestamp 1688980957
transform 1 0 29164 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_312
timestamp 1688980957
transform 1 0 29808 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_327
timestamp 1688980957
transform 1 0 31188 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 1688980957
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_353
timestamp 1688980957
transform 1 0 33580 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_365
timestamp 1688980957
transform 1 0 34684 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_379
timestamp 1688980957
transform 1 0 35972 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_390
timestamp 1688980957
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_393
timestamp 1688980957
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_11
timestamp 1688980957
transform 1 0 2116 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_22
timestamp 1688980957
transform 1 0 3128 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_45
timestamp 1688980957
transform 1 0 5244 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_64
timestamp 1688980957
transform 1 0 6992 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_76
timestamp 1688980957
transform 1 0 8096 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_111
timestamp 1688980957
transform 1 0 11316 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_123
timestamp 1688980957
transform 1 0 12420 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_138
timestamp 1688980957
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_146
timestamp 1688980957
transform 1 0 14536 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_173
timestamp 1688980957
transform 1 0 17020 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_185
timestamp 1688980957
transform 1 0 18124 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_193
timestamp 1688980957
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_209
timestamp 1688980957
transform 1 0 20332 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_217
timestamp 1688980957
transform 1 0 21068 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_227
timestamp 1688980957
transform 1 0 21988 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_247
timestamp 1688980957
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1688980957
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_281
timestamp 1688980957
transform 1 0 26956 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_306
timestamp 1688980957
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_317
timestamp 1688980957
transform 1 0 30268 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_326
timestamp 1688980957
transform 1 0 31096 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_341
timestamp 1688980957
transform 1 0 32476 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_349
timestamp 1688980957
transform 1 0 33212 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_377
timestamp 1688980957
transform 1 0 35788 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_21
timestamp 1688980957
transform 1 0 3036 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_29
timestamp 1688980957
transform 1 0 3772 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_42
timestamp 1688980957
transform 1 0 4968 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_49
timestamp 1688980957
transform 1 0 5612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_70
timestamp 1688980957
transform 1 0 7544 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_74
timestamp 1688980957
transform 1 0 7912 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_98
timestamp 1688980957
transform 1 0 10120 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_110
timestamp 1688980957
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_122
timestamp 1688980957
transform 1 0 12328 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_134
timestamp 1688980957
transform 1 0 13432 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_153
timestamp 1688980957
transform 1 0 15180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_165
timestamp 1688980957
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_176
timestamp 1688980957
transform 1 0 17296 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_195
timestamp 1688980957
transform 1 0 19044 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_205
timestamp 1688980957
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_217
timestamp 1688980957
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1688980957
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_234
timestamp 1688980957
transform 1 0 22632 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_292
timestamp 1688980957
transform 1 0 27968 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_303
timestamp 1688980957
transform 1 0 28980 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_321
timestamp 1688980957
transform 1 0 30636 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_333
timestamp 1688980957
transform 1 0 31740 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_352
timestamp 1688980957
transform 1 0 33488 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_363
timestamp 1688980957
transform 1 0 34500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_375
timestamp 1688980957
transform 1 0 35604 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_381
timestamp 1688980957
transform 1 0 36156 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_389
timestamp 1688980957
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_393
timestamp 1688980957
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_23
timestamp 1688980957
transform 1 0 3220 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_43
timestamp 1688980957
transform 1 0 5060 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_55
timestamp 1688980957
transform 1 0 6164 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_68
timestamp 1688980957
transform 1 0 7360 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_94
timestamp 1688980957
transform 1 0 9752 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_138
timestamp 1688980957
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_148
timestamp 1688980957
transform 1 0 14720 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_156
timestamp 1688980957
transform 1 0 15456 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_165
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_173
timestamp 1688980957
transform 1 0 17020 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_193
timestamp 1688980957
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_201
timestamp 1688980957
transform 1 0 19596 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_216
timestamp 1688980957
transform 1 0 20976 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_228
timestamp 1688980957
transform 1 0 22080 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_240
timestamp 1688980957
transform 1 0 23184 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_259
timestamp 1688980957
transform 1 0 24932 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1688980957
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_277
timestamp 1688980957
transform 1 0 26588 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_283
timestamp 1688980957
transform 1 0 27140 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_287
timestamp 1688980957
transform 1 0 27508 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_299
timestamp 1688980957
transform 1 0 28612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 1688980957
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_309
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_317
timestamp 1688980957
transform 1 0 30268 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_326
timestamp 1688980957
transform 1 0 31096 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_332
timestamp 1688980957
transform 1 0 31648 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_336
timestamp 1688980957
transform 1 0 32016 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_344
timestamp 1688980957
transform 1 0 32752 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_355
timestamp 1688980957
transform 1 0 33764 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_363
timestamp 1688980957
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_377
timestamp 1688980957
transform 1 0 35788 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_381
timestamp 1688980957
transform 1 0 36156 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_394
timestamp 1688980957
transform 1 0 37352 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_400
timestamp 1688980957
transform 1 0 37904 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_9
timestamp 1688980957
transform 1 0 1932 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_21
timestamp 1688980957
transform 1 0 3036 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_67
timestamp 1688980957
transform 1 0 7268 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_79
timestamp 1688980957
transform 1 0 8372 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_91
timestamp 1688980957
transform 1 0 9476 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_103
timestamp 1688980957
transform 1 0 10580 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_153
timestamp 1688980957
transform 1 0 15180 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_157
timestamp 1688980957
transform 1 0 15548 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_166
timestamp 1688980957
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_193
timestamp 1688980957
transform 1 0 18860 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_208
timestamp 1688980957
transform 1 0 20240 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_220
timestamp 1688980957
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_237
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_251
timestamp 1688980957
transform 1 0 24196 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_263
timestamp 1688980957
transform 1 0 25300 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_271
timestamp 1688980957
transform 1 0 26036 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_275
timestamp 1688980957
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1688980957
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1688980957
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_305
timestamp 1688980957
transform 1 0 29164 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_316
timestamp 1688980957
transform 1 0 30176 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_335
timestamp 1688980957
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 1688980957
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_361
timestamp 1688980957
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_373
timestamp 1688980957
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_385
timestamp 1688980957
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 1688980957
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_393
timestamp 1688980957
transform 1 0 37260 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_23
timestamp 1688980957
transform 1 0 3220 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_43
timestamp 1688980957
transform 1 0 5060 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_71
timestamp 1688980957
transform 1 0 7636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_95
timestamp 1688980957
transform 1 0 9844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_107
timestamp 1688980957
transform 1 0 10948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 1688980957
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_147
timestamp 1688980957
transform 1 0 14628 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_159
timestamp 1688980957
transform 1 0 15732 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_166
timestamp 1688980957
transform 1 0 16376 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_190
timestamp 1688980957
transform 1 0 18584 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_209
timestamp 1688980957
transform 1 0 20332 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_217
timestamp 1688980957
transform 1 0 21068 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_225
timestamp 1688980957
transform 1 0 21804 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_235
timestamp 1688980957
transform 1 0 22724 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_243
timestamp 1688980957
transform 1 0 23460 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_268
timestamp 1688980957
transform 1 0 25760 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_273
timestamp 1688980957
transform 1 0 26220 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_280
timestamp 1688980957
transform 1 0 26864 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_291
timestamp 1688980957
transform 1 0 27876 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_305
timestamp 1688980957
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_314
timestamp 1688980957
transform 1 0 29992 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_326
timestamp 1688980957
transform 1 0 31096 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_347
timestamp 1688980957
transform 1 0 33028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_359
timestamp 1688980957
transform 1 0 34132 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_372
timestamp 1688980957
transform 1 0 35328 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_380
timestamp 1688980957
transform 1 0 36064 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_392
timestamp 1688980957
transform 1 0 37168 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_400
timestamp 1688980957
transform 1 0 37904 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_47
timestamp 1688980957
transform 1 0 5428 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_78
timestamp 1688980957
transform 1 0 8280 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_149
timestamp 1688980957
transform 1 0 14812 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_159
timestamp 1688980957
transform 1 0 15732 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_163
timestamp 1688980957
transform 1 0 16100 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1688980957
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 1688980957
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_193
timestamp 1688980957
transform 1 0 18860 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_204
timestamp 1688980957
transform 1 0 19872 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_210
timestamp 1688980957
transform 1 0 20424 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_218
timestamp 1688980957
transform 1 0 21160 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_240
timestamp 1688980957
transform 1 0 23184 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_248
timestamp 1688980957
transform 1 0 23920 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_273
timestamp 1688980957
transform 1 0 26220 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_281
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_297
timestamp 1688980957
transform 1 0 28428 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_305
timestamp 1688980957
transform 1 0 29164 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_324
timestamp 1688980957
transform 1 0 30912 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_334
timestamp 1688980957
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_345
timestamp 1688980957
transform 1 0 32844 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_350
timestamp 1688980957
transform 1 0 33304 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_384
timestamp 1688980957
transform 1 0 36432 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_390
timestamp 1688980957
transform 1 0 36984 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_393
timestamp 1688980957
transform 1 0 37260 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_37
timestamp 1688980957
transform 1 0 4508 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_44
timestamp 1688980957
transform 1 0 5152 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_56
timestamp 1688980957
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_64
timestamp 1688980957
transform 1 0 6992 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_71
timestamp 1688980957
transform 1 0 7636 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_77
timestamp 1688980957
transform 1 0 8188 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_81
timestamp 1688980957
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_94
timestamp 1688980957
transform 1 0 9752 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_106
timestamp 1688980957
transform 1 0 10856 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_157
timestamp 1688980957
transform 1 0 15548 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_164
timestamp 1688980957
transform 1 0 16192 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_176
timestamp 1688980957
transform 1 0 17296 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_188
timestamp 1688980957
transform 1 0 18400 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_211
timestamp 1688980957
transform 1 0 20516 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_223
timestamp 1688980957
transform 1 0 21620 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_239
timestamp 1688980957
transform 1 0 23092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 1688980957
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1688980957
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_277
timestamp 1688980957
transform 1 0 26588 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_283
timestamp 1688980957
transform 1 0 27140 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_287
timestamp 1688980957
transform 1 0 27508 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_299
timestamp 1688980957
transform 1 0 28612 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_333
timestamp 1688980957
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_345
timestamp 1688980957
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_357
timestamp 1688980957
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_363
timestamp 1688980957
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_368
timestamp 1688980957
transform 1 0 34960 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_380
timestamp 1688980957
transform 1 0 36064 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_400
timestamp 1688980957
transform 1 0 37904 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_10
timestamp 1688980957
transform 1 0 2024 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_22
timestamp 1688980957
transform 1 0 3128 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_34
timestamp 1688980957
transform 1 0 4232 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_44
timestamp 1688980957
transform 1 0 5152 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_60
timestamp 1688980957
transform 1 0 6624 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_72
timestamp 1688980957
transform 1 0 7728 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_95
timestamp 1688980957
transform 1 0 9844 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_107
timestamp 1688980957
transform 1 0 10948 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_120
timestamp 1688980957
transform 1 0 12144 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_140
timestamp 1688980957
transform 1 0 13984 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_152
timestamp 1688980957
transform 1 0 15088 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 1688980957
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_180
timestamp 1688980957
transform 1 0 17664 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_188
timestamp 1688980957
transform 1 0 18400 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_194
timestamp 1688980957
transform 1 0 18952 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_206
timestamp 1688980957
transform 1 0 20056 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_218
timestamp 1688980957
transform 1 0 21160 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_225
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_240
timestamp 1688980957
transform 1 0 23184 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_252
timestamp 1688980957
transform 1 0 24288 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_260
timestamp 1688980957
transform 1 0 25024 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_264
timestamp 1688980957
transform 1 0 25392 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_272
timestamp 1688980957
transform 1 0 26128 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_284
timestamp 1688980957
transform 1 0 27232 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_296
timestamp 1688980957
transform 1 0 28336 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_308
timestamp 1688980957
transform 1 0 29440 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_320
timestamp 1688980957
transform 1 0 30544 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_332
timestamp 1688980957
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_348
timestamp 1688980957
transform 1 0 33120 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_384
timestamp 1688980957
transform 1 0 36432 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_393
timestamp 1688980957
transform 1 0 37260 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_7
timestamp 1688980957
transform 1 0 1748 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_43
timestamp 1688980957
transform 1 0 5060 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_69
timestamp 1688980957
transform 1 0 7452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_81
timestamp 1688980957
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 1688980957
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 1688980957
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_121
timestamp 1688980957
transform 1 0 12236 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_132
timestamp 1688980957
transform 1 0 13248 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_168
timestamp 1688980957
transform 1 0 16560 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_172
timestamp 1688980957
transform 1 0 16928 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_207
timestamp 1688980957
transform 1 0 20148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_219
timestamp 1688980957
transform 1 0 21252 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_227
timestamp 1688980957
transform 1 0 21988 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_237
timestamp 1688980957
transform 1 0 22908 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_249
timestamp 1688980957
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_261
timestamp 1688980957
transform 1 0 25116 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_273
timestamp 1688980957
transform 1 0 26220 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_277
timestamp 1688980957
transform 1 0 26588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_293
timestamp 1688980957
transform 1 0 28060 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_305
timestamp 1688980957
transform 1 0 29164 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_315
timestamp 1688980957
transform 1 0 30084 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_321
timestamp 1688980957
transform 1 0 30636 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_325
timestamp 1688980957
transform 1 0 31004 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_334
timestamp 1688980957
transform 1 0 31832 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_340
timestamp 1688980957
transform 1 0 32384 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_350
timestamp 1688980957
transform 1 0 33304 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_362
timestamp 1688980957
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_365
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_369
timestamp 1688980957
transform 1 0 35052 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_391
timestamp 1688980957
transform 1 0 37076 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_399
timestamp 1688980957
transform 1 0 37812 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_7
timestamp 1688980957
transform 1 0 1748 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_11
timestamp 1688980957
transform 1 0 2116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_32
timestamp 1688980957
transform 1 0 4048 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_46
timestamp 1688980957
transform 1 0 5336 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_54
timestamp 1688980957
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_65
timestamp 1688980957
transform 1 0 7084 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_78
timestamp 1688980957
transform 1 0 8280 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_86
timestamp 1688980957
transform 1 0 9016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_107
timestamp 1688980957
transform 1 0 10948 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_121
timestamp 1688980957
transform 1 0 12236 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_135
timestamp 1688980957
transform 1 0 13524 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_147
timestamp 1688980957
transform 1 0 14628 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_159
timestamp 1688980957
transform 1 0 15732 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_164
timestamp 1688980957
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_177
timestamp 1688980957
transform 1 0 17388 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_190
timestamp 1688980957
transform 1 0 18584 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_202
timestamp 1688980957
transform 1 0 19688 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_210
timestamp 1688980957
transform 1 0 20424 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_232
timestamp 1688980957
transform 1 0 22448 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_244
timestamp 1688980957
transform 1 0 23552 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_260
timestamp 1688980957
transform 1 0 25024 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_275
timestamp 1688980957
transform 1 0 26404 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1688980957
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_301
timestamp 1688980957
transform 1 0 28796 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_318
timestamp 1688980957
transform 1 0 30360 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_326
timestamp 1688980957
transform 1 0 31096 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_331
timestamp 1688980957
transform 1 0 31556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 1688980957
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_342
timestamp 1688980957
transform 1 0 32568 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_353
timestamp 1688980957
transform 1 0 33580 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_366
timestamp 1688980957
transform 1 0 34776 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_373
timestamp 1688980957
transform 1 0 35420 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_384
timestamp 1688980957
transform 1 0 36432 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_393
timestamp 1688980957
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_23
timestamp 1688980957
transform 1 0 3220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_45
timestamp 1688980957
transform 1 0 5244 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_57
timestamp 1688980957
transform 1 0 6348 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_63
timestamp 1688980957
transform 1 0 6900 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_96
timestamp 1688980957
transform 1 0 9936 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_107
timestamp 1688980957
transform 1 0 10948 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_111
timestamp 1688980957
transform 1 0 11316 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_117
timestamp 1688980957
transform 1 0 11868 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_125
timestamp 1688980957
transform 1 0 12604 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_135
timestamp 1688980957
transform 1 0 13524 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1688980957
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_148
timestamp 1688980957
transform 1 0 14720 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_169
timestamp 1688980957
transform 1 0 16652 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_181
timestamp 1688980957
transform 1 0 17756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_193
timestamp 1688980957
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_205
timestamp 1688980957
transform 1 0 19964 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_222
timestamp 1688980957
transform 1 0 21528 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_234
timestamp 1688980957
transform 1 0 22632 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_242
timestamp 1688980957
transform 1 0 23368 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_247
timestamp 1688980957
transform 1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 1688980957
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_256
timestamp 1688980957
transform 1 0 24656 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_268
timestamp 1688980957
transform 1 0 25760 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_272
timestamp 1688980957
transform 1 0 26128 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_282
timestamp 1688980957
transform 1 0 27048 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_290
timestamp 1688980957
transform 1 0 27784 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_305
timestamp 1688980957
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_321
timestamp 1688980957
transform 1 0 30636 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_326
timestamp 1688980957
transform 1 0 31096 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_332
timestamp 1688980957
transform 1 0 31648 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_338
timestamp 1688980957
transform 1 0 32200 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_350
timestamp 1688980957
transform 1 0 33304 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_354
timestamp 1688980957
transform 1 0 33672 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_362
timestamp 1688980957
transform 1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_365
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_377
timestamp 1688980957
transform 1 0 35788 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_46
timestamp 1688980957
transform 1 0 5336 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_54
timestamp 1688980957
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_69
timestamp 1688980957
transform 1 0 7452 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_75
timestamp 1688980957
transform 1 0 8004 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_79
timestamp 1688980957
transform 1 0 8372 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_91
timestamp 1688980957
transform 1 0 9476 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_103
timestamp 1688980957
transform 1 0 10580 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1688980957
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 1688980957
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1688980957
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 1688980957
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_181
timestamp 1688980957
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_193
timestamp 1688980957
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_214
timestamp 1688980957
transform 1 0 20792 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_222
timestamp 1688980957
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_256
timestamp 1688980957
transform 1 0 24656 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_268
timestamp 1688980957
transform 1 0 25760 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_281
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_287
timestamp 1688980957
transform 1 0 27508 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_296
timestamp 1688980957
transform 1 0 28336 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_308
timestamp 1688980957
transform 1 0 29440 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_325
timestamp 1688980957
transform 1 0 31004 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_333
timestamp 1688980957
transform 1 0 31740 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_337
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_354
timestamp 1688980957
transform 1 0 33672 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_366
timestamp 1688980957
transform 1 0 34776 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_378
timestamp 1688980957
transform 1 0 35880 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_390
timestamp 1688980957
transform 1 0 36984 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_393
timestamp 1688980957
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_21
timestamp 1688980957
transform 1 0 3036 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_63
timestamp 1688980957
transform 1 0 6900 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_97
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_109
timestamp 1688980957
transform 1 0 11132 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_117
timestamp 1688980957
transform 1 0 11868 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_135
timestamp 1688980957
transform 1 0 13524 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1688980957
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_144
timestamp 1688980957
transform 1 0 14352 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_156
timestamp 1688980957
transform 1 0 15456 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_160
timestamp 1688980957
transform 1 0 15824 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_173
timestamp 1688980957
transform 1 0 17020 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_185
timestamp 1688980957
transform 1 0 18124 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_192
timestamp 1688980957
transform 1 0 18768 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_200
timestamp 1688980957
transform 1 0 19504 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_212
timestamp 1688980957
transform 1 0 20608 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_224
timestamp 1688980957
transform 1 0 21712 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_236
timestamp 1688980957
transform 1 0 22816 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_248
timestamp 1688980957
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_253
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_261
timestamp 1688980957
transform 1 0 25116 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_294
timestamp 1688980957
transform 1 0 28152 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1688980957
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_333
timestamp 1688980957
transform 1 0 31740 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_337
timestamp 1688980957
transform 1 0 32108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_342
timestamp 1688980957
transform 1 0 32568 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_354
timestamp 1688980957
transform 1 0 33672 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_362
timestamp 1688980957
transform 1 0 34408 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_370
timestamp 1688980957
transform 1 0 35144 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_383
timestamp 1688980957
transform 1 0 36340 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_395
timestamp 1688980957
transform 1 0 37444 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_33
timestamp 1688980957
transform 1 0 4140 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_42
timestamp 1688980957
transform 1 0 4968 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1688980957
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_121
timestamp 1688980957
transform 1 0 12236 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_129
timestamp 1688980957
transform 1 0 12972 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_133
timestamp 1688980957
transform 1 0 13340 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_176
timestamp 1688980957
transform 1 0 17296 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_182
timestamp 1688980957
transform 1 0 17848 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_206
timestamp 1688980957
transform 1 0 20056 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_218
timestamp 1688980957
transform 1 0 21160 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_232
timestamp 1688980957
transform 1 0 22448 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_244
timestamp 1688980957
transform 1 0 23552 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_253
timestamp 1688980957
transform 1 0 24380 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_267
timestamp 1688980957
transform 1 0 25668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1688980957
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_286
timestamp 1688980957
transform 1 0 27416 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_293
timestamp 1688980957
transform 1 0 28060 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_305
timestamp 1688980957
transform 1 0 29164 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_331
timestamp 1688980957
transform 1 0 31556 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1688980957
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_368
timestamp 1688980957
transform 1 0 34960 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_386
timestamp 1688980957
transform 1 0 36616 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_393
timestamp 1688980957
transform 1 0 37260 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_49
timestamp 1688980957
transform 1 0 5612 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1688980957
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1688980957
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 1688980957
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_109
timestamp 1688980957
transform 1 0 11132 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_113
timestamp 1688980957
transform 1 0 11500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_120
timestamp 1688980957
transform 1 0 12144 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_132
timestamp 1688980957
transform 1 0 13248 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_152
timestamp 1688980957
transform 1 0 15088 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_167
timestamp 1688980957
transform 1 0 16468 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_179
timestamp 1688980957
transform 1 0 17572 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_190
timestamp 1688980957
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 1688980957
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_227
timestamp 1688980957
transform 1 0 21988 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_238
timestamp 1688980957
transform 1 0 23000 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_243
timestamp 1688980957
transform 1 0 23460 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_261
timestamp 1688980957
transform 1 0 25116 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_270
timestamp 1688980957
transform 1 0 25944 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_282
timestamp 1688980957
transform 1 0 27048 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_288
timestamp 1688980957
transform 1 0 27600 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_293
timestamp 1688980957
transform 1 0 28060 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_305
timestamp 1688980957
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_321
timestamp 1688980957
transform 1 0 30636 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_341
timestamp 1688980957
transform 1 0 32476 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_353
timestamp 1688980957
transform 1 0 33580 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_362
timestamp 1688980957
transform 1 0 34408 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 1688980957
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_377
timestamp 1688980957
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_389
timestamp 1688980957
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 1688980957
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_91
timestamp 1688980957
transform 1 0 9476 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_103
timestamp 1688980957
transform 1 0 10580 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1688980957
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_129
timestamp 1688980957
transform 1 0 12972 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_141
timestamp 1688980957
transform 1 0 14076 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_153
timestamp 1688980957
transform 1 0 15180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_165
timestamp 1688980957
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_181
timestamp 1688980957
transform 1 0 17756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_188
timestamp 1688980957
transform 1 0 18400 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_197
timestamp 1688980957
transform 1 0 19228 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_208
timestamp 1688980957
transform 1 0 20240 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_215
timestamp 1688980957
transform 1 0 20884 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_241
timestamp 1688980957
transform 1 0 23276 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_262
timestamp 1688980957
transform 1 0 25208 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_274
timestamp 1688980957
transform 1 0 26312 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 1688980957
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_305
timestamp 1688980957
transform 1 0 29164 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_309
timestamp 1688980957
transform 1 0 29532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_315
timestamp 1688980957
transform 1 0 30084 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_327
timestamp 1688980957
transform 1 0 31188 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1688980957
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_342
timestamp 1688980957
transform 1 0 32568 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_370
timestamp 1688980957
transform 1 0 35144 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_382
timestamp 1688980957
transform 1 0 36248 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_390
timestamp 1688980957
transform 1 0 36984 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_393
timestamp 1688980957
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1688980957
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_35
timestamp 1688980957
transform 1 0 4324 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_48
timestamp 1688980957
transform 1 0 5520 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_60
timestamp 1688980957
transform 1 0 6624 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_93
timestamp 1688980957
transform 1 0 9660 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_110
timestamp 1688980957
transform 1 0 11224 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_114
timestamp 1688980957
transform 1 0 11592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_118
timestamp 1688980957
transform 1 0 11960 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_126
timestamp 1688980957
transform 1 0 12696 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_130
timestamp 1688980957
transform 1 0 13064 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_138
timestamp 1688980957
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_153
timestamp 1688980957
transform 1 0 15180 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_171
timestamp 1688980957
transform 1 0 16836 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_215
timestamp 1688980957
transform 1 0 20884 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_221
timestamp 1688980957
transform 1 0 21436 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_232
timestamp 1688980957
transform 1 0 22448 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_244
timestamp 1688980957
transform 1 0 23552 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_268
timestamp 1688980957
transform 1 0 25760 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_280
timestamp 1688980957
transform 1 0 26864 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_286
timestamp 1688980957
transform 1 0 27416 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_294
timestamp 1688980957
transform 1 0 28152 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_302
timestamp 1688980957
transform 1 0 28888 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_321
timestamp 1688980957
transform 1 0 30636 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_327
timestamp 1688980957
transform 1 0 31188 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_343
timestamp 1688980957
transform 1 0 32660 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_354
timestamp 1688980957
transform 1 0 33672 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_358
timestamp 1688980957
transform 1 0 34040 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 1688980957
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_372
timestamp 1688980957
transform 1 0 35328 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_384
timestamp 1688980957
transform 1 0 36432 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_396
timestamp 1688980957
transform 1 0 37536 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_31
timestamp 1688980957
transform 1 0 3956 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_84
timestamp 1688980957
transform 1 0 8832 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_108
timestamp 1688980957
transform 1 0 11040 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_121
timestamp 1688980957
transform 1 0 12236 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_166
timestamp 1688980957
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_175
timestamp 1688980957
transform 1 0 17204 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_195
timestamp 1688980957
transform 1 0 19044 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_206
timestamp 1688980957
transform 1 0 20056 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_218
timestamp 1688980957
transform 1 0 21160 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 1688980957
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 1688980957
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_261
timestamp 1688980957
transform 1 0 25116 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_273
timestamp 1688980957
transform 1 0 26220 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 1688980957
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_307
timestamp 1688980957
transform 1 0 29348 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_318
timestamp 1688980957
transform 1 0 30360 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_324
timestamp 1688980957
transform 1 0 30912 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_347
timestamp 1688980957
transform 1 0 33028 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_359
timestamp 1688980957
transform 1 0 34132 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_371
timestamp 1688980957
transform 1 0 35236 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_383
timestamp 1688980957
transform 1 0 36340 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_391
timestamp 1688980957
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_393
timestamp 1688980957
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1688980957
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1688980957
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1688980957
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1688980957
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1688980957
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 1688980957
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1688980957
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_149
timestamp 1688980957
transform 1 0 14812 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_160
timestamp 1688980957
transform 1 0 15824 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_172
timestamp 1688980957
transform 1 0 16928 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_180
timestamp 1688980957
transform 1 0 17664 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_184
timestamp 1688980957
transform 1 0 18032 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_209
timestamp 1688980957
transform 1 0 20332 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_233
timestamp 1688980957
transform 1 0 22540 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_242
timestamp 1688980957
transform 1 0 23368 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_249
timestamp 1688980957
transform 1 0 24012 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_259
timestamp 1688980957
transform 1 0 24932 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_265
timestamp 1688980957
transform 1 0 25484 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_273
timestamp 1688980957
transform 1 0 26220 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_288
timestamp 1688980957
transform 1 0 27600 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_300
timestamp 1688980957
transform 1 0 28704 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 1688980957
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 1688980957
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_345
timestamp 1688980957
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 1688980957
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 1688980957
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 1688980957
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_389
timestamp 1688980957
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1688980957
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1688980957
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1688980957
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_105
timestamp 1688980957
transform 1 0 10764 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_132
timestamp 1688980957
transform 1 0 13248 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_144
timestamp 1688980957
transform 1 0 14352 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_156
timestamp 1688980957
transform 1 0 15456 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_162
timestamp 1688980957
transform 1 0 16008 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_166
timestamp 1688980957
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 1688980957
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_193
timestamp 1688980957
transform 1 0 18860 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_201
timestamp 1688980957
transform 1 0 19596 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_207
timestamp 1688980957
transform 1 0 20148 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_219
timestamp 1688980957
transform 1 0 21252 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 1688980957
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_234
timestamp 1688980957
transform 1 0 22632 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_240
timestamp 1688980957
transform 1 0 23184 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 1688980957
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 1688980957
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1688980957
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 1688980957
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_316
timestamp 1688980957
transform 1 0 30176 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_328
timestamp 1688980957
transform 1 0 31280 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1688980957
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_361
timestamp 1688980957
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_373
timestamp 1688980957
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_385
timestamp 1688980957
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 1688980957
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_393
timestamp 1688980957
transform 1 0 37260 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_7
timestamp 1688980957
transform 1 0 1748 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_19
timestamp 1688980957
transform 1 0 2852 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1688980957
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_88
timestamp 1688980957
transform 1 0 9200 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_99
timestamp 1688980957
transform 1 0 10212 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_150
timestamp 1688980957
transform 1 0 14904 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_154
timestamp 1688980957
transform 1 0 15272 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_174
timestamp 1688980957
transform 1 0 17112 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_182
timestamp 1688980957
transform 1 0 17848 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_186
timestamp 1688980957
transform 1 0 18216 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_192
timestamp 1688980957
transform 1 0 18768 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_214
timestamp 1688980957
transform 1 0 20792 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_219
timestamp 1688980957
transform 1 0 21252 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_238
timestamp 1688980957
transform 1 0 23000 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_250
timestamp 1688980957
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_271
timestamp 1688980957
transform 1 0 26036 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_283
timestamp 1688980957
transform 1 0 27140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_295
timestamp 1688980957
transform 1 0 28244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1688980957
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1688980957
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1688980957
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1688980957
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 1688980957
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 1688980957
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 1688980957
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_389
timestamp 1688980957
transform 1 0 36892 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_393
timestamp 1688980957
transform 1 0 37260 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_397
timestamp 1688980957
transform 1 0 37628 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_100
timestamp 1688980957
transform 1 0 10304 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_129
timestamp 1688980957
transform 1 0 12972 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_133
timestamp 1688980957
transform 1 0 13340 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_141
timestamp 1688980957
transform 1 0 14076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_162
timestamp 1688980957
transform 1 0 16008 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_181
timestamp 1688980957
transform 1 0 17756 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_194
timestamp 1688980957
transform 1 0 18952 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_203
timestamp 1688980957
transform 1 0 19780 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_215
timestamp 1688980957
transform 1 0 20884 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_225
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_231
timestamp 1688980957
transform 1 0 22356 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 1688980957
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_249
timestamp 1688980957
transform 1 0 24012 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_257
timestamp 1688980957
transform 1 0 24748 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_271
timestamp 1688980957
transform 1 0 26036 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1688980957
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1688980957
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 1688980957
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 1688980957
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 1688980957
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 1688980957
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1688980957
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_361
timestamp 1688980957
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_373
timestamp 1688980957
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_385
timestamp 1688980957
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 1688980957
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_393
timestamp 1688980957
transform 1 0 37260 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1688980957
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1688980957
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 1688980957
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1688980957
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_111
timestamp 1688980957
transform 1 0 11316 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_123
timestamp 1688980957
transform 1 0 12420 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_159
timestamp 1688980957
transform 1 0 15732 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_179
timestamp 1688980957
transform 1 0 17572 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_187
timestamp 1688980957
transform 1 0 18308 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_192
timestamp 1688980957
transform 1 0 18768 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_206
timestamp 1688980957
transform 1 0 20056 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_225
timestamp 1688980957
transform 1 0 21804 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_233
timestamp 1688980957
transform 1 0 22540 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_240
timestamp 1688980957
transform 1 0 23184 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_257
timestamp 1688980957
transform 1 0 24748 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_271
timestamp 1688980957
transform 1 0 26036 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_283
timestamp 1688980957
transform 1 0 27140 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_291
timestamp 1688980957
transform 1 0 27876 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_298
timestamp 1688980957
transform 1 0 28520 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_304
timestamp 1688980957
transform 1 0 29072 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1688980957
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_345
timestamp 1688980957
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_357
timestamp 1688980957
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 1688980957
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1688980957
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1688980957
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 1688980957
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1688980957
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1688980957
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1688980957
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1688980957
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1688980957
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 1688980957
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_93
timestamp 1688980957
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 1688980957
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 1688980957
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_117
timestamp 1688980957
transform 1 0 11868 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_148
timestamp 1688980957
transform 1 0 14720 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_160
timestamp 1688980957
transform 1 0 15824 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_181
timestamp 1688980957
transform 1 0 17756 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_206
timestamp 1688980957
transform 1 0 20056 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_212
timestamp 1688980957
transform 1 0 20608 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_222
timestamp 1688980957
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_232
timestamp 1688980957
transform 1 0 22448 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_240
timestamp 1688980957
transform 1 0 23184 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_250
timestamp 1688980957
transform 1 0 24104 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_258
timestamp 1688980957
transform 1 0 24840 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_264
timestamp 1688980957
transform 1 0 25392 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_276
timestamp 1688980957
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 1688980957
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 1688980957
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 1688980957
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 1688980957
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 1688980957
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 1688980957
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 1688980957
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_349
timestamp 1688980957
transform 1 0 33212 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_354
timestamp 1688980957
transform 1 0 33672 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_366
timestamp 1688980957
transform 1 0 34776 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_378
timestamp 1688980957
transform 1 0 35880 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_390
timestamp 1688980957
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_393
timestamp 1688980957
transform 1 0 37260 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_397
timestamp 1688980957
transform 1 0 37628 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1688980957
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 1688980957
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_77
timestamp 1688980957
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 1688980957
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1688980957
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_109
timestamp 1688980957
transform 1 0 11132 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_113
timestamp 1688980957
transform 1 0 11500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_124
timestamp 1688980957
transform 1 0 12512 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_129
timestamp 1688980957
transform 1 0 12972 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_137
timestamp 1688980957
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_153
timestamp 1688980957
transform 1 0 15180 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_161
timestamp 1688980957
transform 1 0 15916 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_167
timestamp 1688980957
transform 1 0 16468 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_179
timestamp 1688980957
transform 1 0 17572 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_191
timestamp 1688980957
transform 1 0 18676 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_195
timestamp 1688980957
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_197
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_218
timestamp 1688980957
transform 1 0 21160 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_230
timestamp 1688980957
transform 1 0 22264 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_242
timestamp 1688980957
transform 1 0 23368 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_250
timestamp 1688980957
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_253
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_259
timestamp 1688980957
transform 1 0 24932 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_270
timestamp 1688980957
transform 1 0 25944 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_282
timestamp 1688980957
transform 1 0 27048 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_294
timestamp 1688980957
transform 1 0 28152 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_306
timestamp 1688980957
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 1688980957
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 1688980957
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_333
timestamp 1688980957
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_345
timestamp 1688980957
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_357
timestamp 1688980957
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 1688980957
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1688980957
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1688980957
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_389
timestamp 1688980957
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_9
timestamp 1688980957
transform 1 0 1932 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_21
timestamp 1688980957
transform 1 0 3036 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_33
timestamp 1688980957
transform 1 0 4140 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_45
timestamp 1688980957
transform 1 0 5244 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_53
timestamp 1688980957
transform 1 0 5980 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_69
timestamp 1688980957
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_81
timestamp 1688980957
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_93
timestamp 1688980957
transform 1 0 9660 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_102
timestamp 1688980957
transform 1 0 10488 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_110
timestamp 1688980957
transform 1 0 11224 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_113
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_125
timestamp 1688980957
transform 1 0 12604 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_132
timestamp 1688980957
transform 1 0 13248 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_144
timestamp 1688980957
transform 1 0 14352 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_156
timestamp 1688980957
transform 1 0 15456 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_178
timestamp 1688980957
transform 1 0 17480 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_188
timestamp 1688980957
transform 1 0 18400 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_200
timestamp 1688980957
transform 1 0 19504 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_218
timestamp 1688980957
transform 1 0 21160 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_225
timestamp 1688980957
transform 1 0 21804 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_229
timestamp 1688980957
transform 1 0 22172 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_242
timestamp 1688980957
transform 1 0 23368 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_250
timestamp 1688980957
transform 1 0 24104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_278
timestamp 1688980957
transform 1 0 26680 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_281
timestamp 1688980957
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_293
timestamp 1688980957
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_305
timestamp 1688980957
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_317
timestamp 1688980957
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_329
timestamp 1688980957
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_335
timestamp 1688980957
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_337
timestamp 1688980957
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_349
timestamp 1688980957
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_361
timestamp 1688980957
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_373
timestamp 1688980957
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_385
timestamp 1688980957
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_391
timestamp 1688980957
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_393
timestamp 1688980957
transform 1 0 37260 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_10
timestamp 1688980957
transform 1 0 2024 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_22
timestamp 1688980957
transform 1 0 3128 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_41
timestamp 1688980957
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_53
timestamp 1688980957
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_65
timestamp 1688980957
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_77
timestamp 1688980957
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_83
timestamp 1688980957
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_97
timestamp 1688980957
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_109
timestamp 1688980957
transform 1 0 11132 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_115
timestamp 1688980957
transform 1 0 11684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_127
timestamp 1688980957
transform 1 0 12788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_139
timestamp 1688980957
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_149
timestamp 1688980957
transform 1 0 14812 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_171
timestamp 1688980957
transform 1 0 16836 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_175
timestamp 1688980957
transform 1 0 17204 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_197
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_201
timestamp 1688980957
transform 1 0 19596 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_222
timestamp 1688980957
transform 1 0 21528 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_245
timestamp 1688980957
transform 1 0 23644 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_273
timestamp 1688980957
transform 1 0 26220 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_285
timestamp 1688980957
transform 1 0 27324 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_297
timestamp 1688980957
transform 1 0 28428 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_305
timestamp 1688980957
transform 1 0 29164 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_309
timestamp 1688980957
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_321
timestamp 1688980957
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_333
timestamp 1688980957
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_345
timestamp 1688980957
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_357
timestamp 1688980957
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_363
timestamp 1688980957
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_365
timestamp 1688980957
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_377
timestamp 1688980957
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_389
timestamp 1688980957
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_15
timestamp 1688980957
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_27
timestamp 1688980957
transform 1 0 3588 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_29
timestamp 1688980957
transform 1 0 3772 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_41
timestamp 1688980957
transform 1 0 4876 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_51
timestamp 1688980957
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 1688980957
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 1688980957
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_81
timestamp 1688980957
transform 1 0 8556 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_85
timestamp 1688980957
transform 1 0 8924 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_93
timestamp 1688980957
transform 1 0 9660 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_100
timestamp 1688980957
transform 1 0 10304 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_113
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_125
timestamp 1688980957
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_137
timestamp 1688980957
transform 1 0 13708 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_141
timestamp 1688980957
transform 1 0 14076 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_149
timestamp 1688980957
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_161
timestamp 1688980957
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_167
timestamp 1688980957
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_169
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_177
timestamp 1688980957
transform 1 0 17388 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_182
timestamp 1688980957
transform 1 0 17848 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_194
timestamp 1688980957
transform 1 0 18952 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_197
timestamp 1688980957
transform 1 0 19228 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_209
timestamp 1688980957
transform 1 0 20332 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_217
timestamp 1688980957
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_223
timestamp 1688980957
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_225
timestamp 1688980957
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_237
timestamp 1688980957
transform 1 0 22908 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_247
timestamp 1688980957
transform 1 0 23828 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_251
timestamp 1688980957
transform 1 0 24196 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_253
timestamp 1688980957
transform 1 0 24380 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_261
timestamp 1688980957
transform 1 0 25116 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_266
timestamp 1688980957
transform 1 0 25576 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_278
timestamp 1688980957
transform 1 0 26680 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_281
timestamp 1688980957
transform 1 0 26956 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_289
timestamp 1688980957
transform 1 0 27692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_301
timestamp 1688980957
transform 1 0 28796 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_307
timestamp 1688980957
transform 1 0 29348 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_309
timestamp 1688980957
transform 1 0 29532 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_321
timestamp 1688980957
transform 1 0 30636 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_333
timestamp 1688980957
transform 1 0 31740 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_343
timestamp 1688980957
transform 1 0 32660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_355
timestamp 1688980957
transform 1 0 33764 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_363
timestamp 1688980957
transform 1 0 34500 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_371
timestamp 1688980957
transform 1 0 35236 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_379
timestamp 1688980957
transform 1 0 35972 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_385
timestamp 1688980957
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_391
timestamp 1688980957
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_393
timestamp 1688980957
transform 1 0 37260 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 4232 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 3404 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 4508 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 4508 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 3588 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 30452 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform -1 0 31556 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform -1 0 31464 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform -1 0 5796 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform -1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform -1 0 21252 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 1688980957
transform 1 0 31004 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1688980957
transform 1 0 37444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12972 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1688980957
transform -1 0 37996 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1688980957
transform 1 0 35512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1688980957
transform -1 0 21068 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1688980957
transform -1 0 37996 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1688980957
transform -1 0 37996 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap1
timestamp 1688980957
transform -1 0 21988 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  max_cap47
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  max_cap48
timestamp 1688980957
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  max_cap49
timestamp 1688980957
transform 1 0 20424 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  max_cap50
timestamp 1688980957
transform -1 0 20884 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap51
timestamp 1688980957
transform 1 0 21344 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  max_cap52
timestamp 1688980957
transform -1 0 18768 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  max_cap53
timestamp 1688980957
transform -1 0 18860 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  max_cap54
timestamp 1688980957
transform 1 0 16008 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  max_cap55
timestamp 1688980957
transform 1 0 15824 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  max_cap57
timestamp 1688980957
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1688980957
transform 1 0 37628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 1688980957
transform 1 0 24564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1688980957
transform 1 0 37628 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1688980957
transform 1 0 25208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1688980957
transform 1 0 27140 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1688980957
transform -1 0 1932 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1688980957
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 1688980957
transform -1 0 1932 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1688980957
transform 1 0 23276 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1688980957
transform 1 0 32108 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1688980957
transform 1 0 37628 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1688980957
transform -1 0 14812 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1688980957
transform -1 0 4508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1688980957
transform -1 0 2576 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1688980957
transform 1 0 1932 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1688980957
transform 1 0 36156 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1688980957
transform -1 0 16100 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1688980957
transform 1 0 37628 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1688980957
transform 1 0 37444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1688980957
transform -1 0 1932 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output33
timestamp 1688980957
transform -1 0 1932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 1688980957
transform -1 0 7084 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1688980957
transform -1 0 1932 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1688980957
transform 1 0 37628 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1688980957
transform 1 0 20056 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform -1 0 1932 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1688980957
transform 1 0 34684 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1688980957
transform -1 0 5796 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output42
timestamp 1688980957
transform -1 0 10304 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output43
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output44
timestamp 1688980957
transform -1 0 1932 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output45
timestamp 1688980957
transform -1 0 1932 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 38272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 38272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 38272 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 38272 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 38272 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 38272 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 38272 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 38272 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 38272 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 38272 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 38272 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 38272 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 38272 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 38272 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 38272 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 38272 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 38272 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 38272 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 38272 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 38272 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 38272 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 38272 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 38272 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 38272 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 38272 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 38272 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 38272 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 38272 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 38272 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 38272 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 38272 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 38272 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 38272 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 38272 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 38272 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 38272 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 38272 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 38272 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 38272 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 38272 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 38272 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 38272 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 38272 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 38272 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 38272 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 38272 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 38272 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 38272 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 38272 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 38272 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 38272 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 38272 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 38272 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 38272 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 38272 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 38272 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 38272 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 38272 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 38272 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 38272 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 38272 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 38272 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 38272 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 38272 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 38272 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 38272 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 38272 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 38272 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1688980957
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1688980957
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1688980957
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1688980957
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1688980957
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1688980957
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1688980957
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1688980957
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1688980957
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1688980957
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1688980957
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1688980957
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1688980957
transform 1 0 3680 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1688980957
transform 1 0 8832 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1688980957
transform 1 0 13984 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1688980957
transform 1 0 19136 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1688980957
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1688980957
transform 1 0 24288 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1688980957
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1688980957
transform 1 0 29440 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1688980957
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1688980957
transform 1 0 34592 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1688980957
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  wire46
timestamp 1688980957
transform -1 0 12788 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  wire56
timestamp 1688980957
transform 1 0 14812 0 -1 16320
box -38 -48 590 592
<< labels >>
flabel metal4 s 4868 2128 5188 39216 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 39216 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 6006 38320 6326 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 36642 38320 36962 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 39216 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 34928 2128 35248 39216 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 5346 38320 5666 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 35982 38320 36302 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 2594 40765 2650 41565 0 FreeSans 224 90 0 0 clk
port 2 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 cs
port 3 nsew signal input
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 gpi[0]
port 4 nsew signal input
flabel metal3 s 0 32648 800 32768 0 FreeSans 480 0 0 0 gpi[10]
port 5 nsew signal input
flabel metal3 s 38621 23808 39421 23928 0 FreeSans 480 0 0 0 gpi[11]
port 6 nsew signal input
flabel metal2 s 16118 40765 16174 41565 0 FreeSans 224 90 0 0 gpi[12]
port 7 nsew signal input
flabel metal2 s 38658 40765 38714 41565 0 FreeSans 224 90 0 0 gpi[13]
port 8 nsew signal input
flabel metal3 s 38621 27888 39421 28008 0 FreeSans 480 0 0 0 gpi[14]
port 9 nsew signal input
flabel metal3 s 38621 6808 39421 6928 0 FreeSans 480 0 0 0 gpi[15]
port 10 nsew signal input
flabel metal3 s 38621 25848 39421 25968 0 FreeSans 480 0 0 0 gpi[16]
port 11 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 gpi[17]
port 12 nsew signal input
flabel metal3 s 38621 9528 39421 9648 0 FreeSans 480 0 0 0 gpi[18]
port 13 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 gpi[19]
port 14 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 gpi[1]
port 15 nsew signal input
flabel metal3 s 38621 4768 39421 4888 0 FreeSans 480 0 0 0 gpi[20]
port 16 nsew signal input
flabel metal2 s 11610 40765 11666 41565 0 FreeSans 224 90 0 0 gpi[21]
port 17 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 gpi[22]
port 18 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 gpi[23]
port 19 nsew signal input
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 gpi[24]
port 20 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 gpi[25]
port 21 nsew signal input
flabel metal3 s 38621 30608 39421 30728 0 FreeSans 480 0 0 0 gpi[26]
port 22 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 gpi[27]
port 23 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 gpi[28]
port 24 nsew signal input
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 gpi[29]
port 25 nsew signal input
flabel metal3 s 38621 32648 39421 32768 0 FreeSans 480 0 0 0 gpi[2]
port 26 nsew signal input
flabel metal3 s 38621 16328 39421 16448 0 FreeSans 480 0 0 0 gpi[30]
port 27 nsew signal input
flabel metal2 s 29642 40765 29698 41565 0 FreeSans 224 90 0 0 gpi[31]
port 28 nsew signal input
flabel metal2 s 7102 40765 7158 41565 0 FreeSans 224 90 0 0 gpi[32]
port 29 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 gpi[33]
port 30 nsew signal input
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 gpi[3]
port 31 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 gpi[4]
port 32 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 gpi[5]
port 33 nsew signal input
flabel metal2 s 20626 40765 20682 41565 0 FreeSans 224 90 0 0 gpi[6]
port 34 nsew signal input
flabel metal3 s 38621 40128 39421 40248 0 FreeSans 480 0 0 0 gpi[7]
port 35 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 gpi[8]
port 36 nsew signal input
flabel metal2 s 18694 40765 18750 41565 0 FreeSans 224 90 0 0 gpi[9]
port 37 nsew signal input
flabel metal3 s 38621 2048 39421 2168 0 FreeSans 480 0 0 0 gpo[0]
port 38 nsew signal tristate
flabel metal3 s 38621 11568 39421 11688 0 FreeSans 480 0 0 0 gpo[10]
port 39 nsew signal tristate
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 gpo[11]
port 40 nsew signal tristate
flabel metal3 s 38621 14288 39421 14408 0 FreeSans 480 0 0 0 gpo[12]
port 41 nsew signal tristate
flabel metal2 s 25134 40765 25190 41565 0 FreeSans 224 90 0 0 gpo[13]
port 42 nsew signal tristate
flabel metal2 s 27066 40765 27122 41565 0 FreeSans 224 90 0 0 gpo[14]
port 43 nsew signal tristate
flabel metal2 s 662 40765 718 41565 0 FreeSans 224 90 0 0 gpo[15]
port 44 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 gpo[16]
port 45 nsew signal tristate
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 gpo[17]
port 46 nsew signal tristate
flabel metal2 s 23202 40765 23258 41565 0 FreeSans 224 90 0 0 gpo[18]
port 47 nsew signal tristate
flabel metal2 s 31574 40765 31630 41565 0 FreeSans 224 90 0 0 gpo[19]
port 48 nsew signal tristate
flabel metal3 s 38621 37408 39421 37528 0 FreeSans 480 0 0 0 gpo[1]
port 49 nsew signal tristate
flabel metal2 s 14186 40765 14242 41565 0 FreeSans 224 90 0 0 gpo[20]
port 50 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 gpo[21]
port 51 nsew signal tristate
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 gpo[22]
port 52 nsew signal tristate
flabel metal3 s 0 39448 800 39568 0 FreeSans 480 0 0 0 gpo[23]
port 53 nsew signal tristate
flabel metal2 s 36082 40765 36138 41565 0 FreeSans 224 90 0 0 gpo[24]
port 54 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 gpo[25]
port 55 nsew signal tristate
flabel metal3 s 38621 35368 39421 35488 0 FreeSans 480 0 0 0 gpo[26]
port 56 nsew signal tristate
flabel metal3 s 38621 8 39421 128 0 FreeSans 480 0 0 0 gpo[27]
port 57 nsew signal tristate
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 gpo[28]
port 58 nsew signal tristate
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 gpo[29]
port 59 nsew signal tristate
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 gpo[2]
port 60 nsew signal tristate
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 gpo[30]
port 61 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 gpo[31]
port 62 nsew signal tristate
flabel metal3 s 38621 21088 39421 21208 0 FreeSans 480 0 0 0 gpo[32]
port 63 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 gpo[33]
port 64 nsew signal tristate
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 gpo[3]
port 65 nsew signal tristate
flabel metal2 s 34150 40765 34206 41565 0 FreeSans 224 90 0 0 gpo[4]
port 66 nsew signal tristate
flabel metal2 s 5170 40765 5226 41565 0 FreeSans 224 90 0 0 gpo[5]
port 67 nsew signal tristate
flabel metal2 s 9678 40765 9734 41565 0 FreeSans 224 90 0 0 gpo[6]
port 68 nsew signal tristate
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 gpo[7]
port 69 nsew signal tristate
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 gpo[8]
port 70 nsew signal tristate
flabel metal3 s 0 37408 800 37528 0 FreeSans 480 0 0 0 gpo[9]
port 71 nsew signal tristate
flabel metal3 s 38621 19048 39421 19168 0 FreeSans 480 0 0 0 nrst
port 72 nsew signal input
rlabel metal1 19688 39168 19688 39168 0 VGND
rlabel metal1 19688 38624 19688 38624 0 VPWR
rlabel metal2 27278 19924 27278 19924 0 ALU.flags_to_alu\[0\]
rlabel metal1 30636 17714 30636 17714 0 ALU.flags_to_alu\[1\]
rlabel metal1 18814 19414 18814 19414 0 ALU.flags_to_alu\[2\]
rlabel metal1 18078 7480 18078 7480 0 ALU.flags_to_alu\[3\]
rlabel metal2 25990 10302 25990 10302 0 ALU.flags_to_alu\[4\]
rlabel metal1 26266 13294 26266 13294 0 ALU.flags_to_alu\[5\]
rlabel metal1 20562 16116 20562 16116 0 ALU.flags_to_alu\[6\]
rlabel metal1 23782 19686 23782 19686 0 ALU.flags_to_alu\[7\]
rlabel via2 19458 21539 19458 21539 0 ALU.immediate\[0\]
rlabel metal1 7636 31314 7636 31314 0 ALU.immediate\[10\]
rlabel metal1 5520 32810 5520 32810 0 ALU.immediate\[11\]
rlabel metal1 8694 32334 8694 32334 0 ALU.immediate\[12\]
rlabel metal1 12650 31280 12650 31280 0 ALU.immediate\[13\]
rlabel metal2 8786 29342 8786 29342 0 ALU.immediate\[14\]
rlabel metal1 19550 27472 19550 27472 0 ALU.immediate\[15\]
rlabel metal2 32430 19601 32430 19601 0 ALU.immediate\[1\]
rlabel metal1 18906 19890 18906 19890 0 ALU.immediate\[2\]
rlabel metal2 3174 20825 3174 20825 0 ALU.immediate\[3\]
rlabel metal1 29854 19856 29854 19856 0 ALU.immediate\[4\]
rlabel metal1 9476 26418 9476 26418 0 ALU.immediate\[5\]
rlabel metal2 19688 20570 19688 20570 0 ALU.immediate\[6\]
rlabel metal1 22540 24922 22540 24922 0 ALU.immediate\[7\]
rlabel metal1 17066 35020 17066 35020 0 ALU.immediate\[8\]
rlabel metal1 7728 32742 7728 32742 0 ALU.immediate\[9\]
rlabel metal1 3772 26418 3772 26418 0 ByteBuffer.counter\[0\]
rlabel metal1 4922 26962 4922 26962 0 ByteBuffer.counter\[1\]
rlabel metal1 6118 17170 6118 17170 0 ByteBuffer.instr\[16\]
rlabel metal1 8326 18870 8326 18870 0 ByteBuffer.instr\[17\]
rlabel metal1 3910 16490 3910 16490 0 ByteBuffer.instr\[18\]
rlabel metal1 18354 21590 18354 21590 0 ByteBuffer.instr\[19\]
rlabel metal1 8418 21964 8418 21964 0 ByteBuffer.instr\[20\]
rlabel metal1 21896 23154 21896 23154 0 ByteBuffer.instr\[21\]
rlabel metal1 14536 23086 14536 23086 0 ByteBuffer.instr\[22\]
rlabel metal2 11546 23868 11546 23868 0 ByteBuffer.instr\[23\]
rlabel metal1 2231 26418 2231 26418 0 ByteBuffer.next_counter\[0\]
rlabel metal2 3450 26452 3450 26452 0 ByteBuffer.next_counter\[1\]
rlabel metal1 3404 29750 3404 29750 0 ByteDecoder.num_bytes\[1\]
rlabel metal2 3450 30736 3450 30736 0 ByteDecoder.num_bytes\[2\]
rlabel metal1 3588 28730 3588 28730 0 ByteDecoder.num_bytes\[3\]
rlabel metal1 4876 30702 4876 30702 0 ByteDecoder.state\[0\]
rlabel metal2 5106 31076 5106 31076 0 ByteDecoder.state\[1\]
rlabel metal1 4554 30906 4554 30906 0 FSM.next_state\[0\]
rlabel metal1 5934 30090 5934 30090 0 FSM.next_state\[1\]
rlabel metal1 2530 23630 2530 23630 0 MemControl.state\[0\]
rlabel metal1 3772 23630 3772 23630 0 MemControl.state\[1\]
rlabel metal1 3772 25330 3772 25330 0 MemControl.state\[2\]
rlabel metal1 21252 36142 21252 36142 0 PC.i_mem_addr\[0\]
rlabel metal1 20470 35020 20470 35020 0 PC.i_mem_addr\[10\]
rlabel metal2 12650 35904 12650 35904 0 PC.i_mem_addr\[11\]
rlabel metal1 12604 32878 12604 32878 0 PC.i_mem_addr\[12\]
rlabel metal1 13294 30804 13294 30804 0 PC.i_mem_addr\[13\]
rlabel metal2 12742 29036 12742 29036 0 PC.i_mem_addr\[14\]
rlabel metal1 13478 27370 13478 27370 0 PC.i_mem_addr\[15\]
rlabel metal1 21160 36074 21160 36074 0 PC.i_mem_addr\[1\]
rlabel metal1 21114 38182 21114 38182 0 PC.i_mem_addr\[2\]
rlabel metal1 22954 35122 22954 35122 0 PC.i_mem_addr\[3\]
rlabel metal1 25944 35734 25944 35734 0 PC.i_mem_addr\[4\]
rlabel metal1 24932 37978 24932 37978 0 PC.i_mem_addr\[5\]
rlabel metal2 21574 37196 21574 37196 0 PC.i_mem_addr\[6\]
rlabel metal1 16928 37978 16928 37978 0 PC.i_mem_addr\[7\]
rlabel metal1 15548 27098 15548 27098 0 PC.i_mem_addr\[8\]
rlabel metal2 12466 34544 12466 34544 0 PC.i_mem_addr\[9\]
rlabel metal1 32338 16762 32338 16762 0 RegFile.A\[0\]
rlabel metal1 30866 3094 30866 3094 0 RegFile.A\[1\]
rlabel metal2 6394 10268 6394 10268 0 RegFile.A\[2\]
rlabel metal1 15318 9996 15318 9996 0 RegFile.A\[3\]
rlabel metal1 12466 2380 12466 2380 0 RegFile.A\[4\]
rlabel metal2 5290 13498 5290 13498 0 RegFile.A\[5\]
rlabel metal1 6762 15606 6762 15606 0 RegFile.A\[6\]
rlabel metal2 18630 3230 18630 3230 0 RegFile.A\[7\]
rlabel metal2 32614 15130 32614 15130 0 RegFile.B\[0\]
rlabel metal1 29854 7820 29854 7820 0 RegFile.B\[1\]
rlabel metal2 8510 10880 8510 10880 0 RegFile.B\[2\]
rlabel metal1 7038 7514 7038 7514 0 RegFile.B\[3\]
rlabel viali 20102 10030 20102 10030 0 RegFile.B\[4\]
rlabel metal1 26652 12818 26652 12818 0 RegFile.B\[5\]
rlabel metal1 6716 14450 6716 14450 0 RegFile.B\[6\]
rlabel metal2 20746 4794 20746 4794 0 RegFile.B\[7\]
rlabel metal1 33580 14246 33580 14246 0 RegFile.C\[0\]
rlabel metal1 32292 5338 32292 5338 0 RegFile.C\[1\]
rlabel metal1 12144 8806 12144 8806 0 RegFile.C\[2\]
rlabel metal1 16284 6766 16284 6766 0 RegFile.C\[3\]
rlabel metal1 27508 9554 27508 9554 0 RegFile.C\[4\]
rlabel metal1 27646 12750 27646 12750 0 RegFile.C\[5\]
rlabel metal2 16514 13498 16514 13498 0 RegFile.C\[6\]
rlabel metal2 22034 8160 22034 8160 0 RegFile.C\[7\]
rlabel metal1 24224 16082 24224 16082 0 RegFile.D\[0\]
rlabel metal1 26450 3366 26450 3366 0 RegFile.D\[1\]
rlabel metal1 8188 9690 8188 9690 0 RegFile.D\[2\]
rlabel metal1 8556 7514 8556 7514 0 RegFile.D\[3\]
rlabel metal2 13938 3230 13938 3230 0 RegFile.D\[4\]
rlabel via1 24702 12818 24702 12818 0 RegFile.D\[5\]
rlabel metal2 8510 13906 8510 13906 0 RegFile.D\[6\]
rlabel metal1 17986 3910 17986 3910 0 RegFile.D\[7\]
rlabel metal2 32522 14314 32522 14314 0 RegFile.E\[0\]
rlabel metal1 30912 5338 30912 5338 0 RegFile.E\[1\]
rlabel metal2 18032 10642 18032 10642 0 RegFile.E\[2\]
rlabel metal1 17710 6426 17710 6426 0 RegFile.E\[3\]
rlabel metal2 28198 10846 28198 10846 0 RegFile.E\[4\]
rlabel metal1 25944 13294 25944 13294 0 RegFile.E\[5\]
rlabel metal1 21344 13906 21344 13906 0 RegFile.E\[6\]
rlabel metal1 21298 8840 21298 8840 0 RegFile.E\[7\]
rlabel metal1 28014 17306 28014 17306 0 RegFile.H\[0\]
rlabel metal1 25714 6800 25714 6800 0 RegFile.H\[1\]
rlabel metal1 19826 11152 19826 11152 0 RegFile.H\[2\]
rlabel via1 18456 7378 18456 7378 0 RegFile.H\[3\]
rlabel metal1 21298 10574 21298 10574 0 RegFile.H\[4\]
rlabel metal1 18722 13158 18722 13158 0 RegFile.H\[5\]
rlabel metal1 9292 14926 9292 14926 0 RegFile.H\[6\]
rlabel metal1 21344 2890 21344 2890 0 RegFile.H\[7\]
rlabel viali 25898 15470 25898 15470 0 RegFile.L\[0\]
rlabel metal1 32246 7242 32246 7242 0 RegFile.L\[1\]
rlabel metal1 17020 9622 17020 9622 0 RegFile.L\[2\]
rlabel metal2 14582 5338 14582 5338 0 RegFile.L\[3\]
rlabel metal1 27278 9520 27278 9520 0 RegFile.L\[4\]
rlabel metal1 27830 12342 27830 12342 0 RegFile.L\[5\]
rlabel metal1 14536 13974 14536 13974 0 RegFile.L\[6\]
rlabel metal1 23874 5134 23874 5134 0 RegFile.L\[7\]
rlabel metal1 3312 23834 3312 23834 0 _0000_
rlabel metal1 2116 24922 2116 24922 0 _0001_
rlabel metal1 1748 23154 1748 23154 0 _0066_
rlabel metal1 2162 28424 2162 28424 0 _0067_
rlabel metal1 3128 30906 3128 30906 0 _0068_
rlabel metal1 1794 29274 1794 29274 0 _0069_
rlabel metal1 5842 33626 5842 33626 0 _0070_
rlabel metal1 7130 33558 7130 33558 0 _0071_
rlabel metal1 6624 31450 6624 31450 0 _0072_
rlabel metal1 4554 33082 4554 33082 0 _0073_
rlabel metal1 8096 32470 8096 32470 0 _0074_
rlabel metal1 7728 30362 7728 30362 0 _0075_
rlabel metal1 7682 29274 7682 29274 0 _0076_
rlabel metal2 8326 27812 8326 27812 0 _0077_
rlabel metal1 4370 17272 4370 17272 0 _0078_
rlabel metal1 5520 17578 5520 17578 0 _0079_
rlabel metal1 2346 16626 2346 16626 0 _0080_
rlabel metal1 3220 21862 3220 21862 0 _0081_
rlabel metal1 6210 21658 6210 21658 0 _0082_
rlabel metal2 8326 25058 8326 25058 0 _0083_
rlabel metal1 1886 18360 1886 18360 0 _0084_
rlabel metal1 9614 24106 9614 24106 0 _0085_
rlabel metal1 4738 21862 4738 21862 0 _0086_
rlabel metal2 6486 20060 6486 20060 0 _0087_
rlabel metal2 4094 19618 4094 19618 0 _0088_
rlabel metal1 1787 21114 1787 21114 0 _0089_
rlabel metal1 6992 23290 6992 23290 0 _0090_
rlabel metal1 9062 27030 9062 27030 0 _0091_
rlabel metal1 1840 19414 1840 19414 0 _0092_
rlabel metal1 11500 24922 11500 24922 0 _0093_
rlabel metal2 25070 19618 25070 19618 0 _0094_
rlabel metal1 28888 17850 28888 17850 0 _0095_
rlabel metal1 17388 19278 17388 19278 0 _0096_
rlabel metal1 12696 7922 12696 7922 0 _0097_
rlabel metal2 30498 9180 30498 9180 0 _0098_
rlabel metal1 30222 11866 30222 11866 0 _0099_
rlabel metal1 19872 18394 19872 18394 0 _0100_
rlabel metal1 22034 19720 22034 19720 0 _0101_
rlabel metal1 33028 16626 33028 16626 0 _0102_
rlabel metal1 32108 6970 32108 6970 0 _0103_
rlabel metal1 12742 9146 12742 9146 0 _0104_
rlabel metal1 13248 4726 13248 4726 0 _0105_
rlabel metal1 34684 9622 34684 9622 0 _0106_
rlabel metal1 33672 13498 33672 13498 0 _0107_
rlabel metal1 13340 12886 13340 12886 0 _0108_
rlabel metal1 24610 4658 24610 4658 0 _0109_
rlabel metal1 27140 17714 27140 17714 0 _0110_
rlabel metal1 27738 4488 27738 4488 0 _0111_
rlabel metal1 9246 9928 9246 9928 0 _0112_
rlabel metal1 9476 7446 9476 7446 0 _0113_
rlabel metal1 14858 3128 14858 3128 0 _0114_
rlabel metal1 9016 5270 9016 5270 0 _0115_
rlabel metal1 7636 15062 7636 15062 0 _0116_
rlabel metal1 20240 3094 20240 3094 0 _0117_
rlabel metal2 31418 14178 31418 14178 0 _0118_
rlabel metal1 29992 5746 29992 5746 0 _0119_
rlabel metal1 12742 11322 12742 11322 0 _0120_
rlabel metal1 12144 5882 12144 5882 0 _0121_
rlabel metal2 31326 10268 31326 10268 0 _0122_
rlabel metal1 32246 12750 32246 12750 0 _0123_
rlabel metal1 19826 12886 19826 12886 0 _0124_
rlabel metal1 22172 3094 22172 3094 0 _0125_
rlabel metal1 23000 14450 23000 14450 0 _0126_
rlabel metal1 26956 2958 26956 2958 0 _0127_
rlabel metal1 6670 9656 6670 9656 0 _0128_
rlabel metal1 7498 7514 7498 7514 0 _0129_
rlabel metal1 12236 3570 12236 3570 0 _0130_
rlabel metal1 7176 5066 7176 5066 0 _0131_
rlabel metal1 7084 13362 7084 13362 0 _0132_
rlabel metal1 16882 4046 16882 4046 0 _0133_
rlabel metal1 33626 15096 33626 15096 0 _0134_
rlabel metal2 31786 5338 31786 5338 0 _0135_
rlabel metal1 10212 9146 10212 9146 0 _0136_
rlabel metal2 15042 4930 15042 4930 0 _0137_
rlabel metal1 32798 8874 32798 8874 0 _0138_
rlabel metal1 34684 11798 34684 11798 0 _0139_
rlabel metal2 15226 13600 15226 13600 0 _0140_
rlabel metal1 21620 4250 21620 4250 0 _0141_
rlabel metal1 30958 15402 30958 15402 0 _0142_
rlabel metal2 28106 4692 28106 4692 0 _0143_
rlabel metal1 7084 11186 7084 11186 0 _0144_
rlabel metal1 5835 6970 5835 6970 0 _0145_
rlabel metal1 10718 5066 10718 5066 0 _0146_
rlabel metal1 5566 11866 5566 11866 0 _0147_
rlabel metal1 5244 14042 5244 14042 0 _0148_
rlabel metal2 19274 5338 19274 5338 0 _0149_
rlabel via1 30951 16762 30951 16762 0 _0150_
rlabel metal1 24656 2958 24656 2958 0 _0151_
rlabel metal1 4685 10234 4685 10234 0 _0152_
rlabel metal2 4922 8228 4922 8228 0 _0153_
rlabel metal1 9752 2890 9752 2890 0 _0154_
rlabel metal2 4554 12716 4554 12716 0 _0155_
rlabel metal1 5060 15538 5060 15538 0 _0156_
rlabel metal1 17618 3128 17618 3128 0 _0157_
rlabel metal1 18492 36346 18492 36346 0 _0158_
rlabel metal1 22218 37978 22218 37978 0 _0159_
rlabel metal1 20056 37978 20056 37978 0 _0160_
rlabel metal2 21022 34408 21022 34408 0 _0161_
rlabel metal1 23690 34170 23690 34170 0 _0162_
rlabel metal1 24610 38386 24610 38386 0 _0163_
rlabel metal2 17618 38658 17618 38658 0 _0164_
rlabel metal1 15456 37978 15456 37978 0 _0165_
rlabel metal1 14582 35258 14582 35258 0 _0166_
rlabel metal1 9936 35802 9936 35802 0 _0167_
rlabel metal1 13110 36856 13110 36856 0 _0168_
rlabel metal2 8970 35428 8970 35428 0 _0169_
rlabel metal2 9798 33320 9798 33320 0 _0170_
rlabel metal1 9706 30906 9706 30906 0 _0171_
rlabel metal1 9568 29206 9568 29206 0 _0172_
rlabel metal1 11546 26418 11546 26418 0 _0173_
rlabel metal2 34454 27710 34454 27710 0 _0174_
rlabel metal1 31234 25466 31234 25466 0 _0175_
rlabel metal1 32062 26010 32062 26010 0 _0176_
rlabel metal2 32982 26724 32982 26724 0 _0177_
rlabel metal1 33718 26996 33718 26996 0 _0178_
rlabel metal1 34638 26826 34638 26826 0 _0179_
rlabel metal1 34454 26350 34454 26350 0 _0180_
rlabel metal2 34730 27506 34730 27506 0 _0181_
rlabel metal1 33166 26520 33166 26520 0 _0182_
rlabel metal1 18860 32538 18860 32538 0 _0183_
rlabel metal1 17894 32912 17894 32912 0 _0184_
rlabel metal2 17802 33354 17802 33354 0 _0185_
rlabel metal1 17802 26486 17802 26486 0 _0186_
rlabel metal4 12972 10324 12972 10324 0 _0187_
rlabel metal1 5244 7854 5244 7854 0 _0188_
rlabel metal1 34960 23834 34960 23834 0 _0189_
rlabel metal1 35512 24242 35512 24242 0 _0190_
rlabel metal1 36754 23562 36754 23562 0 _0191_
rlabel metal1 36478 23732 36478 23732 0 _0192_
rlabel metal2 37122 21046 37122 21046 0 _0193_
rlabel metal1 36892 23086 36892 23086 0 _0194_
rlabel metal1 33304 23698 33304 23698 0 _0195_
rlabel metal1 33626 21862 33626 21862 0 _0196_
rlabel metal1 32890 23494 32890 23494 0 _0197_
rlabel metal2 33166 24038 33166 24038 0 _0198_
rlabel metal1 32890 23800 32890 23800 0 _0199_
rlabel metal1 35604 23086 35604 23086 0 _0200_
rlabel metal1 36386 23290 36386 23290 0 _0201_
rlabel metal2 36294 24072 36294 24072 0 _0202_
rlabel metal1 19780 25670 19780 25670 0 _0203_
rlabel metal2 20470 32640 20470 32640 0 _0204_
rlabel metal1 19826 33524 19826 33524 0 _0205_
rlabel metal1 19872 32878 19872 32878 0 _0206_
rlabel metal1 19734 33014 19734 33014 0 _0207_
rlabel metal1 16100 26282 16100 26282 0 _0208_
rlabel metal2 15778 24480 15778 24480 0 _0209_
rlabel metal1 5198 10642 5198 10642 0 _0210_
rlabel metal1 35558 22032 35558 22032 0 _0211_
rlabel metal2 35926 22474 35926 22474 0 _0212_
rlabel metal1 35374 19482 35374 19482 0 _0213_
rlabel metal2 34822 20944 34822 20944 0 _0214_
rlabel metal1 33304 21114 33304 21114 0 _0215_
rlabel metal1 33948 20026 33948 20026 0 _0216_
rlabel metal1 32890 21964 32890 21964 0 _0217_
rlabel metal1 32246 22202 32246 22202 0 _0218_
rlabel metal1 33074 21998 33074 21998 0 _0219_
rlabel metal1 33580 22066 33580 22066 0 _0220_
rlabel metal1 34684 21998 34684 21998 0 _0221_
rlabel metal1 35512 22202 35512 22202 0 _0222_
rlabel metal1 20102 37230 20102 37230 0 _0223_
rlabel metal1 22911 31654 22911 31654 0 _0224_
rlabel via1 22199 31314 22199 31314 0 _0225_
rlabel metal1 21620 31178 21620 31178 0 _0226_
rlabel metal1 21344 30294 21344 30294 0 _0227_
rlabel metal2 21022 29240 21022 29240 0 _0228_
rlabel metal3 25323 23596 25323 23596 0 _0229_
rlabel metal1 25300 2414 25300 2414 0 _0230_
rlabel metal1 31004 20910 31004 20910 0 _0231_
rlabel metal1 31924 20298 31924 20298 0 _0232_
rlabel metal1 31004 20026 31004 20026 0 _0233_
rlabel metal1 31372 20978 31372 20978 0 _0234_
rlabel metal1 30728 21114 30728 21114 0 _0235_
rlabel metal1 30452 22542 30452 22542 0 _0236_
rlabel metal2 31326 23018 31326 23018 0 _0237_
rlabel metal1 29992 21658 29992 21658 0 _0238_
rlabel metal1 29578 21930 29578 21930 0 _0239_
rlabel metal2 30130 22610 30130 22610 0 _0240_
rlabel metal1 30544 22610 30544 22610 0 _0241_
rlabel metal2 19274 25823 19274 25823 0 _0242_
rlabel metal1 24656 29478 24656 29478 0 _0243_
rlabel metal1 23736 30090 23736 30090 0 _0244_
rlabel metal1 24150 30226 24150 30226 0 _0245_
rlabel metal1 24426 30192 24426 30192 0 _0246_
rlabel metal2 18722 26418 18722 26418 0 _0247_
rlabel metal1 23690 13974 23690 13974 0 _0248_
rlabel metal1 30636 17170 30636 17170 0 _0249_
rlabel metal2 10258 15164 10258 15164 0 _0250_
rlabel metal1 19044 4658 19044 4658 0 _0251_
rlabel metal1 19412 4454 19412 4454 0 _0252_
rlabel metal1 5980 13906 5980 13906 0 _0253_
rlabel metal1 6118 11730 6118 11730 0 _0254_
rlabel metal1 11270 5202 11270 5202 0 _0255_
rlabel metal1 6256 7378 6256 7378 0 _0256_
rlabel metal1 7498 10778 7498 10778 0 _0257_
rlabel metal1 27232 4794 27232 4794 0 _0258_
rlabel metal1 30682 15130 30682 15130 0 _0259_
rlabel metal2 13294 23460 13294 23460 0 _0260_
rlabel metal1 21622 24174 21622 24174 0 _0261_
rlabel metal1 21436 24174 21436 24174 0 _0262_
rlabel metal2 22586 19907 22586 19907 0 _0263_
rlabel metal1 10258 13328 10258 13328 0 _0264_
rlabel metal1 8786 12818 8786 12818 0 _0265_
rlabel metal1 9752 12886 9752 12886 0 _0266_
rlabel metal1 11362 13430 11362 13430 0 _0267_
rlabel metal1 11270 13362 11270 13362 0 _0268_
rlabel metal1 33580 14450 33580 14450 0 _0269_
rlabel metal1 21988 4114 21988 4114 0 _0270_
rlabel metal1 14812 24582 14812 24582 0 _0271_
rlabel metal1 15502 13294 15502 13294 0 _0272_
rlabel metal1 33534 12308 33534 12308 0 _0273_
rlabel metal1 34362 12172 34362 12172 0 _0274_
rlabel metal2 21804 18428 21804 18428 0 _0275_
rlabel metal1 32430 9044 32430 9044 0 _0276_
rlabel metal2 13892 20570 13892 20570 0 _0277_
rlabel metal1 15226 4658 15226 4658 0 _0278_
rlabel metal2 17158 18547 17158 18547 0 _0279_
rlabel metal1 10718 8874 10718 8874 0 _0280_
rlabel metal1 32614 5066 32614 5066 0 _0281_
rlabel metal1 32154 5100 32154 5100 0 _0282_
rlabel metal1 33488 16218 33488 16218 0 _0283_
rlabel metal1 33166 14586 33166 14586 0 _0284_
rlabel metal1 8970 12682 8970 12682 0 _0285_
rlabel metal1 10166 11764 10166 11764 0 _0286_
rlabel metal1 11178 11696 11178 11696 0 _0287_
rlabel metal1 16974 3570 16974 3570 0 _0288_
rlabel metal1 16744 3706 16744 3706 0 _0289_
rlabel metal1 7544 13906 7544 13906 0 _0290_
rlabel metal1 7590 5202 7590 5202 0 _0291_
rlabel metal1 12742 2890 12742 2890 0 _0292_
rlabel metal1 7958 7378 7958 7378 0 _0293_
rlabel metal1 7176 10030 7176 10030 0 _0294_
rlabel metal1 26588 3026 26588 3026 0 _0295_
rlabel metal2 23414 14518 23414 14518 0 _0296_
rlabel metal2 20194 13175 20194 13175 0 _0297_
rlabel metal1 22678 3502 22678 3502 0 _0298_
rlabel metal1 19366 12886 19366 12886 0 _0299_
rlabel metal2 31970 13124 31970 13124 0 _0300_
rlabel metal1 31786 10642 31786 10642 0 _0301_
rlabel metal1 12558 5712 12558 5712 0 _0302_
rlabel metal1 13110 11118 13110 11118 0 _0303_
rlabel metal1 30130 5338 30130 5338 0 _0304_
rlabel metal1 31947 14042 31947 14042 0 _0305_
rlabel metal1 10626 13192 10626 13192 0 _0306_
rlabel metal2 19366 16405 19366 16405 0 _0307_
rlabel metal1 20746 3570 20746 3570 0 _0308_
rlabel metal2 9154 15300 9154 15300 0 _0309_
rlabel metal1 9292 5678 9292 5678 0 _0310_
rlabel metal1 15180 3502 15180 3502 0 _0311_
rlabel metal1 9752 7854 9752 7854 0 _0312_
rlabel metal1 8464 10030 8464 10030 0 _0313_
rlabel metal2 27002 4726 27002 4726 0 _0314_
rlabel metal2 27002 17782 27002 17782 0 _0315_
rlabel metal1 14490 13872 14490 13872 0 _0316_
rlabel metal1 23782 4692 23782 4692 0 _0317_
rlabel metal1 13846 13906 13846 13906 0 _0318_
rlabel metal1 33212 13294 33212 13294 0 _0319_
rlabel metal1 33948 10642 33948 10642 0 _0320_
rlabel metal1 13846 4590 13846 4590 0 _0321_
rlabel metal1 13294 8976 13294 8976 0 _0322_
rlabel metal2 31970 6970 31970 6970 0 _0323_
rlabel metal2 33258 16694 33258 16694 0 _0324_
rlabel metal2 17526 27234 17526 27234 0 _0325_
rlabel metal1 18354 22610 18354 22610 0 _0326_
rlabel metal1 22356 19482 22356 19482 0 _0327_
rlabel metal1 9982 19142 9982 19142 0 _0328_
rlabel metal1 9752 18598 9752 18598 0 _0329_
rlabel metal1 9660 18938 9660 18938 0 _0330_
rlabel metal1 9706 19278 9706 19278 0 _0331_
rlabel metal1 10396 19754 10396 19754 0 _0332_
rlabel metal1 9752 19754 9752 19754 0 _0333_
rlabel metal1 18906 18802 18906 18802 0 _0334_
rlabel metal1 21942 19482 21942 19482 0 _0335_
rlabel metal1 19274 18224 19274 18224 0 _0336_
rlabel via2 18354 26435 18354 26435 0 _0337_
rlabel metal1 17710 25432 17710 25432 0 _0338_
rlabel metal1 17894 25330 17894 25330 0 _0339_
rlabel metal1 18262 25296 18262 25296 0 _0340_
rlabel metal1 17756 25194 17756 25194 0 _0341_
rlabel metal1 18354 20434 18354 20434 0 _0342_
rlabel metal2 19366 18513 19366 18513 0 _0343_
rlabel metal1 19136 18258 19136 18258 0 _0344_
rlabel metal1 19688 28730 19688 28730 0 _0345_
rlabel metal1 19550 27948 19550 27948 0 _0346_
rlabel metal1 33994 29172 33994 29172 0 _0347_
rlabel metal1 35558 29274 35558 29274 0 _0348_
rlabel metal1 36570 22712 36570 22712 0 _0349_
rlabel metal1 37674 22678 37674 22678 0 _0350_
rlabel metal1 34178 22644 34178 22644 0 _0351_
rlabel metal1 36938 22542 36938 22542 0 _0352_
rlabel metal1 37352 22406 37352 22406 0 _0353_
rlabel metal1 37490 29648 37490 29648 0 _0354_
rlabel metal1 32752 30702 32752 30702 0 _0355_
rlabel metal1 32660 30838 32660 30838 0 _0356_
rlabel metal1 32476 23222 32476 23222 0 _0357_
rlabel metal1 35420 30158 35420 30158 0 _0358_
rlabel metal2 21942 29121 21942 29121 0 _0359_
rlabel metal1 22264 28594 22264 28594 0 _0360_
rlabel metal1 16951 29818 16951 29818 0 _0361_
rlabel metal1 20700 29818 20700 29818 0 _0362_
rlabel metal1 20332 29818 20332 29818 0 _0363_
rlabel metal1 21068 29546 21068 29546 0 _0364_
rlabel metal1 21206 29648 21206 29648 0 _0365_
rlabel metal1 24794 29070 24794 29070 0 _0366_
rlabel metal1 29118 29580 29118 29580 0 _0367_
rlabel metal1 24058 29104 24058 29104 0 _0368_
rlabel metal1 24334 29036 24334 29036 0 _0369_
rlabel metal1 21252 29070 21252 29070 0 _0370_
rlabel via1 21490 29206 21490 29206 0 _0371_
rlabel metal2 22218 29240 22218 29240 0 _0372_
rlabel viali 22128 28526 22128 28526 0 _0373_
rlabel metal1 22540 27846 22540 27846 0 _0374_
rlabel via1 22863 28050 22863 28050 0 _0375_
rlabel metal1 32821 27914 32821 27914 0 _0376_
rlabel metal1 22586 27472 22586 27472 0 _0377_
rlabel metal2 22770 27642 22770 27642 0 _0378_
rlabel metal1 19228 24718 19228 24718 0 _0379_
rlabel metal1 20240 24922 20240 24922 0 _0380_
rlabel metal1 20378 25330 20378 25330 0 _0381_
rlabel metal1 21114 25466 21114 25466 0 _0382_
rlabel metal1 21160 26418 21160 26418 0 _0383_
rlabel metal1 21919 26486 21919 26486 0 _0384_
rlabel metal1 22770 26554 22770 26554 0 _0385_
rlabel metal1 23092 26826 23092 26826 0 _0386_
rlabel metal1 17158 20570 17158 20570 0 _0387_
rlabel metal1 17342 19890 17342 19890 0 _0388_
rlabel metal2 17894 19890 17894 19890 0 _0389_
rlabel metal1 29256 17850 29256 17850 0 _0390_
rlabel metal2 25714 33082 25714 33082 0 _0391_
rlabel metal1 24932 32742 24932 32742 0 _0392_
rlabel metal1 27784 28526 27784 28526 0 _0393_
rlabel metal1 25346 22610 25346 22610 0 _0394_
rlabel metal1 26036 22746 26036 22746 0 _0395_
rlabel metal1 27554 28492 27554 28492 0 _0396_
rlabel metal1 24886 28560 24886 28560 0 _0397_
rlabel metal1 24334 28050 24334 28050 0 _0398_
rlabel metal1 19734 27438 19734 27438 0 _0399_
rlabel metal1 19412 27642 19412 27642 0 _0400_
rlabel metal1 19274 28118 19274 28118 0 _0401_
rlabel metal1 23966 27982 23966 27982 0 _0402_
rlabel metal1 18630 23664 18630 23664 0 _0403_
rlabel metal1 24702 19924 24702 19924 0 _0404_
rlabel metal1 25024 19346 25024 19346 0 _0405_
rlabel metal1 7636 32946 7636 32946 0 _0406_
rlabel metal1 4876 26350 4876 26350 0 _0407_
rlabel metal1 4922 19244 4922 19244 0 _0408_
rlabel metal1 2714 24752 2714 24752 0 _0409_
rlabel metal1 4002 23154 4002 23154 0 _0410_
rlabel metal1 4554 24786 4554 24786 0 _0411_
rlabel metal1 4462 24922 4462 24922 0 _0412_
rlabel metal1 3818 30362 3818 30362 0 _0413_
rlabel metal2 4462 30464 4462 30464 0 _0414_
rlabel metal1 4094 30838 4094 30838 0 _0415_
rlabel metal1 12098 24752 12098 24752 0 _0416_
rlabel metal1 10948 25194 10948 25194 0 _0417_
rlabel metal1 5796 28594 5796 28594 0 _0418_
rlabel metal2 7314 27030 7314 27030 0 _0419_
rlabel metal2 9430 26265 9430 26265 0 _0420_
rlabel metal1 7590 32878 7590 32878 0 _0421_
rlabel metal1 7774 26996 7774 26996 0 _0422_
rlabel metal2 8234 27234 8234 27234 0 _0423_
rlabel metal1 5980 27642 5980 27642 0 _0424_
rlabel metal1 5520 18394 5520 18394 0 _0425_
rlabel metal2 5934 26860 5934 26860 0 _0426_
rlabel metal1 5842 27030 5842 27030 0 _0427_
rlabel metal1 4830 18734 4830 18734 0 _0428_
rlabel metal2 5658 27744 5658 27744 0 _0429_
rlabel metal1 4462 29002 4462 29002 0 _0430_
rlabel metal2 5290 28934 5290 28934 0 _0431_
rlabel metal2 6394 27200 6394 27200 0 _0432_
rlabel metal1 6072 28390 6072 28390 0 _0433_
rlabel metal1 5290 19414 5290 19414 0 _0434_
rlabel metal1 6992 20502 6992 20502 0 _0435_
rlabel metal1 7314 28628 7314 28628 0 _0436_
rlabel metal1 5106 29172 5106 29172 0 _0437_
rlabel metal1 4646 30260 4646 30260 0 _0438_
rlabel metal1 4462 23290 4462 23290 0 _0439_
rlabel metal2 3910 23528 3910 23528 0 _0440_
rlabel metal1 14168 36142 14168 36142 0 _0441_
rlabel metal1 34914 18054 34914 18054 0 _0442_
rlabel metal1 31464 3026 31464 3026 0 _0443_
rlabel metal2 2162 11526 2162 11526 0 _0444_
rlabel metal2 4186 5372 4186 5372 0 _0445_
rlabel metal1 11500 2414 11500 2414 0 _0446_
rlabel metal2 1978 14790 1978 14790 0 _0447_
rlabel metal2 37398 18292 37398 18292 0 _0448_
rlabel metal1 19780 2414 19780 2414 0 _0449_
rlabel metal2 14398 25840 14398 25840 0 _0450_
rlabel metal1 12880 33558 12880 33558 0 _0451_
rlabel metal1 16698 2414 16698 2414 0 _0452_
rlabel metal1 13662 26350 13662 26350 0 _0453_
rlabel metal2 14444 36142 14444 36142 0 _0454_
rlabel metal1 19596 35122 19596 35122 0 _0455_
rlabel metal1 19412 33082 19412 33082 0 _0456_
rlabel metal1 20470 37196 20470 37196 0 _0457_
rlabel metal2 23138 33873 23138 33873 0 _0458_
rlabel metal1 23552 26486 23552 26486 0 _0459_
rlabel metal2 25116 31484 25116 31484 0 _0460_
rlabel metal1 25576 37434 25576 37434 0 _0461_
rlabel metal1 26036 37434 26036 37434 0 _0462_
rlabel metal1 16376 37434 16376 37434 0 _0463_
rlabel metal3 14375 4012 14375 4012 0 _0464_
rlabel metal2 12466 3230 12466 3230 0 _0465_
rlabel metal1 13386 29138 13386 29138 0 _0466_
rlabel metal1 2714 29648 2714 29648 0 _0467_
rlabel metal1 20194 34714 20194 34714 0 _0468_
rlabel metal1 14398 36176 14398 36176 0 _0469_
rlabel metal2 12926 33762 12926 33762 0 _0470_
rlabel metal1 13478 30294 13478 30294 0 _0471_
rlabel metal1 13754 28084 13754 28084 0 _0472_
rlabel metal2 13064 37842 13064 37842 0 _0473_
rlabel metal1 2277 38318 2277 38318 0 _0474_
rlabel metal2 12558 2618 12558 2618 0 _0475_
rlabel metal1 19826 36040 19826 36040 0 _0476_
rlabel metal2 36938 3196 36938 3196 0 _0477_
rlabel metal2 37398 36550 37398 36550 0 _0478_
rlabel metal1 8142 3026 8142 3026 0 _0479_
rlabel metal1 10580 15674 10580 15674 0 _0480_
rlabel metal2 28474 36550 28474 36550 0 _0481_
rlabel metal2 11638 37876 11638 37876 0 _0482_
rlabel metal2 12098 37638 12098 37638 0 _0483_
rlabel metal1 25852 3026 25852 3026 0 _0484_
rlabel metal1 1978 23732 1978 23732 0 _0485_
rlabel metal1 2415 29138 2415 29138 0 _0486_
rlabel metal1 5980 33082 5980 33082 0 _0487_
rlabel metal1 6808 33082 6808 33082 0 _0488_
rlabel metal1 6532 31314 6532 31314 0 _0489_
rlabel metal1 4370 21998 4370 21998 0 _0490_
rlabel metal1 4692 32878 4692 32878 0 _0491_
rlabel metal1 8556 32878 8556 32878 0 _0492_
rlabel metal1 8648 30226 8648 30226 0 _0493_
rlabel metal1 8096 29138 8096 29138 0 _0494_
rlabel metal1 8740 27438 8740 27438 0 _0495_
rlabel metal1 4692 25262 4692 25262 0 _0496_
rlabel metal1 5658 18224 5658 18224 0 _0497_
rlabel metal1 4876 17646 4876 17646 0 _0498_
rlabel metal1 6118 18734 6118 18734 0 _0499_
rlabel metal1 3450 17170 3450 17170 0 _0500_
rlabel metal1 3680 21862 3680 21862 0 _0501_
rlabel metal2 6578 21801 6578 21801 0 _0502_
rlabel metal1 7912 25262 7912 25262 0 _0503_
rlabel metal1 2645 18734 2645 18734 0 _0504_
rlabel metal1 9246 24276 9246 24276 0 _0505_
rlabel metal1 5244 21658 5244 21658 0 _0506_
rlabel metal1 6716 20434 6716 20434 0 _0507_
rlabel metal1 4324 19346 4324 19346 0 _0508_
rlabel metal1 2346 21522 2346 21522 0 _0509_
rlabel metal1 7222 23120 7222 23120 0 _0510_
rlabel metal1 8878 26554 8878 26554 0 _0511_
rlabel metal1 2392 19822 2392 19822 0 _0512_
rlabel metal1 11408 24786 11408 24786 0 _0513_
rlabel metal4 13156 10608 13156 10608 0 _0514_
rlabel via3 22333 12580 22333 12580 0 _0515_
rlabel metal2 19366 7174 19366 7174 0 _0516_
rlabel metal1 12236 5338 12236 5338 0 _0517_
rlabel metal1 13478 19414 13478 19414 0 _0518_
rlabel metal2 20746 19652 20746 19652 0 _0519_
rlabel metal2 20194 23698 20194 23698 0 _0520_
rlabel metal1 19734 22542 19734 22542 0 _0521_
rlabel metal2 20240 33388 20240 33388 0 _0522_
rlabel metal1 16836 23086 16836 23086 0 _0523_
rlabel metal1 18170 21590 18170 21590 0 _0524_
rlabel metal2 15870 22746 15870 22746 0 _0525_
rlabel metal1 17480 22066 17480 22066 0 _0526_
rlabel metal2 17618 23222 17618 23222 0 _0527_
rlabel metal2 18354 23324 18354 23324 0 _0528_
rlabel metal1 16514 23120 16514 23120 0 _0529_
rlabel metal1 17664 22202 17664 22202 0 _0530_
rlabel metal1 17618 21658 17618 21658 0 _0531_
rlabel metal1 17250 21998 17250 21998 0 _0532_
rlabel metal1 17020 22202 17020 22202 0 _0533_
rlabel via2 16790 24157 16790 24157 0 _0534_
rlabel metal1 17020 23290 17020 23290 0 _0535_
rlabel metal2 15962 23188 15962 23188 0 _0536_
rlabel metal1 16422 24208 16422 24208 0 _0537_
rlabel metal1 15134 22746 15134 22746 0 _0538_
rlabel metal2 16054 23562 16054 23562 0 _0539_
rlabel metal2 12282 34102 12282 34102 0 _0540_
rlabel metal1 19872 35258 19872 35258 0 _0541_
rlabel metal1 15502 36244 15502 36244 0 _0542_
rlabel metal1 18998 36142 18998 36142 0 _0543_
rlabel metal1 24748 20570 24748 20570 0 _0544_
rlabel via3 25461 21556 25461 21556 0 _0545_
rlabel metal1 23460 36686 23460 36686 0 _0546_
rlabel metal1 23184 36890 23184 36890 0 _0547_
rlabel metal1 22540 37842 22540 37842 0 _0548_
rlabel metal1 21252 36754 21252 36754 0 _0549_
rlabel metal1 21528 36142 21528 36142 0 _0550_
rlabel metal2 22126 36346 22126 36346 0 _0551_
rlabel metal1 21482 36346 21482 36346 0 _0552_
rlabel metal1 20792 36890 20792 36890 0 _0553_
rlabel metal1 20332 37842 20332 37842 0 _0554_
rlabel metal1 21666 34918 21666 34918 0 _0555_
rlabel metal1 22770 35462 22770 35462 0 _0556_
rlabel metal1 22494 35088 22494 35088 0 _0557_
rlabel metal1 22264 34986 22264 34986 0 _0558_
rlabel metal1 22356 34714 22356 34714 0 _0559_
rlabel metal1 21528 34714 21528 34714 0 _0560_
rlabel metal3 25829 34612 25829 34612 0 _0561_
rlabel metal1 25622 35122 25622 35122 0 _0562_
rlabel metal1 25070 34918 25070 34918 0 _0563_
rlabel metal1 24196 33966 24196 33966 0 _0564_
rlabel metal1 25852 19142 25852 19142 0 _0565_
rlabel metal2 25392 33932 25392 33932 0 _0566_
rlabel metal1 19826 35666 19826 35666 0 _0567_
rlabel metal1 25668 36754 25668 36754 0 _0568_
rlabel metal1 25346 36278 25346 36278 0 _0569_
rlabel metal2 24886 37060 24886 37060 0 _0570_
rlabel metal1 24242 37978 24242 37978 0 _0571_
rlabel metal1 18722 35666 18722 35666 0 _0572_
rlabel metal1 16974 35802 16974 35802 0 _0573_
rlabel metal1 18032 35258 18032 35258 0 _0574_
rlabel metal1 18308 35598 18308 35598 0 _0575_
rlabel metal1 18124 35802 18124 35802 0 _0576_
rlabel metal1 17710 37978 17710 37978 0 _0577_
rlabel metal1 19412 33626 19412 33626 0 _0578_
rlabel metal1 16974 36210 16974 36210 0 _0579_
rlabel metal1 16974 36346 16974 36346 0 _0580_
rlabel metal1 15778 37876 15778 37876 0 _0581_
rlabel metal2 16146 35020 16146 35020 0 _0582_
rlabel metal1 16468 34714 16468 34714 0 _0583_
rlabel metal2 16560 35054 16560 35054 0 _0584_
rlabel metal2 12374 25874 12374 25874 0 _0585_
rlabel metal1 15916 35258 15916 35258 0 _0586_
rlabel metal1 14904 35054 14904 35054 0 _0587_
rlabel metal1 12466 35734 12466 35734 0 _0588_
rlabel metal1 11776 35054 11776 35054 0 _0589_
rlabel metal1 11546 35088 11546 35088 0 _0590_
rlabel metal1 11224 35258 11224 35258 0 _0591_
rlabel metal1 10442 35666 10442 35666 0 _0592_
rlabel metal1 13110 35088 13110 35088 0 _0593_
rlabel metal1 13294 35054 13294 35054 0 _0594_
rlabel metal2 13386 35530 13386 35530 0 _0595_
rlabel metal2 12742 37060 12742 37060 0 _0596_
rlabel metal1 12098 31756 12098 31756 0 _0597_
rlabel metal1 11546 34646 11546 34646 0 _0598_
rlabel metal1 11684 34578 11684 34578 0 _0599_
rlabel metal1 10718 34714 10718 34714 0 _0600_
rlabel metal1 9292 35054 9292 35054 0 _0601_
rlabel metal2 11822 33286 11822 33286 0 _0602_
rlabel metal1 12006 33014 12006 33014 0 _0603_
rlabel metal1 11224 32878 11224 32878 0 _0604_
rlabel metal1 10212 32878 10212 32878 0 _0605_
rlabel metal1 11316 30838 11316 30838 0 _0606_
rlabel metal1 11546 31382 11546 31382 0 _0607_
rlabel metal1 11638 31314 11638 31314 0 _0608_
rlabel metal1 10810 30838 10810 30838 0 _0609_
rlabel metal1 10166 30702 10166 30702 0 _0610_
rlabel metal2 11822 28560 11822 28560 0 _0611_
rlabel metal1 11730 29172 11730 29172 0 _0612_
rlabel metal2 11546 29376 11546 29376 0 _0613_
rlabel metal1 10028 29614 10028 29614 0 _0614_
rlabel metal2 12558 27676 12558 27676 0 _0615_
rlabel metal1 12006 27302 12006 27302 0 _0616_
rlabel metal1 11224 27438 11224 27438 0 _0617_
rlabel metal1 13202 24140 13202 24140 0 _0618_
rlabel metal1 8418 21522 8418 21522 0 _0619_
rlabel metal1 9338 18768 9338 18768 0 _0620_
rlabel metal2 13800 21828 13800 21828 0 _0621_
rlabel metal1 8234 17578 8234 17578 0 _0622_
rlabel metal2 15686 20128 15686 20128 0 _0623_
rlabel metal1 4186 18156 4186 18156 0 _0624_
rlabel metal1 10902 23120 10902 23120 0 _0625_
rlabel metal1 13110 16082 13110 16082 0 _0626_
rlabel metal1 5060 29750 5060 29750 0 _0627_
rlabel metal1 15824 20502 15824 20502 0 _0628_
rlabel metal1 28520 19346 28520 19346 0 _0629_
rlabel metal2 9522 13090 9522 13090 0 _0630_
rlabel metal1 21666 24276 21666 24276 0 _0631_
rlabel metal1 9890 21556 9890 21556 0 _0632_
rlabel metal1 12282 16524 12282 16524 0 _0633_
rlabel metal1 14582 17646 14582 17646 0 _0634_
rlabel metal1 14444 20026 14444 20026 0 _0635_
rlabel metal1 15824 19414 15824 19414 0 _0636_
rlabel metal1 14904 17646 14904 17646 0 _0637_
rlabel metal1 17250 9452 17250 9452 0 _0638_
rlabel metal1 8326 18632 8326 18632 0 _0639_
rlabel metal1 16330 17612 16330 17612 0 _0640_
rlabel metal1 8970 16592 8970 16592 0 _0641_
rlabel metal1 9016 17170 9016 17170 0 _0642_
rlabel metal1 7912 16218 7912 16218 0 _0643_
rlabel metal1 16928 17170 16928 17170 0 _0644_
rlabel via1 14927 21522 14927 21522 0 _0645_
rlabel metal2 20470 17238 20470 17238 0 _0646_
rlabel metal1 9890 21998 9890 21998 0 _0647_
rlabel metal1 14306 21522 14306 21522 0 _0648_
rlabel metal1 16284 18326 16284 18326 0 _0649_
rlabel metal1 18722 17068 18722 17068 0 _0650_
rlabel metal2 20838 17476 20838 17476 0 _0651_
rlabel metal1 22126 18870 22126 18870 0 _0652_
rlabel metal1 16100 18734 16100 18734 0 _0653_
rlabel metal1 29854 9010 29854 9010 0 _0654_
rlabel metal1 14582 8500 14582 8500 0 _0655_
rlabel metal2 10994 21896 10994 21896 0 _0656_
rlabel metal1 11178 21012 11178 21012 0 _0657_
rlabel metal2 4738 28526 4738 28526 0 _0658_
rlabel metal2 10350 19737 10350 19737 0 _0659_
rlabel metal1 8970 22032 8970 22032 0 _0660_
rlabel metal1 9522 20434 9522 20434 0 _0661_
rlabel metal1 9798 22678 9798 22678 0 _0662_
rlabel metal1 10166 21454 10166 21454 0 _0663_
rlabel metal2 19458 20587 19458 20587 0 _0664_
rlabel metal2 10718 16626 10718 16626 0 _0665_
rlabel metal2 13110 20128 13110 20128 0 _0666_
rlabel via1 12926 19345 12926 19345 0 _0667_
rlabel metal2 13202 19040 13202 19040 0 _0668_
rlabel metal1 12604 19142 12604 19142 0 _0669_
rlabel metal2 21252 19924 21252 19924 0 _0670_
rlabel metal1 12466 19788 12466 19788 0 _0671_
rlabel metal1 13754 17136 13754 17136 0 _0672_
rlabel metal1 13662 19890 13662 19890 0 _0673_
rlabel metal1 19780 19822 19780 19822 0 _0674_
rlabel metal1 13136 32402 13136 32402 0 _0675_
rlabel metal1 24886 18666 24886 18666 0 _0676_
rlabel metal2 17526 15776 17526 15776 0 _0677_
rlabel metal1 15870 16082 15870 16082 0 _0678_
rlabel metal1 17450 16490 17450 16490 0 _0679_
rlabel metal1 18814 15980 18814 15980 0 _0680_
rlabel metal1 17342 9588 17342 9588 0 _0681_
rlabel metal1 20148 6426 20148 6426 0 _0682_
rlabel metal1 17733 14994 17733 14994 0 _0683_
rlabel metal1 22494 16490 22494 16490 0 _0684_
rlabel metal1 27048 9622 27048 9622 0 _0685_
rlabel metal1 18262 15436 18262 15436 0 _0686_
rlabel metal1 25990 7344 25990 7344 0 _0687_
rlabel metal1 18170 14960 18170 14960 0 _0688_
rlabel metal1 18308 14858 18308 14858 0 _0689_
rlabel metal1 17572 17850 17572 17850 0 _0690_
rlabel metal1 16238 28526 16238 28526 0 _0691_
rlabel metal1 19872 19754 19872 19754 0 _0692_
rlabel metal1 19504 20570 19504 20570 0 _0693_
rlabel metal1 14168 16082 14168 16082 0 _0694_
rlabel metal2 14398 18938 14398 18938 0 _0695_
rlabel metal1 13110 18700 13110 18700 0 _0696_
rlabel metal1 14858 22066 14858 22066 0 _0697_
rlabel metal2 14214 17340 14214 17340 0 _0698_
rlabel metal1 15318 12614 15318 12614 0 _0699_
rlabel metal2 12466 21114 12466 21114 0 _0700_
rlabel metal1 12650 15674 12650 15674 0 _0701_
rlabel metal2 13386 17340 13386 17340 0 _0702_
rlabel metal1 27692 6630 27692 6630 0 _0703_
rlabel metal2 28244 9316 28244 9316 0 _0704_
rlabel metal1 29716 7854 29716 7854 0 _0705_
rlabel metal1 14720 16082 14720 16082 0 _0706_
rlabel metal1 14904 6698 14904 6698 0 _0707_
rlabel metal1 16054 11050 16054 11050 0 _0708_
rlabel metal1 21482 15368 21482 15368 0 _0709_
rlabel metal1 12512 14586 12512 14586 0 _0710_
rlabel metal1 13386 13328 13386 13328 0 _0711_
rlabel metal1 11960 15130 11960 15130 0 _0712_
rlabel metal1 12236 15674 12236 15674 0 _0713_
rlabel metal1 15226 28526 15226 28526 0 _0714_
rlabel metal1 17940 28050 17940 28050 0 _0715_
rlabel metal1 16054 28730 16054 28730 0 _0716_
rlabel metal1 15548 28050 15548 28050 0 _0717_
rlabel metal2 15962 28662 15962 28662 0 _0718_
rlabel metal2 17986 8262 17986 8262 0 _0719_
rlabel metal1 17802 8602 17802 8602 0 _0720_
rlabel metal1 18262 33490 18262 33490 0 _0721_
rlabel metal1 12098 7242 12098 7242 0 _0722_
rlabel metal1 11500 8058 11500 8058 0 _0723_
rlabel metal1 11822 32402 11822 32402 0 _0724_
rlabel metal2 18078 32810 18078 32810 0 _0725_
rlabel via1 17986 32878 17986 32878 0 _0726_
rlabel metal1 18216 11322 18216 11322 0 _0727_
rlabel metal1 18676 11866 18676 11866 0 _0728_
rlabel metal2 18032 17238 18032 17238 0 _0729_
rlabel metal1 12236 10778 12236 10778 0 _0730_
rlabel metal1 11730 10676 11730 10676 0 _0731_
rlabel metal2 12558 30515 12558 30515 0 _0732_
rlabel metal1 18538 30668 18538 30668 0 _0733_
rlabel metal1 19412 31246 19412 31246 0 _0734_
rlabel metal1 19688 31314 19688 31314 0 _0735_
rlabel metal1 18308 31790 18308 31790 0 _0736_
rlabel metal1 20010 32300 20010 32300 0 _0737_
rlabel metal1 25162 7514 25162 7514 0 _0738_
rlabel metal1 24702 8058 24702 8058 0 _0739_
rlabel metal4 22172 18700 22172 18700 0 _0740_
rlabel metal1 28198 8874 28198 8874 0 _0741_
rlabel metal1 29716 7514 29716 7514 0 _0742_
rlabel metal1 29210 8058 29210 8058 0 _0743_
rlabel metal3 29095 9588 29095 9588 0 _0744_
rlabel viali 21390 32401 21390 32401 0 _0745_
rlabel metal1 21758 32470 21758 32470 0 _0746_
rlabel metal2 25070 15980 25070 15980 0 _0747_
rlabel metal1 25162 16218 25162 16218 0 _0748_
rlabel metal1 24472 18938 24472 18938 0 _0749_
rlabel metal1 26082 15028 26082 15028 0 _0750_
rlabel metal1 26496 15130 26496 15130 0 _0751_
rlabel metal2 26910 16099 26910 16099 0 _0752_
rlabel metal1 24012 32198 24012 32198 0 _0753_
rlabel metal1 24380 31450 24380 31450 0 _0754_
rlabel metal1 24242 31858 24242 31858 0 _0755_
rlabel metal1 23276 32266 23276 32266 0 _0756_
rlabel metal2 17802 18122 17802 18122 0 _0757_
rlabel metal2 12190 17476 12190 17476 0 _0758_
rlabel metal1 18814 17714 18814 17714 0 _0759_
rlabel metal1 18630 14382 18630 14382 0 _0760_
rlabel metal1 18124 10642 18124 10642 0 _0761_
rlabel metal2 17434 7990 17434 7990 0 _0762_
rlabel metal2 20838 15878 20838 15878 0 _0763_
rlabel metal2 25806 12954 25806 12954 0 _0764_
rlabel metal2 19458 14892 19458 14892 0 _0765_
rlabel metal1 22770 17170 22770 17170 0 _0766_
rlabel metal2 18722 15878 18722 15878 0 _0767_
rlabel metal1 24840 12682 24840 12682 0 _0768_
rlabel metal1 25714 12716 25714 12716 0 _0769_
rlabel metal2 21896 6766 21896 6766 0 _0770_
rlabel metal2 17250 8942 17250 8942 0 _0771_
rlabel metal1 21482 17544 21482 17544 0 _0772_
rlabel metal1 25760 12818 25760 12818 0 _0773_
rlabel metal2 18676 6766 18676 6766 0 _0774_
rlabel metal1 28152 19822 28152 19822 0 _0775_
rlabel metal1 27186 13396 27186 13396 0 _0776_
rlabel metal1 27048 13294 27048 13294 0 _0777_
rlabel metal1 27922 19788 27922 19788 0 _0778_
rlabel metal1 23000 20842 23000 20842 0 _0779_
rlabel metal2 30130 20519 30130 20519 0 _0780_
rlabel metal1 27922 26350 27922 26350 0 _0781_
rlabel metal1 29210 27404 29210 27404 0 _0782_
rlabel metal2 14950 15708 14950 15708 0 _0783_
rlabel metal1 21252 14382 21252 14382 0 _0784_
rlabel metal2 27186 6494 27186 6494 0 _0785_
rlabel metal2 15824 9452 15824 9452 0 _0786_
rlabel metal1 24978 12308 24978 12308 0 _0787_
rlabel metal2 22862 9316 22862 9316 0 _0788_
rlabel metal2 21160 13906 21160 13906 0 _0789_
rlabel metal1 28566 12954 28566 12954 0 _0790_
rlabel metal1 28198 13430 28198 13430 0 _0791_
rlabel metal1 22264 9350 22264 9350 0 _0792_
rlabel metal1 20102 13906 20102 13906 0 _0793_
rlabel metal1 21988 13906 21988 13906 0 _0794_
rlabel metal1 27186 12410 27186 12410 0 _0795_
rlabel metal2 27922 13124 27922 13124 0 _0796_
rlabel metal2 27830 13498 27830 13498 0 _0797_
rlabel metal1 29946 13328 29946 13328 0 _0798_
rlabel metal1 29486 12784 29486 12784 0 _0799_
rlabel metal2 29394 13056 29394 13056 0 _0800_
rlabel metal1 30130 12954 30130 12954 0 _0801_
rlabel metal1 29724 26282 29724 26282 0 _0802_
rlabel metal1 29762 30158 29762 30158 0 _0803_
rlabel metal1 30498 30260 30498 30260 0 _0804_
rlabel via1 29394 34595 29394 34595 0 _0805_
rlabel metal2 31694 33490 31694 33490 0 _0806_
rlabel metal1 18032 9554 18032 9554 0 _0807_
rlabel metal1 17848 9418 17848 9418 0 _0808_
rlabel metal1 18492 9690 18492 9690 0 _0809_
rlabel metal1 18906 10506 18906 10506 0 _0810_
rlabel metal1 18492 10574 18492 10574 0 _0811_
rlabel metal1 18400 10778 18400 10778 0 _0812_
rlabel metal1 18722 11152 18722 11152 0 _0813_
rlabel metal1 17618 10744 17618 10744 0 _0814_
rlabel metal2 20930 19754 20930 19754 0 _0815_
rlabel metal1 33488 21998 33488 21998 0 _0816_
rlabel metal1 16008 8262 16008 8262 0 _0817_
rlabel metal1 15272 11118 15272 11118 0 _0818_
rlabel metal1 16514 11186 16514 11186 0 _0819_
rlabel viali 15318 10643 15318 10643 0 _0820_
rlabel metal1 15916 10778 15916 10778 0 _0821_
rlabel metal1 16698 10778 16698 10778 0 _0822_
rlabel metal1 16836 11254 16836 11254 0 _0823_
rlabel metal1 16468 12206 16468 12206 0 _0824_
rlabel metal1 14306 10778 14306 10778 0 _0825_
rlabel metal1 14996 11322 14996 11322 0 _0826_
rlabel metal1 16054 12240 16054 12240 0 _0827_
rlabel metal3 17871 19244 17871 19244 0 _0828_
rlabel metal1 19826 19958 19826 19958 0 _0829_
rlabel metal1 20102 21114 20102 21114 0 _0830_
rlabel via2 21206 19771 21206 19771 0 _0831_
rlabel metal1 36570 25296 36570 25296 0 _0832_
rlabel metal2 15410 7820 15410 7820 0 _0833_
rlabel metal1 16284 7514 16284 7514 0 _0834_
rlabel metal1 16146 7208 16146 7208 0 _0835_
rlabel metal1 16054 8058 16054 8058 0 _0836_
rlabel metal1 16376 7854 16376 7854 0 _0837_
rlabel metal2 16790 8772 16790 8772 0 _0838_
rlabel metal1 16330 9588 16330 9588 0 _0839_
rlabel metal1 14628 6766 14628 6766 0 _0840_
rlabel metal1 15548 6630 15548 6630 0 _0841_
rlabel metal1 16100 9146 16100 9146 0 _0842_
rlabel metal3 18768 18020 18768 18020 0 _0843_
rlabel metal1 21620 21590 21620 21590 0 _0844_
rlabel metal2 17802 5916 17802 5916 0 _0845_
rlabel metal1 17664 6154 17664 6154 0 _0846_
rlabel metal1 18308 6426 18308 6426 0 _0847_
rlabel metal2 18446 7038 18446 7038 0 _0848_
rlabel metal1 18768 6834 18768 6834 0 _0849_
rlabel metal1 18216 6970 18216 6970 0 _0850_
rlabel metal1 18446 7514 18446 7514 0 _0851_
rlabel metal1 17710 6630 17710 6630 0 _0852_
rlabel metal1 20792 21998 20792 21998 0 _0853_
rlabel metal1 29302 21658 29302 21658 0 _0854_
rlabel metal1 32522 23630 32522 23630 0 _0855_
rlabel metal1 36340 28186 36340 28186 0 _0856_
rlabel metal1 24794 6222 24794 6222 0 _0857_
rlabel metal1 24886 5882 24886 5882 0 _0858_
rlabel metal2 24886 6562 24886 6562 0 _0859_
rlabel metal1 24978 6732 24978 6732 0 _0860_
rlabel metal1 25530 6086 25530 6086 0 _0861_
rlabel metal2 25070 7514 25070 7514 0 _0862_
rlabel metal1 25714 8398 25714 8398 0 _0863_
rlabel metal1 25990 6970 25990 6970 0 _0864_
rlabel metal1 26036 7242 26036 7242 0 _0865_
rlabel viali 26178 8466 26178 8466 0 _0866_
rlabel via1 34454 20910 34454 20910 0 _0867_
rlabel metal1 35972 19822 35972 19822 0 _0868_
rlabel metal1 33304 18734 33304 18734 0 _0869_
rlabel metal1 27968 8058 27968 8058 0 _0870_
rlabel metal1 28474 8398 28474 8398 0 _0871_
rlabel metal1 28428 6426 28428 6426 0 _0872_
rlabel metal1 28106 6698 28106 6698 0 _0873_
rlabel metal1 28428 6834 28428 6834 0 _0874_
rlabel metal1 28290 6766 28290 6766 0 _0875_
rlabel metal1 29164 8602 29164 8602 0 _0876_
rlabel metal2 29578 7004 29578 7004 0 _0877_
rlabel metal1 30452 7514 30452 7514 0 _0878_
rlabel metal2 30590 8466 30590 8466 0 _0879_
rlabel metal2 30130 9384 30130 9384 0 _0880_
rlabel metal1 35834 19924 35834 19924 0 _0881_
rlabel metal1 37076 20230 37076 20230 0 _0882_
rlabel metal1 33580 20434 33580 20434 0 _0883_
rlabel metal1 33948 19346 33948 19346 0 _0884_
rlabel metal1 20378 21352 20378 21352 0 _0885_
rlabel metal1 26864 14790 26864 14790 0 _0886_
rlabel metal1 27784 15470 27784 15470 0 _0887_
rlabel metal1 28658 15606 28658 15606 0 _0888_
rlabel metal1 28704 15062 28704 15062 0 _0889_
rlabel metal1 28704 15130 28704 15130 0 _0890_
rlabel metal1 28658 15504 28658 15504 0 _0891_
rlabel metal2 29118 15878 29118 15878 0 _0892_
rlabel metal1 30360 15674 30360 15674 0 _0893_
rlabel metal1 30590 15878 30590 15878 0 _0894_
rlabel metal1 29578 16116 29578 16116 0 _0895_
rlabel metal1 31096 19346 31096 19346 0 _0896_
rlabel metal1 25208 15470 25208 15470 0 _0897_
rlabel metal1 26128 15674 26128 15674 0 _0898_
rlabel metal1 25576 17102 25576 17102 0 _0899_
rlabel metal1 24840 17034 24840 17034 0 _0900_
rlabel metal1 25070 17170 25070 17170 0 _0901_
rlabel metal2 24702 17714 24702 17714 0 _0902_
rlabel metal2 26082 19448 26082 19448 0 _0903_
rlabel metal1 26634 16218 26634 16218 0 _0904_
rlabel metal1 26588 16490 26588 16490 0 _0905_
rlabel via1 27178 19414 27178 19414 0 _0906_
rlabel metal2 27002 19958 27002 19958 0 _0907_
rlabel metal1 28474 24242 28474 24242 0 _0908_
rlabel metal1 32752 19822 32752 19822 0 _0909_
rlabel metal1 34178 20332 34178 20332 0 _0910_
rlabel metal1 36846 21012 36846 21012 0 _0911_
rlabel metal2 36938 21284 36938 21284 0 _0912_
rlabel metal1 36064 29070 36064 29070 0 _0913_
rlabel metal1 25990 11152 25990 11152 0 _0914_
rlabel metal1 24794 9690 24794 9690 0 _0915_
rlabel metal1 25760 10234 25760 10234 0 _0916_
rlabel metal1 25760 9418 25760 9418 0 _0917_
rlabel metal1 26266 11186 26266 11186 0 _0918_
rlabel metal1 26450 10778 26450 10778 0 _0919_
rlabel metal1 26772 9418 26772 9418 0 _0920_
rlabel metal1 29716 20434 29716 20434 0 _0921_
rlabel metal1 31602 25840 31602 25840 0 _0922_
rlabel metal1 27968 10982 27968 10982 0 _0923_
rlabel metal1 25760 9350 25760 9350 0 _0924_
rlabel metal1 28290 10234 28290 10234 0 _0925_
rlabel metal1 28934 10608 28934 10608 0 _0926_
rlabel metal1 28152 10506 28152 10506 0 _0927_
rlabel metal1 27784 10778 27784 10778 0 _0928_
rlabel metal1 29762 19720 29762 19720 0 _0929_
rlabel metal1 29394 10234 29394 10234 0 _0930_
rlabel metal2 29854 10948 29854 10948 0 _0931_
rlabel metal1 30084 11186 30084 11186 0 _0932_
rlabel metal1 29532 19822 29532 19822 0 _0933_
rlabel metal2 30728 24106 30728 24106 0 _0934_
rlabel metal1 31786 29648 31786 29648 0 _0935_
rlabel metal1 31700 33490 31700 33490 0 _0936_
rlabel metal1 36018 30702 36018 30702 0 _0937_
rlabel metal1 35374 29138 35374 29138 0 _0938_
rlabel metal1 22448 6290 22448 6290 0 _0939_
rlabel metal2 22126 6579 22126 6579 0 _0940_
rlabel metal1 22310 6358 22310 6358 0 _0941_
rlabel metal1 22218 6358 22218 6358 0 _0942_
rlabel metal1 22816 6086 22816 6086 0 _0943_
rlabel metal1 23322 6324 23322 6324 0 _0944_
rlabel metal2 23230 6902 23230 6902 0 _0945_
rlabel metal2 23506 6647 23506 6647 0 _0946_
rlabel metal2 28750 24446 28750 24446 0 _0947_
rlabel metal2 22494 9622 22494 9622 0 _0948_
rlabel metal1 22862 8942 22862 8942 0 _0949_
rlabel metal1 21666 8398 21666 8398 0 _0950_
rlabel metal1 21620 8874 21620 8874 0 _0951_
rlabel metal1 22586 9044 22586 9044 0 _0952_
rlabel metal1 22448 8602 22448 8602 0 _0953_
rlabel metal1 22770 8806 22770 8806 0 _0954_
rlabel metal2 22126 10591 22126 10591 0 _0955_
rlabel metal1 23506 8058 23506 8058 0 _0956_
rlabel metal1 23046 8500 23046 8500 0 _0957_
rlabel metal1 22632 8602 22632 8602 0 _0958_
rlabel metal1 24932 24786 24932 24786 0 _0959_
rlabel metal1 27278 24820 27278 24820 0 _0960_
rlabel metal1 20056 15062 20056 15062 0 _0961_
rlabel metal1 18308 14586 18308 14586 0 _0962_
rlabel metal1 20010 14960 20010 14960 0 _0963_
rlabel metal1 20102 14960 20102 14960 0 _0964_
rlabel metal2 19642 15164 19642 15164 0 _0965_
rlabel metal1 20010 15130 20010 15130 0 _0966_
rlabel metal1 20194 15980 20194 15980 0 _0967_
rlabel metal1 19826 15572 19826 15572 0 _0968_
rlabel metal2 19734 23766 19734 23766 0 _0969_
rlabel metal2 25806 25976 25806 25976 0 _0970_
rlabel metal1 22264 15674 22264 15674 0 _0971_
rlabel metal1 22126 14382 22126 14382 0 _0972_
rlabel metal1 20608 14042 20608 14042 0 _0973_
rlabel metal1 21850 13974 21850 13974 0 _0974_
rlabel metal1 21896 14042 21896 14042 0 _0975_
rlabel metal1 21666 14314 21666 14314 0 _0976_
rlabel metal1 22172 14246 22172 14246 0 _0977_
rlabel metal1 22494 16218 22494 16218 0 _0978_
rlabel metal1 20700 15470 20700 15470 0 _0979_
rlabel metal1 21712 15674 21712 15674 0 _0980_
rlabel metal1 22356 18394 22356 18394 0 _0981_
rlabel metal1 22862 18802 22862 18802 0 _0982_
rlabel metal1 28014 30668 28014 30668 0 _0983_
rlabel metal1 29394 29036 29394 29036 0 _0984_
rlabel metal1 29578 29138 29578 29138 0 _0985_
rlabel metal1 25806 27030 25806 27030 0 _0986_
rlabel metal1 25898 27098 25898 27098 0 _0987_
rlabel metal1 26726 28186 26726 28186 0 _0988_
rlabel metal1 30222 29036 30222 29036 0 _0989_
rlabel metal1 28060 28730 28060 28730 0 _0990_
rlabel viali 22214 32888 22214 32888 0 _0991_
rlabel metal1 23782 32368 23782 32368 0 _0992_
rlabel metal1 23230 32436 23230 32436 0 _0993_
rlabel metal1 20424 32402 20424 32402 0 _0994_
rlabel metal1 19136 30702 19136 30702 0 _0995_
rlabel metal1 19780 30906 19780 30906 0 _0996_
rlabel metal1 18998 32810 18998 32810 0 _0997_
rlabel metal1 18722 33456 18722 33456 0 _0998_
rlabel metal1 17710 32810 17710 32810 0 _0999_
rlabel metal1 17158 33014 17158 33014 0 _1000_
rlabel metal1 18170 13362 18170 13362 0 _1001_
rlabel metal1 18078 13498 18078 13498 0 _1002_
rlabel metal2 17526 14569 17526 14569 0 _1003_
rlabel metal1 12926 12954 12926 12954 0 _1004_
rlabel metal2 12374 13702 12374 13702 0 _1005_
rlabel metal1 11868 14042 11868 14042 0 _1006_
rlabel metal1 13202 31314 13202 31314 0 _1007_
rlabel metal1 14352 31450 14352 31450 0 _1008_
rlabel metal1 13984 30906 13984 30906 0 _1009_
rlabel metal2 14122 31518 14122 31518 0 _1010_
rlabel metal1 15594 31280 15594 31280 0 _1011_
rlabel metal1 20884 10234 20884 10234 0 _1012_
rlabel metal2 20930 10914 20930 10914 0 _1013_
rlabel metal1 15134 32946 15134 32946 0 _1014_
rlabel metal1 23230 10234 23230 10234 0 _1015_
rlabel metal2 23322 10948 23322 10948 0 _1016_
rlabel metal1 13202 32810 13202 32810 0 _1017_
rlabel metal1 14950 32912 14950 32912 0 _1018_
rlabel metal1 14858 32844 14858 32844 0 _1019_
rlabel metal1 14628 32810 14628 32810 0 _1020_
rlabel metal1 15226 33626 15226 33626 0 _1021_
rlabel metal2 15962 33184 15962 33184 0 _1022_
rlabel metal1 14421 31314 14421 31314 0 _1023_
rlabel metal1 16744 31314 16744 31314 0 _1024_
rlabel metal1 16928 29614 16928 29614 0 _1025_
rlabel metal2 18170 29444 18170 29444 0 _1026_
rlabel metal1 20746 8398 20746 8398 0 _1027_
rlabel metal1 20194 8602 20194 8602 0 _1028_
rlabel metal2 19918 26877 19918 26877 0 _1029_
rlabel metal1 19918 7956 19918 7956 0 _1030_
rlabel metal1 20470 8058 20470 8058 0 _1031_
rlabel via2 21022 9163 21022 9163 0 _1032_
rlabel metal1 19458 27404 19458 27404 0 _1033_
rlabel metal1 20240 28526 20240 28526 0 _1034_
rlabel metal1 19826 28016 19826 28016 0 _1035_
rlabel metal2 19918 28356 19918 28356 0 _1036_
rlabel metal1 18170 28084 18170 28084 0 _1037_
rlabel metal1 18906 27982 18906 27982 0 _1038_
rlabel metal1 15821 21522 15821 21522 0 _1039_
rlabel metal1 14076 21046 14076 21046 0 _1040_
rlabel viali 14490 21522 14490 21522 0 _1041_
rlabel metal1 16146 21556 16146 21556 0 _1042_
rlabel metal1 16468 32946 16468 32946 0 _1043_
rlabel via2 12006 21947 12006 21947 0 _1044_
rlabel metal1 22862 21964 22862 21964 0 _1045_
rlabel metal1 22724 21522 22724 21522 0 _1046_
rlabel metal1 23460 21454 23460 21454 0 _1047_
rlabel metal1 23874 21522 23874 21522 0 _1048_
rlabel metal2 20102 32878 20102 32878 0 _1049_
rlabel metal2 33902 22831 33902 22831 0 _1050_
rlabel metal2 18538 28730 18538 28730 0 _1051_
rlabel metal1 18446 31858 18446 31858 0 _1052_
rlabel metal1 22586 32436 22586 32436 0 _1053_
rlabel metal2 22494 31586 22494 31586 0 _1054_
rlabel metal1 23920 31858 23920 31858 0 _1055_
rlabel metal1 32706 27846 32706 27846 0 _1056_
rlabel metal2 36938 23936 36938 23936 0 _1057_
rlabel metal1 33626 20366 33626 20366 0 _1058_
rlabel metal1 33718 20298 33718 20298 0 _1059_
rlabel metal1 33856 20570 33856 20570 0 _1060_
rlabel metal1 33028 26010 33028 26010 0 _1061_
rlabel metal1 33902 24922 33902 24922 0 _1062_
rlabel metal2 33074 26996 33074 26996 0 _1063_
rlabel metal1 32154 29206 32154 29206 0 _1064_
rlabel metal1 28481 29173 28481 29173 0 _1065_
rlabel metal1 26864 26350 26864 26350 0 _1066_
rlabel metal1 26680 25670 26680 25670 0 _1067_
rlabel metal1 26634 24106 26634 24106 0 _1068_
rlabel metal1 26634 26996 26634 26996 0 _1069_
rlabel metal1 27186 28118 27186 28118 0 _1070_
rlabel metal1 30268 27370 30268 27370 0 _1071_
rlabel metal1 30452 20366 30452 20366 0 _1072_
rlabel metal1 30590 26928 30590 26928 0 _1073_
rlabel metal1 29440 27506 29440 27506 0 _1074_
rlabel metal1 27232 26962 27232 26962 0 _1075_
rlabel metal1 27094 26928 27094 26928 0 _1076_
rlabel metal1 27554 27098 27554 27098 0 _1077_
rlabel metal1 28014 29036 28014 29036 0 _1078_
rlabel metal2 27922 30532 27922 30532 0 _1079_
rlabel metal1 22862 31790 22862 31790 0 _1080_
rlabel metal1 21758 31790 21758 31790 0 _1081_
rlabel metal1 20654 32742 20654 32742 0 _1082_
rlabel metal1 18906 31246 18906 31246 0 _1083_
rlabel metal1 18768 31790 18768 31790 0 _1084_
rlabel metal1 16238 31824 16238 31824 0 _1085_
rlabel metal1 14720 31790 14720 31790 0 _1086_
rlabel metal1 16422 30668 16422 30668 0 _1087_
rlabel metal1 16008 29682 16008 29682 0 _1088_
rlabel metal2 17158 28492 17158 28492 0 _1089_
rlabel metal1 17710 28186 17710 28186 0 _1090_
rlabel metal1 24564 21658 24564 21658 0 _1091_
rlabel metal1 17020 33490 17020 33490 0 _1092_
rlabel metal1 18262 28526 18262 28526 0 _1093_
rlabel metal1 17480 28526 17480 28526 0 _1094_
rlabel metal1 27002 32878 27002 32878 0 _1095_
rlabel metal1 26404 33422 26404 33422 0 _1096_
rlabel metal2 26542 33286 26542 33286 0 _1097_
rlabel metal1 26542 34034 26542 34034 0 _1098_
rlabel metal1 26312 30906 26312 30906 0 _1099_
rlabel metal1 29624 34578 29624 34578 0 _1100_
rlabel metal1 29946 34646 29946 34646 0 _1101_
rlabel metal1 30130 34544 30130 34544 0 _1102_
rlabel metal1 30176 34034 30176 34034 0 _1103_
rlabel metal1 35972 28730 35972 28730 0 _1104_
rlabel metal1 35190 32742 35190 32742 0 _1105_
rlabel metal1 37168 26350 37168 26350 0 _1106_
rlabel metal1 36708 20026 36708 20026 0 _1107_
rlabel metal1 35098 19346 35098 19346 0 _1108_
rlabel metal1 30682 19754 30682 19754 0 _1109_
rlabel metal1 35558 19924 35558 19924 0 _1110_
rlabel metal1 36662 23664 36662 23664 0 _1111_
rlabel metal1 36708 26350 36708 26350 0 _1112_
rlabel metal1 34040 26418 34040 26418 0 _1113_
rlabel via1 36570 27098 36570 27098 0 _1114_
rlabel metal1 36294 30906 36294 30906 0 _1115_
rlabel metal1 34914 32980 34914 32980 0 _1116_
rlabel metal1 34132 32878 34132 32878 0 _1117_
rlabel metal1 33258 32878 33258 32878 0 _1118_
rlabel metal1 31096 33966 31096 33966 0 _1119_
rlabel metal1 29808 33490 29808 33490 0 _1120_
rlabel metal1 26956 33898 26956 33898 0 _1121_
rlabel metal2 25806 22508 25806 22508 0 _1122_
rlabel metal1 31786 20978 31786 20978 0 _1123_
rlabel metal1 34776 22066 34776 22066 0 _1124_
rlabel metal1 26642 33830 26642 33830 0 _1125_
rlabel metal1 27186 33490 27186 33490 0 _1126_
rlabel metal1 31786 28560 31786 28560 0 _1127_
rlabel metal1 29026 30702 29026 30702 0 _1128_
rlabel metal1 27692 31450 27692 31450 0 _1129_
rlabel metal2 28198 33252 28198 33252 0 _1130_
rlabel metal1 29072 30770 29072 30770 0 _1131_
rlabel metal1 32062 31892 32062 31892 0 _1132_
rlabel metal1 31648 28730 31648 28730 0 _1133_
rlabel metal1 33856 31790 33856 31790 0 _1134_
rlabel metal1 32706 29138 32706 29138 0 _1135_
rlabel metal1 33810 29070 33810 29070 0 _1136_
rlabel metal1 35282 24072 35282 24072 0 _1137_
rlabel metal1 34592 19414 34592 19414 0 _1138_
rlabel metal1 34086 20978 34086 20978 0 _1139_
rlabel metal1 30314 20944 30314 20944 0 _1140_
rlabel metal1 31050 20842 31050 20842 0 _1141_
rlabel metal1 34960 21658 34960 21658 0 _1142_
rlabel metal1 34684 24174 34684 24174 0 _1143_
rlabel metal2 34270 25432 34270 25432 0 _1144_
rlabel metal1 35466 27030 35466 27030 0 _1145_
rlabel metal1 34086 26928 34086 26928 0 _1146_
rlabel metal2 33718 32606 33718 32606 0 _1147_
rlabel metal1 29256 32946 29256 32946 0 _1148_
rlabel metal2 28106 32572 28106 32572 0 _1149_
rlabel metal1 16606 20910 16606 20910 0 _1150_
rlabel metal1 16744 20842 16744 20842 0 _1151_
rlabel metal1 27370 33524 27370 33524 0 _1152_
rlabel metal1 26818 29614 26818 29614 0 _1153_
rlabel metal2 31050 30532 31050 30532 0 _1154_
rlabel metal1 27922 30736 27922 30736 0 _1155_
rlabel metal1 27140 30226 27140 30226 0 _1156_
rlabel metal1 26174 29070 26174 29070 0 _1157_
rlabel metal1 26588 29274 26588 29274 0 _1158_
rlabel via1 25814 21658 25814 21658 0 _1159_
rlabel metal2 28290 22304 28290 22304 0 _1160_
rlabel metal2 33810 26639 33810 26639 0 _1161_
rlabel metal1 30912 21930 30912 21930 0 _1162_
rlabel metal1 26358 22678 26358 22678 0 _1163_
rlabel metal1 27278 23086 27278 23086 0 _1164_
rlabel metal1 26634 26316 26634 26316 0 _1165_
rlabel metal2 35190 22039 35190 22039 0 _1166_
rlabel metal2 27646 23664 27646 23664 0 _1167_
rlabel metal2 26634 21869 26634 21869 0 _1168_
rlabel metal1 27646 24242 27646 24242 0 _1169_
rlabel metal1 27278 24378 27278 24378 0 _1170_
rlabel metal1 27324 20910 27324 20910 0 _1171_
rlabel metal1 27416 20774 27416 20774 0 _1172_
rlabel metal1 29210 24208 29210 24208 0 _1173_
rlabel metal1 29072 24378 29072 24378 0 _1174_
rlabel metal1 32016 24174 32016 24174 0 _1175_
rlabel metal1 27922 24684 27922 24684 0 _1176_
rlabel metal2 28198 24548 28198 24548 0 _1177_
rlabel metal1 27646 24378 27646 24378 0 _1178_
rlabel metal2 27002 26656 27002 26656 0 _1179_
rlabel metal1 27324 28730 27324 28730 0 _1180_
rlabel metal2 27554 32419 27554 32419 0 _1181_
rlabel metal1 16146 37400 16146 37400 0 _1182_
rlabel metal1 17020 26486 17020 26486 0 _1183_
rlabel metal2 17618 3689 17618 3689 0 _1184_
rlabel metal1 10235 16558 10235 16558 0 _1185_
rlabel metal2 10626 16320 10626 16320 0 _1186_
rlabel metal1 10304 16490 10304 16490 0 _1187_
rlabel metal1 10074 15504 10074 15504 0 _1188_
rlabel metal2 10258 17612 10258 17612 0 _1189_
rlabel metal2 9798 16558 9798 16558 0 _1190_
rlabel metal2 9798 15776 9798 15776 0 _1191_
rlabel metal1 10902 11730 10902 11730 0 _1192_
rlabel metal1 9982 15402 9982 15402 0 _1193_
rlabel metal1 9246 21658 9246 21658 0 _1194_
rlabel metal1 9568 21862 9568 21862 0 _1195_
rlabel metal1 10442 21420 10442 21420 0 _1196_
rlabel metal2 9798 21012 9798 21012 0 _1197_
rlabel metal1 9706 21556 9706 21556 0 _1198_
rlabel metal2 10718 21590 10718 21590 0 _1199_
rlabel metal1 10074 20910 10074 20910 0 _1200_
rlabel via1 12558 20315 12558 20315 0 _1201_
rlabel metal2 9890 13668 9890 13668 0 _1202_
rlabel metal2 18814 3519 18814 3519 0 _1203_
rlabel metal1 18170 3570 18170 3570 0 _1204_
rlabel metal1 30268 33490 30268 33490 0 _1205_
rlabel metal1 29762 32946 29762 32946 0 _1206_
rlabel metal1 35236 32334 35236 32334 0 _1207_
rlabel metal1 29724 32538 29724 32538 0 _1208_
rlabel metal2 30038 32810 30038 32810 0 _1209_
rlabel metal2 32522 31178 32522 31178 0 _1210_
rlabel metal1 27692 30294 27692 30294 0 _1211_
rlabel metal1 28290 30362 28290 30362 0 _1212_
rlabel metal1 32430 31212 32430 31212 0 _1213_
rlabel via1 28934 24157 28934 24157 0 _1214_
rlabel metal1 27094 26384 27094 26384 0 _1215_
rlabel metal1 27876 26554 27876 26554 0 _1216_
rlabel metal1 27922 26486 27922 26486 0 _1217_
rlabel metal2 28382 29206 28382 29206 0 _1218_
rlabel metal1 29624 31450 29624 31450 0 _1219_
rlabel metal1 29440 33082 29440 33082 0 _1220_
rlabel metal1 18722 24786 18722 24786 0 _1221_
rlabel metal1 15410 29750 15410 29750 0 _1222_
rlabel metal1 15594 29682 15594 29682 0 _1223_
rlabel metal1 15410 27574 15410 27574 0 _1224_
rlabel metal2 8050 14688 8050 14688 0 _1225_
rlabel metal1 5934 16082 5934 16082 0 _1226_
rlabel metal1 34684 30906 34684 30906 0 _1227_
rlabel metal1 34224 32402 34224 32402 0 _1228_
rlabel metal1 32476 31314 32476 31314 0 _1229_
rlabel metal1 29302 26962 29302 26962 0 _1230_
rlabel metal1 30406 26996 30406 26996 0 _1231_
rlabel metal1 30176 26010 30176 26010 0 _1232_
rlabel metal1 31947 31314 31947 31314 0 _1233_
rlabel metal1 33166 31450 33166 31450 0 _1234_
rlabel metal1 32936 32198 32936 32198 0 _1235_
rlabel metal1 35282 32878 35282 32878 0 _1236_
rlabel metal1 33442 32912 33442 32912 0 _1237_
rlabel metal1 33258 32436 33258 32436 0 _1238_
rlabel metal2 17986 25619 17986 25619 0 _1239_
rlabel metal1 15962 31824 15962 31824 0 _1240_
rlabel metal1 16238 31382 16238 31382 0 _1241_
rlabel metal1 15778 32912 15778 32912 0 _1242_
rlabel metal2 15962 32241 15962 32241 0 _1243_
rlabel metal2 16606 30940 16606 30940 0 _1244_
rlabel metal1 16790 30770 16790 30770 0 _1245_
rlabel metal1 14306 29546 14306 29546 0 _1246_
rlabel metal2 6992 14892 6992 14892 0 _1247_
rlabel metal1 4830 13158 4830 13158 0 _1248_
rlabel metal1 34546 31382 34546 31382 0 _1249_
rlabel metal1 36432 28730 36432 28730 0 _1250_
rlabel metal1 35834 29206 35834 29206 0 _1251_
rlabel metal1 34086 29580 34086 29580 0 _1252_
rlabel metal1 32706 25126 32706 25126 0 _1253_
rlabel metal1 32729 22610 32729 22610 0 _1254_
rlabel metal1 29854 21556 29854 21556 0 _1255_
rlabel metal1 32016 24038 32016 24038 0 _1256_
rlabel metal1 32430 29104 32430 29104 0 _1257_
rlabel metal1 32154 25908 32154 25908 0 _1258_
rlabel metal1 32844 25942 32844 25942 0 _1259_
rlabel metal1 31326 24378 31326 24378 0 _1260_
rlabel metal1 31970 27098 31970 27098 0 _1261_
rlabel metal1 33304 28186 33304 28186 0 _1262_
rlabel metal1 34500 29818 34500 29818 0 _1263_
rlabel metal1 35052 31314 35052 31314 0 _1264_
rlabel metal1 21574 24072 21574 24072 0 _1265_
rlabel metal2 16054 33286 16054 33286 0 _1266_
rlabel metal1 16146 33524 16146 33524 0 _1267_
rlabel metal2 15686 33762 15686 33762 0 _1268_
rlabel metal2 15594 3162 15594 3162 0 _1269_
rlabel metal1 10258 3026 10258 3026 0 _1270_
rlabel metal1 36984 26962 36984 26962 0 _1271_
rlabel metal1 36478 26962 36478 26962 0 _1272_
rlabel metal1 35098 26962 35098 26962 0 _1273_
rlabel metal1 34431 26962 34431 26962 0 _1274_
rlabel metal1 36800 27642 36800 27642 0 _1275_
rlabel metal2 2622 39076 2622 39076 0 clk
rlabel metal1 14858 9350 14858 9350 0 clknet_0__0514_
rlabel metal1 23506 12614 23506 12614 0 clknet_0__0515_
rlabel metal1 20930 7412 20930 7412 0 clknet_0__0516_
rlabel metal2 19182 9214 19182 9214 0 clknet_0__0517_
rlabel metal1 12742 33422 12742 33422 0 clknet_0_clk
rlabel metal2 4002 14382 4002 14382 0 clknet_1_0__leaf__0514_
rlabel metal1 19412 18734 19412 18734 0 clknet_1_0__leaf__0515_
rlabel metal1 14674 3978 14674 3978 0 clknet_1_0__leaf__0516_
rlabel metal1 17020 4590 17020 4590 0 clknet_1_0__leaf__0517_
rlabel metal1 9062 3468 9062 3468 0 clknet_1_1__leaf__0514_
rlabel metal1 32154 7854 32154 7854 0 clknet_1_1__leaf__0515_
rlabel metal1 32246 13362 32246 13362 0 clknet_1_1__leaf__0516_
rlabel metal1 31786 5236 31786 5236 0 clknet_1_1__leaf__0517_
rlabel metal2 1426 22032 1426 22032 0 clknet_2_0__leaf_clk
rlabel metal2 2162 26758 2162 26758 0 clknet_2_1__leaf_clk
rlabel metal1 4784 31858 4784 31858 0 clknet_2_2__leaf_clk
rlabel metal2 14214 34612 14214 34612 0 clknet_2_3__leaf_clk
rlabel metal2 30958 1027 30958 1027 0 cs
rlabel metal3 820 34748 820 34748 0 gpi[0]
rlabel metal2 37398 1299 37398 1299 0 gpi[1]
rlabel metal2 12926 1027 12926 1027 0 gpi[23]
rlabel metal1 38134 32878 38134 32878 0 gpi[2]
rlabel metal3 820 18428 820 18428 0 gpi[3]
rlabel metal3 820 4148 820 4148 0 gpi[4]
rlabel metal2 35466 1571 35466 1571 0 gpi[5]
rlabel metal1 20838 38998 20838 38998 0 gpi[6]
rlabel metal1 37536 38998 37536 38998 0 gpi[7]
rlabel metal1 37720 2278 37720 2278 0 gpo[0]
rlabel via2 37858 11611 37858 11611 0 gpo[10]
rlabel metal2 24518 1520 24518 1520 0 gpo[11]
rlabel metal1 38088 14586 38088 14586 0 gpo[12]
rlabel metal1 25300 39066 25300 39066 0 gpo[13]
rlabel metal2 27370 39967 27370 39967 0 gpo[14]
rlabel metal1 1104 39066 1104 39066 0 gpo[15]
rlabel metal2 46 1554 46 1554 0 gpo[16]
rlabel metal3 820 25908 820 25908 0 gpo[17]
rlabel metal1 23368 39066 23368 39066 0 gpo[18]
rlabel via1 31878 39083 31878 39083 0 gpo[19]
rlabel metal2 37858 37553 37858 37553 0 gpo[1]
rlabel metal1 14398 39066 14398 39066 0 gpo[20]
rlabel metal2 3910 959 3910 959 0 gpo[21]
rlabel metal2 1978 959 1978 959 0 gpo[22]
rlabel metal3 912 39508 912 39508 0 gpo[23]
rlabel metal2 36386 39967 36386 39967 0 gpo[24]
rlabel metal2 15502 1554 15502 1554 0 gpo[25]
rlabel via2 37858 35445 37858 35445 0 gpo[26]
rlabel metal3 38326 68 38326 68 0 gpo[27]
rlabel metal3 820 11628 820 11628 0 gpo[28]
rlabel metal3 1096 2108 1096 2108 0 gpo[29]
rlabel metal2 6486 959 6486 959 0 gpo[2]
rlabel metal2 10994 1095 10994 1095 0 gpo[30]
rlabel metal3 820 21148 820 21148 0 gpo[31]
rlabel metal2 37858 21233 37858 21233 0 gpo[32]
rlabel metal2 20010 823 20010 823 0 gpo[33]
rlabel metal3 820 16388 820 16388 0 gpo[3]
rlabel metal1 34546 39066 34546 39066 0 gpo[4]
rlabel metal1 5336 39066 5336 39066 0 gpo[5]
rlabel metal1 9844 39066 9844 39066 0 gpo[6]
rlabel metal2 26450 1520 26450 1520 0 gpo[7]
rlabel metal3 1096 13668 1096 13668 0 gpo[8]
rlabel metal3 820 37468 820 37468 0 gpo[9]
rlabel metal1 31188 2482 31188 2482 0 net1
rlabel metal1 36294 38964 36294 38964 0 net10
rlabel metal1 30958 10030 30958 10030 0 net100
rlabel metal1 32154 12852 32154 12852 0 net101
rlabel metal2 19688 12750 19688 12750 0 net102
rlabel metal1 21850 3060 21850 3060 0 net103
rlabel metal1 22586 14042 22586 14042 0 net104
rlabel metal1 27002 3060 27002 3060 0 net105
rlabel metal1 6394 9588 6394 9588 0 net106
rlabel metal1 6946 7854 6946 7854 0 net107
rlabel metal1 11914 3638 11914 3638 0 net108
rlabel metal1 6670 5746 6670 5746 0 net109
rlabel metal1 36478 17238 36478 17238 0 net11
rlabel metal1 6670 13294 6670 13294 0 net110
rlabel metal2 16698 4250 16698 4250 0 net111
rlabel metal2 33350 15130 33350 15130 0 net112
rlabel metal1 31602 5338 31602 5338 0 net113
rlabel metal1 9614 9588 9614 9588 0 net114
rlabel metal2 14766 5610 14766 5610 0 net115
rlabel metal1 32798 8602 32798 8602 0 net116
rlabel metal1 35098 11798 35098 11798 0 net117
rlabel metal1 14766 13940 14766 13940 0 net118
rlabel metal1 21022 4658 21022 4658 0 net119
rlabel metal1 37352 2414 37352 2414 0 net12
rlabel metal1 30958 15130 30958 15130 0 net120
rlabel metal2 27830 4522 27830 4522 0 net121
rlabel metal1 6670 11118 6670 11118 0 net122
rlabel metal1 5382 6766 5382 6766 0 net123
rlabel metal1 10304 5746 10304 5746 0 net124
rlabel metal1 5106 12206 5106 12206 0 net125
rlabel metal1 4738 14042 4738 14042 0 net126
rlabel metal1 18998 5236 18998 5236 0 net127
rlabel metal1 30590 16558 30590 16558 0 net128
rlabel metal1 4140 30022 4140 30022 0 net129
rlabel metal2 37674 12019 37674 12019 0 net13
rlabel metal1 5106 31450 5106 31450 0 net130
rlabel metal1 3542 30804 3542 30804 0 net131
rlabel metal1 3450 26316 3450 26316 0 net132
rlabel metal1 4508 28526 4508 28526 0 net133
rlabel metal1 3358 24922 3358 24922 0 net134
rlabel metal1 2254 23596 2254 23596 0 net135
rlabel metal1 4968 23630 4968 23630 0 net136
rlabel metal1 29026 17680 29026 17680 0 net137
rlabel metal1 29670 9520 29670 9520 0 net138
rlabel metal1 29578 11764 29578 11764 0 net139
rlabel via3 24725 2652 24725 2652 0 net14
rlabel metal1 5152 30294 5152 30294 0 net140
rlabel metal1 14030 8058 14030 8058 0 net141
rlabel metal1 20010 18326 20010 18326 0 net142
rlabel metal2 20746 16626 20746 16626 0 net143
rlabel metal2 37628 18292 37628 18292 0 net15
rlabel metal2 25254 38454 25254 38454 0 net16
rlabel metal1 26956 37978 26956 37978 0 net17
rlabel metal2 1794 38284 1794 38284 0 net18
rlabel metal1 1886 2414 1886 2414 0 net19
rlabel metal1 13570 24072 13570 24072 0 net2
rlabel metal2 1794 26894 1794 26894 0 net20
rlabel metal2 23414 37094 23414 37094 0 net21
rlabel metal2 14858 37604 14858 37604 0 net22
rlabel metal1 37628 36890 37628 36890 0 net23
rlabel metal2 14766 36550 14766 36550 0 net24
rlabel metal1 4370 2448 4370 2448 0 net25
rlabel metal1 2438 2516 2438 2516 0 net26
rlabel metal1 2024 38522 2024 38522 0 net27
rlabel metal1 36202 38862 36202 38862 0 net28
rlabel metal1 16629 2278 16629 2278 0 net29
rlabel metal3 26611 8092 26611 8092 0 net3
rlabel metal1 37628 35258 37628 35258 0 net30
rlabel metal1 34730 3094 34730 3094 0 net31
rlabel metal1 1794 11832 1794 11832 0 net32
rlabel metal2 1794 4046 1794 4046 0 net33
rlabel metal1 6900 2822 6900 2822 0 net34
rlabel metal1 11362 2346 11362 2346 0 net35
rlabel metal2 1794 18326 1794 18326 0 net36
rlabel metal1 37628 18938 37628 18938 0 net37
rlabel metal1 20102 2346 20102 2346 0 net38
rlabel metal1 1794 16184 1794 16184 0 net39
rlabel metal2 12374 23970 12374 23970 0 net4
rlabel metal2 33626 37910 33626 37910 0 net40
rlabel metal1 10580 38522 10580 38522 0 net41
rlabel metal1 10212 37978 10212 37978 0 net42
rlabel metal1 26910 2414 26910 2414 0 net43
rlabel metal2 6486 16048 6486 16048 0 net44
rlabel metal2 20010 37570 20010 37570 0 net45
rlabel metal2 21298 36788 21298 36788 0 net46
rlabel metal2 12466 10608 12466 10608 0 net47
rlabel metal1 19826 3536 19826 3536 0 net48
rlabel metal1 29578 22039 29578 22039 0 net49
rlabel metal1 33350 32300 33350 32300 0 net5
rlabel via1 19813 14994 19813 14994 0 net50
rlabel metal1 21873 17782 21873 17782 0 net51
rlabel metal1 25714 7276 25714 7276 0 net52
rlabel metal1 18170 8432 18170 8432 0 net53
rlabel metal1 22954 8024 22954 8024 0 net54
rlabel metal1 16146 11832 16146 11832 0 net55
rlabel metal1 15594 14994 15594 14994 0 net56
rlabel metal1 21850 18054 21850 18054 0 net57
rlabel metal1 13754 11662 13754 11662 0 net58
rlabel metal2 18354 19584 18354 19584 0 net59
rlabel metal1 1702 18870 1702 18870 0 net6
rlabel metal1 21206 2985 21206 2985 0 net60
rlabel metal1 33771 12818 33771 12818 0 net61
rlabel metal1 12505 25262 12505 25262 0 net62
rlabel metal1 15785 35734 15785 35734 0 net63
rlabel metal2 19090 19618 19090 19618 0 net64
rlabel metal1 23874 3060 23874 3060 0 net65
rlabel metal1 4278 10030 4278 10030 0 net66
rlabel metal1 4186 8500 4186 8500 0 net67
rlabel metal1 9246 3502 9246 3502 0 net68
rlabel metal1 3542 12852 3542 12852 0 net69
rlabel metal2 20746 24497 20746 24497 0 net7
rlabel metal1 4646 15470 4646 15470 0 net70
rlabel metal1 17158 3026 17158 3026 0 net71
rlabel metal1 25346 19482 25346 19482 0 net72
rlabel metal1 28750 18292 28750 18292 0 net73
rlabel metal1 17066 19380 17066 19380 0 net74
rlabel metal1 12282 7514 12282 7514 0 net75
rlabel metal1 30314 8602 30314 8602 0 net76
rlabel metal1 29946 12206 29946 12206 0 net77
rlabel metal1 19642 18734 19642 18734 0 net78
rlabel metal1 21896 19890 21896 19890 0 net79
rlabel metal2 35742 2329 35742 2329 0 net8
rlabel metal1 32798 16218 32798 16218 0 net80
rlabel metal1 32154 7412 32154 7412 0 net81
rlabel metal1 12006 9588 12006 9588 0 net82
rlabel metal2 12834 5338 12834 5338 0 net83
rlabel metal2 35098 9690 35098 9690 0 net84
rlabel metal1 35420 13906 35420 13906 0 net85
rlabel metal1 13018 12852 13018 12852 0 net86
rlabel metal1 24288 4658 24288 4658 0 net87
rlabel metal1 26818 17714 26818 17714 0 net88
rlabel via1 27462 4573 27462 4573 0 net89
rlabel metal2 13984 35700 13984 35700 0 net9
rlabel metal1 8970 9996 8970 9996 0 net90
rlabel metal1 9154 7412 9154 7412 0 net91
rlabel metal1 14582 3060 14582 3060 0 net92
rlabel metal2 8694 5610 8694 5610 0 net93
rlabel metal2 7222 15130 7222 15130 0 net94
rlabel metal1 19826 3094 19826 3094 0 net95
rlabel metal1 31050 14382 31050 14382 0 net96
rlabel metal1 29762 5338 29762 5338 0 net97
rlabel metal2 12466 11934 12466 11934 0 net98
rlabel metal1 11638 6324 11638 6324 0 net99
rlabel metal1 38134 19346 38134 19346 0 nrst
<< properties >>
string FIXED_BBOX 0 0 39421 41565
<< end >>
