// This is the unpowered netlist.
module stopwatch (clk,
    nrst,
    pb_0,
    pb_1,
    time_done,
    out_0,
    out_1,
    out_2,
    out_3);
 input clk;
 input nrst;
 input pb_0;
 input pb_1;
 output time_done;
 output [6:0] out_0;
 output [6:0] out_1;
 output [6:0] out_2;
 output [6:0] out_3;

 wire \CLKDIV.count[0] ;
 wire \CLKDIV.count[10] ;
 wire \CLKDIV.count[11] ;
 wire \CLKDIV.count[12] ;
 wire \CLKDIV.count[13] ;
 wire \CLKDIV.count[14] ;
 wire \CLKDIV.count[15] ;
 wire \CLKDIV.count[16] ;
 wire \CLKDIV.count[17] ;
 wire \CLKDIV.count[18] ;
 wire \CLKDIV.count[19] ;
 wire \CLKDIV.count[1] ;
 wire \CLKDIV.count[20] ;
 wire \CLKDIV.count[21] ;
 wire \CLKDIV.count[22] ;
 wire \CLKDIV.count[23] ;
 wire \CLKDIV.count[2] ;
 wire \CLKDIV.count[3] ;
 wire \CLKDIV.count[4] ;
 wire \CLKDIV.count[5] ;
 wire \CLKDIV.count[6] ;
 wire \CLKDIV.count[7] ;
 wire \CLKDIV.count[8] ;
 wire \CLKDIV.count[9] ;
 wire \CLKDIV.secpulse ;
 wire \CTR.minutes ;
 wire \CTR.time_out[0] ;
 wire \CTR.time_out[10] ;
 wire \CTR.time_out[11] ;
 wire \CTR.time_out[1] ;
 wire \CTR.time_out[2] ;
 wire \CTR.time_out[3] ;
 wire \CTR.time_out[4] ;
 wire \CTR.time_out[5] ;
 wire \CTR.time_out[6] ;
 wire \CTR.time_out[7] ;
 wire \CTR.time_out[8] ;
 wire \CTR.time_out[9] ;
 wire \FSM.next_state[0] ;
 wire \FSM.next_state[1] ;
 wire \FSM.next_state[2] ;
 wire \FSM.next_state[3] ;
 wire \FSM.state[0] ;
 wire \FSM.state[1] ;
 wire \FSM.state[2] ;
 wire \FSM.state[3] ;
 wire \MEM.addr[0] ;
 wire \MEM.addr[1] ;
 wire \MEM.addr[2] ;
 wire \MEM.mem1[0] ;
 wire \MEM.mem1[10] ;
 wire \MEM.mem1[11] ;
 wire \MEM.mem1[1] ;
 wire \MEM.mem1[2] ;
 wire \MEM.mem1[3] ;
 wire \MEM.mem1[4] ;
 wire \MEM.mem1[5] ;
 wire \MEM.mem1[6] ;
 wire \MEM.mem1[7] ;
 wire \MEM.mem1[8] ;
 wire \MEM.mem1[9] ;
 wire \MEM.mem2[0] ;
 wire \MEM.mem2[10] ;
 wire \MEM.mem2[11] ;
 wire \MEM.mem2[1] ;
 wire \MEM.mem2[2] ;
 wire \MEM.mem2[3] ;
 wire \MEM.mem2[4] ;
 wire \MEM.mem2[5] ;
 wire \MEM.mem2[6] ;
 wire \MEM.mem2[7] ;
 wire \MEM.mem2[8] ;
 wire \MEM.mem2[9] ;
 wire \MEM.mem3[0] ;
 wire \MEM.mem3[10] ;
 wire \MEM.mem3[11] ;
 wire \MEM.mem3[1] ;
 wire \MEM.mem3[2] ;
 wire \MEM.mem3[3] ;
 wire \MEM.mem3[4] ;
 wire \MEM.mem3[5] ;
 wire \MEM.mem3[6] ;
 wire \MEM.mem3[7] ;
 wire \MEM.mem3[8] ;
 wire \MEM.mem3[9] ;
 wire \MEM.mem4[0] ;
 wire \MEM.mem4[10] ;
 wire \MEM.mem4[11] ;
 wire \MEM.mem4[1] ;
 wire \MEM.mem4[2] ;
 wire \MEM.mem4[3] ;
 wire \MEM.mem4[4] ;
 wire \MEM.mem4[5] ;
 wire \MEM.mem4[6] ;
 wire \MEM.mem4[7] ;
 wire \MEM.mem4[8] ;
 wire \MEM.mem4[9] ;
 wire \MEM.mem5[0] ;
 wire \MEM.mem5[10] ;
 wire \MEM.mem5[11] ;
 wire \MEM.mem5[1] ;
 wire \MEM.mem5[2] ;
 wire \MEM.mem5[3] ;
 wire \MEM.mem5[4] ;
 wire \MEM.mem5[5] ;
 wire \MEM.mem5[6] ;
 wire \MEM.mem5[7] ;
 wire \MEM.mem5[8] ;
 wire \MEM.mem5[9] ;
 wire \MEM.next_mem1[0] ;
 wire \MEM.next_mem1[10] ;
 wire \MEM.next_mem1[11] ;
 wire \MEM.next_mem1[1] ;
 wire \MEM.next_mem1[2] ;
 wire \MEM.next_mem1[3] ;
 wire \MEM.next_mem1[4] ;
 wire \MEM.next_mem1[5] ;
 wire \MEM.next_mem1[6] ;
 wire \MEM.next_mem1[7] ;
 wire \MEM.next_mem1[8] ;
 wire \MEM.next_mem1[9] ;
 wire \MEM.next_mem2[0] ;
 wire \MEM.next_mem2[10] ;
 wire \MEM.next_mem2[11] ;
 wire \MEM.next_mem2[1] ;
 wire \MEM.next_mem2[2] ;
 wire \MEM.next_mem2[3] ;
 wire \MEM.next_mem2[4] ;
 wire \MEM.next_mem2[5] ;
 wire \MEM.next_mem2[6] ;
 wire \MEM.next_mem2[7] ;
 wire \MEM.next_mem2[8] ;
 wire \MEM.next_mem2[9] ;
 wire \MEM.next_mem3[0] ;
 wire \MEM.next_mem3[10] ;
 wire \MEM.next_mem3[11] ;
 wire \MEM.next_mem3[1] ;
 wire \MEM.next_mem3[2] ;
 wire \MEM.next_mem3[3] ;
 wire \MEM.next_mem3[4] ;
 wire \MEM.next_mem3[5] ;
 wire \MEM.next_mem3[6] ;
 wire \MEM.next_mem3[7] ;
 wire \MEM.next_mem3[8] ;
 wire \MEM.next_mem3[9] ;
 wire \MEM.next_mem4[0] ;
 wire \MEM.next_mem4[10] ;
 wire \MEM.next_mem4[11] ;
 wire \MEM.next_mem4[1] ;
 wire \MEM.next_mem4[2] ;
 wire \MEM.next_mem4[3] ;
 wire \MEM.next_mem4[4] ;
 wire \MEM.next_mem4[5] ;
 wire \MEM.next_mem4[6] ;
 wire \MEM.next_mem4[7] ;
 wire \MEM.next_mem4[8] ;
 wire \MEM.next_mem4[9] ;
 wire \MEM.next_mem5[0] ;
 wire \MEM.next_mem5[10] ;
 wire \MEM.next_mem5[11] ;
 wire \MEM.next_mem5[1] ;
 wire \MEM.next_mem5[2] ;
 wire \MEM.next_mem5[3] ;
 wire \MEM.next_mem5[4] ;
 wire \MEM.next_mem5[5] ;
 wire \MEM.next_mem5[6] ;
 wire \MEM.next_mem5[7] ;
 wire \MEM.next_mem5[8] ;
 wire \MEM.next_mem5[9] ;
 wire \MEM.raddr[0] ;
 wire \MEM.raddr[1] ;
 wire \MEM.raddr[2] ;
 wire \TIM.cnt[0] ;
 wire \TIM.cnt[10] ;
 wire \TIM.cnt[11] ;
 wire \TIM.cnt[1] ;
 wire \TIM.cnt[2] ;
 wire \TIM.cnt[3] ;
 wire \TIM.cnt[4] ;
 wire \TIM.cnt[5] ;
 wire \TIM.cnt[6] ;
 wire \TIM.cnt[7] ;
 wire \TIM.cnt[8] ;
 wire \TIM.cnt[9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire \e1.edge_d ;
 wire \e1.intermediate ;
 wire \e1.sync ;
 wire \e2.edge_d ;
 wire \e2.intermediate ;
 wire \e2.sync ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net6));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_99 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__or4b_1 _0462_ (.A(\CLKDIV.count[5] ),
    .B(\CLKDIV.count[4] ),
    .C(\CLKDIV.count[6] ),
    .D_N(\CLKDIV.count[7] ),
    .X(_0057_));
 sky130_fd_sc_hd__or2_1 _0463_ (.A(\CLKDIV.count[1] ),
    .B(\CLKDIV.count[0] ),
    .X(_0058_));
 sky130_fd_sc_hd__or4_1 _0464_ (.A(\CLKDIV.count[3] ),
    .B(\CLKDIV.count[2] ),
    .C(_0057_),
    .D(_0058_),
    .X(_0059_));
 sky130_fd_sc_hd__or4bb_1 _0465_ (.A(\CLKDIV.count[13] ),
    .B(\CLKDIV.count[14] ),
    .C_N(\CLKDIV.count[15] ),
    .D_N(\CLKDIV.count[12] ),
    .X(_0060_));
 sky130_fd_sc_hd__or4bb_1 _0466_ (.A(\CLKDIV.count[8] ),
    .B(\CLKDIV.count[11] ),
    .C_N(\CLKDIV.count[10] ),
    .D_N(\CLKDIV.count[9] ),
    .X(_0061_));
 sky130_fd_sc_hd__or4bb_1 _0467_ (.A(\CLKDIV.count[21] ),
    .B(\CLKDIV.count[22] ),
    .C_N(\CLKDIV.count[23] ),
    .D_N(\CLKDIV.count[20] ),
    .X(_0062_));
 sky130_fd_sc_hd__or4b_1 _0468_ (.A(\CLKDIV.count[17] ),
    .B(\CLKDIV.count[16] ),
    .C(\CLKDIV.count[18] ),
    .D_N(\CLKDIV.count[19] ),
    .X(_0063_));
 sky130_fd_sc_hd__or4_1 _0469_ (.A(_0060_),
    .B(_0061_),
    .C(_0062_),
    .D(_0063_),
    .X(_0064_));
 sky130_fd_sc_hd__or2_2 _0470_ (.A(_0059_),
    .B(_0064_),
    .X(_0065_));
 sky130_fd_sc_hd__inv_2 _0471_ (.A(_0065_),
    .Y(_0024_));
 sky130_fd_sc_hd__buf_4 _0472_ (.A(\FSM.state[0] ),
    .X(_0066_));
 sky130_fd_sc_hd__or4bb_4 _0473_ (.A(\FSM.state[3] ),
    .B(_0066_),
    .C_N(\FSM.state[1] ),
    .D_N(\FSM.state[2] ),
    .X(_0067_));
 sky130_fd_sc_hd__or4bb_4 _0474_ (.A(\FSM.state[3] ),
    .B(\FSM.state[1] ),
    .C_N(_0066_),
    .D_N(\FSM.state[2] ),
    .X(_0068_));
 sky130_fd_sc_hd__nand2_8 _0475_ (.A(_0067_),
    .B(_0068_),
    .Y(_0069_));
 sky130_fd_sc_hd__buf_6 _0476_ (.A(\MEM.raddr[2] ),
    .X(_0070_));
 sky130_fd_sc_hd__clkinv_4 _0477_ (.A(_0070_),
    .Y(_0071_));
 sky130_fd_sc_hd__buf_4 _0478_ (.A(\MEM.raddr[1] ),
    .X(_0072_));
 sky130_fd_sc_hd__clkbuf_8 _0479_ (.A(\MEM.raddr[0] ),
    .X(_0073_));
 sky130_fd_sc_hd__and2_1 _0480_ (.A(_0072_),
    .B(_0073_),
    .X(_0074_));
 sky130_fd_sc_hd__buf_4 _0481_ (.A(_0074_),
    .X(_0075_));
 sky130_fd_sc_hd__nor2_4 _0482_ (.A(_0072_),
    .B(_0073_),
    .Y(_0076_));
 sky130_fd_sc_hd__a221o_1 _0483_ (.A1(\MEM.mem5[11] ),
    .A2(_0075_),
    .B1(_0076_),
    .B2(\MEM.mem2[11] ),
    .C1(_0070_),
    .X(_0077_));
 sky130_fd_sc_hd__nor3b_4 _0484_ (.A(_0073_),
    .B(_0070_),
    .C_N(_0072_),
    .Y(_0078_));
 sky130_fd_sc_hd__nor3b_2 _0485_ (.A(_0072_),
    .B(_0070_),
    .C_N(_0073_),
    .Y(_0079_));
 sky130_fd_sc_hd__a22o_1 _0486_ (.A1(\MEM.mem4[11] ),
    .A2(_0078_),
    .B1(net33),
    .B2(\MEM.mem3[11] ),
    .X(_0080_));
 sky130_fd_sc_hd__o22a_1 _0487_ (.A1(_0071_),
    .A2(\MEM.mem1[11] ),
    .B1(_0077_),
    .B2(_0080_),
    .X(_0081_));
 sky130_fd_sc_hd__nand4b_4 _0488_ (.A_N(\FSM.state[3] ),
    .B(\FSM.state[1] ),
    .C(_0066_),
    .D(\FSM.state[2] ),
    .Y(_0082_));
 sky130_fd_sc_hd__or4b_1 _0489_ (.A(\FSM.state[2] ),
    .B(\FSM.state[1] ),
    .C(_0066_),
    .D_N(\FSM.state[3] ),
    .X(_0083_));
 sky130_fd_sc_hd__clkbuf_4 _0490_ (.A(_0083_),
    .X(_0084_));
 sky130_fd_sc_hd__nand2_8 _0491_ (.A(_0082_),
    .B(_0084_),
    .Y(_0085_));
 sky130_fd_sc_hd__nor3b_4 _0492_ (.A(\FSM.state[2] ),
    .B(\FSM.state[3] ),
    .C_N(\FSM.state[1] ),
    .Y(_0086_));
 sky130_fd_sc_hd__a22o_1 _0493_ (.A1(\TIM.cnt[11] ),
    .A2(_0085_),
    .B1(_0086_),
    .B2(\CTR.time_out[11] ),
    .X(_0087_));
 sky130_fd_sc_hd__a21oi_4 _0494_ (.A1(_0069_),
    .A2(_0081_),
    .B1(_0087_),
    .Y(_0088_));
 sky130_fd_sc_hd__a221o_1 _0495_ (.A1(\MEM.mem5[9] ),
    .A2(_0075_),
    .B1(_0076_),
    .B2(\MEM.mem2[9] ),
    .C1(_0070_),
    .X(_0089_));
 sky130_fd_sc_hd__a22o_1 _0496_ (.A1(\MEM.mem4[9] ),
    .A2(_0078_),
    .B1(net33),
    .B2(\MEM.mem3[9] ),
    .X(_0090_));
 sky130_fd_sc_hd__or2_1 _0497_ (.A(_0071_),
    .B(\MEM.mem1[9] ),
    .X(_0091_));
 sky130_fd_sc_hd__o211ai_2 _0498_ (.A1(_0089_),
    .A2(_0090_),
    .B1(_0091_),
    .C1(_0069_),
    .Y(_0092_));
 sky130_fd_sc_hd__a22oi_2 _0499_ (.A1(\TIM.cnt[9] ),
    .A2(_0085_),
    .B1(_0086_),
    .B2(\CTR.time_out[9] ),
    .Y(_0093_));
 sky130_fd_sc_hd__and4bb_1 _0500_ (.A_N(_0072_),
    .B_N(\MEM.raddr[2] ),
    .C(\MEM.mem3[10] ),
    .D(_0073_),
    .X(_0094_));
 sky130_fd_sc_hd__nor3b_1 _0501_ (.A(_0072_),
    .B(_0073_),
    .C_N(\MEM.mem2[10] ),
    .Y(_0095_));
 sky130_fd_sc_hd__and4bb_1 _0502_ (.A_N(_0073_),
    .B_N(\MEM.raddr[2] ),
    .C(\MEM.mem4[10] ),
    .D(_0072_),
    .X(_0096_));
 sky130_fd_sc_hd__a31o_1 _0503_ (.A1(_0072_),
    .A2(_0073_),
    .A3(\MEM.mem5[10] ),
    .B1(_0070_),
    .X(_0097_));
 sky130_fd_sc_hd__or4_2 _0504_ (.A(_0094_),
    .B(_0095_),
    .C(_0096_),
    .D(_0097_),
    .X(_0098_));
 sky130_fd_sc_hd__o2bb2a_1 _0505_ (.A1_N(_0067_),
    .A2_N(_0068_),
    .B1(_0071_),
    .B2(\MEM.mem1[10] ),
    .X(_0099_));
 sky130_fd_sc_hd__and2_1 _0506_ (.A(\CTR.time_out[10] ),
    .B(_0086_),
    .X(_0100_));
 sky130_fd_sc_hd__a221oi_1 _0507_ (.A1(\TIM.cnt[10] ),
    .A2(_0085_),
    .B1(_0098_),
    .B2(_0099_),
    .C1(_0100_),
    .Y(_0101_));
 sky130_fd_sc_hd__a21o_1 _0508_ (.A1(_0092_),
    .A2(_0093_),
    .B1(_0101_),
    .X(_0102_));
 sky130_fd_sc_hd__a221o_2 _0509_ (.A1(\TIM.cnt[10] ),
    .A2(_0085_),
    .B1(_0098_),
    .B2(_0099_),
    .C1(_0100_),
    .X(_0103_));
 sky130_fd_sc_hd__and4bb_1 _0510_ (.A_N(_0072_),
    .B_N(\MEM.raddr[2] ),
    .C(\MEM.mem3[8] ),
    .D(_0073_),
    .X(_0104_));
 sky130_fd_sc_hd__nor3b_1 _0511_ (.A(_0072_),
    .B(_0073_),
    .C_N(\MEM.mem2[8] ),
    .Y(_0105_));
 sky130_fd_sc_hd__and4bb_1 _0512_ (.A_N(_0073_),
    .B_N(\MEM.raddr[2] ),
    .C(\MEM.mem4[8] ),
    .D(_0072_),
    .X(_0106_));
 sky130_fd_sc_hd__a31o_1 _0513_ (.A1(_0072_),
    .A2(_0073_),
    .A3(\MEM.mem5[8] ),
    .B1(\MEM.raddr[2] ),
    .X(_0107_));
 sky130_fd_sc_hd__or4_1 _0514_ (.A(_0104_),
    .B(_0105_),
    .C(_0106_),
    .D(_0107_),
    .X(_0108_));
 sky130_fd_sc_hd__o2bb2a_1 _0515_ (.A1_N(_0067_),
    .A2_N(_0068_),
    .B1(_0071_),
    .B2(\MEM.mem1[8] ),
    .X(_0109_));
 sky130_fd_sc_hd__and2_1 _0516_ (.A(\CTR.time_out[8] ),
    .B(_0086_),
    .X(_0110_));
 sky130_fd_sc_hd__a221o_2 _0517_ (.A1(\TIM.cnt[8] ),
    .A2(_0085_),
    .B1(_0108_),
    .B2(_0109_),
    .C1(_0110_),
    .X(_0111_));
 sky130_fd_sc_hd__nand2_1 _0518_ (.A(_0103_),
    .B(_0111_),
    .Y(_0112_));
 sky130_fd_sc_hd__nand3_2 _0519_ (.A(_0088_),
    .B(_0102_),
    .C(_0112_),
    .Y(net31));
 sky130_fd_sc_hd__nand2_2 _0520_ (.A(_0092_),
    .B(_0093_),
    .Y(_0113_));
 sky130_fd_sc_hd__and4bb_1 _0521_ (.A_N(_0072_),
    .B_N(_0070_),
    .C(\MEM.mem3[7] ),
    .D(_0073_),
    .X(_0114_));
 sky130_fd_sc_hd__nor3b_1 _0522_ (.A(_0072_),
    .B(_0073_),
    .C_N(\MEM.mem2[7] ),
    .Y(_0115_));
 sky130_fd_sc_hd__and4bb_1 _0523_ (.A_N(_0073_),
    .B_N(_0070_),
    .C(\MEM.mem4[7] ),
    .D(_0072_),
    .X(_0116_));
 sky130_fd_sc_hd__a31o_1 _0524_ (.A1(_0072_),
    .A2(_0073_),
    .A3(\MEM.mem5[7] ),
    .B1(_0070_),
    .X(_0117_));
 sky130_fd_sc_hd__or4_1 _0525_ (.A(_0114_),
    .B(_0115_),
    .C(_0116_),
    .D(_0117_),
    .X(_0118_));
 sky130_fd_sc_hd__o2bb2a_1 _0526_ (.A1_N(_0067_),
    .A2_N(_0068_),
    .B1(_0071_),
    .B2(\MEM.mem1[7] ),
    .X(_0119_));
 sky130_fd_sc_hd__and2_1 _0527_ (.A(\CTR.time_out[7] ),
    .B(_0086_),
    .X(_0120_));
 sky130_fd_sc_hd__a221o_2 _0528_ (.A1(\TIM.cnt[7] ),
    .A2(_0085_),
    .B1(_0118_),
    .B2(_0119_),
    .C1(_0120_),
    .X(_0121_));
 sky130_fd_sc_hd__or2_2 _0529_ (.A(_0111_),
    .B(_0121_),
    .X(_0122_));
 sky130_fd_sc_hd__a21oi_1 _0530_ (.A1(_0113_),
    .A2(_0122_),
    .B1(_0103_),
    .Y(_0123_));
 sky130_fd_sc_hd__nand2_1 _0531_ (.A(_0111_),
    .B(_0121_),
    .Y(_0124_));
 sky130_fd_sc_hd__o21a_1 _0532_ (.A1(_0102_),
    .A2(_0124_),
    .B1(_0088_),
    .X(_0125_));
 sky130_fd_sc_hd__o21a_1 _0533_ (.A1(net31),
    .A2(_0123_),
    .B1(_0125_),
    .X(_0126_));
 sky130_fd_sc_hd__nor2_1 _0534_ (.A(_0103_),
    .B(_0113_),
    .Y(_0127_));
 sky130_fd_sc_hd__nor2_1 _0535_ (.A(_0088_),
    .B(_0127_),
    .Y(_0128_));
 sky130_fd_sc_hd__or2_1 _0536_ (.A(_0088_),
    .B(_0101_),
    .X(_0129_));
 sky130_fd_sc_hd__o21bai_4 _0537_ (.A1(_0113_),
    .A2(_0122_),
    .B1_N(_0129_),
    .Y(net26));
 sky130_fd_sc_hd__o21ai_1 _0538_ (.A1(_0126_),
    .A2(_0128_),
    .B1(net26),
    .Y(_0130_));
 sky130_fd_sc_hd__or3b_2 _0539_ (.A(_0088_),
    .B(_0102_),
    .C_N(_0111_),
    .X(_0131_));
 sky130_fd_sc_hd__or2b_1 _0540_ (.A(_0126_),
    .B_N(_0131_),
    .X(_0132_));
 sky130_fd_sc_hd__clkbuf_2 _0541_ (.A(_0132_),
    .X(net29));
 sky130_fd_sc_hd__a21o_1 _0542_ (.A1(net31),
    .A2(_0130_),
    .B1(net29),
    .X(net25));
 sky130_fd_sc_hd__inv_2 _0543_ (.A(net31),
    .Y(_0133_));
 sky130_fd_sc_hd__nand2_1 _0544_ (.A(_0131_),
    .B(_0130_),
    .Y(_0134_));
 sky130_fd_sc_hd__or3b_1 _0545_ (.A(_0133_),
    .B(_0128_),
    .C_N(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__buf_1 _0546_ (.A(_0135_),
    .X(net27));
 sky130_fd_sc_hd__a21o_1 _0547_ (.A1(net31),
    .A2(_0130_),
    .B1(net29),
    .X(net28));
 sky130_fd_sc_hd__a31o_1 _0548_ (.A1(_0133_),
    .A2(_0126_),
    .A3(net26),
    .B1(_0128_),
    .X(net30));
 sky130_fd_sc_hd__nor2_1 _0549_ (.A(net114),
    .B(_0024_),
    .Y(_0000_));
 sky130_fd_sc_hd__nand2_1 _0550_ (.A(\CLKDIV.count[1] ),
    .B(\CLKDIV.count[0] ),
    .Y(_0136_));
 sky130_fd_sc_hd__and2_1 _0551_ (.A(_0058_),
    .B(_0136_),
    .X(_0137_));
 sky130_fd_sc_hd__clkbuf_1 _0552_ (.A(_0137_),
    .X(_0011_));
 sky130_fd_sc_hd__a21oi_1 _0553_ (.A1(\CLKDIV.count[1] ),
    .A2(net114),
    .B1(net125),
    .Y(_0138_));
 sky130_fd_sc_hd__and3_1 _0554_ (.A(\CLKDIV.count[1] ),
    .B(\CLKDIV.count[0] ),
    .C(\CLKDIV.count[2] ),
    .X(_0139_));
 sky130_fd_sc_hd__nor2_1 _0555_ (.A(net126),
    .B(_0139_),
    .Y(_0016_));
 sky130_fd_sc_hd__and4_1 _0556_ (.A(\CLKDIV.count[1] ),
    .B(\CLKDIV.count[0] ),
    .C(\CLKDIV.count[3] ),
    .D(\CLKDIV.count[2] ),
    .X(_0140_));
 sky130_fd_sc_hd__nor2_1 _0557_ (.A(net121),
    .B(_0139_),
    .Y(_0141_));
 sky130_fd_sc_hd__nor2_1 _0558_ (.A(_0140_),
    .B(_0141_),
    .Y(_0017_));
 sky130_fd_sc_hd__nand2_1 _0559_ (.A(\CLKDIV.count[4] ),
    .B(_0140_),
    .Y(_0142_));
 sky130_fd_sc_hd__or2_1 _0560_ (.A(\CLKDIV.count[4] ),
    .B(_0140_),
    .X(_0143_));
 sky130_fd_sc_hd__and2_1 _0561_ (.A(_0142_),
    .B(_0143_),
    .X(_0144_));
 sky130_fd_sc_hd__clkbuf_1 _0562_ (.A(_0144_),
    .X(_0018_));
 sky130_fd_sc_hd__xnor2_1 _0563_ (.A(net122),
    .B(_0142_),
    .Y(_0019_));
 sky130_fd_sc_hd__and4_1 _0564_ (.A(\CLKDIV.count[5] ),
    .B(\CLKDIV.count[4] ),
    .C(\CLKDIV.count[6] ),
    .D(_0140_),
    .X(_0145_));
 sky130_fd_sc_hd__a31o_1 _0565_ (.A1(\CLKDIV.count[5] ),
    .A2(\CLKDIV.count[4] ),
    .A3(_0140_),
    .B1(\CLKDIV.count[6] ),
    .X(_0146_));
 sky130_fd_sc_hd__and2b_1 _0566_ (.A_N(_0145_),
    .B(_0146_),
    .X(_0147_));
 sky130_fd_sc_hd__clkbuf_1 _0567_ (.A(_0147_),
    .X(_0020_));
 sky130_fd_sc_hd__or2_1 _0568_ (.A(\CLKDIV.count[7] ),
    .B(_0145_),
    .X(_0148_));
 sky130_fd_sc_hd__nand2_1 _0569_ (.A(\CLKDIV.count[7] ),
    .B(_0145_),
    .Y(_0149_));
 sky130_fd_sc_hd__and3_1 _0570_ (.A(_0065_),
    .B(_0148_),
    .C(_0149_),
    .X(_0150_));
 sky130_fd_sc_hd__clkbuf_1 _0571_ (.A(_0150_),
    .X(_0021_));
 sky130_fd_sc_hd__and3_1 _0572_ (.A(\CLKDIV.count[7] ),
    .B(\CLKDIV.count[8] ),
    .C(_0145_),
    .X(_0151_));
 sky130_fd_sc_hd__a21oi_1 _0573_ (.A1(\CLKDIV.count[7] ),
    .A2(_0145_),
    .B1(net119),
    .Y(_0152_));
 sky130_fd_sc_hd__nor2_1 _0574_ (.A(_0151_),
    .B(net120),
    .Y(_0022_));
 sky130_fd_sc_hd__and2_1 _0575_ (.A(\CLKDIV.count[9] ),
    .B(_0151_),
    .X(_0153_));
 sky130_fd_sc_hd__nor2_1 _0576_ (.A(_0024_),
    .B(_0153_),
    .Y(_0154_));
 sky130_fd_sc_hd__o21a_1 _0577_ (.A1(net113),
    .A2(_0151_),
    .B1(_0154_),
    .X(_0023_));
 sky130_fd_sc_hd__or2_1 _0578_ (.A(\CLKDIV.count[10] ),
    .B(_0153_),
    .X(_0155_));
 sky130_fd_sc_hd__nand2_1 _0579_ (.A(\CLKDIV.count[10] ),
    .B(_0153_),
    .Y(_0156_));
 sky130_fd_sc_hd__and3_1 _0580_ (.A(_0065_),
    .B(_0155_),
    .C(_0156_),
    .X(_0157_));
 sky130_fd_sc_hd__clkbuf_1 _0581_ (.A(_0157_),
    .X(_0001_));
 sky130_fd_sc_hd__xnor2_1 _0582_ (.A(net116),
    .B(_0156_),
    .Y(_0002_));
 sky130_fd_sc_hd__and4_1 _0583_ (.A(\CLKDIV.count[11] ),
    .B(\CLKDIV.count[10] ),
    .C(\CLKDIV.count[12] ),
    .D(_0153_),
    .X(_0158_));
 sky130_fd_sc_hd__buf_1 _0584_ (.A(_0158_),
    .X(_0159_));
 sky130_fd_sc_hd__a31o_1 _0585_ (.A1(\CLKDIV.count[11] ),
    .A2(\CLKDIV.count[10] ),
    .A3(_0153_),
    .B1(\CLKDIV.count[12] ),
    .X(_0160_));
 sky130_fd_sc_hd__nor3b_1 _0586_ (.A(_0024_),
    .B(_0159_),
    .C_N(_0160_),
    .Y(_0003_));
 sky130_fd_sc_hd__xor2_1 _0587_ (.A(net111),
    .B(_0159_),
    .X(_0004_));
 sky130_fd_sc_hd__and3_1 _0588_ (.A(\CLKDIV.count[13] ),
    .B(\CLKDIV.count[14] ),
    .C(_0159_),
    .X(_0161_));
 sky130_fd_sc_hd__a21oi_1 _0589_ (.A1(\CLKDIV.count[13] ),
    .A2(_0159_),
    .B1(net105),
    .Y(_0162_));
 sky130_fd_sc_hd__nor2_1 _0590_ (.A(_0161_),
    .B(net106),
    .Y(_0005_));
 sky130_fd_sc_hd__and2_1 _0591_ (.A(\CLKDIV.count[15] ),
    .B(_0161_),
    .X(_0163_));
 sky130_fd_sc_hd__nor2_1 _0592_ (.A(_0024_),
    .B(_0163_),
    .Y(_0164_));
 sky130_fd_sc_hd__o21a_1 _0593_ (.A1(net109),
    .A2(_0161_),
    .B1(_0164_),
    .X(_0006_));
 sky130_fd_sc_hd__nand2_1 _0594_ (.A(\CLKDIV.count[16] ),
    .B(_0163_),
    .Y(_0165_));
 sky130_fd_sc_hd__or2_1 _0595_ (.A(\CLKDIV.count[16] ),
    .B(_0163_),
    .X(_0166_));
 sky130_fd_sc_hd__and2_1 _0596_ (.A(_0165_),
    .B(_0166_),
    .X(_0167_));
 sky130_fd_sc_hd__clkbuf_1 _0597_ (.A(_0167_),
    .X(_0007_));
 sky130_fd_sc_hd__xnor2_1 _0598_ (.A(net115),
    .B(_0165_),
    .Y(_0008_));
 sky130_fd_sc_hd__and4_1 _0599_ (.A(\CLKDIV.count[17] ),
    .B(\CLKDIV.count[16] ),
    .C(\CLKDIV.count[18] ),
    .D(_0163_),
    .X(_0168_));
 sky130_fd_sc_hd__a31o_1 _0600_ (.A1(\CLKDIV.count[17] ),
    .A2(\CLKDIV.count[16] ),
    .A3(_0163_),
    .B1(\CLKDIV.count[18] ),
    .X(_0169_));
 sky130_fd_sc_hd__and2b_1 _0601_ (.A_N(_0168_),
    .B(_0169_),
    .X(_0170_));
 sky130_fd_sc_hd__clkbuf_1 _0602_ (.A(_0170_),
    .X(_0009_));
 sky130_fd_sc_hd__o21ai_1 _0603_ (.A1(net102),
    .A2(_0168_),
    .B1(_0065_),
    .Y(_0171_));
 sky130_fd_sc_hd__a21oi_1 _0604_ (.A1(net102),
    .A2(_0168_),
    .B1(_0171_),
    .Y(_0010_));
 sky130_fd_sc_hd__a21oi_1 _0605_ (.A1(\CLKDIV.count[19] ),
    .A2(_0168_),
    .B1(net131),
    .Y(_0172_));
 sky130_fd_sc_hd__and3_1 _0606_ (.A(\CLKDIV.count[19] ),
    .B(\CLKDIV.count[20] ),
    .C(_0168_),
    .X(_0173_));
 sky130_fd_sc_hd__nor3_1 _0607_ (.A(_0024_),
    .B(_0172_),
    .C(_0173_),
    .Y(_0012_));
 sky130_fd_sc_hd__and2_1 _0608_ (.A(\CLKDIV.count[21] ),
    .B(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__nor2_1 _0609_ (.A(net124),
    .B(_0173_),
    .Y(_0175_));
 sky130_fd_sc_hd__nor2_1 _0610_ (.A(_0174_),
    .B(_0175_),
    .Y(_0013_));
 sky130_fd_sc_hd__xor2_1 _0611_ (.A(net123),
    .B(_0174_),
    .X(_0014_));
 sky130_fd_sc_hd__nand3_1 _0612_ (.A(\CLKDIV.count[22] ),
    .B(\CLKDIV.count[23] ),
    .C(_0174_),
    .Y(_0176_));
 sky130_fd_sc_hd__a31o_1 _0613_ (.A1(\CLKDIV.count[21] ),
    .A2(\CLKDIV.count[22] ),
    .A3(_0173_),
    .B1(\CLKDIV.count[23] ),
    .X(_0177_));
 sky130_fd_sc_hd__and3_1 _0614_ (.A(_0065_),
    .B(_0176_),
    .C(_0177_),
    .X(_0178_));
 sky130_fd_sc_hd__clkbuf_1 _0615_ (.A(_0178_),
    .X(_0015_));
 sky130_fd_sc_hd__a221o_1 _0616_ (.A1(\MEM.mem5[4] ),
    .A2(_0075_),
    .B1(_0076_),
    .B2(\MEM.mem2[4] ),
    .C1(_0070_),
    .X(_0179_));
 sky130_fd_sc_hd__a221o_1 _0617_ (.A1(\MEM.mem4[4] ),
    .A2(_0078_),
    .B1(_0079_),
    .B2(\MEM.mem3[4] ),
    .C1(_0179_),
    .X(_0180_));
 sky130_fd_sc_hd__or2_1 _0618_ (.A(_0071_),
    .B(\MEM.mem1[4] ),
    .X(_0181_));
 sky130_fd_sc_hd__a22o_1 _0619_ (.A1(\TIM.cnt[4] ),
    .A2(_0085_),
    .B1(net34),
    .B2(\CTR.time_out[4] ),
    .X(_0182_));
 sky130_fd_sc_hd__a31o_2 _0620_ (.A1(_0069_),
    .A2(_0180_),
    .A3(_0181_),
    .B1(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__inv_2 _0621_ (.A(_0073_),
    .Y(_0184_));
 sky130_fd_sc_hd__a31o_1 _0622_ (.A1(_0072_),
    .A2(_0184_),
    .A3(\MEM.mem4[3] ),
    .B1(_0070_),
    .X(_0185_));
 sky130_fd_sc_hd__a22o_1 _0623_ (.A1(\MEM.mem5[3] ),
    .A2(_0075_),
    .B1(_0076_),
    .B2(\MEM.mem2[3] ),
    .X(_0186_));
 sky130_fd_sc_hd__a211o_1 _0624_ (.A1(\MEM.mem3[3] ),
    .A2(_0079_),
    .B1(_0185_),
    .C1(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__or2_1 _0625_ (.A(_0071_),
    .B(\MEM.mem1[3] ),
    .X(_0188_));
 sky130_fd_sc_hd__clkbuf_4 _0626_ (.A(\CTR.time_out[3] ),
    .X(_0189_));
 sky130_fd_sc_hd__a22o_1 _0627_ (.A1(\TIM.cnt[3] ),
    .A2(_0085_),
    .B1(net34),
    .B2(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__a31o_4 _0628_ (.A1(_0069_),
    .A2(_0187_),
    .A3(_0188_),
    .B1(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__a221o_1 _0629_ (.A1(\MEM.mem5[2] ),
    .A2(_0075_),
    .B1(_0076_),
    .B2(\MEM.mem2[2] ),
    .C1(_0070_),
    .X(_0192_));
 sky130_fd_sc_hd__a221o_1 _0630_ (.A1(\MEM.mem4[2] ),
    .A2(_0078_),
    .B1(net33),
    .B2(\MEM.mem3[2] ),
    .C1(_0192_),
    .X(_0193_));
 sky130_fd_sc_hd__or2_1 _0631_ (.A(_0071_),
    .B(\MEM.mem1[2] ),
    .X(_0194_));
 sky130_fd_sc_hd__a22o_1 _0632_ (.A1(\TIM.cnt[2] ),
    .A2(_0085_),
    .B1(net34),
    .B2(\CTR.time_out[2] ),
    .X(_0195_));
 sky130_fd_sc_hd__a31oi_4 _0633_ (.A1(_0069_),
    .A2(_0193_),
    .A3(_0194_),
    .B1(_0195_),
    .Y(_0196_));
 sky130_fd_sc_hd__a221o_1 _0634_ (.A1(\MEM.mem5[1] ),
    .A2(_0075_),
    .B1(_0076_),
    .B2(\MEM.mem2[1] ),
    .C1(_0070_),
    .X(_0197_));
 sky130_fd_sc_hd__a221o_1 _0635_ (.A1(\MEM.mem4[1] ),
    .A2(_0078_),
    .B1(net33),
    .B2(\MEM.mem3[1] ),
    .C1(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__o21a_1 _0636_ (.A1(_0071_),
    .A2(\MEM.mem1[1] ),
    .B1(_0069_),
    .X(_0199_));
 sky130_fd_sc_hd__clkbuf_4 _0637_ (.A(\CTR.time_out[1] ),
    .X(_0200_));
 sky130_fd_sc_hd__a22o_1 _0638_ (.A1(\TIM.cnt[1] ),
    .A2(_0085_),
    .B1(net34),
    .B2(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__a21oi_4 _0639_ (.A1(_0198_),
    .A2(_0199_),
    .B1(_0201_),
    .Y(_0202_));
 sky130_fd_sc_hd__nor2_2 _0640_ (.A(_0196_),
    .B(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__a221o_1 _0641_ (.A1(\MEM.mem5[5] ),
    .A2(_0075_),
    .B1(_0076_),
    .B2(\MEM.mem2[5] ),
    .C1(_0070_),
    .X(_0204_));
 sky130_fd_sc_hd__a221o_1 _0642_ (.A1(\MEM.mem4[5] ),
    .A2(_0078_),
    .B1(_0079_),
    .B2(\MEM.mem3[5] ),
    .C1(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__or2_1 _0643_ (.A(_0071_),
    .B(\MEM.mem1[5] ),
    .X(_0206_));
 sky130_fd_sc_hd__a22o_1 _0644_ (.A1(\TIM.cnt[5] ),
    .A2(_0085_),
    .B1(net34),
    .B2(\CTR.time_out[5] ),
    .X(_0207_));
 sky130_fd_sc_hd__a31o_2 _0645_ (.A1(_0069_),
    .A2(_0205_),
    .A3(_0206_),
    .B1(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__a31oi_4 _0646_ (.A1(_0183_),
    .A2(_0191_),
    .A3(_0203_),
    .B1(_0208_),
    .Y(_0209_));
 sky130_fd_sc_hd__inv_2 _0647_ (.A(_0183_),
    .Y(_0210_));
 sky130_fd_sc_hd__a21bo_1 _0648_ (.A1(_0196_),
    .A2(_0202_),
    .B1_N(_0191_),
    .X(_0211_));
 sky130_fd_sc_hd__a31o_1 _0649_ (.A1(_0069_),
    .A2(_0193_),
    .A3(_0194_),
    .B1(_0195_),
    .X(_0212_));
 sky130_fd_sc_hd__o21a_1 _0650_ (.A1(_0191_),
    .A2(_0212_),
    .B1(_0183_),
    .X(_0213_));
 sky130_fd_sc_hd__a21o_1 _0651_ (.A1(_0210_),
    .A2(_0211_),
    .B1(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__and2_1 _0652_ (.A(_0209_),
    .B(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__nand2_1 _0653_ (.A(_0196_),
    .B(_0202_),
    .Y(_0216_));
 sky130_fd_sc_hd__and2_1 _0654_ (.A(_0208_),
    .B(_0183_),
    .X(_0217_));
 sky130_fd_sc_hd__o21ai_2 _0655_ (.A1(_0191_),
    .A2(_0216_),
    .B1(_0217_),
    .Y(net12));
 sky130_fd_sc_hd__o21a_1 _0656_ (.A1(_0183_),
    .A2(_0191_),
    .B1(_0208_),
    .X(_0218_));
 sky130_fd_sc_hd__a21o_1 _0657_ (.A1(_0209_),
    .A2(_0214_),
    .B1(_0218_),
    .X(_0219_));
 sky130_fd_sc_hd__nor2_2 _0658_ (.A(_0208_),
    .B(_0213_),
    .Y(_0220_));
 sky130_fd_sc_hd__a21oi_1 _0659_ (.A1(net12),
    .A2(_0219_),
    .B1(_0220_),
    .Y(_0221_));
 sky130_fd_sc_hd__or2_1 _0660_ (.A(_0215_),
    .B(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__clkbuf_1 _0661_ (.A(_0222_),
    .X(net11));
 sky130_fd_sc_hd__and2_1 _0662_ (.A(_0191_),
    .B(_0212_),
    .X(_0223_));
 sky130_fd_sc_hd__and2_1 _0663_ (.A(_0217_),
    .B(_0223_),
    .X(_0224_));
 sky130_fd_sc_hd__a21o_1 _0664_ (.A1(net12),
    .A2(_0219_),
    .B1(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__or3b_2 _0665_ (.A(_0218_),
    .B(_0220_),
    .C_N(_0225_),
    .X(_0226_));
 sky130_fd_sc_hd__clkbuf_1 _0666_ (.A(_0226_),
    .X(net13));
 sky130_fd_sc_hd__or2_1 _0667_ (.A(_0215_),
    .B(_0221_),
    .X(_0227_));
 sky130_fd_sc_hd__clkbuf_1 _0668_ (.A(_0227_),
    .X(net14));
 sky130_fd_sc_hd__or2_1 _0669_ (.A(_0215_),
    .B(_0224_),
    .X(_0228_));
 sky130_fd_sc_hd__clkbuf_1 _0670_ (.A(_0228_),
    .X(net15));
 sky130_fd_sc_hd__a31o_1 _0671_ (.A1(_0215_),
    .A2(net12),
    .A3(_0220_),
    .B1(_0218_),
    .X(net16));
 sky130_fd_sc_hd__inv_2 _0672_ (.A(_0220_),
    .Y(net17));
 sky130_fd_sc_hd__buf_4 _0673_ (.A(\CTR.time_out[0] ),
    .X(_0229_));
 sky130_fd_sc_hd__inv_2 _0674_ (.A(\MEM.addr[2] ),
    .Y(_0230_));
 sky130_fd_sc_hd__nor3b_4 _0675_ (.A(\FSM.state[3] ),
    .B(\FSM.state[1] ),
    .C_N(\FSM.state[2] ),
    .Y(_0231_));
 sky130_fd_sc_hd__nand2b_4 _0676_ (.A_N(_0066_),
    .B(_0231_),
    .Y(_0232_));
 sky130_fd_sc_hd__nor2_8 _0677_ (.A(_0230_),
    .B(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__nor2_1 _0678_ (.A(\FSM.state[2] ),
    .B(\FSM.state[3] ),
    .Y(_0234_));
 sky130_fd_sc_hd__and2b_1 _0679_ (.A_N(\FSM.state[1] ),
    .B(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__buf_8 _0680_ (.A(_0235_),
    .X(_0236_));
 sky130_fd_sc_hd__nor2_4 _0681_ (.A(_0233_),
    .B(_0236_),
    .Y(_0237_));
 sky130_fd_sc_hd__a22o_1 _0682_ (.A1(_0229_),
    .A2(_0233_),
    .B1(_0237_),
    .B2(net57),
    .X(\MEM.next_mem1[0] ));
 sky130_fd_sc_hd__a22o_1 _0683_ (.A1(_0200_),
    .A2(_0233_),
    .B1(_0237_),
    .B2(net87),
    .X(\MEM.next_mem1[1] ));
 sky130_fd_sc_hd__a22o_1 _0684_ (.A1(\CTR.time_out[2] ),
    .A2(_0233_),
    .B1(_0237_),
    .B2(net50),
    .X(\MEM.next_mem1[2] ));
 sky130_fd_sc_hd__a22o_1 _0685_ (.A1(_0189_),
    .A2(_0233_),
    .B1(_0237_),
    .B2(net47),
    .X(\MEM.next_mem1[3] ));
 sky130_fd_sc_hd__a22o_1 _0686_ (.A1(\CTR.time_out[4] ),
    .A2(_0233_),
    .B1(_0237_),
    .B2(net48),
    .X(\MEM.next_mem1[4] ));
 sky130_fd_sc_hd__a22o_1 _0687_ (.A1(\CTR.time_out[5] ),
    .A2(_0233_),
    .B1(_0237_),
    .B2(net46),
    .X(\MEM.next_mem1[5] ));
 sky130_fd_sc_hd__a22o_1 _0688_ (.A1(\CTR.time_out[6] ),
    .A2(_0233_),
    .B1(_0237_),
    .B2(net55),
    .X(\MEM.next_mem1[6] ));
 sky130_fd_sc_hd__a22o_1 _0689_ (.A1(\CTR.time_out[7] ),
    .A2(_0233_),
    .B1(_0237_),
    .B2(net52),
    .X(\MEM.next_mem1[7] ));
 sky130_fd_sc_hd__a22o_1 _0690_ (.A1(\CTR.time_out[8] ),
    .A2(_0233_),
    .B1(_0237_),
    .B2(net49),
    .X(\MEM.next_mem1[8] ));
 sky130_fd_sc_hd__a22o_1 _0691_ (.A1(\CTR.time_out[9] ),
    .A2(_0233_),
    .B1(_0237_),
    .B2(net51),
    .X(\MEM.next_mem1[9] ));
 sky130_fd_sc_hd__a22o_1 _0692_ (.A1(\CTR.time_out[10] ),
    .A2(_0233_),
    .B1(_0237_),
    .B2(net64),
    .X(\MEM.next_mem1[10] ));
 sky130_fd_sc_hd__a22o_1 _0693_ (.A1(\CTR.time_out[11] ),
    .A2(_0233_),
    .B1(_0237_),
    .B2(net78),
    .X(\MEM.next_mem1[11] ));
 sky130_fd_sc_hd__or3_4 _0694_ (.A(\FSM.state[2] ),
    .B(\FSM.state[3] ),
    .C(\FSM.state[1] ),
    .X(_0238_));
 sky130_fd_sc_hd__o41a_1 _0695_ (.A1(\MEM.addr[0] ),
    .A2(\MEM.addr[1] ),
    .A3(\MEM.addr[2] ),
    .A4(_0232_),
    .B1(_0238_),
    .X(_0239_));
 sky130_fd_sc_hd__buf_4 _0696_ (.A(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__inv_2 _0697_ (.A(\MEM.addr[1] ),
    .Y(_0241_));
 sky130_fd_sc_hd__nor2b_2 _0698_ (.A(_0066_),
    .B_N(_0231_),
    .Y(_0242_));
 sky130_fd_sc_hd__and4b_1 _0699_ (.A_N(\MEM.addr[0] ),
    .B(_0241_),
    .C(_0230_),
    .D(_0242_),
    .X(_0243_));
 sky130_fd_sc_hd__buf_4 _0700_ (.A(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__a22o_1 _0701_ (.A1(net99),
    .A2(_0240_),
    .B1(_0244_),
    .B2(_0229_),
    .X(\MEM.next_mem2[0] ));
 sky130_fd_sc_hd__a22o_1 _0702_ (.A1(net93),
    .A2(_0240_),
    .B1(_0244_),
    .B2(_0200_),
    .X(\MEM.next_mem2[1] ));
 sky130_fd_sc_hd__a22o_1 _0703_ (.A1(net100),
    .A2(_0240_),
    .B1(_0244_),
    .B2(\CTR.time_out[2] ),
    .X(\MEM.next_mem2[2] ));
 sky130_fd_sc_hd__a22o_1 _0704_ (.A1(net90),
    .A2(_0240_),
    .B1(_0244_),
    .B2(_0189_),
    .X(\MEM.next_mem2[3] ));
 sky130_fd_sc_hd__a22o_1 _0705_ (.A1(net96),
    .A2(_0240_),
    .B1(_0244_),
    .B2(\CTR.time_out[4] ),
    .X(\MEM.next_mem2[4] ));
 sky130_fd_sc_hd__a22o_1 _0706_ (.A1(net94),
    .A2(_0240_),
    .B1(_0244_),
    .B2(\CTR.time_out[5] ),
    .X(\MEM.next_mem2[5] ));
 sky130_fd_sc_hd__a22o_1 _0707_ (.A1(net91),
    .A2(_0240_),
    .B1(_0244_),
    .B2(\CTR.time_out[6] ),
    .X(\MEM.next_mem2[6] ));
 sky130_fd_sc_hd__a22o_1 _0708_ (.A1(net58),
    .A2(_0240_),
    .B1(_0244_),
    .B2(\CTR.time_out[7] ),
    .X(\MEM.next_mem2[7] ));
 sky130_fd_sc_hd__a22o_1 _0709_ (.A1(net73),
    .A2(_0240_),
    .B1(_0244_),
    .B2(\CTR.time_out[8] ),
    .X(\MEM.next_mem2[8] ));
 sky130_fd_sc_hd__a22o_1 _0710_ (.A1(net108),
    .A2(_0240_),
    .B1(_0244_),
    .B2(\CTR.time_out[9] ),
    .X(\MEM.next_mem2[9] ));
 sky130_fd_sc_hd__a22o_1 _0711_ (.A1(net83),
    .A2(_0240_),
    .B1(_0244_),
    .B2(\CTR.time_out[10] ),
    .X(\MEM.next_mem2[10] ));
 sky130_fd_sc_hd__a22o_1 _0712_ (.A1(net98),
    .A2(_0240_),
    .B1(_0244_),
    .B2(\CTR.time_out[11] ),
    .X(\MEM.next_mem2[11] ));
 sky130_fd_sc_hd__and4_1 _0713_ (.A(\MEM.addr[0] ),
    .B(_0241_),
    .C(_0230_),
    .D(_0242_),
    .X(_0245_));
 sky130_fd_sc_hd__buf_4 _0714_ (.A(_0245_),
    .X(_0246_));
 sky130_fd_sc_hd__nor2_4 _0715_ (.A(_0236_),
    .B(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__a22o_1 _0716_ (.A1(_0229_),
    .A2(_0246_),
    .B1(_0247_),
    .B2(net80),
    .X(\MEM.next_mem3[0] ));
 sky130_fd_sc_hd__a22o_1 _0717_ (.A1(_0200_),
    .A2(_0246_),
    .B1(_0247_),
    .B2(net92),
    .X(\MEM.next_mem3[1] ));
 sky130_fd_sc_hd__a22o_1 _0718_ (.A1(\CTR.time_out[2] ),
    .A2(_0246_),
    .B1(_0247_),
    .B2(net76),
    .X(\MEM.next_mem3[2] ));
 sky130_fd_sc_hd__a22o_1 _0719_ (.A1(_0189_),
    .A2(_0246_),
    .B1(_0247_),
    .B2(net77),
    .X(\MEM.next_mem3[3] ));
 sky130_fd_sc_hd__a22o_1 _0720_ (.A1(\CTR.time_out[4] ),
    .A2(_0246_),
    .B1(_0247_),
    .B2(net65),
    .X(\MEM.next_mem3[4] ));
 sky130_fd_sc_hd__a22o_1 _0721_ (.A1(\CTR.time_out[5] ),
    .A2(_0246_),
    .B1(_0247_),
    .B2(net59),
    .X(\MEM.next_mem3[5] ));
 sky130_fd_sc_hd__a22o_1 _0722_ (.A1(\CTR.time_out[6] ),
    .A2(_0246_),
    .B1(_0247_),
    .B2(net62),
    .X(\MEM.next_mem3[6] ));
 sky130_fd_sc_hd__a22o_1 _0723_ (.A1(\CTR.time_out[7] ),
    .A2(_0246_),
    .B1(_0247_),
    .B2(net54),
    .X(\MEM.next_mem3[7] ));
 sky130_fd_sc_hd__a22o_1 _0724_ (.A1(\CTR.time_out[8] ),
    .A2(_0246_),
    .B1(_0247_),
    .B2(net56),
    .X(\MEM.next_mem3[8] ));
 sky130_fd_sc_hd__a22o_1 _0725_ (.A1(\CTR.time_out[9] ),
    .A2(_0246_),
    .B1(_0247_),
    .B2(net68),
    .X(\MEM.next_mem3[9] ));
 sky130_fd_sc_hd__a22o_1 _0726_ (.A1(\CTR.time_out[10] ),
    .A2(_0246_),
    .B1(_0247_),
    .B2(net84),
    .X(\MEM.next_mem3[10] ));
 sky130_fd_sc_hd__a22o_1 _0727_ (.A1(\CTR.time_out[11] ),
    .A2(_0246_),
    .B1(_0247_),
    .B2(net66),
    .X(\MEM.next_mem3[11] ));
 sky130_fd_sc_hd__and4b_1 _0728_ (.A_N(\MEM.addr[0] ),
    .B(\MEM.addr[1] ),
    .C(_0230_),
    .D(_0242_),
    .X(_0248_));
 sky130_fd_sc_hd__buf_4 _0729_ (.A(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__nor2_4 _0730_ (.A(_0236_),
    .B(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hd__a22o_1 _0731_ (.A1(_0229_),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net72),
    .X(\MEM.next_mem4[0] ));
 sky130_fd_sc_hd__a22o_1 _0732_ (.A1(_0200_),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net85),
    .X(\MEM.next_mem4[1] ));
 sky130_fd_sc_hd__a22o_1 _0733_ (.A1(\CTR.time_out[2] ),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net63),
    .X(\MEM.next_mem4[2] ));
 sky130_fd_sc_hd__a22o_1 _0734_ (.A1(_0189_),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net104),
    .X(\MEM.next_mem4[3] ));
 sky130_fd_sc_hd__a22o_1 _0735_ (.A1(\CTR.time_out[4] ),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net107),
    .X(\MEM.next_mem4[4] ));
 sky130_fd_sc_hd__a22o_1 _0736_ (.A1(\CTR.time_out[5] ),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net70),
    .X(\MEM.next_mem4[5] ));
 sky130_fd_sc_hd__a22o_1 _0737_ (.A1(\CTR.time_out[6] ),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net74),
    .X(\MEM.next_mem4[6] ));
 sky130_fd_sc_hd__a22o_1 _0738_ (.A1(\CTR.time_out[7] ),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net79),
    .X(\MEM.next_mem4[7] ));
 sky130_fd_sc_hd__a22o_1 _0739_ (.A1(\CTR.time_out[8] ),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net67),
    .X(\MEM.next_mem4[8] ));
 sky130_fd_sc_hd__a22o_1 _0740_ (.A1(\CTR.time_out[9] ),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net69),
    .X(\MEM.next_mem4[9] ));
 sky130_fd_sc_hd__a22o_1 _0741_ (.A1(\CTR.time_out[10] ),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net81),
    .X(\MEM.next_mem4[10] ));
 sky130_fd_sc_hd__a22o_1 _0742_ (.A1(\CTR.time_out[11] ),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net53),
    .X(\MEM.next_mem4[11] ));
 sky130_fd_sc_hd__nand2_1 _0743_ (.A(\MEM.addr[0] ),
    .B(\MEM.addr[1] ),
    .Y(_0251_));
 sky130_fd_sc_hd__and3b_1 _0744_ (.A_N(_0251_),
    .B(_0230_),
    .C(_0242_),
    .X(_0252_));
 sky130_fd_sc_hd__buf_4 _0745_ (.A(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__nor2_4 _0746_ (.A(_0236_),
    .B(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__a22o_1 _0747_ (.A1(_0229_),
    .A2(_0253_),
    .B1(_0254_),
    .B2(net60),
    .X(\MEM.next_mem5[0] ));
 sky130_fd_sc_hd__a22o_1 _0748_ (.A1(_0200_),
    .A2(_0253_),
    .B1(_0254_),
    .B2(net103),
    .X(\MEM.next_mem5[1] ));
 sky130_fd_sc_hd__a22o_1 _0749_ (.A1(\CTR.time_out[2] ),
    .A2(_0253_),
    .B1(_0254_),
    .B2(net86),
    .X(\MEM.next_mem5[2] ));
 sky130_fd_sc_hd__a22o_1 _0750_ (.A1(_0189_),
    .A2(_0253_),
    .B1(_0254_),
    .B2(net95),
    .X(\MEM.next_mem5[3] ));
 sky130_fd_sc_hd__a22o_1 _0751_ (.A1(\CTR.time_out[4] ),
    .A2(_0253_),
    .B1(_0254_),
    .B2(net89),
    .X(\MEM.next_mem5[4] ));
 sky130_fd_sc_hd__a22o_1 _0752_ (.A1(\CTR.time_out[5] ),
    .A2(_0253_),
    .B1(_0254_),
    .B2(net75),
    .X(\MEM.next_mem5[5] ));
 sky130_fd_sc_hd__a22o_1 _0753_ (.A1(\CTR.time_out[6] ),
    .A2(_0253_),
    .B1(_0254_),
    .B2(net112),
    .X(\MEM.next_mem5[6] ));
 sky130_fd_sc_hd__a22o_1 _0754_ (.A1(\CTR.time_out[7] ),
    .A2(_0253_),
    .B1(_0254_),
    .B2(net82),
    .X(\MEM.next_mem5[7] ));
 sky130_fd_sc_hd__a22o_1 _0755_ (.A1(\CTR.time_out[8] ),
    .A2(_0253_),
    .B1(_0254_),
    .B2(net110),
    .X(\MEM.next_mem5[8] ));
 sky130_fd_sc_hd__a22o_1 _0756_ (.A1(\CTR.time_out[9] ),
    .A2(_0253_),
    .B1(_0254_),
    .B2(net61),
    .X(\MEM.next_mem5[9] ));
 sky130_fd_sc_hd__a22o_1 _0757_ (.A1(\CTR.time_out[10] ),
    .A2(_0253_),
    .B1(_0254_),
    .B2(net88),
    .X(\MEM.next_mem5[10] ));
 sky130_fd_sc_hd__a22o_1 _0758_ (.A1(\CTR.time_out[11] ),
    .A2(_0253_),
    .B1(_0254_),
    .B2(net71),
    .X(\MEM.next_mem5[11] ));
 sky130_fd_sc_hd__a221o_1 _0759_ (.A1(\MEM.mem5[0] ),
    .A2(_0075_),
    .B1(_0076_),
    .B2(\MEM.mem2[0] ),
    .C1(_0070_),
    .X(_0255_));
 sky130_fd_sc_hd__a221o_1 _0760_ (.A1(\MEM.mem4[0] ),
    .A2(_0078_),
    .B1(net33),
    .B2(\MEM.mem3[0] ),
    .C1(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__o211a_1 _0761_ (.A1(_0071_),
    .A2(\MEM.mem1[0] ),
    .B1(_0069_),
    .C1(_0256_),
    .X(_0257_));
 sky130_fd_sc_hd__a221o_2 _0762_ (.A1(\TIM.cnt[0] ),
    .A2(_0085_),
    .B1(net34),
    .B2(_0229_),
    .C1(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__inv_2 _0763_ (.A(_0258_),
    .Y(_0259_));
 sky130_fd_sc_hd__xnor2_2 _0764_ (.A(_0202_),
    .B(_0225_),
    .Y(_0260_));
 sky130_fd_sc_hd__and2_1 _0765_ (.A(_0259_),
    .B(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__o21ai_1 _0766_ (.A1(_0183_),
    .A2(_0191_),
    .B1(_0208_),
    .Y(_0262_));
 sky130_fd_sc_hd__a21o_1 _0767_ (.A1(_0196_),
    .A2(net12),
    .B1(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__and2_1 _0768_ (.A(_0210_),
    .B(_0211_),
    .X(_0264_));
 sky130_fd_sc_hd__nor2_1 _0769_ (.A(_0210_),
    .B(_0211_),
    .Y(_0265_));
 sky130_fd_sc_hd__o21ai_1 _0770_ (.A1(_0264_),
    .A2(_0265_),
    .B1(_0212_),
    .Y(_0266_));
 sky130_fd_sc_hd__and2b_1 _0771_ (.A_N(_0203_),
    .B(_0216_),
    .X(_0267_));
 sky130_fd_sc_hd__o31a_1 _0772_ (.A1(_0264_),
    .A2(_0265_),
    .A3(_0267_),
    .B1(_0220_),
    .X(_0268_));
 sky130_fd_sc_hd__a22o_1 _0773_ (.A1(_0212_),
    .A2(net17),
    .B1(_0266_),
    .B2(_0268_),
    .X(_0269_));
 sky130_fd_sc_hd__nor2_1 _0774_ (.A(_0209_),
    .B(_0267_),
    .Y(_0270_));
 sky130_fd_sc_hd__a211o_1 _0775_ (.A1(_0209_),
    .A2(_0269_),
    .B1(_0270_),
    .C1(_0218_),
    .X(_0271_));
 sky130_fd_sc_hd__o21a_1 _0776_ (.A1(_0223_),
    .A2(_0267_),
    .B1(_0217_),
    .X(_0272_));
 sky130_fd_sc_hd__a21oi_4 _0777_ (.A1(_0263_),
    .A2(_0271_),
    .B1(_0272_),
    .Y(_0273_));
 sky130_fd_sc_hd__nand2_1 _0778_ (.A(_0261_),
    .B(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__or3b_1 _0779_ (.A(_0259_),
    .B(_0273_),
    .C_N(_0260_),
    .X(_0275_));
 sky130_fd_sc_hd__nor2_1 _0780_ (.A(_0191_),
    .B(_0212_),
    .Y(_0276_));
 sky130_fd_sc_hd__nor2_1 _0781_ (.A(_0191_),
    .B(_0216_),
    .Y(_0277_));
 sky130_fd_sc_hd__a21oi_1 _0782_ (.A1(_0210_),
    .A2(_0216_),
    .B1(_0277_),
    .Y(_0278_));
 sky130_fd_sc_hd__o311a_1 _0783_ (.A1(_0276_),
    .A2(_0220_),
    .A3(_0223_),
    .B1(_0278_),
    .C1(_0209_),
    .X(_0279_));
 sky130_fd_sc_hd__nand2_1 _0784_ (.A(_0191_),
    .B(_0203_),
    .Y(_0280_));
 sky130_fd_sc_hd__or2_1 _0785_ (.A(_0191_),
    .B(_0203_),
    .X(_0281_));
 sky130_fd_sc_hd__and3_1 _0786_ (.A(_0208_),
    .B(_0280_),
    .C(_0281_),
    .X(_0282_));
 sky130_fd_sc_hd__o32a_1 _0787_ (.A1(_0217_),
    .A2(_0279_),
    .A3(_0282_),
    .B1(_0277_),
    .B2(_0262_),
    .X(_0283_));
 sky130_fd_sc_hd__a21oi_1 _0788_ (.A1(_0208_),
    .A2(_0265_),
    .B1(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__nor2_1 _0789_ (.A(_0224_),
    .B(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__a21o_1 _0790_ (.A1(_0274_),
    .A2(_0275_),
    .B1(_0285_),
    .X(net4));
 sky130_fd_sc_hd__xnor2_1 _0791_ (.A(_0258_),
    .B(_0260_),
    .Y(_0286_));
 sky130_fd_sc_hd__nand2_1 _0792_ (.A(_0273_),
    .B(_0286_),
    .Y(net5));
 sky130_fd_sc_hd__nor2_1 _0793_ (.A(_0260_),
    .B(_0273_),
    .Y(_0287_));
 sky130_fd_sc_hd__nand2_2 _0794_ (.A(_0259_),
    .B(_0287_),
    .Y(net6));
 sky130_fd_sc_hd__or2b_1 _0795_ (.A(_0286_),
    .B_N(_0273_),
    .X(_0288_));
 sky130_fd_sc_hd__a21o_1 _0796_ (.A1(_0275_),
    .A2(_0288_),
    .B1(_0285_),
    .X(net7));
 sky130_fd_sc_hd__a21oi_1 _0797_ (.A1(_0260_),
    .A2(_0273_),
    .B1(_0258_),
    .Y(net8));
 sky130_fd_sc_hd__or2_1 _0798_ (.A(_0259_),
    .B(_0260_),
    .X(_0289_));
 sky130_fd_sc_hd__a211o_1 _0799_ (.A1(_0273_),
    .A2(_0289_),
    .B1(_0285_),
    .C1(_0261_),
    .X(net9));
 sky130_fd_sc_hd__a211o_1 _0800_ (.A1(_0273_),
    .A2(_0289_),
    .B1(_0287_),
    .C1(_0285_),
    .X(net10));
 sky130_fd_sc_hd__nand2_1 _0801_ (.A(_0124_),
    .B(_0122_),
    .Y(_0290_));
 sky130_fd_sc_hd__or2_1 _0802_ (.A(_0103_),
    .B(_0111_),
    .X(_0291_));
 sky130_fd_sc_hd__o21ai_1 _0803_ (.A1(_0127_),
    .A2(_0290_),
    .B1(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__mux2_1 _0804_ (.A0(_0111_),
    .A1(_0292_),
    .S(_0133_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _0805_ (.A0(_0290_),
    .A1(_0293_),
    .S(_0125_),
    .X(_0294_));
 sky130_fd_sc_hd__nand2_1 _0806_ (.A(_0111_),
    .B(_0128_),
    .Y(_0295_));
 sky130_fd_sc_hd__o211ai_1 _0807_ (.A1(_0128_),
    .A2(_0294_),
    .B1(_0295_),
    .C1(net26),
    .Y(_0296_));
 sky130_fd_sc_hd__o211a_1 _0808_ (.A1(_0129_),
    .A2(_0290_),
    .B1(_0296_),
    .C1(_0131_),
    .X(_0297_));
 sky130_fd_sc_hd__xnor2_2 _0809_ (.A(_0121_),
    .B(_0134_),
    .Y(_0298_));
 sky130_fd_sc_hd__nor2_1 _0810_ (.A(_0297_),
    .B(_0298_),
    .Y(_0299_));
 sky130_fd_sc_hd__and3b_1 _0811_ (.A_N(_0129_),
    .B(_0122_),
    .C(_0113_),
    .X(_0300_));
 sky130_fd_sc_hd__a21oi_1 _0812_ (.A1(_0112_),
    .A2(_0291_),
    .B1(_0121_),
    .Y(_0301_));
 sky130_fd_sc_hd__and3_1 _0813_ (.A(_0088_),
    .B(_0113_),
    .C(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__nor2_1 _0814_ (.A(_0103_),
    .B(_0111_),
    .Y(_0303_));
 sky130_fd_sc_hd__a21oi_1 _0815_ (.A1(_0088_),
    .A2(_0111_),
    .B1(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__nand2_1 _0816_ (.A(_0121_),
    .B(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__a21oi_1 _0817_ (.A1(_0129_),
    .A2(_0305_),
    .B1(_0113_),
    .Y(_0306_));
 sky130_fd_sc_hd__o21a_1 _0818_ (.A1(_0302_),
    .A2(_0306_),
    .B1(net26),
    .X(_0307_));
 sky130_fd_sc_hd__o21a_1 _0819_ (.A1(_0300_),
    .A2(_0307_),
    .B1(_0131_),
    .X(_0308_));
 sky130_fd_sc_hd__a221o_1 _0820_ (.A1(\MEM.mem5[6] ),
    .A2(_0075_),
    .B1(_0076_),
    .B2(\MEM.mem2[6] ),
    .C1(_0070_),
    .X(_0309_));
 sky130_fd_sc_hd__a221o_1 _0821_ (.A1(\MEM.mem4[6] ),
    .A2(_0078_),
    .B1(_0079_),
    .B2(\MEM.mem3[6] ),
    .C1(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__o211a_1 _0822_ (.A1(_0071_),
    .A2(\MEM.mem1[6] ),
    .B1(_0069_),
    .C1(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__a221o_1 _0823_ (.A1(\TIM.cnt[6] ),
    .A2(_0085_),
    .B1(_0086_),
    .B2(\CTR.time_out[6] ),
    .C1(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__nor2_1 _0824_ (.A(_0298_),
    .B(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__nor2_1 _0825_ (.A(_0308_),
    .B(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__or4b_1 _0826_ (.A(_0297_),
    .B(_0298_),
    .C(_0308_),
    .D_N(_0312_),
    .X(_0315_));
 sky130_fd_sc_hd__o21a_1 _0827_ (.A1(_0299_),
    .A2(_0314_),
    .B1(_0315_),
    .X(net18));
 sky130_fd_sc_hd__nand2_1 _0828_ (.A(_0298_),
    .B(_0312_),
    .Y(_0316_));
 sky130_fd_sc_hd__and2b_1 _0829_ (.A_N(_0313_),
    .B(_0316_),
    .X(_0317_));
 sky130_fd_sc_hd__nand2_1 _0830_ (.A(_0297_),
    .B(_0317_),
    .Y(net19));
 sky130_fd_sc_hd__or3b_2 _0831_ (.A(_0297_),
    .B(_0312_),
    .C_N(_0298_),
    .X(_0318_));
 sky130_fd_sc_hd__clkbuf_1 _0832_ (.A(_0318_),
    .X(net20));
 sky130_fd_sc_hd__inv_2 _0833_ (.A(_0297_),
    .Y(_0319_));
 sky130_fd_sc_hd__o21a_1 _0834_ (.A1(_0319_),
    .A2(_0317_),
    .B1(_0315_),
    .X(net21));
 sky130_fd_sc_hd__o21ba_1 _0835_ (.A1(_0319_),
    .A2(_0298_),
    .B1_N(_0312_),
    .X(net22));
 sky130_fd_sc_hd__a211o_1 _0836_ (.A1(_0297_),
    .A2(_0316_),
    .B1(_0313_),
    .C1(_0308_),
    .X(net23));
 sky130_fd_sc_hd__inv_2 _0837_ (.A(_0308_),
    .Y(_0320_));
 sky130_fd_sc_hd__o2bb2a_2 _0838_ (.A1_N(_0299_),
    .A2_N(_0320_),
    .B1(_0316_),
    .B2(_0319_),
    .X(net24));
 sky130_fd_sc_hd__or2b_2 _0839_ (.A(\e2.edge_d ),
    .B_N(\e2.sync ),
    .X(_0321_));
 sky130_fd_sc_hd__and2b_1 _0840_ (.A_N(_0082_),
    .B(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__or2_1 _0841_ (.A(_0066_),
    .B(_0321_),
    .X(_0323_));
 sky130_fd_sc_hd__nor2_1 _0842_ (.A(_0238_),
    .B(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__a21o_1 _0843_ (.A1(_0066_),
    .A2(net34),
    .B1(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__or3b_2 _0844_ (.A(\FSM.state[2] ),
    .B(\FSM.state[1] ),
    .C_N(\FSM.state[3] ),
    .X(_0326_));
 sky130_fd_sc_hd__nor2_4 _0845_ (.A(_0066_),
    .B(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__nand2b_2 _0846_ (.A_N(\e1.edge_d ),
    .B(\e1.sync ),
    .Y(_0328_));
 sky130_fd_sc_hd__nor2_1 _0847_ (.A(_0066_),
    .B(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__and2b_1 _0848_ (.A_N(\e1.edge_d ),
    .B(\e1.sync ),
    .X(_0330_));
 sky130_fd_sc_hd__nor3b_1 _0849_ (.A(_0330_),
    .B(_0326_),
    .C_N(_0066_),
    .Y(_0331_));
 sky130_fd_sc_hd__a221o_1 _0850_ (.A1(net32),
    .A2(_0327_),
    .B1(_0234_),
    .B2(_0329_),
    .C1(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__or3_1 _0851_ (.A(_0067_),
    .B(_0321_),
    .C(_0330_),
    .X(_0333_));
 sky130_fd_sc_hd__or4b_1 _0852_ (.A(_0322_),
    .B(_0325_),
    .C(_0332_),
    .D_N(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__clkbuf_1 _0853_ (.A(_0334_),
    .X(\FSM.next_state[0] ));
 sky130_fd_sc_hd__or2b_2 _0854_ (.A(_0066_),
    .B_N(_0086_),
    .X(_0335_));
 sky130_fd_sc_hd__inv_2 _0855_ (.A(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__nor2_1 _0856_ (.A(_0067_),
    .B(_0330_),
    .Y(_0337_));
 sky130_fd_sc_hd__o22a_1 _0857_ (.A1(_0321_),
    .A2(_0330_),
    .B1(_0336_),
    .B2(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__a211o_1 _0858_ (.A1(_0066_),
    .A2(_0236_),
    .B1(_0322_),
    .C1(_0231_),
    .X(_0339_));
 sky130_fd_sc_hd__a211o_1 _0859_ (.A1(_0328_),
    .A2(_0325_),
    .B1(_0338_),
    .C1(_0339_),
    .X(\FSM.next_state[1] ));
 sky130_fd_sc_hd__and2_2 _0860_ (.A(_0066_),
    .B(_0231_),
    .X(_0340_));
 sky130_fd_sc_hd__or2_1 _0861_ (.A(_0066_),
    .B(_0328_),
    .X(_0341_));
 sky130_fd_sc_hd__nand2_1 _0862_ (.A(_0328_),
    .B(_0323_),
    .Y(_0342_));
 sky130_fd_sc_hd__a32o_1 _0863_ (.A1(net34),
    .A2(_0341_),
    .A3(_0342_),
    .B1(_0324_),
    .B2(_0328_),
    .X(_0343_));
 sky130_fd_sc_hd__or4_1 _0864_ (.A(_0340_),
    .B(_0322_),
    .C(_0337_),
    .D(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_1 _0865_ (.A(_0344_),
    .X(\FSM.next_state[2] ));
 sky130_fd_sc_hd__nor2_1 _0866_ (.A(_0082_),
    .B(_0321_),
    .Y(_0345_));
 sky130_fd_sc_hd__or3_1 _0867_ (.A(_0327_),
    .B(_0331_),
    .C(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__clkbuf_1 _0868_ (.A(_0346_),
    .X(\FSM.next_state[3] ));
 sky130_fd_sc_hd__nor2_1 _0869_ (.A(\TIM.cnt[6] ),
    .B(_0234_),
    .Y(_0347_));
 sky130_fd_sc_hd__a41o_1 _0870_ (.A1(\TIM.cnt[1] ),
    .A2(\TIM.cnt[3] ),
    .A3(\TIM.cnt[2] ),
    .A4(\TIM.cnt[4] ),
    .B1(\TIM.cnt[5] ),
    .X(_0348_));
 sky130_fd_sc_hd__inv_2 _0871_ (.A(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__or2_1 _0872_ (.A(\TIM.cnt[1] ),
    .B(\TIM.cnt[2] ),
    .X(_0350_));
 sky130_fd_sc_hd__or2_1 _0873_ (.A(\TIM.cnt[3] ),
    .B(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__or2_1 _0874_ (.A(\TIM.cnt[4] ),
    .B(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__nor3_1 _0875_ (.A(\TIM.cnt[0] ),
    .B(\TIM.cnt[5] ),
    .C(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hd__nand2_2 _0876_ (.A(_0327_),
    .B(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__or4_1 _0877_ (.A(\TIM.cnt[9] ),
    .B(\TIM.cnt[8] ),
    .C(\TIM.cnt[11] ),
    .D(\TIM.cnt[10] ),
    .X(_0355_));
 sky130_fd_sc_hd__or4_1 _0878_ (.A(\TIM.cnt[7] ),
    .B(\TIM.cnt[6] ),
    .C(_0354_),
    .D(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__o221a_1 _0879_ (.A1(_0085_),
    .A2(_0236_),
    .B1(_0330_),
    .B2(_0082_),
    .C1(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__o21ai_4 _0880_ (.A1(\CLKDIV.secpulse ),
    .A2(_0354_),
    .B1(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__a31o_1 _0881_ (.A1(_0084_),
    .A2(_0238_),
    .A3(_0349_),
    .B1(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__or2_2 _0882_ (.A(_0084_),
    .B(_0353_),
    .X(_0360_));
 sky130_fd_sc_hd__or2b_1 _0883_ (.A(_0359_),
    .B_N(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__buf_2 _0884_ (.A(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _0885_ (.A0(_0347_),
    .A1(\TIM.cnt[6] ),
    .S(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__clkbuf_1 _0886_ (.A(_0363_),
    .X(_0025_));
 sky130_fd_sc_hd__nor2_1 _0887_ (.A(_0236_),
    .B(_0362_),
    .Y(_0364_));
 sky130_fd_sc_hd__or2_1 _0888_ (.A(\TIM.cnt[7] ),
    .B(_0327_),
    .X(_0365_));
 sky130_fd_sc_hd__nand2_1 _0889_ (.A(\TIM.cnt[7] ),
    .B(_0327_),
    .Y(_0366_));
 sky130_fd_sc_hd__a21o_1 _0890_ (.A1(_0365_),
    .A2(_0366_),
    .B1(\TIM.cnt[6] ),
    .X(_0367_));
 sky130_fd_sc_hd__nand3_1 _0891_ (.A(\TIM.cnt[6] ),
    .B(_0365_),
    .C(_0366_),
    .Y(_0368_));
 sky130_fd_sc_hd__a32o_1 _0892_ (.A1(_0364_),
    .A2(_0367_),
    .A3(_0368_),
    .B1(_0362_),
    .B2(net134),
    .X(_0026_));
 sky130_fd_sc_hd__nor2_1 _0893_ (.A(\TIM.cnt[8] ),
    .B(_0327_),
    .Y(_0369_));
 sky130_fd_sc_hd__and2_1 _0894_ (.A(\TIM.cnt[8] ),
    .B(_0327_),
    .X(_0370_));
 sky130_fd_sc_hd__o211a_1 _0895_ (.A1(_0369_),
    .A2(_0370_),
    .B1(_0366_),
    .C1(_0368_),
    .X(_0371_));
 sky130_fd_sc_hd__a211oi_1 _0896_ (.A1(_0366_),
    .A2(_0368_),
    .B1(_0369_),
    .C1(_0370_),
    .Y(_0372_));
 sky130_fd_sc_hd__nor2_1 _0897_ (.A(_0371_),
    .B(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__a22o_1 _0898_ (.A1(net136),
    .A2(_0362_),
    .B1(_0364_),
    .B2(_0373_),
    .X(_0027_));
 sky130_fd_sc_hd__nor2_1 _0899_ (.A(\TIM.cnt[9] ),
    .B(_0327_),
    .Y(_0374_));
 sky130_fd_sc_hd__and2_1 _0900_ (.A(\TIM.cnt[9] ),
    .B(_0327_),
    .X(_0375_));
 sky130_fd_sc_hd__or2_1 _0901_ (.A(_0370_),
    .B(_0372_),
    .X(_0376_));
 sky130_fd_sc_hd__o21bai_1 _0902_ (.A1(_0374_),
    .A2(_0375_),
    .B1_N(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__or3b_1 _0903_ (.A(_0374_),
    .B(_0375_),
    .C_N(_0376_),
    .X(_0378_));
 sky130_fd_sc_hd__a32o_1 _0904_ (.A1(_0364_),
    .A2(_0377_),
    .A3(_0378_),
    .B1(_0362_),
    .B2(net127),
    .X(_0028_));
 sky130_fd_sc_hd__and2b_1 _0905_ (.A_N(_0374_),
    .B(_0376_),
    .X(_0379_));
 sky130_fd_sc_hd__or2_1 _0906_ (.A(\TIM.cnt[10] ),
    .B(_0327_),
    .X(_0380_));
 sky130_fd_sc_hd__nand2_2 _0907_ (.A(\TIM.cnt[10] ),
    .B(_0327_),
    .Y(_0381_));
 sky130_fd_sc_hd__o211ai_2 _0908_ (.A1(_0375_),
    .A2(_0379_),
    .B1(_0380_),
    .C1(_0381_),
    .Y(_0382_));
 sky130_fd_sc_hd__a211o_1 _0909_ (.A1(_0381_),
    .A2(_0380_),
    .B1(_0379_),
    .C1(_0375_),
    .X(_0383_));
 sky130_fd_sc_hd__a32o_1 _0910_ (.A1(_0364_),
    .A2(_0382_),
    .A3(_0383_),
    .B1(_0362_),
    .B2(net128),
    .X(_0029_));
 sky130_fd_sc_hd__xor2_1 _0911_ (.A(\TIM.cnt[11] ),
    .B(_0084_),
    .X(_0384_));
 sky130_fd_sc_hd__a21oi_1 _0912_ (.A1(_0381_),
    .A2(_0382_),
    .B1(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__a311o_1 _0913_ (.A1(_0381_),
    .A2(_0382_),
    .A3(_0384_),
    .B1(_0362_),
    .C1(_0236_),
    .X(_0386_));
 sky130_fd_sc_hd__a2bb2o_1 _0914_ (.A1_N(_0385_),
    .A2_N(_0386_),
    .B1(net133),
    .B2(_0362_),
    .X(_0030_));
 sky130_fd_sc_hd__and4_1 _0915_ (.A(_0189_),
    .B(\CTR.time_out[2] ),
    .C(\CTR.time_out[5] ),
    .D(\CTR.time_out[4] ),
    .X(_0387_));
 sky130_fd_sc_hd__nor3b_1 _0916_ (.A(_0200_),
    .B(_0229_),
    .C_N(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__nor2_2 _0917_ (.A(_0335_),
    .B(_0387_),
    .Y(_0389_));
 sky130_fd_sc_hd__nor2_1 _0918_ (.A(_0236_),
    .B(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__o21a_1 _0919_ (.A1(net118),
    .A2(_0388_),
    .B1(_0390_),
    .X(_0031_));
 sky130_fd_sc_hd__and2_1 _0920_ (.A(\CTR.minutes ),
    .B(_0336_),
    .X(_0391_));
 sky130_fd_sc_hd__nor2_1 _0921_ (.A(_0236_),
    .B(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__mux2_1 _0922_ (.A0(_0391_),
    .A1(_0392_),
    .S(\CTR.time_out[6] ),
    .X(_0393_));
 sky130_fd_sc_hd__clkbuf_1 _0923_ (.A(_0393_),
    .X(_0032_));
 sky130_fd_sc_hd__or2_1 _0924_ (.A(\CTR.time_out[7] ),
    .B(\CTR.time_out[6] ),
    .X(_0394_));
 sky130_fd_sc_hd__nand2_1 _0925_ (.A(\CTR.time_out[7] ),
    .B(\CTR.time_out[6] ),
    .Y(_0395_));
 sky130_fd_sc_hd__a32o_1 _0926_ (.A1(_0391_),
    .A2(_0394_),
    .A3(_0395_),
    .B1(_0392_),
    .B2(\CTR.time_out[7] ),
    .X(_0033_));
 sky130_fd_sc_hd__or2_1 _0927_ (.A(_0236_),
    .B(_0391_),
    .X(_0396_));
 sky130_fd_sc_hd__a31o_1 _0928_ (.A1(\CTR.time_out[7] ),
    .A2(\CTR.time_out[6] ),
    .A3(_0396_),
    .B1(\CTR.time_out[8] ),
    .X(_0397_));
 sky130_fd_sc_hd__and4_1 _0929_ (.A(\CTR.time_out[7] ),
    .B(\CTR.time_out[6] ),
    .C(\CTR.time_out[8] ),
    .D(_0396_),
    .X(_0398_));
 sky130_fd_sc_hd__inv_2 _0930_ (.A(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__and3_1 _0931_ (.A(_0238_),
    .B(_0397_),
    .C(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__clkbuf_1 _0932_ (.A(_0400_),
    .X(_0034_));
 sky130_fd_sc_hd__and2_1 _0933_ (.A(\CTR.time_out[9] ),
    .B(_0398_),
    .X(_0401_));
 sky130_fd_sc_hd__nor2_1 _0934_ (.A(_0236_),
    .B(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__o21a_1 _0935_ (.A1(\CTR.time_out[9] ),
    .A2(_0398_),
    .B1(_0402_),
    .X(_0035_));
 sky130_fd_sc_hd__and3_1 _0936_ (.A(\CTR.time_out[10] ),
    .B(\CTR.time_out[9] ),
    .C(_0398_),
    .X(_0403_));
 sky130_fd_sc_hd__nor2_1 _0937_ (.A(_0236_),
    .B(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__o21a_1 _0938_ (.A1(\CTR.time_out[10] ),
    .A2(_0401_),
    .B1(_0404_),
    .X(_0036_));
 sky130_fd_sc_hd__o21ai_1 _0939_ (.A1(\CTR.time_out[11] ),
    .A2(_0403_),
    .B1(_0238_),
    .Y(_0405_));
 sky130_fd_sc_hd__a21oi_1 _0940_ (.A1(net130),
    .A2(_0403_),
    .B1(_0405_),
    .Y(_0037_));
 sky130_fd_sc_hd__nor2_2 _0941_ (.A(_0236_),
    .B(_0358_),
    .Y(_0406_));
 sky130_fd_sc_hd__inv_2 _0942_ (.A(\CLKDIV.secpulse ),
    .Y(_0407_));
 sky130_fd_sc_hd__o21a_1 _0943_ (.A1(\TIM.cnt[0] ),
    .A2(_0407_),
    .B1(\TIM.cnt[1] ),
    .X(_0408_));
 sky130_fd_sc_hd__or3_1 _0944_ (.A(\TIM.cnt[0] ),
    .B(\TIM.cnt[1] ),
    .C(_0407_),
    .X(_0409_));
 sky130_fd_sc_hd__or3b_1 _0945_ (.A(_0360_),
    .B(_0408_),
    .C_N(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__o21ai_1 _0946_ (.A1(\TIM.cnt[1] ),
    .A2(\TIM.cnt[5] ),
    .B1(_0084_),
    .Y(_0411_));
 sky130_fd_sc_hd__a32o_1 _0947_ (.A1(_0406_),
    .A2(_0410_),
    .A3(_0411_),
    .B1(_0358_),
    .B2(net137),
    .X(_0038_));
 sky130_fd_sc_hd__nand2_1 _0948_ (.A(\TIM.cnt[1] ),
    .B(\TIM.cnt[2] ),
    .Y(_0412_));
 sky130_fd_sc_hd__a21o_1 _0949_ (.A1(_0350_),
    .A2(_0412_),
    .B1(_0348_),
    .X(_0413_));
 sky130_fd_sc_hd__nand2_1 _0950_ (.A(\TIM.cnt[2] ),
    .B(_0409_),
    .Y(_0414_));
 sky130_fd_sc_hd__or2_1 _0951_ (.A(\TIM.cnt[2] ),
    .B(_0409_),
    .X(_0415_));
 sky130_fd_sc_hd__and3_1 _0952_ (.A(_0327_),
    .B(_0414_),
    .C(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__a21oi_1 _0953_ (.A1(_0084_),
    .A2(_0413_),
    .B1(_0416_),
    .Y(_0417_));
 sky130_fd_sc_hd__a32o_1 _0954_ (.A1(_0354_),
    .A2(_0406_),
    .A3(_0417_),
    .B1(_0358_),
    .B2(net132),
    .X(_0039_));
 sky130_fd_sc_hd__a21oi_1 _0955_ (.A1(\TIM.cnt[3] ),
    .A2(_0415_),
    .B1(_0360_),
    .Y(_0418_));
 sky130_fd_sc_hd__o21ai_1 _0956_ (.A1(\TIM.cnt[3] ),
    .A2(_0415_),
    .B1(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__nand2_1 _0957_ (.A(\TIM.cnt[3] ),
    .B(_0350_),
    .Y(_0420_));
 sky130_fd_sc_hd__a21o_1 _0958_ (.A1(_0351_),
    .A2(_0420_),
    .B1(_0348_),
    .X(_0421_));
 sky130_fd_sc_hd__nand2_1 _0959_ (.A(_0084_),
    .B(_0421_),
    .Y(_0422_));
 sky130_fd_sc_hd__a32o_1 _0960_ (.A1(_0406_),
    .A2(_0419_),
    .A3(_0422_),
    .B1(_0358_),
    .B2(\TIM.cnt[3] ),
    .X(_0040_));
 sky130_fd_sc_hd__or3_1 _0961_ (.A(\TIM.cnt[3] ),
    .B(\TIM.cnt[4] ),
    .C(_0415_),
    .X(_0423_));
 sky130_fd_sc_hd__inv_2 _0962_ (.A(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__o21a_1 _0963_ (.A1(\TIM.cnt[3] ),
    .A2(_0415_),
    .B1(\TIM.cnt[4] ),
    .X(_0425_));
 sky130_fd_sc_hd__nand2_1 _0964_ (.A(\TIM.cnt[4] ),
    .B(_0351_),
    .Y(_0426_));
 sky130_fd_sc_hd__a21oi_1 _0965_ (.A1(_0352_),
    .A2(_0426_),
    .B1(_0348_),
    .Y(_0427_));
 sky130_fd_sc_hd__o32a_1 _0966_ (.A1(_0360_),
    .A2(_0424_),
    .A3(_0425_),
    .B1(_0427_),
    .B2(_0327_),
    .X(_0428_));
 sky130_fd_sc_hd__a22o_1 _0967_ (.A1(\TIM.cnt[4] ),
    .A2(_0358_),
    .B1(_0406_),
    .B2(_0428_),
    .X(_0041_));
 sky130_fd_sc_hd__a21o_1 _0968_ (.A1(\TIM.cnt[5] ),
    .A2(_0423_),
    .B1(_0360_),
    .X(_0429_));
 sky130_fd_sc_hd__a21o_1 _0969_ (.A1(_0352_),
    .A2(_0349_),
    .B1(_0327_),
    .X(_0430_));
 sky130_fd_sc_hd__a32o_1 _0970_ (.A1(_0406_),
    .A2(_0429_),
    .A3(_0430_),
    .B1(_0358_),
    .B2(net129),
    .X(_0042_));
 sky130_fd_sc_hd__a21bo_1 _0971_ (.A1(net117),
    .A2(_0238_),
    .B1_N(_0356_),
    .X(_0043_));
 sky130_fd_sc_hd__or2_1 _0972_ (.A(\FSM.state[3] ),
    .B(\FSM.state[1] ),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _0973_ (.A0(_0231_),
    .A1(_0431_),
    .S(_0073_),
    .X(_0432_));
 sky130_fd_sc_hd__a41o_1 _0974_ (.A1(_0070_),
    .A2(\MEM.addr[0] ),
    .A3(_0340_),
    .A4(_0075_),
    .B1(_0432_),
    .X(_0044_));
 sky130_fd_sc_hd__nand2_1 _0975_ (.A(_0070_),
    .B(_0075_),
    .Y(_0433_));
 sky130_fd_sc_hd__o221a_1 _0976_ (.A1(\MEM.addr[1] ),
    .A2(_0433_),
    .B1(_0076_),
    .B2(_0075_),
    .C1(_0340_),
    .X(_0434_));
 sky130_fd_sc_hd__nor3_1 _0977_ (.A(_0075_),
    .B(_0076_),
    .C(_0232_),
    .Y(_0435_));
 sky130_fd_sc_hd__a211o_1 _0978_ (.A1(_0072_),
    .A2(_0431_),
    .B1(_0434_),
    .C1(_0435_),
    .X(_0045_));
 sky130_fd_sc_hd__or2_1 _0979_ (.A(_0070_),
    .B(_0075_),
    .X(_0436_));
 sky130_fd_sc_hd__a21oi_1 _0980_ (.A1(_0230_),
    .A2(_0075_),
    .B1(_0076_),
    .Y(_0437_));
 sky130_fd_sc_hd__a21o_1 _0981_ (.A1(_0340_),
    .A2(_0437_),
    .B1(_0431_),
    .X(_0438_));
 sky130_fd_sc_hd__a32o_1 _0982_ (.A1(_0433_),
    .A2(_0436_),
    .A3(_0242_),
    .B1(_0438_),
    .B2(_0070_),
    .X(_0439_));
 sky130_fd_sc_hd__a31o_1 _0983_ (.A1(_0071_),
    .A2(_0340_),
    .A3(_0076_),
    .B1(_0439_),
    .X(_0046_));
 sky130_fd_sc_hd__xor2_1 _0984_ (.A(\TIM.cnt[0] ),
    .B(\CLKDIV.secpulse ),
    .X(_0440_));
 sky130_fd_sc_hd__o21a_1 _0985_ (.A1(_0353_),
    .A2(_0440_),
    .B1(_0327_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _0986_ (.A0(_0441_),
    .A1(\TIM.cnt[0] ),
    .S(_0359_),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_1 _0987_ (.A(_0442_),
    .X(_0047_));
 sky130_fd_sc_hd__nor2_1 _0988_ (.A(_0242_),
    .B(_0236_),
    .Y(_0443_));
 sky130_fd_sc_hd__nor2_1 _0989_ (.A(\MEM.addr[0] ),
    .B(_0232_),
    .Y(_0444_));
 sky130_fd_sc_hd__a21o_1 _0990_ (.A1(net135),
    .A2(_0443_),
    .B1(_0444_),
    .X(_0048_));
 sky130_fd_sc_hd__o21a_1 _0991_ (.A1(_0443_),
    .A2(_0444_),
    .B1(\MEM.addr[1] ),
    .X(_0445_));
 sky130_fd_sc_hd__a31o_1 _0992_ (.A1(\MEM.addr[0] ),
    .A2(_0241_),
    .A3(_0242_),
    .B1(_0445_),
    .X(_0049_));
 sky130_fd_sc_hd__xnor2_1 _0993_ (.A(\MEM.addr[2] ),
    .B(_0251_),
    .Y(_0446_));
 sky130_fd_sc_hd__a22o_1 _0994_ (.A1(\MEM.addr[2] ),
    .A2(_0443_),
    .B1(_0446_),
    .B2(_0242_),
    .X(_0050_));
 sky130_fd_sc_hd__or2_1 _0995_ (.A(_0229_),
    .B(\CLKDIV.secpulse ),
    .X(_0447_));
 sky130_fd_sc_hd__nand2_1 _0996_ (.A(_0229_),
    .B(\CLKDIV.secpulse ),
    .Y(_0448_));
 sky130_fd_sc_hd__a32o_1 _0997_ (.A1(_0389_),
    .A2(_0447_),
    .A3(_0448_),
    .B1(_0390_),
    .B2(_0229_),
    .X(_0051_));
 sky130_fd_sc_hd__a21o_1 _0998_ (.A1(_0229_),
    .A2(\CLKDIV.secpulse ),
    .B1(_0200_),
    .X(_0449_));
 sky130_fd_sc_hd__nand3_1 _0999_ (.A(_0200_),
    .B(_0229_),
    .C(\CLKDIV.secpulse ),
    .Y(_0450_));
 sky130_fd_sc_hd__a32o_1 _1000_ (.A1(_0389_),
    .A2(_0449_),
    .A3(_0450_),
    .B1(_0390_),
    .B2(_0200_),
    .X(_0052_));
 sky130_fd_sc_hd__a31o_1 _1001_ (.A1(_0200_),
    .A2(_0229_),
    .A3(\CLKDIV.secpulse ),
    .B1(\CTR.time_out[2] ),
    .X(_0451_));
 sky130_fd_sc_hd__and4_1 _1002_ (.A(_0200_),
    .B(_0229_),
    .C(\CTR.time_out[2] ),
    .D(\CLKDIV.secpulse ),
    .X(_0452_));
 sky130_fd_sc_hd__inv_2 _1003_ (.A(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__and2b_1 _1004_ (.A_N(_0388_),
    .B(_0390_),
    .X(_0454_));
 sky130_fd_sc_hd__a32o_1 _1005_ (.A1(_0389_),
    .A2(_0451_),
    .A3(_0453_),
    .B1(_0454_),
    .B2(\CTR.time_out[2] ),
    .X(_0053_));
 sky130_fd_sc_hd__or2_1 _1006_ (.A(_0189_),
    .B(_0452_),
    .X(_0455_));
 sky130_fd_sc_hd__nand2_1 _1007_ (.A(_0189_),
    .B(_0452_),
    .Y(_0456_));
 sky130_fd_sc_hd__a32o_1 _1008_ (.A1(_0389_),
    .A2(_0455_),
    .A3(_0456_),
    .B1(_0454_),
    .B2(_0189_),
    .X(_0054_));
 sky130_fd_sc_hd__nand3_1 _1009_ (.A(_0189_),
    .B(\CTR.time_out[4] ),
    .C(_0452_),
    .Y(_0457_));
 sky130_fd_sc_hd__a21o_1 _1010_ (.A1(_0389_),
    .A2(_0457_),
    .B1(_0454_),
    .X(_0458_));
 sky130_fd_sc_hd__or4_1 _1011_ (.A(\CTR.time_out[4] ),
    .B(_0335_),
    .C(_0387_),
    .D(_0456_),
    .X(_0459_));
 sky130_fd_sc_hd__a21bo_1 _1012_ (.A1(\CTR.time_out[4] ),
    .A2(_0458_),
    .B1_N(_0459_),
    .X(_0055_));
 sky130_fd_sc_hd__nor2_1 _1013_ (.A(_0335_),
    .B(_0457_),
    .Y(_0460_));
 sky130_fd_sc_hd__mux2_1 _1014_ (.A0(_0460_),
    .A1(_0458_),
    .S(\CTR.time_out[5] ),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_1 _1015_ (.A(_0461_),
    .X(_0056_));
 sky130_fd_sc_hd__dfrtp_1 _1016_ (.CLK(clknet_4_1_0_clk),
    .D(net42),
    .RESET_B(net35),
    .Q(\e1.sync ));
 sky130_fd_sc_hd__dfrtp_1 _1017_ (.CLK(clknet_4_8_0_clk),
    .D(net45),
    .RESET_B(net40),
    .Q(\e1.edge_d ));
 sky130_fd_sc_hd__dfrtp_1 _1018_ (.CLK(clknet_4_1_0_clk),
    .D(net2),
    .RESET_B(net35),
    .Q(\e1.intermediate ));
 sky130_fd_sc_hd__dfrtp_1 _1019_ (.CLK(clknet_4_5_0_clk),
    .D(net43),
    .RESET_B(net37),
    .Q(\e2.sync ));
 sky130_fd_sc_hd__dfrtp_1 _1020_ (.CLK(clknet_4_5_0_clk),
    .D(net44),
    .RESET_B(net38),
    .Q(\e2.edge_d ));
 sky130_fd_sc_hd__dfrtp_1 _1021_ (.CLK(clknet_4_5_0_clk),
    .D(net3),
    .RESET_B(net37),
    .Q(\e2.intermediate ));
 sky130_fd_sc_hd__dfrtp_4 _1022_ (.CLK(clknet_4_15_0_clk),
    .D(_0024_),
    .RESET_B(net39),
    .Q(\CLKDIV.secpulse ));
 sky130_fd_sc_hd__dfrtp_1 _1023_ (.CLK(clknet_4_7_0_clk),
    .D(_0000_),
    .RESET_B(net37),
    .Q(\CLKDIV.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1024_ (.CLK(clknet_4_5_0_clk),
    .D(_0011_),
    .RESET_B(net37),
    .Q(\CLKDIV.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1025_ (.CLK(clknet_4_5_0_clk),
    .D(_0016_),
    .RESET_B(net37),
    .Q(\CLKDIV.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1026_ (.CLK(clknet_4_5_0_clk),
    .D(_0017_),
    .RESET_B(net37),
    .Q(\CLKDIV.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1027_ (.CLK(clknet_4_5_0_clk),
    .D(_0018_),
    .RESET_B(net37),
    .Q(\CLKDIV.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1028_ (.CLK(clknet_4_5_0_clk),
    .D(_0019_),
    .RESET_B(net37),
    .Q(\CLKDIV.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1029_ (.CLK(clknet_4_5_0_clk),
    .D(_0020_),
    .RESET_B(net37),
    .Q(\CLKDIV.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1030_ (.CLK(clknet_4_5_0_clk),
    .D(_0021_),
    .RESET_B(net37),
    .Q(\CLKDIV.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1031_ (.CLK(clknet_4_5_0_clk),
    .D(_0022_),
    .RESET_B(net41),
    .Q(\CLKDIV.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1032_ (.CLK(clknet_4_5_0_clk),
    .D(_0023_),
    .RESET_B(net38),
    .Q(\CLKDIV.count[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1033_ (.CLK(clknet_4_7_0_clk),
    .D(_0001_),
    .RESET_B(net38),
    .Q(\CLKDIV.count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1034_ (.CLK(clknet_4_13_0_clk),
    .D(_0002_),
    .RESET_B(net38),
    .Q(\CLKDIV.count[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1035_ (.CLK(clknet_4_7_0_clk),
    .D(_0003_),
    .RESET_B(net38),
    .Q(\CLKDIV.count[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1036_ (.CLK(clknet_4_7_0_clk),
    .D(_0004_),
    .RESET_B(net38),
    .Q(\CLKDIV.count[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1037_ (.CLK(clknet_4_13_0_clk),
    .D(_0005_),
    .RESET_B(net38),
    .Q(\CLKDIV.count[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1038_ (.CLK(clknet_4_13_0_clk),
    .D(_0006_),
    .RESET_B(net38),
    .Q(\CLKDIV.count[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1039_ (.CLK(clknet_4_14_0_clk),
    .D(_0007_),
    .RESET_B(net39),
    .Q(\CLKDIV.count[16] ));
 sky130_fd_sc_hd__dfrtp_1 _1040_ (.CLK(clknet_4_14_0_clk),
    .D(_0008_),
    .RESET_B(net39),
    .Q(\CLKDIV.count[17] ));
 sky130_fd_sc_hd__dfrtp_1 _1041_ (.CLK(clknet_4_14_0_clk),
    .D(_0009_),
    .RESET_B(net39),
    .Q(\CLKDIV.count[18] ));
 sky130_fd_sc_hd__dfrtp_1 _1042_ (.CLK(clknet_4_15_0_clk),
    .D(_0010_),
    .RESET_B(net39),
    .Q(\CLKDIV.count[19] ));
 sky130_fd_sc_hd__dfrtp_1 _1043_ (.CLK(clknet_4_15_0_clk),
    .D(_0012_),
    .RESET_B(net39),
    .Q(\CLKDIV.count[20] ));
 sky130_fd_sc_hd__dfrtp_1 _1044_ (.CLK(clknet_4_15_0_clk),
    .D(_0013_),
    .RESET_B(net39),
    .Q(\CLKDIV.count[21] ));
 sky130_fd_sc_hd__dfrtp_1 _1045_ (.CLK(clknet_4_15_0_clk),
    .D(_0014_),
    .RESET_B(net41),
    .Q(\CLKDIV.count[22] ));
 sky130_fd_sc_hd__dfrtp_1 _1046_ (.CLK(clknet_4_15_0_clk),
    .D(_0015_),
    .RESET_B(net39),
    .Q(\CLKDIV.count[23] ));
 sky130_fd_sc_hd__dfrtp_2 _1047_ (.CLK(clknet_4_10_0_clk),
    .D(_0025_),
    .RESET_B(net40),
    .Q(\TIM.cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1048_ (.CLK(clknet_4_10_0_clk),
    .D(_0026_),
    .RESET_B(net40),
    .Q(\TIM.cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1049_ (.CLK(clknet_4_10_0_clk),
    .D(_0027_),
    .RESET_B(net40),
    .Q(\TIM.cnt[8] ));
 sky130_fd_sc_hd__dfrtp_2 _1050_ (.CLK(clknet_4_10_0_clk),
    .D(_0028_),
    .RESET_B(net40),
    .Q(\TIM.cnt[9] ));
 sky130_fd_sc_hd__dfrtp_2 _1051_ (.CLK(clknet_4_10_0_clk),
    .D(_0029_),
    .RESET_B(net40),
    .Q(\TIM.cnt[10] ));
 sky130_fd_sc_hd__dfrtp_2 _1052_ (.CLK(clknet_4_10_0_clk),
    .D(_0030_),
    .RESET_B(net40),
    .Q(\TIM.cnt[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1053_ (.CLK(clknet_4_12_0_clk),
    .D(_0031_),
    .RESET_B(net39),
    .Q(\CTR.minutes ));
 sky130_fd_sc_hd__dfrtp_4 _1054_ (.CLK(clknet_4_1_0_clk),
    .D(_0032_),
    .RESET_B(net35),
    .Q(\CTR.time_out[6] ));
 sky130_fd_sc_hd__dfrtp_4 _1055_ (.CLK(clknet_4_1_0_clk),
    .D(_0033_),
    .RESET_B(net35),
    .Q(\CTR.time_out[7] ));
 sky130_fd_sc_hd__dfrtp_4 _1056_ (.CLK(clknet_4_2_0_clk),
    .D(_0034_),
    .RESET_B(net36),
    .Q(\CTR.time_out[8] ));
 sky130_fd_sc_hd__dfrtp_4 _1057_ (.CLK(clknet_4_2_0_clk),
    .D(_0035_),
    .RESET_B(net36),
    .Q(\CTR.time_out[9] ));
 sky130_fd_sc_hd__dfrtp_4 _1058_ (.CLK(clknet_4_2_0_clk),
    .D(_0036_),
    .RESET_B(net36),
    .Q(\CTR.time_out[10] ));
 sky130_fd_sc_hd__dfrtp_4 _1059_ (.CLK(clknet_4_2_0_clk),
    .D(_0037_),
    .RESET_B(net36),
    .Q(\CTR.time_out[11] ));
 sky130_fd_sc_hd__dfrtp_4 _1060_ (.CLK(clknet_4_11_0_clk),
    .D(_0038_),
    .RESET_B(net41),
    .Q(\TIM.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1061_ (.CLK(clknet_4_11_0_clk),
    .D(_0039_),
    .RESET_B(net40),
    .Q(\TIM.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1062_ (.CLK(clknet_4_11_0_clk),
    .D(_0040_),
    .RESET_B(net40),
    .Q(\TIM.cnt[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1063_ (.CLK(clknet_4_11_0_clk),
    .D(_0041_),
    .RESET_B(net41),
    .Q(\TIM.cnt[4] ));
 sky130_fd_sc_hd__dfrtp_2 _1064_ (.CLK(clknet_4_11_0_clk),
    .D(_0042_),
    .RESET_B(net41),
    .Q(\TIM.cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1065_ (.CLK(clknet_4_11_0_clk),
    .D(_0043_),
    .RESET_B(net40),
    .Q(net32));
 sky130_fd_sc_hd__dfstp_1 _1066_ (.CLK(clknet_4_2_0_clk),
    .D(_0044_),
    .SET_B(net36),
    .Q(\MEM.raddr[0] ));
 sky130_fd_sc_hd__dfstp_1 _1067_ (.CLK(clknet_4_2_0_clk),
    .D(_0045_),
    .SET_B(net36),
    .Q(\MEM.raddr[1] ));
 sky130_fd_sc_hd__dfstp_1 _1068_ (.CLK(clknet_4_2_0_clk),
    .D(_0046_),
    .SET_B(net35),
    .Q(\MEM.raddr[2] ));
 sky130_fd_sc_hd__dfrtp_2 _1069_ (.CLK(clknet_4_9_0_clk),
    .D(_0047_),
    .RESET_B(net39),
    .Q(\TIM.cnt[0] ));
 sky130_fd_sc_hd__dfstp_2 _1070_ (.CLK(clknet_4_2_0_clk),
    .D(_0048_),
    .SET_B(net36),
    .Q(\MEM.addr[0] ));
 sky130_fd_sc_hd__dfstp_2 _1071_ (.CLK(clknet_4_2_0_clk),
    .D(_0049_),
    .SET_B(net36),
    .Q(\MEM.addr[1] ));
 sky130_fd_sc_hd__dfstp_1 _1072_ (.CLK(clknet_4_2_0_clk),
    .D(_0050_),
    .SET_B(net36),
    .Q(\MEM.addr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1073_ (.CLK(clknet_4_14_0_clk),
    .D(_0051_),
    .RESET_B(net39),
    .Q(\CTR.time_out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1074_ (.CLK(clknet_4_15_0_clk),
    .D(_0052_),
    .RESET_B(net39),
    .Q(\CTR.time_out[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1075_ (.CLK(clknet_4_14_0_clk),
    .D(_0053_),
    .RESET_B(net39),
    .Q(\CTR.time_out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1076_ (.CLK(clknet_4_13_0_clk),
    .D(_0054_),
    .RESET_B(net39),
    .Q(\CTR.time_out[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1077_ (.CLK(clknet_4_13_0_clk),
    .D(_0055_),
    .RESET_B(net38),
    .Q(\CTR.time_out[4] ));
 sky130_fd_sc_hd__dfrtp_4 _1078_ (.CLK(clknet_4_7_0_clk),
    .D(_0056_),
    .RESET_B(net41),
    .Q(\CTR.time_out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1079_ (.CLK(clknet_4_6_0_clk),
    .D(\MEM.next_mem5[0] ),
    .RESET_B(net38),
    .Q(\MEM.mem5[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1080_ (.CLK(clknet_4_7_0_clk),
    .D(\MEM.next_mem5[1] ),
    .RESET_B(net41),
    .Q(\MEM.mem5[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1081_ (.CLK(clknet_4_6_0_clk),
    .D(\MEM.next_mem5[2] ),
    .RESET_B(net38),
    .Q(\MEM.mem5[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1082_ (.CLK(clknet_4_4_0_clk),
    .D(\MEM.next_mem5[3] ),
    .RESET_B(net37),
    .Q(\MEM.mem5[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1083_ (.CLK(clknet_4_4_0_clk),
    .D(\MEM.next_mem5[4] ),
    .RESET_B(net37),
    .Q(\MEM.mem5[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1084_ (.CLK(clknet_4_4_0_clk),
    .D(\MEM.next_mem5[5] ),
    .RESET_B(net37),
    .Q(\MEM.mem5[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1085_ (.CLK(clknet_4_1_0_clk),
    .D(\MEM.next_mem5[6] ),
    .RESET_B(net35),
    .Q(\MEM.mem5[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1086_ (.CLK(clknet_4_0_0_clk),
    .D(\MEM.next_mem5[7] ),
    .RESET_B(net35),
    .Q(\MEM.mem5[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1087_ (.CLK(clknet_4_0_0_clk),
    .D(\MEM.next_mem5[8] ),
    .RESET_B(net35),
    .Q(\MEM.mem5[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1088_ (.CLK(clknet_4_3_0_clk),
    .D(\MEM.next_mem5[9] ),
    .RESET_B(net36),
    .Q(\MEM.mem5[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1089_ (.CLK(clknet_4_0_0_clk),
    .D(\MEM.next_mem5[10] ),
    .RESET_B(net35),
    .Q(\MEM.mem5[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1090_ (.CLK(clknet_4_3_0_clk),
    .D(\MEM.next_mem5[11] ),
    .RESET_B(net36),
    .Q(\MEM.mem5[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1091_ (.CLK(clknet_4_9_0_clk),
    .D(\MEM.next_mem4[0] ),
    .RESET_B(net38),
    .Q(\MEM.mem4[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1092_ (.CLK(clknet_4_12_0_clk),
    .D(\MEM.next_mem4[1] ),
    .RESET_B(net38),
    .Q(\MEM.mem4[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1093_ (.CLK(clknet_4_6_0_clk),
    .D(\MEM.next_mem4[2] ),
    .RESET_B(net38),
    .Q(\MEM.mem4[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1094_ (.CLK(clknet_4_1_0_clk),
    .D(\MEM.next_mem4[3] ),
    .RESET_B(net35),
    .Q(\MEM.mem4[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1095_ (.CLK(clknet_4_4_0_clk),
    .D(\MEM.next_mem4[4] ),
    .RESET_B(net37),
    .Q(\MEM.mem4[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1096_ (.CLK(clknet_4_6_0_clk),
    .D(\MEM.next_mem4[5] ),
    .RESET_B(net38),
    .Q(\MEM.mem4[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1097_ (.CLK(clknet_4_1_0_clk),
    .D(\MEM.next_mem4[6] ),
    .RESET_B(net35),
    .Q(\MEM.mem4[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1098_ (.CLK(clknet_4_0_0_clk),
    .D(\MEM.next_mem4[7] ),
    .RESET_B(net35),
    .Q(\MEM.mem4[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1099_ (.CLK(clknet_4_0_0_clk),
    .D(\MEM.next_mem4[8] ),
    .RESET_B(net35),
    .Q(\MEM.mem4[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1100_ (.CLK(clknet_4_3_0_clk),
    .D(\MEM.next_mem4[9] ),
    .RESET_B(net36),
    .Q(\MEM.mem4[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1101_ (.CLK(clknet_4_0_0_clk),
    .D(\MEM.next_mem4[10] ),
    .RESET_B(net35),
    .Q(\MEM.mem4[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1102_ (.CLK(clknet_4_3_0_clk),
    .D(\MEM.next_mem4[11] ),
    .RESET_B(net36),
    .Q(\MEM.mem4[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1103_ (.CLK(clknet_4_6_0_clk),
    .D(\MEM.next_mem3[0] ),
    .RESET_B(net38),
    .Q(\MEM.mem3[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1104_ (.CLK(clknet_4_6_0_clk),
    .D(\MEM.next_mem3[1] ),
    .RESET_B(net38),
    .Q(\MEM.mem3[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1105_ (.CLK(clknet_4_6_0_clk),
    .D(\MEM.next_mem3[2] ),
    .RESET_B(net38),
    .Q(\MEM.mem3[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1106_ (.CLK(clknet_4_4_0_clk),
    .D(\MEM.next_mem3[3] ),
    .RESET_B(net37),
    .Q(\MEM.mem3[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1107_ (.CLK(clknet_4_4_0_clk),
    .D(\MEM.next_mem3[4] ),
    .RESET_B(net37),
    .Q(\MEM.mem3[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1108_ (.CLK(clknet_4_4_0_clk),
    .D(\MEM.next_mem3[5] ),
    .RESET_B(net37),
    .Q(\MEM.mem3[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1109_ (.CLK(clknet_4_1_0_clk),
    .D(\MEM.next_mem3[6] ),
    .RESET_B(net35),
    .Q(\MEM.mem3[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1110_ (.CLK(clknet_4_0_0_clk),
    .D(\MEM.next_mem3[7] ),
    .RESET_B(net35),
    .Q(\MEM.mem3[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1111_ (.CLK(clknet_4_0_0_clk),
    .D(\MEM.next_mem3[8] ),
    .RESET_B(net35),
    .Q(\MEM.mem3[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1112_ (.CLK(clknet_4_3_0_clk),
    .D(\MEM.next_mem3[9] ),
    .RESET_B(net36),
    .Q(\MEM.mem3[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1113_ (.CLK(clknet_4_0_0_clk),
    .D(\MEM.next_mem3[10] ),
    .RESET_B(net35),
    .Q(\MEM.mem3[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1114_ (.CLK(clknet_4_3_0_clk),
    .D(\MEM.next_mem3[11] ),
    .RESET_B(net36),
    .Q(\MEM.mem3[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1115_ (.CLK(clknet_4_6_0_clk),
    .D(\MEM.next_mem2[0] ),
    .RESET_B(net38),
    .Q(\MEM.mem2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1116_ (.CLK(clknet_4_7_0_clk),
    .D(\MEM.next_mem2[1] ),
    .RESET_B(net41),
    .Q(\MEM.mem2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1117_ (.CLK(clknet_4_7_0_clk),
    .D(net101),
    .RESET_B(net38),
    .Q(\MEM.mem2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1118_ (.CLK(clknet_4_4_0_clk),
    .D(\MEM.next_mem2[3] ),
    .RESET_B(net37),
    .Q(\MEM.mem2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1119_ (.CLK(clknet_4_4_0_clk),
    .D(net97),
    .RESET_B(net37),
    .Q(\MEM.mem2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1120_ (.CLK(clknet_4_6_0_clk),
    .D(\MEM.next_mem2[5] ),
    .RESET_B(net37),
    .Q(\MEM.mem2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1121_ (.CLK(clknet_4_1_0_clk),
    .D(\MEM.next_mem2[6] ),
    .RESET_B(net36),
    .Q(\MEM.mem2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1122_ (.CLK(clknet_4_1_0_clk),
    .D(\MEM.next_mem2[7] ),
    .RESET_B(net36),
    .Q(\MEM.mem2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1123_ (.CLK(clknet_4_0_0_clk),
    .D(\MEM.next_mem2[8] ),
    .RESET_B(net35),
    .Q(\MEM.mem2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1124_ (.CLK(clknet_4_3_0_clk),
    .D(\MEM.next_mem2[9] ),
    .RESET_B(net36),
    .Q(\MEM.mem2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1125_ (.CLK(clknet_4_0_0_clk),
    .D(\MEM.next_mem2[10] ),
    .RESET_B(net35),
    .Q(\MEM.mem2[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1126_ (.CLK(clknet_4_3_0_clk),
    .D(\MEM.next_mem2[11] ),
    .RESET_B(net36),
    .Q(\MEM.mem2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1127_ (.CLK(clknet_4_12_0_clk),
    .D(\MEM.next_mem1[0] ),
    .RESET_B(net39),
    .Q(\MEM.mem1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1128_ (.CLK(clknet_4_12_0_clk),
    .D(\MEM.next_mem1[1] ),
    .RESET_B(net39),
    .Q(\MEM.mem1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1129_ (.CLK(clknet_4_12_0_clk),
    .D(\MEM.next_mem1[2] ),
    .RESET_B(net39),
    .Q(\MEM.mem1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1130_ (.CLK(clknet_4_9_0_clk),
    .D(\MEM.next_mem1[3] ),
    .RESET_B(net39),
    .Q(\MEM.mem1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1131_ (.CLK(clknet_4_12_0_clk),
    .D(\MEM.next_mem1[4] ),
    .RESET_B(net39),
    .Q(\MEM.mem1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1132_ (.CLK(clknet_4_12_0_clk),
    .D(\MEM.next_mem1[5] ),
    .RESET_B(net39),
    .Q(\MEM.mem1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1133_ (.CLK(clknet_4_8_0_clk),
    .D(\MEM.next_mem1[6] ),
    .RESET_B(net40),
    .Q(\MEM.mem1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1134_ (.CLK(clknet_4_8_0_clk),
    .D(\MEM.next_mem1[7] ),
    .RESET_B(net40),
    .Q(\MEM.mem1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1135_ (.CLK(clknet_4_8_0_clk),
    .D(\MEM.next_mem1[8] ),
    .RESET_B(net40),
    .Q(\MEM.mem1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1136_ (.CLK(clknet_4_8_0_clk),
    .D(\MEM.next_mem1[9] ),
    .RESET_B(net40),
    .Q(\MEM.mem1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1137_ (.CLK(clknet_4_10_0_clk),
    .D(\MEM.next_mem1[10] ),
    .RESET_B(net40),
    .Q(\MEM.mem1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1138_ (.CLK(clknet_4_8_0_clk),
    .D(\MEM.next_mem1[11] ),
    .RESET_B(net40),
    .Q(\MEM.mem1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1139_ (.CLK(clknet_4_9_0_clk),
    .D(\FSM.next_state[0] ),
    .RESET_B(net40),
    .Q(\FSM.state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1140_ (.CLK(clknet_4_8_0_clk),
    .D(\FSM.next_state[1] ),
    .RESET_B(net40),
    .Q(\FSM.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1141_ (.CLK(clknet_4_10_0_clk),
    .D(\FSM.next_state[2] ),
    .RESET_B(net40),
    .Q(\FSM.state[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1142_ (.CLK(clknet_4_10_0_clk),
    .D(\FSM.next_state[3] ),
    .RESET_B(net40),
    .Q(\FSM.state[3] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__buf_6 fanout35 (.A(net36),
    .X(net35));
 sky130_fd_sc_hd__buf_6 fanout36 (.A(net41),
    .X(net36));
 sky130_fd_sc_hd__buf_6 fanout37 (.A(net41),
    .X(net37));
 sky130_fd_sc_hd__buf_6 fanout38 (.A(net41),
    .X(net38));
 sky130_fd_sc_hd__buf_6 fanout39 (.A(net41),
    .X(net39));
 sky130_fd_sc_hd__buf_8 fanout40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__buf_6 fanout41 (.A(net1),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\e1.intermediate ),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\MEM.mem1[9] ),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\MEM.mem1[7] ),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\MEM.mem4[11] ),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\MEM.mem3[7] ),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\MEM.mem1[6] ),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\MEM.mem3[8] ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\MEM.mem1[0] ),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\MEM.mem2[7] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\MEM.mem3[5] ),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\MEM.mem5[0] ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\e2.intermediate ),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\MEM.mem5[9] ),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\MEM.mem3[6] ),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\MEM.mem4[2] ),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\MEM.mem1[10] ),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\MEM.mem3[4] ),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\MEM.mem3[11] ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\MEM.mem4[8] ),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\MEM.mem3[9] ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\MEM.mem4[9] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\MEM.mem4[5] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\e2.sync ),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\MEM.mem5[11] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\MEM.mem4[0] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\MEM.mem2[8] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\MEM.mem4[6] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\MEM.mem5[5] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\MEM.mem3[2] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\MEM.mem3[3] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\MEM.mem1[11] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\MEM.mem4[7] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\MEM.mem3[0] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\e1.sync ),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\MEM.mem4[10] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\MEM.mem5[7] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\MEM.mem2[10] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\MEM.mem3[10] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\MEM.mem4[1] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\MEM.mem5[2] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\MEM.mem1[1] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\MEM.mem5[10] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\MEM.mem5[4] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\MEM.mem2[3] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\MEM.mem1[5] ),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\MEM.mem2[6] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\MEM.mem3[1] ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\MEM.mem2[1] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\MEM.mem2[5] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\MEM.mem5[3] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\MEM.mem2[4] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\MEM.next_mem2[4] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\MEM.mem2[11] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\MEM.mem2[0] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\MEM.mem2[2] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\MEM.mem1[3] ),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\MEM.next_mem2[2] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\CLKDIV.count[19] ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\MEM.mem5[1] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\MEM.mem4[3] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\CLKDIV.count[14] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_0162_),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\MEM.mem4[4] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\MEM.mem2[9] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\CLKDIV.count[15] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\MEM.mem5[8] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\MEM.mem1[4] ),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\CLKDIV.count[13] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\MEM.mem5[6] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\CLKDIV.count[9] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\CLKDIV.count[0] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\CLKDIV.count[17] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\CLKDIV.count[11] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net32),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\CTR.minutes ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\CLKDIV.count[8] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_0152_),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\MEM.mem1[8] ),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\CLKDIV.count[3] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\CLKDIV.count[5] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\CLKDIV.count[22] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\CLKDIV.count[21] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\CLKDIV.count[2] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(_0138_),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\TIM.cnt[9] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\TIM.cnt[10] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\TIM.cnt[5] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\CTR.time_out[11] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\MEM.mem1[2] ),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\CLKDIV.count[20] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\TIM.cnt[2] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\TIM.cnt[11] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\TIM.cnt[7] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\MEM.addr[0] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\TIM.cnt[8] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\TIM.cnt[1] ),
    .X(net137));
 sky130_fd_sc_hd__buf_1 input1 (.A(nrst),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(pb_0),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(pb_1),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 max_cap33 (.A(_0079_),
    .X(net33));
 sky130_fd_sc_hd__buf_4 max_cap34 (.A(_0086_),
    .X(net34));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(out_0[6]));
 sky130_fd_sc_hd__clkbuf_4 output11 (.A(net11),
    .X(out_1[0]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(out_1[1]));
 sky130_fd_sc_hd__clkbuf_4 output13 (.A(net13),
    .X(out_1[2]));
 sky130_fd_sc_hd__clkbuf_4 output14 (.A(net14),
    .X(out_1[3]));
 sky130_fd_sc_hd__clkbuf_4 output15 (.A(net15),
    .X(out_1[4]));
 sky130_fd_sc_hd__clkbuf_4 output16 (.A(net16),
    .X(out_1[5]));
 sky130_fd_sc_hd__clkbuf_4 output17 (.A(net17),
    .X(out_1[6]));
 sky130_fd_sc_hd__clkbuf_4 output18 (.A(net18),
    .X(out_2[0]));
 sky130_fd_sc_hd__clkbuf_4 output19 (.A(net19),
    .X(out_2[1]));
 sky130_fd_sc_hd__clkbuf_4 output20 (.A(net20),
    .X(out_2[2]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(out_2[3]));
 sky130_fd_sc_hd__clkbuf_4 output22 (.A(net22),
    .X(out_2[4]));
 sky130_fd_sc_hd__clkbuf_4 output23 (.A(net23),
    .X(out_2[5]));
 sky130_fd_sc_hd__clkbuf_4 output24 (.A(net24),
    .X(out_2[6]));
 sky130_fd_sc_hd__clkbuf_4 output25 (.A(net25),
    .X(out_3[0]));
 sky130_fd_sc_hd__clkbuf_4 output26 (.A(net26),
    .X(out_3[1]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(out_3[2]));
 sky130_fd_sc_hd__clkbuf_4 output28 (.A(net28),
    .X(out_3[3]));
 sky130_fd_sc_hd__clkbuf_4 output29 (.A(net29),
    .X(out_3[4]));
 sky130_fd_sc_hd__clkbuf_4 output30 (.A(net30),
    .X(out_3[5]));
 sky130_fd_sc_hd__clkbuf_4 output31 (.A(net31),
    .X(out_3[6]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(time_done));
 sky130_fd_sc_hd__clkbuf_4 output4 (.A(net4),
    .X(out_0[0]));
 sky130_fd_sc_hd__clkbuf_4 output5 (.A(net5),
    .X(out_0[1]));
 sky130_fd_sc_hd__clkbuf_4 output6 (.A(net6),
    .X(out_0[2]));
 sky130_fd_sc_hd__clkbuf_4 output7 (.A(net7),
    .X(out_0[3]));
 sky130_fd_sc_hd__clkbuf_4 output8 (.A(net8),
    .X(out_0[4]));
 sky130_fd_sc_hd__clkbuf_4 output9 (.A(net9),
    .X(out_0[5]));
endmodule

