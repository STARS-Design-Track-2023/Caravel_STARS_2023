magic
tech sky130A
magscale 1 2
timestamp 1693189295
<< viali >>
rect 1593 42313 1627 42347
rect 35081 42313 35115 42347
rect 9229 42245 9263 42279
rect 1501 42177 1535 42211
rect 17509 42177 17543 42211
rect 19717 42177 19751 42211
rect 31033 42177 31067 42211
rect 34989 42177 35023 42211
rect 35633 42177 35667 42211
rect 38761 42177 38795 42211
rect 31309 42109 31343 42143
rect 38945 42109 38979 42143
rect 9321 41973 9355 42007
rect 17325 41973 17359 42007
rect 19533 41973 19567 42007
rect 17128 41769 17162 41803
rect 10149 41633 10183 41667
rect 14105 41633 14139 41667
rect 16865 41633 16899 41667
rect 19349 41633 19383 41667
rect 19625 41633 19659 41667
rect 21373 41633 21407 41667
rect 9873 41565 9907 41599
rect 11805 41565 11839 41599
rect 16129 41565 16163 41599
rect 18889 41565 18923 41599
rect 22201 41565 22235 41599
rect 12081 41497 12115 41531
rect 13829 41497 13863 41531
rect 14381 41497 14415 41531
rect 22477 41497 22511 41531
rect 24225 41497 24259 41531
rect 11621 41429 11655 41463
rect 12357 41225 12391 41259
rect 14289 41225 14323 41259
rect 16865 41225 16899 41259
rect 19441 41225 19475 41259
rect 19809 41225 19843 41259
rect 21557 41225 21591 41259
rect 1685 41157 1719 41191
rect 12725 41157 12759 41191
rect 14933 41157 14967 41191
rect 12265 41089 12299 41123
rect 12449 41089 12483 41123
rect 12633 41089 12667 41123
rect 12817 41089 12851 41123
rect 14105 41089 14139 41123
rect 14289 41089 14323 41123
rect 14841 41089 14875 41123
rect 15025 41089 15059 41123
rect 17233 41089 17267 41123
rect 21373 41089 21407 41123
rect 21649 41089 21683 41123
rect 40785 41089 40819 41123
rect 1409 41021 1443 41055
rect 3433 41021 3467 41055
rect 3801 41021 3835 41055
rect 4077 41021 4111 41055
rect 5825 41021 5859 41055
rect 10517 41021 10551 41055
rect 17325 41021 17359 41055
rect 17509 41021 17543 41055
rect 19901 41021 19935 41055
rect 20085 41021 20119 41055
rect 21833 41021 21867 41055
rect 22109 41021 22143 41055
rect 23857 41021 23891 41055
rect 21189 40953 21223 40987
rect 11069 40885 11103 40919
rect 40969 40885 41003 40919
rect 2053 40681 2087 40715
rect 4261 40681 4295 40715
rect 11069 40681 11103 40715
rect 17049 40681 17083 40715
rect 22477 40681 22511 40715
rect 2513 40613 2547 40647
rect 15669 40613 15703 40647
rect 16037 40613 16071 40647
rect 17969 40613 18003 40647
rect 3157 40545 3191 40579
rect 5273 40545 5307 40579
rect 14381 40545 14415 40579
rect 14933 40545 14967 40579
rect 16221 40545 16255 40579
rect 16405 40545 16439 40579
rect 17693 40545 17727 40579
rect 18797 40545 18831 40579
rect 18889 40545 18923 40579
rect 19441 40545 19475 40579
rect 2237 40477 2271 40511
rect 2881 40477 2915 40511
rect 4445 40477 4479 40511
rect 4997 40477 5031 40511
rect 10425 40477 10459 40511
rect 10573 40477 10607 40511
rect 10890 40477 10924 40511
rect 11253 40477 11287 40511
rect 11437 40477 11471 40511
rect 14289 40477 14323 40511
rect 14473 40477 14507 40511
rect 14565 40477 14599 40511
rect 14749 40477 14783 40511
rect 14841 40477 14875 40511
rect 15025 40477 15059 40511
rect 15301 40477 15335 40511
rect 15485 40477 15519 40511
rect 16497 40477 16531 40511
rect 17877 40477 17911 40511
rect 22385 40477 22419 40511
rect 22569 40477 22603 40511
rect 22661 40477 22695 40511
rect 22845 40477 22879 40511
rect 2973 40409 3007 40443
rect 8033 40409 8067 40443
rect 10701 40409 10735 40443
rect 10793 40409 10827 40443
rect 14657 40409 14691 40443
rect 15761 40409 15795 40443
rect 19717 40409 19751 40443
rect 21465 40409 21499 40443
rect 22753 40409 22787 40443
rect 4629 40341 4663 40375
rect 5089 40341 5123 40375
rect 8309 40341 8343 40375
rect 11345 40341 11379 40375
rect 16865 40341 16899 40375
rect 17417 40341 17451 40375
rect 17509 40341 17543 40375
rect 18337 40341 18371 40375
rect 18705 40341 18739 40375
rect 10354 40137 10388 40171
rect 10517 40137 10551 40171
rect 17049 40137 17083 40171
rect 19257 40137 19291 40171
rect 22937 40137 22971 40171
rect 24961 40137 24995 40171
rect 7481 40069 7515 40103
rect 8677 40069 8711 40103
rect 10175 40069 10209 40103
rect 15393 40069 15427 40103
rect 16221 40069 16255 40103
rect 19993 40069 20027 40103
rect 23489 40069 23523 40103
rect 8493 40001 8527 40035
rect 9873 40001 9907 40035
rect 10057 40001 10091 40035
rect 10609 40001 10643 40035
rect 10793 40001 10827 40035
rect 11161 40001 11195 40035
rect 11345 40001 11379 40035
rect 11713 40001 11747 40035
rect 15301 40001 15335 40035
rect 15485 40001 15519 40035
rect 15669 40001 15703 40035
rect 15761 40001 15795 40035
rect 16865 40001 16899 40035
rect 18889 40001 18923 40035
rect 22017 40001 22051 40035
rect 23121 40001 23155 40035
rect 8217 39933 8251 39967
rect 10977 39933 11011 39967
rect 11253 39933 11287 39967
rect 11529 39933 11563 39967
rect 11897 39933 11931 39967
rect 12909 39933 12943 39967
rect 13185 39933 13219 39967
rect 14933 39933 14967 39967
rect 16681 39933 16715 39967
rect 18797 39933 18831 39967
rect 20729 39933 20763 39967
rect 23213 39933 23247 39967
rect 15853 39865 15887 39899
rect 8861 39797 8895 39831
rect 9965 39797 9999 39831
rect 10333 39797 10367 39831
rect 15117 39797 15151 39831
rect 16221 39797 16255 39831
rect 16405 39797 16439 39831
rect 21833 39797 21867 39831
rect 8217 39593 8251 39627
rect 11069 39593 11103 39627
rect 13461 39593 13495 39627
rect 15117 39593 15151 39627
rect 15761 39593 15795 39627
rect 23029 39593 23063 39627
rect 11805 39525 11839 39559
rect 3801 39457 3835 39491
rect 7389 39457 7423 39491
rect 8953 39457 8987 39491
rect 9229 39457 9263 39491
rect 21465 39457 21499 39491
rect 23489 39457 23523 39491
rect 23581 39457 23615 39491
rect 25881 39457 25915 39491
rect 7573 39389 7607 39423
rect 7849 39389 7883 39423
rect 11253 39389 11287 39423
rect 11437 39389 11471 39423
rect 11621 39389 11655 39423
rect 11713 39389 11747 39423
rect 11805 39389 11839 39423
rect 12081 39389 12115 39423
rect 12817 39389 12851 39423
rect 12910 39389 12944 39423
rect 13282 39389 13316 39423
rect 14749 39389 14783 39423
rect 14933 39389 14967 39423
rect 16221 39389 16255 39423
rect 18061 39389 18095 39423
rect 21189 39389 21223 39423
rect 23397 39389 23431 39423
rect 8217 39321 8251 39355
rect 10977 39321 11011 39355
rect 11345 39321 11379 39355
rect 11989 39321 12023 39355
rect 13093 39321 13127 39355
rect 13185 39321 13219 39355
rect 15393 39321 15427 39355
rect 15577 39321 15611 39355
rect 15853 39321 15887 39355
rect 16037 39321 16071 39355
rect 26157 39321 26191 39355
rect 4445 39253 4479 39287
rect 7757 39253 7791 39287
rect 8401 39253 8435 39287
rect 17877 39253 17911 39287
rect 22937 39253 22971 39287
rect 27629 39253 27663 39287
rect 4077 39049 4111 39083
rect 9045 39049 9079 39083
rect 11253 39049 11287 39083
rect 17233 39049 17267 39083
rect 17601 39049 17635 39083
rect 21649 39049 21683 39083
rect 26157 39049 26191 39083
rect 4445 38981 4479 39015
rect 7205 38981 7239 39015
rect 8769 38981 8803 39015
rect 17693 38981 17727 39015
rect 18337 38981 18371 39015
rect 21189 38981 21223 39015
rect 25881 38981 25915 39015
rect 27629 38981 27663 39015
rect 7021 38913 7055 38947
rect 7297 38913 7331 38947
rect 7573 38913 7607 38947
rect 8401 38913 8435 38947
rect 8494 38913 8528 38947
rect 8677 38913 8711 38947
rect 8866 38913 8900 38947
rect 10885 38913 10919 38947
rect 11069 38913 11103 38947
rect 11713 38913 11747 38947
rect 12633 38913 12667 38947
rect 18061 38913 18095 38947
rect 22109 38913 22143 38947
rect 22753 38913 22787 38947
rect 22937 38913 22971 38947
rect 25605 38913 25639 38947
rect 25789 38913 25823 38947
rect 25973 38913 26007 38947
rect 27077 38913 27111 38947
rect 2329 38845 2363 38879
rect 2605 38845 2639 38879
rect 4169 38845 4203 38879
rect 6193 38845 6227 38879
rect 7665 38845 7699 38879
rect 7941 38845 7975 38879
rect 11805 38845 11839 38879
rect 12909 38845 12943 38879
rect 14657 38845 14691 38879
rect 14841 38845 14875 38879
rect 17785 38845 17819 38879
rect 20085 38845 20119 38879
rect 22661 38845 22695 38879
rect 12081 38777 12115 38811
rect 21557 38777 21591 38811
rect 6837 38709 6871 38743
rect 15393 38709 15427 38743
rect 23029 38709 23063 38743
rect 3433 38505 3467 38539
rect 4721 38505 4755 38539
rect 6561 38505 6595 38539
rect 7573 38505 7607 38539
rect 11345 38505 11379 38539
rect 12633 38505 12667 38539
rect 18061 38505 18095 38539
rect 22017 38505 22051 38539
rect 5273 38437 5307 38471
rect 7849 38437 7883 38471
rect 11253 38437 11287 38471
rect 4445 38369 4479 38403
rect 5917 38369 5951 38403
rect 7113 38369 7147 38403
rect 7205 38369 7239 38403
rect 10885 38369 10919 38403
rect 24685 38369 24719 38403
rect 3617 38301 3651 38335
rect 4169 38301 4203 38335
rect 4905 38301 4939 38335
rect 6285 38301 6319 38335
rect 6653 38301 6687 38335
rect 7297 38301 7331 38335
rect 7389 38301 7423 38335
rect 7849 38301 7883 38335
rect 8033 38301 8067 38335
rect 11069 38301 11103 38335
rect 11345 38301 11379 38335
rect 11529 38301 11563 38335
rect 11989 38301 12023 38335
rect 12082 38301 12116 38335
rect 12495 38301 12529 38335
rect 17049 38301 17083 38335
rect 17141 38301 17175 38335
rect 17509 38301 17543 38335
rect 17877 38301 17911 38335
rect 20269 38301 20303 38335
rect 27629 38301 27663 38335
rect 5641 38233 5675 38267
rect 12265 38233 12299 38267
rect 12357 38233 12391 38267
rect 17693 38233 17727 38267
rect 17785 38233 17819 38267
rect 20545 38233 20579 38267
rect 24961 38233 24995 38267
rect 27905 38233 27939 38267
rect 3801 38165 3835 38199
rect 4261 38165 4295 38199
rect 5733 38165 5767 38199
rect 6837 38165 6871 38199
rect 6929 38165 6963 38199
rect 17325 38165 17359 38199
rect 26433 38165 26467 38199
rect 29377 38165 29411 38199
rect 6469 37961 6503 37995
rect 9321 37961 9355 37995
rect 9505 37961 9539 37995
rect 10977 37961 11011 37995
rect 11621 37961 11655 37995
rect 16129 37961 16163 37995
rect 18061 37961 18095 37995
rect 18153 37961 18187 37995
rect 7849 37893 7883 37927
rect 18889 37893 18923 37927
rect 19809 37893 19843 37927
rect 25973 37893 26007 37927
rect 6377 37825 6411 37859
rect 6561 37825 6595 37859
rect 6929 37825 6963 37859
rect 7113 37825 7147 37859
rect 7481 37825 7515 37859
rect 8953 37825 8987 37859
rect 9413 37825 9447 37859
rect 9597 37825 9631 37859
rect 10793 37825 10827 37859
rect 11529 37825 11563 37859
rect 11713 37825 11747 37859
rect 14565 37825 14599 37859
rect 14749 37825 14783 37859
rect 15945 37825 15979 37859
rect 17785 37825 17819 37859
rect 18337 37825 18371 37859
rect 18613 37825 18647 37859
rect 19625 37825 19659 37859
rect 20821 37825 20855 37859
rect 21925 37825 21959 37859
rect 22017 37825 22051 37859
rect 22661 37825 22695 37859
rect 23121 37825 23155 37859
rect 23305 37825 23339 37859
rect 23397 37825 23431 37859
rect 23489 37825 23523 37859
rect 23765 37825 23799 37859
rect 7205 37757 7239 37791
rect 7297 37757 7331 37791
rect 9045 37757 9079 37791
rect 18061 37757 18095 37791
rect 19441 37757 19475 37791
rect 24041 37757 24075 37791
rect 25789 37757 25823 37791
rect 26985 37757 27019 37791
rect 27261 37757 27295 37791
rect 17877 37689 17911 37723
rect 18429 37689 18463 37723
rect 18521 37689 18555 37723
rect 19257 37689 19291 37723
rect 22109 37689 22143 37723
rect 23673 37689 23707 37723
rect 6745 37621 6779 37655
rect 7665 37621 7699 37655
rect 8125 37621 8159 37655
rect 14657 37621 14691 37655
rect 19349 37621 19383 37655
rect 20913 37621 20947 37655
rect 22477 37621 22511 37655
rect 26065 37621 26099 37655
rect 28733 37621 28767 37655
rect 6837 37417 6871 37451
rect 10701 37417 10735 37451
rect 11161 37417 11195 37451
rect 14657 37417 14691 37451
rect 18429 37417 18463 37451
rect 19625 37417 19659 37451
rect 26525 37417 26559 37451
rect 27905 37417 27939 37451
rect 31953 37417 31987 37451
rect 15301 37349 15335 37383
rect 24961 37349 24995 37383
rect 29561 37349 29595 37383
rect 7021 37281 7055 37315
rect 10333 37281 10367 37315
rect 13093 37281 13127 37315
rect 14841 37281 14875 37315
rect 17049 37281 17083 37315
rect 22293 37281 22327 37315
rect 25421 37281 25455 37315
rect 6745 37213 6779 37247
rect 10425 37213 10459 37247
rect 11161 37213 11195 37247
rect 11345 37213 11379 37247
rect 12909 37213 12943 37247
rect 13737 37213 13771 37247
rect 13921 37213 13955 37247
rect 14473 37213 14507 37247
rect 14749 37213 14783 37247
rect 14933 37213 14967 37247
rect 15025 37213 15059 37247
rect 15485 37213 15519 37247
rect 15945 37213 15979 37247
rect 16221 37213 16255 37247
rect 16405 37213 16439 37247
rect 16957 37213 16991 37247
rect 18613 37213 18647 37247
rect 18981 37213 19015 37247
rect 19073 37213 19107 37247
rect 22017 37213 22051 37247
rect 24409 37213 24443 37247
rect 24685 37213 24719 37247
rect 24777 37213 24811 37247
rect 25973 37213 26007 37247
rect 26341 37213 26375 37247
rect 27353 37213 27387 37247
rect 27721 37213 27755 37247
rect 29745 37213 29779 37247
rect 29837 37213 29871 37247
rect 30205 37213 30239 37247
rect 40785 37213 40819 37247
rect 14289 37145 14323 37179
rect 18705 37145 18739 37179
rect 18797 37145 18831 37179
rect 19257 37145 19291 37179
rect 19441 37145 19475 37179
rect 24593 37145 24627 37179
rect 25145 37145 25179 37179
rect 26157 37145 26191 37179
rect 26249 37145 26283 37179
rect 27537 37145 27571 37179
rect 27629 37145 27663 37179
rect 31861 37145 31895 37179
rect 7021 37077 7055 37111
rect 12449 37077 12483 37111
rect 12817 37077 12851 37111
rect 13921 37077 13955 37111
rect 23765 37077 23799 37111
rect 31631 37077 31665 37111
rect 40969 37077 41003 37111
rect 8033 36873 8067 36907
rect 10333 36873 10367 36907
rect 22201 36873 22235 36907
rect 27813 36873 27847 36907
rect 3801 36805 3835 36839
rect 14105 36805 14139 36839
rect 21649 36805 21683 36839
rect 1777 36737 1811 36771
rect 6653 36737 6687 36771
rect 6837 36737 6871 36771
rect 6929 36737 6963 36771
rect 7298 36737 7332 36771
rect 7665 36737 7699 36771
rect 7757 36737 7791 36771
rect 9965 36737 9999 36771
rect 11989 36737 12023 36771
rect 14565 36737 14599 36771
rect 15117 36737 15151 36771
rect 16037 36737 16071 36771
rect 16865 36737 16899 36771
rect 17049 36737 17083 36771
rect 17233 36737 17267 36771
rect 17417 36737 17451 36771
rect 18061 36737 18095 36771
rect 18153 36737 18187 36771
rect 18337 36737 18371 36771
rect 18429 36737 18463 36771
rect 18705 36737 18739 36771
rect 19165 36737 19199 36771
rect 19625 36737 19659 36771
rect 22569 36737 22603 36771
rect 27261 36737 27295 36771
rect 27445 36737 27479 36771
rect 27537 36737 27571 36771
rect 27629 36737 27663 36771
rect 30021 36737 30055 36771
rect 30205 36737 30239 36771
rect 2053 36669 2087 36703
rect 4353 36669 4387 36703
rect 4629 36669 4663 36703
rect 7021 36669 7055 36703
rect 7205 36669 7239 36703
rect 7389 36669 7423 36703
rect 7481 36669 7515 36703
rect 10057 36669 10091 36703
rect 12081 36669 12115 36703
rect 12357 36669 12391 36703
rect 14657 36669 14691 36703
rect 16129 36669 16163 36703
rect 17141 36669 17175 36703
rect 18613 36669 18647 36703
rect 19257 36669 19291 36703
rect 19901 36669 19935 36703
rect 22661 36669 22695 36703
rect 22845 36669 22879 36703
rect 27905 36669 27939 36703
rect 28181 36669 28215 36703
rect 29929 36669 29963 36703
rect 16405 36601 16439 36635
rect 30297 36601 30331 36635
rect 6101 36533 6135 36567
rect 6469 36533 6503 36567
rect 7665 36533 7699 36567
rect 11805 36533 11839 36567
rect 14841 36533 14875 36567
rect 15209 36533 15243 36567
rect 16681 36533 16715 36567
rect 17325 36533 17359 36567
rect 18429 36533 18463 36567
rect 18889 36533 18923 36567
rect 19533 36533 19567 36567
rect 2329 36329 2363 36363
rect 6929 36329 6963 36363
rect 8125 36329 8159 36363
rect 9873 36329 9907 36363
rect 10793 36329 10827 36363
rect 13185 36329 13219 36363
rect 15393 36329 15427 36363
rect 16589 36329 16623 36363
rect 18797 36329 18831 36363
rect 19349 36329 19383 36363
rect 28273 36329 28307 36363
rect 28457 36329 28491 36363
rect 28733 36329 28767 36363
rect 29745 36329 29779 36363
rect 15301 36261 15335 36295
rect 18521 36261 18555 36295
rect 27261 36261 27295 36295
rect 3433 36193 3467 36227
rect 3801 36193 3835 36227
rect 6653 36193 6687 36227
rect 9689 36193 9723 36227
rect 10885 36193 10919 36227
rect 12725 36193 12759 36227
rect 13645 36193 13679 36227
rect 13737 36193 13771 36227
rect 15485 36193 15519 36227
rect 16221 36193 16255 36227
rect 18153 36193 18187 36227
rect 27813 36193 27847 36227
rect 33609 36193 33643 36227
rect 2513 36125 2547 36159
rect 6561 36125 6595 36159
rect 7573 36125 7607 36159
rect 7941 36125 7975 36159
rect 9597 36125 9631 36159
rect 9781 36125 9815 36159
rect 10149 36125 10183 36159
rect 10241 36125 10275 36159
rect 10333 36125 10367 36159
rect 10517 36125 10551 36159
rect 10609 36125 10643 36159
rect 10701 36125 10735 36159
rect 12633 36125 12667 36159
rect 15209 36125 15243 36159
rect 16405 36125 16439 36159
rect 18337 36125 18371 36159
rect 18797 36125 18831 36159
rect 18981 36125 19015 36159
rect 19257 36125 19291 36159
rect 19441 36125 19475 36159
rect 27721 36125 27755 36159
rect 28089 36125 28123 36159
rect 28273 36125 28307 36159
rect 29561 36125 29595 36159
rect 29653 36125 29687 36159
rect 29837 36125 29871 36159
rect 29929 36125 29963 36159
rect 30389 36125 30423 36159
rect 31861 36125 31895 36159
rect 31953 36125 31987 36159
rect 33793 36125 33827 36159
rect 3157 36057 3191 36091
rect 4077 36057 4111 36091
rect 7757 36057 7791 36091
rect 7849 36057 7883 36091
rect 13553 36057 13587 36091
rect 25697 36057 25731 36091
rect 28641 36057 28675 36091
rect 2789 35989 2823 36023
rect 3249 35989 3283 36023
rect 5549 35989 5583 36023
rect 13001 35989 13035 36023
rect 25789 35989 25823 36023
rect 27629 35989 27663 36023
rect 30113 35989 30147 36023
rect 30481 35989 30515 36023
rect 32137 35989 32171 36023
rect 33977 35989 34011 36023
rect 4261 35785 4295 35819
rect 7021 35785 7055 35819
rect 15669 35785 15703 35819
rect 17233 35785 17267 35819
rect 19993 35785 20027 35819
rect 25605 35785 25639 35819
rect 26065 35785 26099 35819
rect 31953 35785 31987 35819
rect 23581 35717 23615 35751
rect 25237 35717 25271 35751
rect 31309 35717 31343 35751
rect 32229 35717 32263 35751
rect 33149 35717 33183 35751
rect 4445 35649 4479 35683
rect 5089 35649 5123 35683
rect 5181 35649 5215 35683
rect 6837 35649 6871 35683
rect 7113 35649 7147 35683
rect 10149 35649 10183 35683
rect 10701 35649 10735 35683
rect 15569 35649 15603 35683
rect 17174 35649 17208 35683
rect 19809 35649 19843 35683
rect 22017 35649 22051 35683
rect 22293 35649 22327 35683
rect 22477 35649 22511 35683
rect 23213 35649 23247 35683
rect 23305 35649 23339 35683
rect 24041 35649 24075 35683
rect 24133 35649 24167 35683
rect 24317 35649 24351 35683
rect 24409 35649 24443 35683
rect 24685 35649 24719 35683
rect 25145 35649 25179 35683
rect 25421 35649 25455 35683
rect 25697 35649 25731 35683
rect 29929 35649 29963 35683
rect 30021 35649 30055 35683
rect 30134 35649 30168 35683
rect 30297 35649 30331 35683
rect 30941 35649 30975 35683
rect 31116 35649 31150 35683
rect 31217 35649 31251 35683
rect 31401 35649 31435 35683
rect 32781 35649 32815 35683
rect 33517 35649 33551 35683
rect 34161 35649 34195 35683
rect 34713 35649 34747 35683
rect 5365 35581 5399 35615
rect 10057 35581 10091 35615
rect 10241 35581 10275 35615
rect 10333 35581 10367 35615
rect 10517 35581 10551 35615
rect 14473 35581 14507 35615
rect 17693 35581 17727 35615
rect 22569 35581 22603 35615
rect 24501 35581 24535 35615
rect 24777 35581 24811 35615
rect 24869 35581 24903 35615
rect 24961 35581 24995 35615
rect 25789 35581 25823 35615
rect 31493 35581 31527 35615
rect 34621 35581 34655 35615
rect 34897 35581 34931 35615
rect 4721 35513 4755 35547
rect 17049 35513 17083 35547
rect 29653 35513 29687 35547
rect 31861 35513 31895 35547
rect 33793 35513 33827 35547
rect 6653 35445 6687 35479
rect 9873 35445 9907 35479
rect 10885 35445 10919 35479
rect 15117 35445 15151 35479
rect 17601 35445 17635 35479
rect 21833 35445 21867 35479
rect 23857 35445 23891 35479
rect 25697 35445 25731 35479
rect 31033 35445 31067 35479
rect 32321 35445 32355 35479
rect 33977 35445 34011 35479
rect 34345 35445 34379 35479
rect 7205 35241 7239 35275
rect 8677 35241 8711 35275
rect 9781 35241 9815 35275
rect 15945 35241 15979 35275
rect 16773 35241 16807 35275
rect 23213 35241 23247 35275
rect 23489 35241 23523 35275
rect 23857 35241 23891 35275
rect 25789 35241 25823 35275
rect 26433 35241 26467 35275
rect 26801 35241 26835 35275
rect 27077 35241 27111 35275
rect 27169 35241 27203 35275
rect 29193 35241 29227 35275
rect 32137 35241 32171 35275
rect 33517 35241 33551 35275
rect 36093 35241 36127 35275
rect 9965 35173 9999 35207
rect 27537 35173 27571 35207
rect 34253 35173 34287 35207
rect 7021 35105 7055 35139
rect 8401 35105 8435 35139
rect 14197 35105 14231 35139
rect 16405 35105 16439 35139
rect 20821 35105 20855 35139
rect 21097 35105 21131 35139
rect 23949 35105 23983 35139
rect 26065 35105 26099 35139
rect 26709 35105 26743 35139
rect 31033 35105 31067 35139
rect 32045 35105 32079 35139
rect 33885 35105 33919 35139
rect 6929 35037 6963 35071
rect 8309 35037 8343 35071
rect 10057 35037 10091 35071
rect 10149 35037 10183 35071
rect 10425 35037 10459 35071
rect 11069 35037 11103 35071
rect 11345 35037 11379 35071
rect 11713 35037 11747 35071
rect 11897 35037 11931 35071
rect 16497 35037 16531 35071
rect 19901 35037 19935 35071
rect 20085 35037 20119 35071
rect 23121 35037 23155 35071
rect 23213 35037 23247 35071
rect 23673 35037 23707 35071
rect 24409 35037 24443 35071
rect 24557 35037 24591 35071
rect 24685 35037 24719 35071
rect 24915 35037 24949 35071
rect 25145 35037 25179 35071
rect 25293 35037 25327 35071
rect 25421 35037 25455 35071
rect 25513 35037 25547 35071
rect 25651 35037 25685 35071
rect 26249 35037 26283 35071
rect 26525 35037 26559 35071
rect 26893 35037 26927 35071
rect 27353 35037 27387 35071
rect 27629 35037 27663 35071
rect 28917 35037 28951 35071
rect 29101 35037 29135 35071
rect 30849 35037 30883 35071
rect 30941 35037 30975 35071
rect 31217 35037 31251 35071
rect 31401 35037 31435 35071
rect 31953 35037 31987 35071
rect 33425 35037 33459 35071
rect 36001 35037 36035 35071
rect 9597 34969 9631 35003
rect 10885 34969 10919 35003
rect 14473 34969 14507 35003
rect 22937 34969 22971 35003
rect 24777 34969 24811 35003
rect 26617 34969 26651 35003
rect 31677 34969 31711 35003
rect 9797 34901 9831 34935
rect 10241 34901 10275 34935
rect 10333 34901 10367 34935
rect 11253 34901 11287 34935
rect 11897 34901 11931 34935
rect 20269 34901 20303 34935
rect 22569 34901 22603 34935
rect 23397 34901 23431 34935
rect 25053 34901 25087 34935
rect 31125 34901 31159 34935
rect 32321 34901 32355 34935
rect 34345 34901 34379 34935
rect 36461 34901 36495 34935
rect 2053 34697 2087 34731
rect 8769 34697 8803 34731
rect 9689 34697 9723 34731
rect 10977 34697 11011 34731
rect 11897 34697 11931 34731
rect 11989 34697 12023 34731
rect 13185 34697 13219 34731
rect 19717 34697 19751 34731
rect 20085 34697 20119 34731
rect 20637 34697 20671 34731
rect 22569 34697 22603 34731
rect 23397 34697 23431 34731
rect 26801 34697 26835 34731
rect 27629 34697 27663 34731
rect 29863 34697 29897 34731
rect 31125 34697 31159 34731
rect 35357 34697 35391 34731
rect 7021 34629 7055 34663
rect 9229 34629 9263 34663
rect 11529 34629 11563 34663
rect 11745 34629 11779 34663
rect 14473 34629 14507 34663
rect 14565 34629 14599 34663
rect 17325 34629 17359 34663
rect 20453 34629 20487 34663
rect 24961 34629 24995 34663
rect 29653 34629 29687 34663
rect 32321 34629 32355 34663
rect 32873 34629 32907 34663
rect 1869 34561 1903 34595
rect 6837 34561 6871 34595
rect 7297 34561 7331 34595
rect 7481 34561 7515 34595
rect 9137 34561 9171 34595
rect 9597 34561 9631 34595
rect 9781 34561 9815 34595
rect 10885 34561 10919 34595
rect 11069 34561 11103 34595
rect 12173 34561 12207 34595
rect 12357 34561 12391 34595
rect 12449 34561 12483 34595
rect 12725 34561 12759 34595
rect 13093 34561 13127 34595
rect 13277 34561 13311 34595
rect 14197 34561 14231 34595
rect 14290 34561 14324 34595
rect 14662 34561 14696 34595
rect 17141 34561 17175 34595
rect 17233 34561 17267 34595
rect 17443 34561 17477 34595
rect 17693 34561 17727 34595
rect 17877 34561 17911 34595
rect 19165 34561 19199 34595
rect 19901 34561 19935 34595
rect 20177 34561 20211 34595
rect 20269 34561 20303 34595
rect 22845 34561 22879 34595
rect 23121 34561 23155 34595
rect 23305 34561 23339 34595
rect 23581 34561 23615 34595
rect 23857 34561 23891 34595
rect 24777 34561 24811 34595
rect 26249 34561 26283 34595
rect 26433 34561 26467 34595
rect 26525 34561 26559 34595
rect 26617 34561 26651 34595
rect 26985 34561 27019 34595
rect 27133 34561 27167 34595
rect 27261 34561 27295 34595
rect 27350 34561 27384 34595
rect 27491 34561 27525 34595
rect 29101 34561 29135 34595
rect 29377 34561 29411 34595
rect 29561 34561 29595 34595
rect 31033 34561 31067 34595
rect 32689 34561 32723 34595
rect 32781 34561 32815 34595
rect 33149 34561 33183 34595
rect 35265 34561 35299 34595
rect 35449 34561 35483 34595
rect 36277 34561 36311 34595
rect 9321 34493 9355 34527
rect 12909 34493 12943 34527
rect 13001 34493 13035 34527
rect 17601 34493 17635 34527
rect 19625 34493 19659 34527
rect 23029 34493 23063 34527
rect 23765 34493 23799 34527
rect 25145 34493 25179 34527
rect 32229 34493 32263 34527
rect 33425 34493 33459 34527
rect 35633 34493 35667 34527
rect 36461 34493 36495 34527
rect 12541 34425 12575 34459
rect 14841 34425 14875 34459
rect 19533 34425 19567 34459
rect 23673 34425 23707 34459
rect 29193 34425 29227 34459
rect 29285 34425 29319 34459
rect 30021 34425 30055 34459
rect 35081 34425 35115 34459
rect 7205 34357 7239 34391
rect 7389 34357 7423 34391
rect 11735 34357 11769 34391
rect 16957 34357 16991 34391
rect 18061 34357 18095 34391
rect 22937 34357 22971 34391
rect 28917 34357 28951 34391
rect 29837 34357 29871 34391
rect 5181 34153 5215 34187
rect 8309 34153 8343 34187
rect 9781 34153 9815 34187
rect 11621 34153 11655 34187
rect 12909 34153 12943 34187
rect 13737 34153 13771 34187
rect 19901 34153 19935 34187
rect 20453 34153 20487 34187
rect 20821 34153 20855 34187
rect 24041 34153 24075 34187
rect 30849 34153 30883 34187
rect 36921 34153 36955 34187
rect 37473 34153 37507 34187
rect 4813 34085 4847 34119
rect 11989 34085 12023 34119
rect 24869 34085 24903 34119
rect 27721 34085 27755 34119
rect 31493 34085 31527 34119
rect 4077 34017 4111 34051
rect 5365 34017 5399 34051
rect 7297 34017 7331 34051
rect 7573 34017 7607 34051
rect 7665 34017 7699 34051
rect 12081 34017 12115 34051
rect 13461 34017 13495 34051
rect 14105 34017 14139 34051
rect 16957 34017 16991 34051
rect 19809 34017 19843 34051
rect 20361 34017 20395 34051
rect 21189 34017 21223 34051
rect 21465 34017 21499 34051
rect 21557 34017 21591 34051
rect 23949 34017 23983 34051
rect 24409 34017 24443 34051
rect 30297 34017 30331 34051
rect 31677 34017 31711 34051
rect 32045 34017 32079 34051
rect 33149 34017 33183 34051
rect 35357 34017 35391 34051
rect 36277 34017 36311 34051
rect 3985 33949 4019 33983
rect 4537 33949 4571 33983
rect 4721 33949 4755 33983
rect 4813 33949 4847 33983
rect 5089 33949 5123 33983
rect 5457 33949 5491 33983
rect 5733 33949 5767 33983
rect 5825 33949 5859 33983
rect 6285 33949 6319 33983
rect 6929 33949 6963 33983
rect 7021 33949 7055 33983
rect 7481 33949 7515 33983
rect 7757 33949 7791 33983
rect 8033 33949 8067 33983
rect 9689 33949 9723 33983
rect 9873 33951 9907 33985
rect 11437 33949 11471 33983
rect 11805 33949 11839 33983
rect 11897 33949 11931 33983
rect 13093 33949 13127 33983
rect 13277 33949 13311 33983
rect 13369 33949 13403 33983
rect 13737 33949 13771 33983
rect 13921 33949 13955 33983
rect 14289 33949 14323 33983
rect 14473 33949 14507 33983
rect 14565 33949 14599 33983
rect 16589 33949 16623 33983
rect 16865 33949 16899 33983
rect 19349 33949 19383 33983
rect 20085 33949 20119 33983
rect 20269 33949 20303 33983
rect 20453 33949 20487 33983
rect 20637 33949 20671 33983
rect 21373 33949 21407 33983
rect 21649 33949 21683 33983
rect 22293 33949 22327 33983
rect 22441 33949 22475 33983
rect 22569 33949 22603 33983
rect 22661 33949 22695 33983
rect 22799 33949 22833 33983
rect 24041 33949 24075 33983
rect 24593 33949 24627 33983
rect 24685 33949 24719 33983
rect 24961 33949 24995 33983
rect 26709 33949 26743 33983
rect 26801 33949 26835 33983
rect 26985 33949 27019 33983
rect 27077 33949 27111 33983
rect 27169 33949 27203 33983
rect 27353 33949 27387 33983
rect 27537 33949 27571 33983
rect 28549 33949 28583 33983
rect 28642 33949 28676 33983
rect 28825 33949 28859 33983
rect 29014 33949 29048 33983
rect 29561 33949 29595 33983
rect 29654 33949 29688 33983
rect 29929 33949 29963 33983
rect 30026 33949 30060 33983
rect 30481 33949 30515 33983
rect 30573 33949 30607 33983
rect 30665 33949 30699 33983
rect 32873 33949 32907 33983
rect 33425 33949 33459 33983
rect 34069 33949 34103 33983
rect 34345 33949 34379 33983
rect 34713 33949 34747 33983
rect 34897 33949 34931 33983
rect 36645 33949 36679 33983
rect 38117 33949 38151 33983
rect 5917 33881 5951 33915
rect 6101 33881 6135 33915
rect 6561 33881 6595 33915
rect 11253 33881 11287 33915
rect 16405 33881 16439 33915
rect 17233 33881 17267 33915
rect 18981 33881 19015 33915
rect 23765 33881 23799 33915
rect 27445 33881 27479 33915
rect 27905 33881 27939 33915
rect 28917 33881 28951 33915
rect 29837 33881 29871 33915
rect 31125 33881 31159 33915
rect 31953 33881 31987 33915
rect 32162 33881 32196 33915
rect 35909 33881 35943 33915
rect 36093 33881 36127 33915
rect 36553 33881 36587 33915
rect 36737 33881 36771 33915
rect 37381 33881 37415 33915
rect 37933 33881 37967 33915
rect 4353 33813 4387 33847
rect 4629 33813 4663 33847
rect 4997 33813 5031 33847
rect 7205 33813 7239 33847
rect 16773 33813 16807 33847
rect 19349 33813 19383 33847
rect 22937 33813 22971 33847
rect 24225 33813 24259 33847
rect 26525 33813 26559 33847
rect 27997 33813 28031 33847
rect 29193 33813 29227 33847
rect 30205 33813 30239 33847
rect 31585 33813 31619 33847
rect 32321 33813 32355 33847
rect 35081 33813 35115 33847
rect 35541 33813 35575 33847
rect 36001 33813 36035 33847
rect 6561 33609 6595 33643
rect 9873 33609 9907 33643
rect 11627 33609 11661 33643
rect 12633 33609 12667 33643
rect 13277 33609 13311 33643
rect 14663 33609 14697 33643
rect 14749 33609 14783 33643
rect 16497 33609 16531 33643
rect 17693 33609 17727 33643
rect 23949 33609 23983 33643
rect 33241 33609 33275 33643
rect 34345 33609 34379 33643
rect 35541 33609 35575 33643
rect 36737 33609 36771 33643
rect 4353 33541 4387 33575
rect 4537 33541 4571 33575
rect 6377 33541 6411 33575
rect 7849 33541 7883 33575
rect 11529 33541 11563 33575
rect 14131 33541 14165 33575
rect 14321 33541 14355 33575
rect 4261 33473 4295 33507
rect 4445 33473 4479 33507
rect 4813 33473 4847 33507
rect 5273 33473 5307 33507
rect 6653 33473 6687 33507
rect 8677 33473 8711 33507
rect 9505 33473 9539 33507
rect 9689 33473 9723 33507
rect 9965 33473 9999 33507
rect 10149 33473 10183 33507
rect 10241 33473 10275 33507
rect 11713 33473 11747 33507
rect 11805 33473 11839 33507
rect 12173 33473 12207 33507
rect 12909 33473 12943 33507
rect 13093 33473 13127 33507
rect 14565 33473 14599 33507
rect 14841 33473 14875 33507
rect 16129 33473 16163 33507
rect 16773 33473 16807 33507
rect 17325 33473 17359 33507
rect 17601 33473 17635 33507
rect 17785 33473 17819 33507
rect 19533 33473 19567 33507
rect 21925 33473 21959 33507
rect 22293 33473 22327 33507
rect 24133 33473 24167 33507
rect 25513 33473 25547 33507
rect 25789 33473 25823 33507
rect 27261 33473 27295 33507
rect 32321 33473 32355 33507
rect 32505 33473 32539 33507
rect 33057 33473 33091 33507
rect 33977 33473 34011 33507
rect 34186 33473 34220 33507
rect 35357 33473 35391 33507
rect 35725 33473 35759 33507
rect 35872 33473 35906 33507
rect 36553 33473 36587 33507
rect 37289 33473 37323 33507
rect 37933 33473 37967 33507
rect 38301 33473 38335 33507
rect 38669 33473 38703 33507
rect 4721 33405 4755 33439
rect 5089 33405 5123 33439
rect 16037 33405 16071 33439
rect 17233 33405 17267 33439
rect 19625 33405 19659 33439
rect 24409 33405 24443 33439
rect 32597 33405 32631 33439
rect 33425 33405 33459 33439
rect 33701 33405 33735 33439
rect 34069 33405 34103 33439
rect 36093 33405 36127 33439
rect 37565 33405 37599 33439
rect 39221 33405 39255 33439
rect 39497 33405 39531 33439
rect 5457 33337 5491 33371
rect 6377 33337 6411 33371
rect 14473 33337 14507 33371
rect 24317 33337 24351 33371
rect 25605 33337 25639 33371
rect 25697 33337 25731 33371
rect 36185 33337 36219 33371
rect 4537 33269 4571 33303
rect 4997 33269 5031 33303
rect 10241 33269 10275 33303
rect 10425 33269 10459 33303
rect 12357 33269 12391 33303
rect 14289 33269 14323 33303
rect 19349 33269 19383 33303
rect 19882 33269 19916 33303
rect 21373 33269 21407 33303
rect 25329 33269 25363 33303
rect 27445 33269 27479 33303
rect 32137 33269 32171 33303
rect 33425 33269 33459 33303
rect 36001 33269 36035 33303
rect 40969 33269 41003 33303
rect 7297 33065 7331 33099
rect 12081 33065 12115 33099
rect 15853 33065 15887 33099
rect 15945 33065 15979 33099
rect 17601 33065 17635 33099
rect 19533 33065 19567 33099
rect 22661 33065 22695 33099
rect 26065 33065 26099 33099
rect 30665 33065 30699 33099
rect 36461 33065 36495 33099
rect 37749 33065 37783 33099
rect 38301 33065 38335 33099
rect 38853 33065 38887 33099
rect 41061 33065 41095 33099
rect 12265 32997 12299 33031
rect 24501 32997 24535 33031
rect 34161 32997 34195 33031
rect 16037 32929 16071 32963
rect 16497 32929 16531 32963
rect 20177 32929 20211 32963
rect 24685 32929 24719 32963
rect 37105 32929 37139 32963
rect 39405 32929 39439 32963
rect 7205 32861 7239 32895
rect 11621 32861 11655 32895
rect 11713 32861 11747 32895
rect 12081 32861 12115 32895
rect 15761 32861 15795 32895
rect 16147 32861 16181 32895
rect 17509 32861 17543 32895
rect 19901 32861 19935 32895
rect 20821 32861 20855 32895
rect 21097 32861 21131 32895
rect 22845 32861 22879 32895
rect 24501 32861 24535 32895
rect 24777 32861 24811 32895
rect 25789 32861 25823 32895
rect 25973 32861 26007 32895
rect 26065 32861 26099 32895
rect 30573 32861 30607 32895
rect 33885 32861 33919 32895
rect 33977 32861 34011 32895
rect 34713 32861 34747 32895
rect 34897 32861 34931 32895
rect 36369 32861 36403 32895
rect 36737 32861 36771 32895
rect 36829 32861 36863 32895
rect 37590 32861 37624 32895
rect 37933 32861 37967 32895
rect 38025 32861 38059 32895
rect 38393 32861 38427 32895
rect 39221 32861 39255 32895
rect 39865 32861 39899 32895
rect 40509 32861 40543 32895
rect 16313 32793 16347 32827
rect 22569 32793 22603 32827
rect 22753 32793 22787 32827
rect 24869 32793 24903 32827
rect 37381 32793 37415 32827
rect 38761 32793 38795 32827
rect 7665 32725 7699 32759
rect 19993 32725 20027 32759
rect 26249 32725 26283 32759
rect 35081 32725 35115 32759
rect 37013 32725 37047 32759
rect 37473 32725 37507 32759
rect 38577 32725 38611 32759
rect 39957 32725 39991 32759
rect 6929 32521 6963 32555
rect 7941 32521 7975 32555
rect 10333 32521 10367 32555
rect 11989 32521 12023 32555
rect 13553 32521 13587 32555
rect 13829 32521 13863 32555
rect 14749 32521 14783 32555
rect 16037 32521 16071 32555
rect 18153 32521 18187 32555
rect 24685 32521 24719 32555
rect 26985 32521 27019 32555
rect 30757 32521 30791 32555
rect 32597 32521 32631 32555
rect 32873 32521 32907 32555
rect 36185 32521 36219 32555
rect 38301 32521 38335 32555
rect 40601 32521 40635 32555
rect 40969 32521 41003 32555
rect 5089 32453 5123 32487
rect 9321 32453 9355 32487
rect 18061 32453 18095 32487
rect 22661 32453 22695 32487
rect 24225 32453 24259 32487
rect 28365 32453 28399 32487
rect 28457 32453 28491 32487
rect 30113 32453 30147 32487
rect 4813 32385 4847 32419
rect 6009 32385 6043 32419
rect 6193 32385 6227 32419
rect 6561 32385 6595 32419
rect 7205 32385 7239 32419
rect 9045 32385 9079 32419
rect 9138 32385 9172 32419
rect 9413 32385 9447 32419
rect 9510 32385 9544 32419
rect 9965 32385 9999 32419
rect 11805 32385 11839 32419
rect 11989 32385 12023 32419
rect 13461 32385 13495 32419
rect 13645 32385 13679 32419
rect 14013 32385 14047 32419
rect 14565 32385 14599 32419
rect 15853 32385 15887 32419
rect 16037 32385 16071 32419
rect 22017 32385 22051 32419
rect 22385 32385 22419 32419
rect 24501 32385 24535 32419
rect 26525 32385 26559 32419
rect 26709 32385 26743 32419
rect 26801 32385 26835 32419
rect 27537 32385 27571 32419
rect 27721 32385 27755 32419
rect 28181 32385 28215 32419
rect 28549 32385 28583 32419
rect 29029 32385 29063 32419
rect 29193 32385 29227 32419
rect 29285 32385 29319 32419
rect 29377 32385 29411 32419
rect 29745 32385 29779 32419
rect 30389 32385 30423 32419
rect 31033 32385 31067 32419
rect 31493 32385 31527 32419
rect 32137 32385 32171 32419
rect 32413 32385 32447 32419
rect 32689 32385 32723 32419
rect 32965 32385 32999 32419
rect 36369 32385 36403 32419
rect 36645 32385 36679 32419
rect 37749 32385 37783 32419
rect 38117 32385 38151 32419
rect 38853 32385 38887 32419
rect 40785 32385 40819 32419
rect 5089 32317 5123 32351
rect 6469 32317 6503 32351
rect 8309 32317 8343 32351
rect 8401 32317 8435 32351
rect 9873 32317 9907 32351
rect 14289 32317 14323 32351
rect 14381 32317 14415 32351
rect 22293 32317 22327 32351
rect 24409 32317 24443 32351
rect 27261 32317 27295 32351
rect 30573 32317 30607 32351
rect 30665 32317 30699 32351
rect 31217 32317 31251 32351
rect 32229 32317 32263 32351
rect 37657 32317 37691 32351
rect 39129 32317 39163 32351
rect 26341 32249 26375 32283
rect 27445 32249 27479 32283
rect 29561 32249 29595 32283
rect 32689 32249 32723 32283
rect 4905 32181 4939 32215
rect 6009 32181 6043 32215
rect 7757 32181 7791 32215
rect 8585 32181 8619 32215
rect 9689 32181 9723 32215
rect 14197 32181 14231 32215
rect 21833 32181 21867 32215
rect 22201 32181 22235 32215
rect 24501 32181 24535 32215
rect 27353 32181 27387 32215
rect 28733 32181 28767 32215
rect 30205 32181 30239 32215
rect 31125 32181 31159 32215
rect 31309 32181 31343 32215
rect 32137 32181 32171 32215
rect 38025 32181 38059 32215
rect 5181 31977 5215 32011
rect 12633 31977 12667 32011
rect 15209 31977 15243 32011
rect 22569 31977 22603 32011
rect 23673 31977 23707 32011
rect 23857 31977 23891 32011
rect 24409 31977 24443 32011
rect 25329 31977 25363 32011
rect 26525 31977 26559 32011
rect 26709 31977 26743 32011
rect 27261 31977 27295 32011
rect 27905 31977 27939 32011
rect 34897 31977 34931 32011
rect 36645 31977 36679 32011
rect 37289 31977 37323 32011
rect 38669 31977 38703 32011
rect 5825 31909 5859 31943
rect 5917 31909 5951 31943
rect 16037 31909 16071 31943
rect 16865 31909 16899 31943
rect 27169 31909 27203 31943
rect 27629 31909 27663 31943
rect 29193 31909 29227 31943
rect 31861 31909 31895 31943
rect 35081 31909 35115 31943
rect 37841 31909 37875 31943
rect 4905 31841 4939 31875
rect 5365 31841 5399 31875
rect 6469 31841 6503 31875
rect 9229 31841 9263 31875
rect 12725 31841 12759 31875
rect 14841 31841 14875 31875
rect 14932 31841 14966 31875
rect 16405 31841 16439 31875
rect 18705 31841 18739 31875
rect 23305 31841 23339 31875
rect 23765 31841 23799 31875
rect 24501 31841 24535 31875
rect 26801 31841 26835 31875
rect 29929 31841 29963 31875
rect 31585 31841 31619 31875
rect 2973 31773 3007 31807
rect 4813 31773 4847 31807
rect 5457 31773 5491 31807
rect 5917 31773 5951 31807
rect 6101 31773 6135 31807
rect 6193 31773 6227 31807
rect 6561 31773 6595 31807
rect 7021 31773 7055 31807
rect 7114 31773 7148 31807
rect 7297 31773 7331 31807
rect 7402 31773 7436 31807
rect 7527 31773 7561 31807
rect 8953 31773 8987 31807
rect 12449 31773 12483 31807
rect 12541 31773 12575 31807
rect 14657 31773 14691 31807
rect 14749 31773 14783 31807
rect 15117 31773 15151 31807
rect 15209 31773 15243 31807
rect 15393 31773 15427 31807
rect 15485 31773 15519 31807
rect 15761 31773 15795 31807
rect 15853 31773 15887 31807
rect 16575 31773 16609 31807
rect 17877 31773 17911 31807
rect 21465 31773 21499 31807
rect 21558 31773 21592 31807
rect 21741 31773 21775 31807
rect 21930 31773 21964 31807
rect 22753 31773 22787 31807
rect 23029 31773 23063 31807
rect 23581 31773 23615 31807
rect 24041 31773 24075 31807
rect 24409 31773 24443 31807
rect 24685 31773 24719 31807
rect 26985 31773 27019 31807
rect 27261 31773 27295 31807
rect 27445 31773 27479 31807
rect 27721 31773 27755 31807
rect 27813 31773 27847 31807
rect 28457 31773 28491 31807
rect 28641 31773 28675 31807
rect 29009 31773 29043 31807
rect 30849 31773 30883 31807
rect 31033 31773 31067 31807
rect 31309 31773 31343 31807
rect 31861 31773 31895 31807
rect 33517 31773 33551 31807
rect 33977 31773 34011 31807
rect 34161 31773 34195 31807
rect 34345 31773 34379 31807
rect 34437 31773 34471 31807
rect 34713 31773 34747 31807
rect 34897 31773 34931 31807
rect 35633 31773 35667 31807
rect 36001 31773 36035 31807
rect 36369 31773 36403 31807
rect 36553 31773 36587 31807
rect 37565 31773 37599 31807
rect 37657 31773 37691 31807
rect 37933 31773 37967 31807
rect 38577 31773 38611 31807
rect 15669 31705 15703 31739
rect 21833 31705 21867 31739
rect 24961 31705 24995 31739
rect 25145 31705 25179 31739
rect 26341 31705 26375 31739
rect 28825 31705 28859 31739
rect 29561 31705 29595 31739
rect 29745 31705 29779 31739
rect 33333 31705 33367 31739
rect 34069 31705 34103 31739
rect 37197 31705 37231 31739
rect 38209 31705 38243 31739
rect 2789 31637 2823 31671
rect 6929 31637 6963 31671
rect 7665 31637 7699 31671
rect 10701 31637 10735 31671
rect 14473 31637 14507 31671
rect 22109 31637 22143 31671
rect 24869 31637 24903 31671
rect 26551 31637 26585 31671
rect 28089 31637 28123 31671
rect 30849 31637 30883 31671
rect 33701 31637 33735 31671
rect 33793 31637 33827 31671
rect 16221 31433 16255 31467
rect 16773 31433 16807 31467
rect 23121 31433 23155 31467
rect 24317 31433 24351 31467
rect 26985 31433 27019 31467
rect 27629 31433 27663 31467
rect 29745 31433 29779 31467
rect 32505 31433 32539 31467
rect 35081 31433 35115 31467
rect 2513 31365 2547 31399
rect 15301 31365 15335 31399
rect 15853 31365 15887 31399
rect 16037 31365 16071 31399
rect 23949 31365 23983 31399
rect 24777 31365 24811 31399
rect 26709 31365 26743 31399
rect 33149 31365 33183 31399
rect 33655 31365 33689 31399
rect 37749 31365 37783 31399
rect 2053 31297 2087 31331
rect 2237 31297 2271 31331
rect 4905 31297 4939 31331
rect 4997 31297 5031 31331
rect 6653 31297 6687 31331
rect 8953 31297 8987 31331
rect 11529 31297 11563 31331
rect 14381 31297 14415 31331
rect 15485 31297 15519 31331
rect 16313 31297 16347 31331
rect 16681 31297 16715 31331
rect 16865 31297 16899 31331
rect 21373 31297 21407 31331
rect 21557 31297 21591 31331
rect 21833 31297 21867 31331
rect 22293 31297 22327 31331
rect 23029 31297 23063 31331
rect 23673 31297 23707 31331
rect 23821 31297 23855 31331
rect 24041 31297 24075 31331
rect 24138 31297 24172 31331
rect 24593 31297 24627 31331
rect 25421 31297 25455 31331
rect 25513 31297 25547 31331
rect 25697 31297 25731 31331
rect 25789 31297 25823 31331
rect 25881 31297 25915 31331
rect 27353 31297 27387 31331
rect 27721 31297 27755 31331
rect 29285 31297 29319 31331
rect 29653 31297 29687 31331
rect 29929 31297 29963 31331
rect 31493 31297 31527 31331
rect 31677 31297 31711 31331
rect 32137 31297 32171 31331
rect 32597 31297 32631 31331
rect 33333 31297 33367 31331
rect 33425 31297 33459 31331
rect 33517 31297 33551 31331
rect 34897 31297 34931 31331
rect 38025 31297 38059 31331
rect 38485 31297 38519 31331
rect 38761 31297 38795 31331
rect 4261 31229 4295 31263
rect 6929 31229 6963 31263
rect 8861 31229 8895 31263
rect 9321 31229 9355 31263
rect 11805 31229 11839 31263
rect 13553 31229 13587 31263
rect 14473 31229 14507 31263
rect 16957 31229 16991 31263
rect 17233 31229 17267 31263
rect 18797 31229 18831 31263
rect 19073 31229 19107 31263
rect 20637 31229 20671 31263
rect 21925 31229 21959 31263
rect 22385 31229 22419 31263
rect 22569 31229 22603 31263
rect 24409 31229 24443 31263
rect 27445 31229 27479 31263
rect 29561 31229 29595 31263
rect 30389 31229 30423 31263
rect 32229 31229 32263 31263
rect 33793 31229 33827 31263
rect 34253 31229 34287 31263
rect 34345 31229 34379 31263
rect 34437 31229 34471 31263
rect 34529 31229 34563 31263
rect 34713 31229 34747 31263
rect 38301 31229 38335 31263
rect 39313 31229 39347 31263
rect 39589 31229 39623 31263
rect 5273 31161 5307 31195
rect 15669 31161 15703 31195
rect 25237 31161 25271 31195
rect 34069 31161 34103 31195
rect 38945 31161 38979 31195
rect 1869 31093 1903 31127
rect 5089 31093 5123 31127
rect 8401 31093 8435 31127
rect 14749 31093 14783 31127
rect 16405 31093 16439 31127
rect 18705 31093 18739 31127
rect 20545 31093 20579 31127
rect 21281 31093 21315 31127
rect 21373 31093 21407 31127
rect 22017 31093 22051 31127
rect 22201 31093 22235 31127
rect 22293 31093 22327 31127
rect 27261 31093 27295 31127
rect 29101 31093 29135 31127
rect 29469 31093 29503 31127
rect 30113 31093 30147 31127
rect 31861 31093 31895 31127
rect 32137 31093 32171 31127
rect 32689 31093 32723 31127
rect 37841 31093 37875 31127
rect 38485 31093 38519 31127
rect 38669 31093 38703 31127
rect 41061 31093 41095 31127
rect 3801 30889 3835 30923
rect 12909 30889 12943 30923
rect 17601 30889 17635 30923
rect 20545 30889 20579 30923
rect 22201 30889 22235 30923
rect 24409 30889 24443 30923
rect 26065 30889 26099 30923
rect 32229 30889 32263 30923
rect 38209 30889 38243 30923
rect 38761 30889 38795 30923
rect 39865 30889 39899 30923
rect 12357 30821 12391 30855
rect 24961 30821 24995 30855
rect 36001 30821 36035 30855
rect 37197 30821 37231 30855
rect 39497 30821 39531 30855
rect 1685 30753 1719 30787
rect 4353 30753 4387 30787
rect 10977 30753 11011 30787
rect 12633 30753 12667 30787
rect 17785 30753 17819 30787
rect 18153 30753 18187 30787
rect 19901 30753 19935 30787
rect 24777 30753 24811 30787
rect 28273 30753 28307 30787
rect 28733 30753 28767 30787
rect 31401 30753 31435 30787
rect 36737 30753 36771 30787
rect 37289 30753 37323 30787
rect 1409 30685 1443 30719
rect 4261 30685 4295 30719
rect 11253 30685 11287 30719
rect 11713 30685 11747 30719
rect 12173 30685 12207 30719
rect 12541 30685 12575 30719
rect 12725 30685 12759 30719
rect 12817 30685 12851 30719
rect 13001 30685 13035 30719
rect 17877 30685 17911 30719
rect 18337 30685 18371 30719
rect 19257 30685 19291 30719
rect 19993 30685 20027 30719
rect 20269 30685 20303 30719
rect 20361 30685 20395 30719
rect 21005 30685 21039 30719
rect 21189 30685 21223 30719
rect 21557 30685 21591 30719
rect 21650 30685 21684 30719
rect 21833 30685 21867 30719
rect 22063 30685 22097 30719
rect 24685 30685 24719 30719
rect 24869 30685 24903 30719
rect 25145 30685 25179 30719
rect 25329 30685 25363 30719
rect 25421 30685 25455 30719
rect 26249 30685 26283 30719
rect 26433 30685 26467 30719
rect 26709 30685 26743 30719
rect 26893 30685 26927 30719
rect 28641 30685 28675 30719
rect 28917 30685 28951 30719
rect 31217 30685 31251 30719
rect 31309 30685 31343 30719
rect 31493 30685 31527 30719
rect 32137 30685 32171 30719
rect 32229 30685 32263 30719
rect 33793 30685 33827 30719
rect 33977 30685 34011 30719
rect 35725 30685 35759 30719
rect 36001 30685 36035 30719
rect 36829 30685 36863 30719
rect 37841 30685 37875 30719
rect 37933 30685 37967 30719
rect 38301 30685 38335 30719
rect 38853 30685 38887 30719
rect 39037 30685 39071 30719
rect 39313 30685 39347 30719
rect 40049 30685 40083 30719
rect 3433 30617 3467 30651
rect 10609 30617 10643 30651
rect 10793 30617 10827 30651
rect 11069 30617 11103 30651
rect 11437 30617 11471 30651
rect 11529 30617 11563 30651
rect 18245 30617 18279 30651
rect 18822 30617 18856 30651
rect 20177 30617 20211 30651
rect 21925 30617 21959 30651
rect 25789 30617 25823 30651
rect 25973 30617 26007 30651
rect 26617 30617 26651 30651
rect 31769 30617 31803 30651
rect 38577 30617 38611 30651
rect 4169 30549 4203 30583
rect 11805 30549 11839 30583
rect 18613 30549 18647 30583
rect 18705 30549 18739 30583
rect 18981 30549 19015 30583
rect 21373 30549 21407 30583
rect 25605 30549 25639 30583
rect 26801 30549 26835 30583
rect 31033 30549 31067 30583
rect 32413 30549 32447 30583
rect 33885 30549 33919 30583
rect 37565 30549 37599 30583
rect 38485 30549 38519 30583
rect 39221 30549 39255 30583
rect 2421 30345 2455 30379
rect 2789 30345 2823 30379
rect 18521 30345 18555 30379
rect 18889 30345 18923 30379
rect 27537 30345 27571 30379
rect 30113 30345 30147 30379
rect 32873 30345 32907 30379
rect 9597 30277 9631 30311
rect 9689 30277 9723 30311
rect 19901 30277 19935 30311
rect 20729 30277 20763 30311
rect 37381 30277 37415 30311
rect 8033 30209 8067 30243
rect 8126 30209 8160 30243
rect 8309 30209 8343 30243
rect 8401 30209 8435 30243
rect 8539 30209 8573 30243
rect 9321 30209 9355 30243
rect 9469 30209 9503 30243
rect 9827 30209 9861 30243
rect 17969 30209 18003 30243
rect 18337 30209 18371 30243
rect 18705 30209 18739 30243
rect 18889 30209 18923 30243
rect 20085 30209 20119 30243
rect 20545 30209 20579 30243
rect 21373 30209 21407 30243
rect 27721 30209 27755 30243
rect 29469 30209 29503 30243
rect 29617 30209 29651 30243
rect 29745 30209 29779 30243
rect 29837 30209 29871 30243
rect 29934 30209 29968 30243
rect 32229 30209 32263 30243
rect 32413 30209 32447 30243
rect 32873 30209 32907 30243
rect 32965 30209 32999 30243
rect 35265 30209 35299 30243
rect 35357 30209 35391 30243
rect 35725 30209 35759 30243
rect 35817 30209 35851 30243
rect 36093 30209 36127 30243
rect 36369 30209 36403 30243
rect 37933 30209 37967 30243
rect 38577 30209 38611 30243
rect 38945 30209 38979 30243
rect 2881 30141 2915 30175
rect 3065 30141 3099 30175
rect 20361 30141 20395 30175
rect 20913 30141 20947 30175
rect 21097 30141 21131 30175
rect 21649 30141 21683 30175
rect 27997 30141 28031 30175
rect 35909 30141 35943 30175
rect 38485 30141 38519 30175
rect 39313 30141 39347 30175
rect 39589 30141 39623 30175
rect 8677 30073 8711 30107
rect 21557 30073 21591 30107
rect 27905 30073 27939 30107
rect 35449 30073 35483 30107
rect 36369 30073 36403 30107
rect 37565 30073 37599 30107
rect 9965 30005 9999 30039
rect 18061 30005 18095 30039
rect 20177 30005 20211 30039
rect 32229 30005 32263 30039
rect 38025 30005 38059 30039
rect 38853 30005 38887 30039
rect 39129 30005 39163 30039
rect 41061 30005 41095 30039
rect 6009 29801 6043 29835
rect 6745 29801 6779 29835
rect 7849 29801 7883 29835
rect 13829 29801 13863 29835
rect 14749 29801 14783 29835
rect 17049 29801 17083 29835
rect 22477 29801 22511 29835
rect 25789 29801 25823 29835
rect 26157 29801 26191 29835
rect 26525 29801 26559 29835
rect 29561 29801 29595 29835
rect 33333 29801 33367 29835
rect 38853 29801 38887 29835
rect 39865 29801 39899 29835
rect 5089 29733 5123 29767
rect 15853 29733 15887 29767
rect 26709 29733 26743 29767
rect 30941 29733 30975 29767
rect 31401 29733 31435 29767
rect 33425 29733 33459 29767
rect 39405 29733 39439 29767
rect 5273 29665 5307 29699
rect 23765 29665 23799 29699
rect 26617 29665 26651 29699
rect 29285 29665 29319 29699
rect 30205 29665 30239 29699
rect 36277 29665 36311 29699
rect 2697 29597 2731 29631
rect 5365 29597 5399 29631
rect 5458 29597 5492 29631
rect 5733 29597 5767 29631
rect 5830 29597 5864 29631
rect 6101 29597 6135 29631
rect 6194 29597 6228 29631
rect 6469 29597 6503 29631
rect 6607 29597 6641 29631
rect 7205 29597 7239 29631
rect 7353 29597 7387 29631
rect 7711 29597 7745 29631
rect 8033 29597 8067 29631
rect 8126 29597 8160 29631
rect 8539 29597 8573 29631
rect 9505 29597 9539 29631
rect 9598 29597 9632 29631
rect 10011 29597 10045 29631
rect 12265 29597 12299 29631
rect 13185 29597 13219 29631
rect 13278 29597 13312 29631
rect 13461 29597 13495 29631
rect 13650 29597 13684 29631
rect 14105 29597 14139 29631
rect 14198 29597 14232 29631
rect 14611 29597 14645 29631
rect 14933 29597 14967 29631
rect 15209 29597 15243 29631
rect 15301 29597 15335 29631
rect 17785 29597 17819 29631
rect 23213 29597 23247 29631
rect 23489 29597 23523 29631
rect 23581 29597 23615 29631
rect 25789 29597 25823 29631
rect 25973 29597 26007 29631
rect 26341 29597 26375 29631
rect 26709 29597 26743 29631
rect 26893 29597 26927 29631
rect 29193 29597 29227 29631
rect 29377 29597 29411 29631
rect 29745 29597 29779 29631
rect 29837 29597 29871 29631
rect 30757 29597 30791 29631
rect 30849 29597 30883 29631
rect 31033 29597 31067 29631
rect 31217 29597 31251 29631
rect 31585 29597 31619 29631
rect 31677 29597 31711 29631
rect 32965 29597 32999 29631
rect 33057 29597 33091 29631
rect 33425 29597 33459 29631
rect 33793 29597 33827 29631
rect 34345 29597 34379 29631
rect 34713 29597 34747 29631
rect 34989 29597 35023 29631
rect 35633 29597 35667 29631
rect 36093 29597 36127 29631
rect 36737 29597 36771 29631
rect 36921 29597 36955 29631
rect 37749 29597 37783 29631
rect 38393 29597 38427 29631
rect 38485 29597 38519 29631
rect 38853 29597 38887 29631
rect 40049 29597 40083 29631
rect 4813 29529 4847 29563
rect 5641 29529 5675 29563
rect 6377 29529 6411 29563
rect 7481 29529 7515 29563
rect 7573 29529 7607 29563
rect 8309 29529 8343 29563
rect 8401 29529 8435 29563
rect 9781 29529 9815 29563
rect 9873 29529 9907 29563
rect 12449 29529 12483 29563
rect 13553 29529 13587 29563
rect 14381 29529 14415 29563
rect 14473 29529 14507 29563
rect 15117 29529 15151 29563
rect 15669 29529 15703 29563
rect 16957 29529 16991 29563
rect 17969 29529 18003 29563
rect 22293 29529 22327 29563
rect 30113 29529 30147 29563
rect 31401 29529 31435 29563
rect 38025 29529 38059 29563
rect 39221 29529 39255 29563
rect 2513 29461 2547 29495
rect 8677 29461 8711 29495
rect 10149 29461 10183 29495
rect 12633 29461 12667 29495
rect 15485 29461 15519 29495
rect 18153 29461 18187 29495
rect 22477 29461 22511 29495
rect 22661 29461 22695 29495
rect 23397 29461 23431 29495
rect 23765 29461 23799 29495
rect 30481 29461 30515 29495
rect 33149 29461 33183 29495
rect 34069 29461 34103 29495
rect 35909 29461 35943 29495
rect 37013 29461 37047 29495
rect 39037 29461 39071 29495
rect 2973 29257 3007 29291
rect 4629 29257 4663 29291
rect 6009 29257 6043 29291
rect 10609 29257 10643 29291
rect 12633 29257 12667 29291
rect 13461 29257 13495 29291
rect 13645 29257 13679 29291
rect 13921 29257 13955 29291
rect 14197 29257 14231 29291
rect 15945 29257 15979 29291
rect 17601 29257 17635 29291
rect 20821 29257 20855 29291
rect 23121 29257 23155 29291
rect 24133 29257 24167 29291
rect 30021 29257 30055 29291
rect 31493 29257 31527 29291
rect 2605 29189 2639 29223
rect 3341 29189 3375 29223
rect 4169 29189 4203 29223
rect 4905 29189 4939 29223
rect 4997 29189 5031 29223
rect 8217 29189 8251 29223
rect 8677 29189 8711 29223
rect 9505 29189 9539 29223
rect 9965 29189 9999 29223
rect 10057 29189 10091 29223
rect 12357 29189 12391 29223
rect 13093 29189 13127 29223
rect 16037 29189 16071 29223
rect 17325 29189 17359 29223
rect 33701 29189 33735 29223
rect 2053 29121 2087 29155
rect 2513 29121 2547 29155
rect 3433 29121 3467 29155
rect 4721 29121 4755 29155
rect 5089 29121 5123 29155
rect 5365 29121 5399 29155
rect 5458 29121 5492 29155
rect 5641 29121 5675 29155
rect 5733 29121 5767 29155
rect 5830 29121 5864 29155
rect 6377 29121 6411 29155
rect 6561 29121 6595 29155
rect 6653 29121 6687 29155
rect 6745 29121 6779 29155
rect 7297 29121 7331 29155
rect 7481 29121 7515 29155
rect 7573 29121 7607 29155
rect 7665 29121 7699 29155
rect 7941 29121 7975 29155
rect 8089 29121 8123 29155
rect 8309 29121 8343 29155
rect 8447 29121 8481 29155
rect 9413 29121 9447 29155
rect 9597 29121 9631 29155
rect 9689 29121 9723 29155
rect 9837 29121 9871 29155
rect 10195 29121 10229 29155
rect 10609 29121 10643 29155
rect 11977 29121 12011 29155
rect 12137 29121 12171 29155
rect 12265 29121 12299 29155
rect 12454 29121 12488 29155
rect 12817 29121 12851 29155
rect 12965 29121 12999 29155
rect 13185 29121 13219 29155
rect 13282 29121 13316 29155
rect 13553 29121 13587 29155
rect 13737 29121 13771 29155
rect 13829 29121 13863 29155
rect 14013 29121 14047 29155
rect 14289 29121 14323 29155
rect 14841 29121 14875 29155
rect 15301 29121 15335 29155
rect 15394 29121 15428 29155
rect 15577 29121 15611 29155
rect 15669 29121 15703 29155
rect 15766 29121 15800 29155
rect 16221 29121 16255 29155
rect 16405 29121 16439 29155
rect 16681 29121 16715 29155
rect 17233 29121 17267 29155
rect 17417 29121 17451 29155
rect 17969 29121 18003 29155
rect 18245 29121 18279 29155
rect 18521 29121 18555 29155
rect 18797 29121 18831 29155
rect 19257 29121 19291 29155
rect 20453 29121 20487 29155
rect 20545 29121 20579 29155
rect 21097 29121 21131 29155
rect 22201 29121 22235 29155
rect 22293 29121 22327 29155
rect 22477 29121 22511 29155
rect 23489 29121 23523 29155
rect 23949 29121 23983 29155
rect 24225 29121 24259 29155
rect 24869 29121 24903 29155
rect 25237 29121 25271 29155
rect 25421 29121 25455 29155
rect 29561 29121 29595 29155
rect 29745 29121 29779 29155
rect 29837 29121 29871 29155
rect 30941 29121 30975 29155
rect 31125 29121 31159 29155
rect 31217 29121 31251 29155
rect 31493 29121 31527 29155
rect 31861 29121 31895 29155
rect 32321 29121 32355 29155
rect 32543 29121 32577 29155
rect 33241 29121 33275 29155
rect 33425 29121 33459 29155
rect 34069 29121 34103 29155
rect 34437 29121 34471 29155
rect 34713 29121 34747 29155
rect 37289 29121 37323 29155
rect 37565 29121 37599 29155
rect 38393 29121 38427 29155
rect 2789 29053 2823 29087
rect 3617 29053 3651 29087
rect 9137 29053 9171 29087
rect 15025 29053 15059 29087
rect 19625 29053 19659 29087
rect 21281 29053 21315 29087
rect 21373 29053 21407 29087
rect 22385 29053 22419 29087
rect 23857 29053 23891 29087
rect 24777 29053 24811 29087
rect 31309 29053 31343 29087
rect 32781 29053 32815 29087
rect 32873 29053 32907 29087
rect 34897 29053 34931 29087
rect 35173 29053 35207 29087
rect 2145 28985 2179 29019
rect 4537 28985 4571 29019
rect 5273 28985 5307 29019
rect 6929 28985 6963 29019
rect 8585 28985 8619 29019
rect 8953 28985 8987 29019
rect 11069 28985 11103 29019
rect 16313 28985 16347 29019
rect 16865 28985 16899 29019
rect 17049 28985 17083 29019
rect 17693 28985 17727 29019
rect 18705 28985 18739 29019
rect 20913 28985 20947 29019
rect 22017 28985 22051 29019
rect 37565 28985 37599 29019
rect 1869 28917 1903 28951
rect 7849 28917 7883 28951
rect 10333 28917 10367 28951
rect 16405 28917 16439 28951
rect 17785 28917 17819 28951
rect 20637 28917 20671 28951
rect 23949 28917 23983 28951
rect 29561 28917 29595 28951
rect 38577 28917 38611 28951
rect 5457 28713 5491 28747
rect 11069 28713 11103 28747
rect 12081 28713 12115 28747
rect 15577 28713 15611 28747
rect 15853 28713 15887 28747
rect 16313 28713 16347 28747
rect 18153 28713 18187 28747
rect 19441 28713 19475 28747
rect 20453 28713 20487 28747
rect 20729 28713 20763 28747
rect 21649 28713 21683 28747
rect 21833 28713 21867 28747
rect 22845 28713 22879 28747
rect 23305 28713 23339 28747
rect 24961 28713 24995 28747
rect 25881 28713 25915 28747
rect 26065 28713 26099 28747
rect 27905 28713 27939 28747
rect 28457 28713 28491 28747
rect 28825 28713 28859 28747
rect 36921 28713 36955 28747
rect 5273 28645 5307 28679
rect 19625 28645 19659 28679
rect 19993 28645 20027 28679
rect 23581 28645 23615 28679
rect 32321 28645 32355 28679
rect 34713 28645 34747 28679
rect 1869 28577 1903 28611
rect 4997 28577 5031 28611
rect 7757 28577 7791 28611
rect 14933 28577 14967 28611
rect 15209 28577 15243 28611
rect 15761 28577 15795 28611
rect 20177 28577 20211 28611
rect 21195 28577 21229 28611
rect 22201 28577 22235 28611
rect 27997 28577 28031 28611
rect 35265 28577 35299 28611
rect 1593 28509 1627 28543
rect 5549 28509 5583 28543
rect 5733 28509 5767 28543
rect 5917 28509 5951 28543
rect 9873 28509 9907 28543
rect 10057 28509 10091 28543
rect 10149 28509 10183 28543
rect 10241 28509 10275 28543
rect 10701 28509 10735 28543
rect 11069 28509 11103 28543
rect 11529 28509 11563 28543
rect 11713 28509 11747 28543
rect 11897 28509 11931 28543
rect 12541 28509 12575 28543
rect 12817 28509 12851 28543
rect 12909 28509 12943 28543
rect 13093 28509 13127 28543
rect 13277 28509 13311 28543
rect 14657 28509 14691 28543
rect 14749 28509 14783 28543
rect 15025 28509 15059 28543
rect 15117 28509 15151 28543
rect 15301 28509 15335 28543
rect 15945 28509 15979 28543
rect 16221 28509 16255 28543
rect 16405 28509 16439 28543
rect 17233 28509 17267 28543
rect 18153 28509 18187 28543
rect 18337 28509 18371 28543
rect 19901 28509 19935 28543
rect 20269 28509 20303 28543
rect 20453 28509 20487 28543
rect 20913 28509 20947 28543
rect 21097 28509 21131 28543
rect 21465 28509 21499 28543
rect 21741 28509 21775 28543
rect 22017 28509 22051 28543
rect 22293 28509 22327 28543
rect 22845 28509 22879 28543
rect 23029 28509 23063 28543
rect 23121 28509 23155 28543
rect 23397 28509 23431 28543
rect 23489 28509 23523 28543
rect 23673 28509 23707 28543
rect 23765 28509 23799 28543
rect 23857 28509 23891 28543
rect 24041 28503 24075 28537
rect 24409 28509 24443 28543
rect 24777 28509 24811 28543
rect 25421 28509 25455 28543
rect 25513 28509 25547 28543
rect 25605 28509 25639 28543
rect 26157 28509 26191 28543
rect 26433 28509 26467 28543
rect 26525 28509 26559 28543
rect 26801 28509 26835 28543
rect 26985 28509 27019 28543
rect 27077 28509 27111 28543
rect 27169 28509 27203 28543
rect 27537 28509 27571 28543
rect 27721 28509 27755 28543
rect 28111 28522 28145 28556
rect 28457 28509 28491 28543
rect 28641 28509 28675 28543
rect 29198 28509 29232 28543
rect 31033 28509 31067 28543
rect 31493 28509 31527 28543
rect 31677 28509 31711 28543
rect 32597 28509 32631 28543
rect 33517 28509 33551 28543
rect 33793 28509 33827 28543
rect 34897 28509 34931 28543
rect 34989 28509 35023 28543
rect 35725 28509 35759 28543
rect 35909 28509 35943 28543
rect 36921 28509 36955 28543
rect 37105 28509 37139 28543
rect 3617 28441 3651 28475
rect 5825 28441 5859 28475
rect 7849 28441 7883 28475
rect 11805 28441 11839 28475
rect 13185 28441 13219 28475
rect 15577 28441 15611 28475
rect 17049 28441 17083 28475
rect 17509 28441 17543 28475
rect 17693 28441 17727 28475
rect 19257 28441 19291 28475
rect 19473 28441 19507 28475
rect 21281 28441 21315 28475
rect 23949 28441 23983 28475
rect 24593 28441 24627 28475
rect 24685 28441 24719 28475
rect 25697 28441 25731 28475
rect 26341 28441 26375 28475
rect 28825 28441 28859 28475
rect 29009 28441 29043 28475
rect 29101 28441 29135 28475
rect 32321 28441 32355 28475
rect 35357 28441 35391 28475
rect 36093 28441 36127 28475
rect 6101 28373 6135 28407
rect 7279 28373 7313 28407
rect 7757 28373 7791 28407
rect 10425 28373 10459 28407
rect 11253 28373 11287 28407
rect 12357 28373 12391 28407
rect 12725 28373 12759 28407
rect 13461 28373 13495 28407
rect 14473 28373 14507 28407
rect 17417 28373 17451 28407
rect 17785 28373 17819 28407
rect 20177 28373 20211 28407
rect 20637 28373 20671 28407
rect 25897 28373 25931 28407
rect 26709 28373 26743 28407
rect 27353 28373 27387 28407
rect 28273 28373 28307 28407
rect 31309 28373 31343 28407
rect 31585 28373 31619 28407
rect 32505 28373 32539 28407
rect 33609 28373 33643 28407
rect 10977 28169 11011 28203
rect 12633 28169 12667 28203
rect 28365 28169 28399 28203
rect 37657 28169 37691 28203
rect 38301 28169 38335 28203
rect 1685 28101 1719 28135
rect 5733 28101 5767 28135
rect 5917 28101 5951 28135
rect 10885 28101 10919 28135
rect 28089 28101 28123 28135
rect 28457 28101 28491 28135
rect 33793 28101 33827 28135
rect 35725 28101 35759 28135
rect 41061 28101 41095 28135
rect 1409 28033 1443 28067
rect 12173 28033 12207 28067
rect 12357 28033 12391 28067
rect 12449 28033 12483 28067
rect 12541 28033 12575 28067
rect 12725 28033 12759 28067
rect 20821 28033 20855 28067
rect 21005 28033 21039 28067
rect 21097 28033 21131 28067
rect 26249 28033 26283 28067
rect 26433 28033 26467 28067
rect 26985 28033 27019 28067
rect 27169 28033 27203 28067
rect 27813 28033 27847 28067
rect 27997 28033 28031 28067
rect 28181 28033 28215 28067
rect 28825 28033 28859 28067
rect 28917 28033 28951 28067
rect 34069 28033 34103 28067
rect 34897 28033 34931 28067
rect 36001 28033 36035 28067
rect 37933 28033 37967 28067
rect 38301 28033 38335 28067
rect 38485 28033 38519 28067
rect 39044 28033 39078 28067
rect 3433 27965 3467 27999
rect 6009 27965 6043 27999
rect 33977 27965 34011 27999
rect 36093 27965 36127 27999
rect 36369 27965 36403 27999
rect 36553 27965 36587 27999
rect 36737 27965 36771 27999
rect 37473 27965 37507 27999
rect 37565 27965 37599 27999
rect 37841 27965 37875 27999
rect 39313 27965 39347 27999
rect 20913 27897 20947 27931
rect 29101 27897 29135 27931
rect 34253 27897 34287 27931
rect 5457 27829 5491 27863
rect 11989 27829 12023 27863
rect 20637 27829 20671 27863
rect 26249 27829 26283 27863
rect 27353 27829 27387 27863
rect 28733 27829 28767 27863
rect 33793 27829 33827 27863
rect 37289 27829 37323 27863
rect 8217 27625 8251 27659
rect 9505 27625 9539 27659
rect 10517 27625 10551 27659
rect 13553 27625 13587 27659
rect 16589 27625 16623 27659
rect 19533 27625 19567 27659
rect 26893 27625 26927 27659
rect 27261 27625 27295 27659
rect 30665 27625 30699 27659
rect 37197 27625 37231 27659
rect 37657 27625 37691 27659
rect 39865 27625 39899 27659
rect 4905 27557 4939 27591
rect 15761 27557 15795 27591
rect 19257 27557 19291 27591
rect 19441 27557 19475 27591
rect 22753 27557 22787 27591
rect 24961 27557 24995 27591
rect 26617 27557 26651 27591
rect 30941 27557 30975 27591
rect 31769 27557 31803 27591
rect 38301 27557 38335 27591
rect 6653 27489 6687 27523
rect 10517 27489 10551 27523
rect 15301 27489 15335 27523
rect 15853 27489 15887 27523
rect 25053 27489 25087 27523
rect 27353 27489 27387 27523
rect 31125 27489 31159 27523
rect 37933 27489 37967 27523
rect 5917 27421 5951 27455
rect 6035 27421 6069 27455
rect 6193 27421 6227 27455
rect 7757 27421 7791 27455
rect 7849 27421 7883 27455
rect 8033 27421 8067 27455
rect 8125 27421 8159 27455
rect 8401 27421 8435 27455
rect 8493 27421 8527 27455
rect 8677 27421 8711 27455
rect 8769 27421 8803 27455
rect 9689 27421 9723 27455
rect 9781 27421 9815 27455
rect 9965 27421 9999 27455
rect 10057 27421 10091 27455
rect 10425 27421 10459 27455
rect 13461 27421 13495 27455
rect 13645 27421 13679 27455
rect 15669 27421 15703 27455
rect 16221 27421 16255 27455
rect 16497 27421 16531 27455
rect 16773 27421 16807 27455
rect 17601 27421 17635 27455
rect 17785 27421 17819 27455
rect 18429 27421 18463 27455
rect 19625 27421 19659 27455
rect 22293 27421 22327 27455
rect 22661 27421 22695 27455
rect 22845 27421 22879 27455
rect 24777 27421 24811 27455
rect 25145 27421 25179 27455
rect 25789 27421 25823 27455
rect 26157 27421 26191 27455
rect 26525 27421 26559 27455
rect 27077 27421 27111 27455
rect 31033 27421 31067 27455
rect 31217 27421 31251 27455
rect 31401 27421 31435 27455
rect 31677 27421 31711 27455
rect 31861 27421 31895 27455
rect 31953 27421 31987 27455
rect 32137 27421 32171 27455
rect 32321 27421 32355 27455
rect 33333 27421 33367 27455
rect 33609 27421 33643 27455
rect 33977 27421 34011 27455
rect 34161 27421 34195 27455
rect 34713 27421 34747 27455
rect 34897 27421 34931 27455
rect 35449 27421 35483 27455
rect 35633 27421 35667 27455
rect 37565 27421 37599 27455
rect 38025 27421 38059 27455
rect 38577 27421 38611 27455
rect 39589 27421 39623 27455
rect 40049 27421 40083 27455
rect 5181 27353 5215 27387
rect 5365 27353 5399 27387
rect 5457 27353 5491 27387
rect 7573 27353 7607 27387
rect 10149 27353 10183 27387
rect 15117 27353 15151 27387
rect 18061 27353 18095 27387
rect 18245 27353 18279 27387
rect 19257 27353 19291 27387
rect 24593 27353 24627 27387
rect 34437 27353 34471 27387
rect 37105 27353 37139 27387
rect 38301 27353 38335 27387
rect 10241 27285 10275 27319
rect 17601 27285 17635 27319
rect 22109 27285 22143 27319
rect 31493 27285 31527 27319
rect 32229 27285 32263 27319
rect 34805 27285 34839 27319
rect 35541 27285 35575 27319
rect 38209 27285 38243 27319
rect 38485 27285 38519 27319
rect 39405 27285 39439 27319
rect 6009 27081 6043 27115
rect 6929 27081 6963 27115
rect 8677 27081 8711 27115
rect 9045 27081 9079 27115
rect 9873 27081 9907 27115
rect 10609 27081 10643 27115
rect 12357 27081 12391 27115
rect 12633 27081 12667 27115
rect 14381 27081 14415 27115
rect 14933 27081 14967 27115
rect 15761 27081 15795 27115
rect 16865 27081 16899 27115
rect 18245 27081 18279 27115
rect 19073 27081 19107 27115
rect 23121 27081 23155 27115
rect 31125 27081 31159 27115
rect 31585 27081 31619 27115
rect 33701 27081 33735 27115
rect 40785 27081 40819 27115
rect 5825 27013 5859 27047
rect 6745 27013 6779 27047
rect 8217 27013 8251 27047
rect 9597 27013 9631 27047
rect 10241 27013 10275 27047
rect 13277 27013 13311 27047
rect 14749 27013 14783 27047
rect 18362 27013 18396 27047
rect 19993 27013 20027 27047
rect 25421 27013 25455 27047
rect 39313 27013 39347 27047
rect 7481 26945 7515 26979
rect 7573 26945 7607 26979
rect 7757 26945 7791 26979
rect 7849 26945 7883 26979
rect 7941 26945 7975 26979
rect 8089 26945 8123 26979
rect 8309 26945 8343 26979
rect 8447 26945 8481 26979
rect 8861 26945 8895 26979
rect 9137 26945 9171 26979
rect 9229 26945 9263 26979
rect 9377 26945 9411 26979
rect 9505 26945 9539 26979
rect 9733 26945 9767 26979
rect 9965 26945 9999 26979
rect 10058 26945 10092 26979
rect 10333 26945 10367 26979
rect 10430 26945 10464 26979
rect 12449 26945 12483 26979
rect 12725 26945 12759 26979
rect 12909 26945 12943 26979
rect 13057 26945 13091 26979
rect 13185 26945 13219 26979
rect 13415 26945 13449 26979
rect 13921 26945 13955 26979
rect 14197 26945 14231 26979
rect 14289 26945 14323 26979
rect 14841 26945 14875 26979
rect 15025 26945 15059 26979
rect 15117 26945 15151 26979
rect 15265 26945 15299 26979
rect 15393 26945 15427 26979
rect 15485 26945 15519 26979
rect 15582 26945 15616 26979
rect 16037 26945 16071 26979
rect 16405 26945 16439 26979
rect 16681 26945 16715 26979
rect 17509 26945 17543 26979
rect 17693 26945 17727 26979
rect 17877 26945 17911 26979
rect 18705 26945 18739 26979
rect 19349 26945 19383 26979
rect 19717 26945 19751 26979
rect 22017 26945 22051 26979
rect 22293 26945 22327 26979
rect 22661 26945 22695 26979
rect 22937 26945 22971 26979
rect 23213 26945 23247 26979
rect 23857 26945 23891 26979
rect 24317 26945 24351 26979
rect 25605 26945 25639 26979
rect 25881 26945 25915 26979
rect 29469 26945 29503 26979
rect 31401 26945 31435 26979
rect 33885 26945 33919 26979
rect 34161 26945 34195 26979
rect 34437 26945 34471 26979
rect 34621 26945 34655 26979
rect 34805 26945 34839 26979
rect 34897 26945 34931 26979
rect 37565 26945 37599 26979
rect 37749 26945 37783 26979
rect 38025 26945 38059 26979
rect 38209 26945 38243 26979
rect 1501 26877 1535 26911
rect 1777 26877 1811 26911
rect 6101 26877 6135 26911
rect 7021 26877 7055 26911
rect 11897 26877 11931 26911
rect 14657 26877 14691 26911
rect 15853 26877 15887 26911
rect 17325 26877 17359 26911
rect 18153 26877 18187 26911
rect 18797 26877 18831 26911
rect 19625 26877 19659 26911
rect 21833 26877 21867 26911
rect 22753 26877 22787 26911
rect 23489 26877 23523 26911
rect 23673 26877 23707 26911
rect 24593 26877 24627 26911
rect 26985 26877 27019 26911
rect 29745 26877 29779 26911
rect 31309 26877 31343 26911
rect 31677 26877 31711 26911
rect 31769 26877 31803 26911
rect 39037 26877 39071 26911
rect 5549 26809 5583 26843
rect 8585 26809 8619 26843
rect 12265 26809 12299 26843
rect 12449 26809 12483 26843
rect 13553 26809 13587 26843
rect 14105 26809 14139 26843
rect 16313 26809 16347 26843
rect 19165 26809 19199 26843
rect 21925 26809 21959 26843
rect 23397 26809 23431 26843
rect 27353 26809 27387 26843
rect 34989 26809 35023 26843
rect 3249 26741 3283 26775
rect 6469 26741 6503 26775
rect 7297 26741 7331 26775
rect 13737 26741 13771 26775
rect 14565 26741 14599 26775
rect 18521 26741 18555 26775
rect 18889 26741 18923 26775
rect 19533 26741 19567 26775
rect 23305 26741 23339 26775
rect 24041 26741 24075 26775
rect 24409 26741 24443 26775
rect 24501 26741 24535 26775
rect 25789 26741 25823 26775
rect 27445 26741 27479 26775
rect 29285 26741 29319 26775
rect 29653 26741 29687 26775
rect 34437 26741 34471 26775
rect 37565 26741 37599 26775
rect 38025 26741 38059 26775
rect 2145 26537 2179 26571
rect 5549 26537 5583 26571
rect 8493 26537 8527 26571
rect 9597 26537 9631 26571
rect 11897 26537 11931 26571
rect 13553 26537 13587 26571
rect 16681 26537 16715 26571
rect 18797 26537 18831 26571
rect 19349 26537 19383 26571
rect 20729 26537 20763 26571
rect 22661 26537 22695 26571
rect 23949 26537 23983 26571
rect 25329 26537 25363 26571
rect 29561 26537 29595 26571
rect 30021 26537 30055 26571
rect 31861 26537 31895 26571
rect 32045 26537 32079 26571
rect 38945 26537 38979 26571
rect 2881 26469 2915 26503
rect 5825 26469 5859 26503
rect 18981 26469 19015 26503
rect 19809 26469 19843 26503
rect 21557 26469 21591 26503
rect 23305 26469 23339 26503
rect 24133 26469 24167 26503
rect 25513 26469 25547 26503
rect 30205 26469 30239 26503
rect 30481 26469 30515 26503
rect 33517 26469 33551 26503
rect 35909 26469 35943 26503
rect 3433 26401 3467 26435
rect 23857 26401 23891 26435
rect 25789 26401 25823 26435
rect 29653 26401 29687 26435
rect 2329 26333 2363 26367
rect 3341 26333 3375 26367
rect 3801 26333 3835 26367
rect 7849 26333 7883 26367
rect 7997 26333 8031 26367
rect 8217 26333 8251 26367
rect 8355 26333 8389 26367
rect 8953 26333 8987 26367
rect 9101 26333 9135 26367
rect 9459 26333 9493 26367
rect 10517 26333 10551 26367
rect 10701 26333 10735 26367
rect 11253 26333 11287 26367
rect 11401 26333 11435 26367
rect 11529 26333 11563 26367
rect 11621 26333 11655 26367
rect 11759 26333 11793 26367
rect 12081 26333 12115 26367
rect 12265 26333 12299 26367
rect 12449 26333 12483 26367
rect 13277 26333 13311 26367
rect 13369 26333 13403 26367
rect 13645 26333 13679 26367
rect 16129 26333 16163 26367
rect 16405 26333 16439 26367
rect 16497 26333 16531 26367
rect 17785 26333 17819 26367
rect 18155 26333 18189 26367
rect 18337 26333 18371 26367
rect 19257 26333 19291 26367
rect 19625 26333 19659 26367
rect 20729 26333 20763 26367
rect 20913 26333 20947 26367
rect 21741 26333 21775 26367
rect 21833 26333 21867 26367
rect 22109 26333 22143 26367
rect 22201 26333 22235 26367
rect 22569 26333 22603 26367
rect 22753 26333 22787 26367
rect 23581 26333 23615 26367
rect 23765 26333 23799 26367
rect 24409 26333 24443 26367
rect 24777 26333 24811 26367
rect 24869 26333 24903 26367
rect 25145 26333 25179 26367
rect 25237 26333 25271 26367
rect 25973 26333 26007 26367
rect 26341 26333 26375 26367
rect 26712 26333 26746 26367
rect 26985 26333 27019 26367
rect 27537 26333 27571 26367
rect 27629 26333 27663 26367
rect 27813 26333 27847 26367
rect 27905 26333 27939 26367
rect 29009 26333 29043 26367
rect 29837 26333 29871 26367
rect 30389 26333 30423 26367
rect 30573 26333 30607 26367
rect 30665 26333 30699 26367
rect 32229 26333 32263 26367
rect 32689 26333 32723 26367
rect 32873 26333 32907 26367
rect 33241 26333 33275 26367
rect 33977 26333 34011 26367
rect 34161 26333 34195 26367
rect 35909 26333 35943 26367
rect 36093 26333 36127 26367
rect 36185 26333 36219 26367
rect 36369 26333 36403 26367
rect 38853 26333 38887 26367
rect 39681 26333 39715 26367
rect 4077 26265 4111 26299
rect 6101 26265 6135 26299
rect 6285 26265 6319 26299
rect 6377 26265 6411 26299
rect 8125 26265 8159 26299
rect 9229 26265 9263 26299
rect 9321 26265 9355 26299
rect 12725 26265 12759 26299
rect 13093 26265 13127 26299
rect 16313 26265 16347 26299
rect 17693 26265 17727 26299
rect 18245 26265 18279 26299
rect 18613 26265 18647 26299
rect 18797 26265 18831 26299
rect 21925 26265 21959 26299
rect 23305 26265 23339 26299
rect 25053 26265 25087 26299
rect 26525 26265 26559 26299
rect 29193 26265 29227 26299
rect 29377 26265 29411 26299
rect 29561 26265 29595 26299
rect 31677 26265 31711 26299
rect 31877 26265 31911 26299
rect 39313 26265 39347 26299
rect 39497 26265 39531 26299
rect 40693 26265 40727 26299
rect 3249 26197 3283 26231
rect 10701 26197 10735 26231
rect 23489 26197 23523 26231
rect 25973 26197 26007 26231
rect 26893 26197 26927 26231
rect 27353 26197 27387 26231
rect 33793 26197 33827 26231
rect 36277 26197 36311 26231
rect 40785 26197 40819 26231
rect 4629 25993 4663 26027
rect 8401 25993 8435 26027
rect 10977 25993 11011 26027
rect 21373 25993 21407 26027
rect 25053 25993 25087 26027
rect 28089 25993 28123 26027
rect 28641 25993 28675 26027
rect 37565 25993 37599 26027
rect 41061 25993 41095 26027
rect 3801 25925 3835 25959
rect 10701 25925 10735 25959
rect 18797 25925 18831 25959
rect 19349 25925 19383 25959
rect 35265 25925 35299 25959
rect 38577 25925 38611 25959
rect 2973 25857 3007 25891
rect 4537 25857 4571 25891
rect 7849 25857 7883 25891
rect 8033 25857 8067 25891
rect 8125 25857 8159 25891
rect 8217 25857 8251 25891
rect 10425 25857 10459 25891
rect 10609 25857 10643 25891
rect 10793 25857 10827 25891
rect 15209 25857 15243 25891
rect 16957 25857 16991 25891
rect 17417 25857 17451 25891
rect 19257 25857 19291 25891
rect 19441 25857 19475 25891
rect 20821 25857 20855 25891
rect 21005 25857 21039 25891
rect 21097 25857 21131 25891
rect 21189 25857 21223 25891
rect 21373 25857 21407 25891
rect 25237 25857 25271 25891
rect 25329 25857 25363 25891
rect 25421 25857 25455 25891
rect 25559 25857 25593 25891
rect 26065 25857 26099 25891
rect 26249 25857 26283 25891
rect 26341 25857 26375 25891
rect 26985 25857 27019 25891
rect 27169 25857 27203 25891
rect 27721 25857 27755 25891
rect 27905 25857 27939 25891
rect 28181 25857 28215 25891
rect 28457 25857 28491 25891
rect 29377 25857 29411 25891
rect 29929 25857 29963 25891
rect 30205 25857 30239 25891
rect 30757 25857 30791 25891
rect 35449 25857 35483 25891
rect 35541 25857 35575 25891
rect 37289 25857 37323 25891
rect 37749 25857 37783 25891
rect 38117 25857 38151 25891
rect 4813 25789 4847 25823
rect 25697 25789 25731 25823
rect 28273 25789 28307 25823
rect 30389 25789 30423 25823
rect 38853 25789 38887 25823
rect 39313 25789 39347 25823
rect 39589 25789 39623 25823
rect 27261 25721 27295 25755
rect 34897 25721 34931 25755
rect 4169 25653 4203 25687
rect 15025 25653 15059 25687
rect 16773 25653 16807 25687
rect 19073 25653 19107 25687
rect 20637 25653 20671 25687
rect 27445 25653 27479 25687
rect 27813 25653 27847 25687
rect 35541 25653 35575 25687
rect 38301 25653 38335 25687
rect 3801 25449 3835 25483
rect 9781 25449 9815 25483
rect 14289 25449 14323 25483
rect 25421 25449 25455 25483
rect 27905 25449 27939 25483
rect 29561 25449 29595 25483
rect 30297 25449 30331 25483
rect 31125 25449 31159 25483
rect 31493 25449 31527 25483
rect 32781 25449 32815 25483
rect 33793 25449 33827 25483
rect 34989 25449 35023 25483
rect 37841 25449 37875 25483
rect 39865 25449 39899 25483
rect 40785 25449 40819 25483
rect 7757 25381 7791 25415
rect 11805 25381 11839 25415
rect 13737 25381 13771 25415
rect 24961 25381 24995 25415
rect 31953 25381 31987 25415
rect 33149 25381 33183 25415
rect 37657 25381 37691 25415
rect 38945 25381 38979 25415
rect 1409 25313 1443 25347
rect 7205 25313 7239 25347
rect 10793 25313 10827 25347
rect 10885 25313 10919 25347
rect 12265 25313 12299 25347
rect 13369 25313 13403 25347
rect 14749 25313 14783 25347
rect 15025 25313 15059 25347
rect 20545 25313 20579 25347
rect 21189 25313 21223 25347
rect 21833 25313 21867 25347
rect 30573 25313 30607 25347
rect 31217 25313 31251 25347
rect 34069 25313 34103 25347
rect 35357 25313 35391 25347
rect 35817 25313 35851 25347
rect 37841 25313 37875 25347
rect 3985 25245 4019 25279
rect 9229 25245 9263 25279
rect 9413 25245 9447 25279
rect 9505 25245 9539 25279
rect 9597 25245 9631 25279
rect 10517 25245 10551 25279
rect 10609 25245 10643 25279
rect 11253 25245 11287 25279
rect 11437 25245 11471 25279
rect 11529 25245 11563 25279
rect 11989 25245 12023 25279
rect 12081 25245 12115 25279
rect 12173 25245 12207 25279
rect 12449 25245 12483 25279
rect 17049 25245 17083 25279
rect 17969 25245 18003 25279
rect 18061 25245 18095 25279
rect 19993 25245 20027 25279
rect 20177 25245 20211 25279
rect 21281 25245 21315 25279
rect 21649 25245 21683 25279
rect 25145 25245 25179 25279
rect 25237 25245 25271 25279
rect 25513 25245 25547 25279
rect 27353 25245 27387 25279
rect 27629 25245 27663 25279
rect 27721 25245 27755 25279
rect 29745 25245 29779 25279
rect 29837 25245 29871 25279
rect 29929 25245 29963 25279
rect 30021 25245 30055 25279
rect 30481 25245 30515 25279
rect 30665 25245 30699 25279
rect 30757 25245 30791 25279
rect 31125 25245 31159 25279
rect 31953 25245 31987 25279
rect 32229 25245 32263 25279
rect 32965 25245 32999 25279
rect 33057 25245 33091 25279
rect 33241 25245 33275 25279
rect 33425 25245 33459 25279
rect 34161 25245 34195 25279
rect 35541 25245 35575 25279
rect 35725 25245 35759 25279
rect 35927 25245 35961 25279
rect 36087 25245 36121 25279
rect 37013 25245 37047 25279
rect 37197 25245 37231 25279
rect 37289 25245 37323 25279
rect 37473 25245 37507 25279
rect 37749 25245 37783 25279
rect 38761 25245 38795 25279
rect 40049 25245 40083 25279
rect 1685 25177 1719 25211
rect 7021 25177 7055 25211
rect 7573 25177 7607 25211
rect 14197 25177 14231 25211
rect 16681 25177 16715 25211
rect 18245 25177 18279 25211
rect 20637 25177 20671 25211
rect 27537 25177 27571 25211
rect 32137 25177 32171 25211
rect 33701 25177 33735 25211
rect 40693 25177 40727 25211
rect 3157 25109 3191 25143
rect 6653 25109 6687 25143
rect 7113 25109 7147 25143
rect 10333 25109 10367 25143
rect 11069 25109 11103 25143
rect 13829 25109 13863 25143
rect 16497 25109 16531 25143
rect 17969 25109 18003 25143
rect 20177 25109 20211 25143
rect 34345 25109 34379 25143
rect 37105 25109 37139 25143
rect 38117 25109 38151 25143
rect 1869 24905 1903 24939
rect 2881 24905 2915 24939
rect 2973 24905 3007 24939
rect 5181 24905 5215 24939
rect 5825 24905 5859 24939
rect 8125 24905 8159 24939
rect 9781 24905 9815 24939
rect 10977 24905 11011 24939
rect 11253 24905 11287 24939
rect 14013 24905 14047 24939
rect 15117 24905 15151 24939
rect 18429 24905 18463 24939
rect 19901 24905 19935 24939
rect 22017 24905 22051 24939
rect 26985 24905 27019 24939
rect 33333 24905 33367 24939
rect 15485 24837 15519 24871
rect 15577 24837 15611 24871
rect 19533 24837 19567 24871
rect 19738 24837 19772 24871
rect 21833 24837 21867 24871
rect 22109 24837 22143 24871
rect 22201 24837 22235 24871
rect 22845 24837 22879 24871
rect 27261 24837 27295 24871
rect 2053 24769 2087 24803
rect 4353 24769 4387 24803
rect 4537 24769 4571 24803
rect 4629 24769 4663 24803
rect 4905 24769 4939 24803
rect 5365 24769 5399 24803
rect 5549 24769 5583 24803
rect 6193 24769 6227 24803
rect 6377 24769 6411 24803
rect 8217 24769 8251 24803
rect 8585 24769 8619 24803
rect 8677 24769 8711 24803
rect 9505 24769 9539 24803
rect 10793 24769 10827 24803
rect 10885 24769 10919 24803
rect 11253 24769 11287 24803
rect 12173 24769 12207 24803
rect 13001 24769 13035 24803
rect 13185 24769 13219 24803
rect 13277 24769 13311 24803
rect 13415 24769 13449 24803
rect 13737 24769 13771 24803
rect 13829 24769 13863 24803
rect 14473 24769 14507 24803
rect 14657 24769 14691 24803
rect 14749 24769 14783 24803
rect 14841 24769 14875 24803
rect 17325 24769 17359 24803
rect 17509 24769 17543 24803
rect 17785 24769 17819 24803
rect 19073 24769 19107 24803
rect 19257 24769 19291 24803
rect 20637 24769 20671 24803
rect 21005 24769 21039 24803
rect 21373 24769 21407 24803
rect 22569 24769 22603 24803
rect 22662 24769 22696 24803
rect 22937 24769 22971 24803
rect 23034 24769 23068 24803
rect 26985 24769 27019 24803
rect 28181 24769 28215 24803
rect 28273 24769 28307 24803
rect 28457 24769 28491 24803
rect 28549 24769 28583 24803
rect 32137 24769 32171 24803
rect 32321 24769 32355 24803
rect 32597 24769 32631 24803
rect 33057 24769 33091 24803
rect 33241 24769 33275 24803
rect 34161 24769 34195 24803
rect 35347 24769 35381 24803
rect 35541 24769 35575 24803
rect 3157 24701 3191 24735
rect 4721 24701 4755 24735
rect 5273 24701 5307 24735
rect 5917 24701 5951 24735
rect 6653 24701 6687 24735
rect 9321 24701 9355 24735
rect 9873 24701 9907 24735
rect 15761 24701 15795 24735
rect 17601 24701 17635 24735
rect 19165 24701 19199 24735
rect 19349 24701 19383 24735
rect 22385 24701 22419 24735
rect 27997 24701 28031 24735
rect 32689 24701 32723 24735
rect 33977 24701 34011 24735
rect 39313 24701 39347 24735
rect 39589 24701 39623 24735
rect 41061 24701 41095 24735
rect 2513 24633 2547 24667
rect 6009 24633 6043 24667
rect 12357 24633 12391 24667
rect 17969 24633 18003 24667
rect 18061 24633 18095 24667
rect 18889 24633 18923 24667
rect 21281 24633 21315 24667
rect 27077 24633 27111 24667
rect 4353 24565 4387 24599
rect 8861 24565 8895 24599
rect 11161 24565 11195 24599
rect 13553 24565 13587 24599
rect 15025 24565 15059 24599
rect 17325 24565 17359 24599
rect 18429 24565 18463 24599
rect 18613 24565 18647 24599
rect 19717 24565 19751 24599
rect 23213 24565 23247 24599
rect 32137 24565 32171 24599
rect 32597 24565 32631 24599
rect 32965 24565 32999 24599
rect 34345 24565 34379 24599
rect 35449 24565 35483 24599
rect 4905 24361 4939 24395
rect 5641 24361 5675 24395
rect 8309 24361 8343 24395
rect 9505 24361 9539 24395
rect 14565 24361 14599 24395
rect 22385 24361 22419 24395
rect 23857 24361 23891 24395
rect 24409 24361 24443 24395
rect 24961 24361 24995 24395
rect 25697 24361 25731 24395
rect 27905 24361 27939 24395
rect 28733 24361 28767 24395
rect 29929 24361 29963 24395
rect 31493 24361 31527 24395
rect 31769 24361 31803 24395
rect 40141 24361 40175 24395
rect 3801 24293 3835 24327
rect 5273 24293 5307 24327
rect 7389 24293 7423 24327
rect 12909 24293 12943 24327
rect 24041 24293 24075 24327
rect 25881 24293 25915 24327
rect 27353 24293 27387 24327
rect 28181 24293 28215 24327
rect 30297 24293 30331 24327
rect 30941 24293 30975 24327
rect 33517 24293 33551 24327
rect 34069 24293 34103 24327
rect 4353 24225 4387 24259
rect 7021 24225 7055 24259
rect 7941 24225 7975 24259
rect 12817 24225 12851 24259
rect 17049 24225 17083 24259
rect 18245 24225 18279 24259
rect 19901 24225 19935 24259
rect 23305 24225 23339 24259
rect 24593 24225 24627 24259
rect 25329 24225 25363 24259
rect 25421 24225 25455 24259
rect 27261 24225 27295 24259
rect 29101 24225 29135 24259
rect 33333 24225 33367 24259
rect 34253 24225 34287 24259
rect 37565 24225 37599 24259
rect 2973 24157 3007 24191
rect 4169 24157 4203 24191
rect 4905 24157 4939 24191
rect 5089 24157 5123 24191
rect 5181 24157 5215 24191
rect 5549 24157 5583 24191
rect 5917 24157 5951 24191
rect 6745 24157 6779 24191
rect 8493 24157 8527 24191
rect 8585 24157 8619 24191
rect 8953 24157 8987 24191
rect 9137 24157 9171 24191
rect 9229 24157 9263 24191
rect 9321 24157 9355 24191
rect 11529 24157 11563 24191
rect 11989 24157 12023 24191
rect 12357 24157 12391 24191
rect 13093 24157 13127 24191
rect 13415 24157 13449 24191
rect 13553 24157 13587 24191
rect 15485 24157 15519 24191
rect 15669 24157 15703 24191
rect 15945 24157 15979 24191
rect 17233 24157 17267 24191
rect 17785 24157 17819 24191
rect 18337 24157 18371 24191
rect 18705 24157 18739 24191
rect 20085 24157 20119 24191
rect 22569 24157 22603 24191
rect 22661 24157 22695 24191
rect 22845 24157 22879 24191
rect 22937 24157 22971 24191
rect 23121 24157 23155 24191
rect 24685 24157 24719 24191
rect 25145 24157 25179 24191
rect 27169 24157 27203 24191
rect 27434 24157 27468 24191
rect 27629 24157 27663 24191
rect 28089 24157 28123 24191
rect 28273 24157 28307 24191
rect 28365 24157 28399 24191
rect 28917 24157 28951 24191
rect 29193 24157 29227 24191
rect 30021 24157 30055 24191
rect 30113 24157 30147 24191
rect 30757 24157 30791 24191
rect 31033 24157 31067 24191
rect 31493 24157 31527 24191
rect 31585 24157 31619 24191
rect 33517 24157 33551 24191
rect 33977 24157 34011 24191
rect 34897 24157 34931 24191
rect 35081 24157 35115 24191
rect 37657 24157 37691 24191
rect 38301 24157 38335 24191
rect 38485 24157 38519 24191
rect 40325 24157 40359 24191
rect 5273 24089 5307 24123
rect 5641 24089 5675 24123
rect 7665 24089 7699 24123
rect 7849 24089 7883 24123
rect 8309 24089 8343 24123
rect 14473 24089 14507 24123
rect 17417 24089 17451 24123
rect 23673 24089 23707 24123
rect 24409 24089 24443 24123
rect 25513 24089 25547 24123
rect 25713 24089 25747 24123
rect 29837 24089 29871 24123
rect 31309 24089 31343 24123
rect 33885 24089 33919 24123
rect 34253 24089 34287 24123
rect 37933 24089 37967 24123
rect 38025 24089 38059 24123
rect 2789 24021 2823 24055
rect 4261 24021 4295 24055
rect 5457 24021 5491 24055
rect 5825 24021 5859 24055
rect 13737 24021 13771 24055
rect 15853 24021 15887 24055
rect 17601 24021 17635 24055
rect 18889 24021 18923 24055
rect 20269 24021 20303 24055
rect 23873 24021 23907 24055
rect 24869 24021 24903 24055
rect 26985 24021 27019 24055
rect 27721 24021 27755 24055
rect 30573 24021 30607 24055
rect 34989 24021 35023 24055
rect 37381 24021 37415 24055
rect 38393 24021 38427 24055
rect 7205 23817 7239 23851
rect 10057 23817 10091 23851
rect 12633 23817 12667 23851
rect 18337 23817 18371 23851
rect 20637 23817 20671 23851
rect 20729 23817 20763 23851
rect 26525 23817 26559 23851
rect 30021 23817 30055 23851
rect 31493 23817 31527 23851
rect 2697 23749 2731 23783
rect 14565 23749 14599 23783
rect 16957 23749 16991 23783
rect 17509 23749 17543 23783
rect 18245 23749 18279 23783
rect 20913 23749 20947 23783
rect 26249 23749 26283 23783
rect 35725 23749 35759 23783
rect 38761 23749 38795 23783
rect 39497 23749 39531 23783
rect 7389 23681 7423 23715
rect 7573 23681 7607 23715
rect 7665 23681 7699 23715
rect 9045 23681 9079 23715
rect 9138 23681 9172 23715
rect 9321 23681 9355 23715
rect 9413 23681 9447 23715
rect 9551 23681 9585 23715
rect 10241 23681 10275 23715
rect 10425 23681 10459 23715
rect 10793 23681 10827 23715
rect 10977 23681 11011 23715
rect 12817 23681 12851 23715
rect 13001 23681 13035 23715
rect 13105 23681 13139 23715
rect 14473 23681 14507 23715
rect 14657 23681 14691 23715
rect 15117 23681 15151 23715
rect 15485 23681 15519 23715
rect 15853 23681 15887 23715
rect 16681 23681 16715 23715
rect 16865 23681 16899 23715
rect 17049 23681 17083 23715
rect 20269 23681 20303 23715
rect 21097 23681 21131 23715
rect 21189 23681 21223 23715
rect 21373 23681 21407 23715
rect 21465 23681 21499 23715
rect 22017 23681 22051 23715
rect 22201 23681 22235 23715
rect 24593 23681 24627 23715
rect 24686 23681 24720 23715
rect 24869 23681 24903 23715
rect 24961 23681 24995 23715
rect 25058 23681 25092 23715
rect 26065 23681 26099 23715
rect 26341 23681 26375 23715
rect 26433 23681 26467 23715
rect 26617 23681 26651 23715
rect 28733 23681 28767 23715
rect 29009 23681 29043 23715
rect 29561 23681 29595 23715
rect 29745 23681 29779 23715
rect 29837 23681 29871 23715
rect 31033 23681 31067 23715
rect 31217 23681 31251 23715
rect 31309 23681 31343 23715
rect 32965 23681 32999 23715
rect 33517 23681 33551 23715
rect 33977 23681 34011 23715
rect 35081 23681 35115 23715
rect 35173 23681 35207 23715
rect 36921 23681 36955 23715
rect 37105 23681 37139 23715
rect 37289 23681 37323 23715
rect 37565 23681 37599 23715
rect 37749 23681 37783 23715
rect 37933 23681 37967 23715
rect 38577 23681 38611 23715
rect 38853 23681 38887 23715
rect 38945 23681 38979 23715
rect 39221 23681 39255 23715
rect 39405 23681 39439 23715
rect 39589 23681 39623 23715
rect 2421 23613 2455 23647
rect 4169 23613 4203 23647
rect 9965 23613 9999 23647
rect 20528 23613 20562 23647
rect 20821 23613 20855 23647
rect 22477 23613 22511 23647
rect 28825 23613 28859 23647
rect 35357 23613 35391 23647
rect 36461 23613 36495 23647
rect 7481 23545 7515 23579
rect 9689 23545 9723 23579
rect 17785 23545 17819 23579
rect 17969 23545 18003 23579
rect 26065 23545 26099 23579
rect 28917 23545 28951 23579
rect 33057 23545 33091 23579
rect 37565 23545 37599 23579
rect 39129 23545 39163 23579
rect 17233 23477 17267 23511
rect 20269 23477 20303 23511
rect 22385 23477 22419 23511
rect 25237 23477 25271 23511
rect 28549 23477 28583 23511
rect 29745 23477 29779 23511
rect 31309 23477 31343 23511
rect 36921 23477 36955 23511
rect 37749 23477 37783 23511
rect 39773 23477 39807 23511
rect 7757 23273 7791 23307
rect 11989 23273 12023 23307
rect 14841 23273 14875 23307
rect 23581 23273 23615 23307
rect 28273 23273 28307 23307
rect 40325 23273 40359 23307
rect 3157 23205 3191 23239
rect 9597 23205 9631 23239
rect 10241 23205 10275 23239
rect 1409 23137 1443 23171
rect 10701 23137 10735 23171
rect 14473 23137 14507 23171
rect 15577 23137 15611 23171
rect 15853 23137 15887 23171
rect 21097 23137 21131 23171
rect 21189 23137 21223 23171
rect 22845 23137 22879 23171
rect 25697 23137 25731 23171
rect 32781 23137 32815 23171
rect 36185 23137 36219 23171
rect 5089 23069 5123 23103
rect 5273 23069 5307 23103
rect 5365 23069 5399 23103
rect 5457 23069 5491 23103
rect 7205 23069 7239 23103
rect 7389 23069 7423 23103
rect 7481 23069 7515 23103
rect 7573 23069 7607 23103
rect 8953 23069 8987 23103
rect 9046 23069 9080 23103
rect 9321 23069 9355 23103
rect 9418 23069 9452 23103
rect 9965 23069 9999 23103
rect 10885 23069 10919 23103
rect 11253 23069 11287 23103
rect 11805 23069 11839 23103
rect 11897 23069 11931 23103
rect 12081 23069 12115 23103
rect 14381 23069 14415 23103
rect 14565 23069 14599 23103
rect 14657 23069 14691 23103
rect 15025 23069 15059 23103
rect 15761 23069 15795 23103
rect 15945 23069 15979 23103
rect 16037 23069 16071 23103
rect 17417 23069 17451 23103
rect 20913 23069 20947 23103
rect 23213 23069 23247 23103
rect 23397 23069 23431 23103
rect 25881 23069 25915 23103
rect 26065 23069 26099 23103
rect 26709 23069 26743 23103
rect 26893 23069 26927 23103
rect 27261 23069 27295 23103
rect 27905 23069 27939 23103
rect 28273 23069 28307 23103
rect 28457 23069 28491 23103
rect 31493 23069 31527 23103
rect 31677 23069 31711 23103
rect 31769 23069 31803 23103
rect 31953 23069 31987 23103
rect 32505 23069 32539 23103
rect 32689 23069 32723 23103
rect 34253 23069 34287 23103
rect 34437 23069 34471 23103
rect 36277 23069 36311 23103
rect 38669 23069 38703 23103
rect 38945 23069 38979 23103
rect 39037 23069 39071 23103
rect 1685 23001 1719 23035
rect 9229 23001 9263 23035
rect 15301 23001 15335 23035
rect 17969 23001 18003 23035
rect 21281 23001 21315 23035
rect 36553 23001 36587 23035
rect 36645 23001 36679 23035
rect 38853 23001 38887 23035
rect 39957 23001 39991 23035
rect 40141 23001 40175 23035
rect 5641 22933 5675 22967
rect 16129 22933 16163 22967
rect 17509 22933 17543 22967
rect 18061 22933 18095 22967
rect 20729 22933 20763 22967
rect 28089 22933 28123 22967
rect 31585 22933 31619 22967
rect 31861 22933 31895 22967
rect 34345 22933 34379 22967
rect 36001 22933 36035 22967
rect 39221 22933 39255 22967
rect 1869 22729 1903 22763
rect 2881 22729 2915 22763
rect 2973 22729 3007 22763
rect 5917 22729 5951 22763
rect 8309 22729 8343 22763
rect 8861 22729 8895 22763
rect 16497 22729 16531 22763
rect 34805 22729 34839 22763
rect 39865 22729 39899 22763
rect 8769 22661 8803 22695
rect 10241 22661 10275 22695
rect 12817 22661 12851 22695
rect 15577 22661 15611 22695
rect 18638 22661 18672 22695
rect 23857 22661 23891 22695
rect 24317 22661 24351 22695
rect 28457 22661 28491 22695
rect 31309 22661 31343 22695
rect 36211 22661 36245 22695
rect 38761 22661 38795 22695
rect 38853 22661 38887 22695
rect 2053 22593 2087 22627
rect 6561 22593 6595 22627
rect 9965 22593 9999 22627
rect 10149 22593 10183 22627
rect 10333 22593 10367 22627
rect 11529 22593 11563 22627
rect 12173 22593 12207 22627
rect 12541 22593 12575 22627
rect 12725 22593 12759 22627
rect 12909 22593 12943 22627
rect 13737 22593 13771 22627
rect 14657 22593 14691 22627
rect 14749 22593 14783 22627
rect 15301 22593 15335 22627
rect 15393 22593 15427 22627
rect 15669 22593 15703 22627
rect 15945 22593 15979 22627
rect 16129 22593 16163 22627
rect 16865 22593 16899 22627
rect 16958 22593 16992 22627
rect 17141 22593 17175 22627
rect 17233 22593 17267 22627
rect 17371 22593 17405 22627
rect 22293 22593 22327 22627
rect 22385 22593 22419 22627
rect 22569 22593 22603 22627
rect 22661 22593 22695 22627
rect 23673 22593 23707 22627
rect 23949 22593 23983 22627
rect 24041 22593 24075 22627
rect 28089 22593 28123 22627
rect 28273 22593 28307 22627
rect 29653 22593 29687 22627
rect 29929 22593 29963 22627
rect 30297 22593 30331 22627
rect 30573 22593 30607 22627
rect 30849 22593 30883 22627
rect 31493 22593 31527 22627
rect 31585 22593 31619 22627
rect 32505 22593 32539 22627
rect 32689 22593 32723 22627
rect 34713 22593 34747 22627
rect 34897 22593 34931 22627
rect 35909 22593 35943 22627
rect 36001 22593 36035 22627
rect 36093 22593 36127 22627
rect 36369 22593 36403 22627
rect 38485 22593 38519 22627
rect 38578 22593 38612 22627
rect 38991 22593 39025 22627
rect 39405 22593 39439 22627
rect 39681 22593 39715 22627
rect 3157 22525 3191 22559
rect 4169 22525 4203 22559
rect 4445 22525 4479 22559
rect 6837 22525 6871 22559
rect 9045 22525 9079 22559
rect 16221 22525 16255 22559
rect 18153 22525 18187 22559
rect 18429 22525 18463 22559
rect 18521 22525 18555 22559
rect 25053 22525 25087 22559
rect 29469 22525 29503 22559
rect 29745 22525 29779 22559
rect 39497 22525 39531 22559
rect 2513 22457 2547 22491
rect 11805 22457 11839 22491
rect 14841 22457 14875 22491
rect 29837 22457 29871 22491
rect 30389 22457 30423 22491
rect 30481 22457 30515 22491
rect 8401 22389 8435 22423
rect 10517 22389 10551 22423
rect 13093 22389 13127 22423
rect 14013 22389 14047 22423
rect 16221 22389 16255 22423
rect 17509 22389 17543 22423
rect 18797 22389 18831 22423
rect 22109 22389 22143 22423
rect 24225 22389 24259 22423
rect 30113 22389 30147 22423
rect 30941 22389 30975 22423
rect 31309 22389 31343 22423
rect 32505 22389 32539 22423
rect 35725 22389 35759 22423
rect 39129 22389 39163 22423
rect 39405 22389 39439 22423
rect 4537 22185 4571 22219
rect 5825 22185 5859 22219
rect 7205 22185 7239 22219
rect 13645 22185 13679 22219
rect 14749 22185 14783 22219
rect 26157 22185 26191 22219
rect 29929 22185 29963 22219
rect 13369 22117 13403 22151
rect 22845 22117 22879 22151
rect 22937 22117 22971 22151
rect 24685 22117 24719 22151
rect 25329 22117 25363 22151
rect 25605 22117 25639 22151
rect 30113 22117 30147 22151
rect 3065 22049 3099 22083
rect 5457 22049 5491 22083
rect 9873 22049 9907 22083
rect 17417 22049 17451 22083
rect 19809 22049 19843 22083
rect 20453 22049 20487 22083
rect 22753 22049 22787 22083
rect 24777 22049 24811 22083
rect 26801 22049 26835 22083
rect 28733 22049 28767 22083
rect 33701 22049 33735 22083
rect 4721 21981 4755 22015
rect 5273 21981 5307 22015
rect 7389 21981 7423 22015
rect 9045 21981 9079 22015
rect 9193 21981 9227 22015
rect 9321 21981 9355 22015
rect 9551 21981 9585 22015
rect 9781 21981 9815 22015
rect 10057 21981 10091 22015
rect 10241 21981 10275 22015
rect 10609 21981 10643 22015
rect 10793 21981 10827 22015
rect 10885 21981 10919 22015
rect 10978 21981 11012 22015
rect 11350 21981 11384 22015
rect 11989 21981 12023 22015
rect 12137 21981 12171 22015
rect 12265 21981 12299 22015
rect 12454 21981 12488 22015
rect 12725 21981 12759 22015
rect 12818 21981 12852 22015
rect 13190 21981 13224 22015
rect 13461 21981 13495 22015
rect 14105 21981 14139 22015
rect 14198 21981 14232 22015
rect 14611 21981 14645 22015
rect 17785 21981 17819 22015
rect 17969 21981 18003 22015
rect 18061 21981 18095 22015
rect 18337 21981 18371 22015
rect 18521 21981 18555 22015
rect 18889 21981 18923 22015
rect 18981 21981 19015 22015
rect 19993 21981 20027 22015
rect 20085 21981 20119 22015
rect 20315 21981 20349 22015
rect 20729 21981 20763 22015
rect 20822 21981 20856 22015
rect 20959 21981 20993 22015
rect 21213 21981 21247 22015
rect 21465 21981 21499 22015
rect 22109 21981 22143 22015
rect 22293 21981 22327 22015
rect 22385 21981 22419 22015
rect 23029 21981 23063 22015
rect 23213 21981 23247 22015
rect 23949 21981 23983 22015
rect 24593 21981 24627 22015
rect 24869 21981 24903 22015
rect 25513 21981 25547 22015
rect 25697 21981 25731 22015
rect 25789 21981 25823 22015
rect 25973 21981 26007 22015
rect 26709 21981 26743 22015
rect 27077 21981 27111 22015
rect 27169 21981 27203 22015
rect 27537 21981 27571 22015
rect 27905 21981 27939 22015
rect 27997 21981 28031 22015
rect 28273 21981 28307 22015
rect 28549 21981 28583 22015
rect 28641 21981 28675 22015
rect 28825 21981 28859 22015
rect 29561 21981 29595 22015
rect 29837 21981 29871 22015
rect 30021 21981 30055 22015
rect 30297 21981 30331 22015
rect 31401 21981 31435 22015
rect 31585 21981 31619 22015
rect 31677 21981 31711 22015
rect 31861 21981 31895 22015
rect 33885 21981 33919 22015
rect 34345 21981 34379 22015
rect 5733 21913 5767 21947
rect 9413 21913 9447 21947
rect 11161 21913 11195 21947
rect 11253 21913 11287 21947
rect 12357 21913 12391 21947
rect 13001 21913 13035 21947
rect 13093 21913 13127 21947
rect 14381 21913 14415 21947
rect 14473 21913 14507 21947
rect 18153 21913 18187 21947
rect 20177 21913 20211 21947
rect 21097 21913 21131 21947
rect 23765 21913 23799 21947
rect 27629 21913 27663 21947
rect 27721 21913 27755 21947
rect 31769 21913 31803 21947
rect 33977 21913 34011 21947
rect 34069 21913 34103 21947
rect 34207 21913 34241 21947
rect 2513 21845 2547 21879
rect 2881 21845 2915 21879
rect 2973 21845 3007 21879
rect 4813 21845 4847 21879
rect 5181 21845 5215 21879
rect 9689 21845 9723 21879
rect 11529 21845 11563 21879
rect 12633 21845 12667 21879
rect 13921 21845 13955 21879
rect 17509 21845 17543 21879
rect 21373 21845 21407 21879
rect 21649 21845 21683 21879
rect 21925 21845 21959 21879
rect 22477 21845 22511 21879
rect 24133 21845 24167 21879
rect 24409 21845 24443 21879
rect 27353 21845 27387 21879
rect 28089 21845 28123 21879
rect 28457 21845 28491 21879
rect 31493 21845 31527 21879
rect 7205 21641 7239 21675
rect 9505 21641 9539 21675
rect 10793 21641 10827 21675
rect 15393 21641 15427 21675
rect 17417 21641 17451 21675
rect 18889 21641 18923 21675
rect 22477 21641 22511 21675
rect 28365 21641 28399 21675
rect 33977 21641 34011 21675
rect 40877 21641 40911 21675
rect 9137 21573 9171 21607
rect 15025 21573 15059 21607
rect 15241 21573 15275 21607
rect 15853 21573 15887 21607
rect 18429 21573 18463 21607
rect 20545 21573 20579 21607
rect 22109 21573 22143 21607
rect 25881 21573 25915 21607
rect 27905 21573 27939 21607
rect 35357 21573 35391 21607
rect 35567 21573 35601 21607
rect 37289 21573 37323 21607
rect 2053 21505 2087 21539
rect 2605 21505 2639 21539
rect 6561 21505 6595 21539
rect 7113 21505 7147 21539
rect 8861 21505 8895 21539
rect 8954 21505 8988 21539
rect 9229 21505 9263 21539
rect 9367 21505 9401 21539
rect 10149 21505 10183 21539
rect 10297 21505 10331 21539
rect 10425 21505 10459 21539
rect 10517 21505 10551 21539
rect 10655 21505 10689 21539
rect 13461 21505 13495 21539
rect 17325 21505 17359 21539
rect 17693 21505 17727 21539
rect 18981 21505 19015 21539
rect 19165 21505 19199 21539
rect 20269 21505 20303 21539
rect 20361 21505 20395 21539
rect 20913 21505 20947 21539
rect 21078 21505 21112 21539
rect 21189 21505 21223 21539
rect 21281 21505 21315 21539
rect 21833 21505 21867 21539
rect 21926 21505 21960 21539
rect 22201 21505 22235 21539
rect 22339 21505 22373 21539
rect 24041 21505 24075 21539
rect 25697 21505 25731 21539
rect 25969 21495 26003 21529
rect 26065 21505 26099 21539
rect 27445 21505 27479 21539
rect 28089 21505 28123 21539
rect 28181 21505 28215 21539
rect 28457 21505 28491 21539
rect 28733 21505 28767 21539
rect 29193 21505 29227 21539
rect 33701 21505 33735 21539
rect 35265 21505 35299 21539
rect 35449 21505 35483 21539
rect 35725 21505 35759 21539
rect 37565 21505 37599 21539
rect 38945 21505 38979 21539
rect 39037 21505 39071 21539
rect 41061 21505 41095 21539
rect 2697 21437 2731 21471
rect 2973 21437 3007 21471
rect 7389 21437 7423 21471
rect 15485 21437 15519 21471
rect 15761 21437 15795 21471
rect 15970 21437 16004 21471
rect 17877 21437 17911 21471
rect 24133 21437 24167 21471
rect 37381 21437 37415 21471
rect 2421 21369 2455 21403
rect 4445 21369 4479 21403
rect 6745 21369 6779 21403
rect 13645 21369 13679 21403
rect 18797 21369 18831 21403
rect 25697 21369 25731 21403
rect 28825 21369 28859 21403
rect 35081 21369 35115 21403
rect 1869 21301 1903 21335
rect 6377 21301 6411 21335
rect 15209 21301 15243 21335
rect 16129 21301 16163 21335
rect 19165 21301 19199 21335
rect 19349 21301 19383 21335
rect 20729 21301 20763 21335
rect 24225 21301 24259 21335
rect 24409 21301 24443 21335
rect 26157 21301 26191 21335
rect 27537 21301 27571 21335
rect 27905 21301 27939 21335
rect 28917 21301 28951 21335
rect 29009 21301 29043 21335
rect 37289 21301 37323 21335
rect 37749 21301 37783 21335
rect 38945 21301 38979 21335
rect 39313 21301 39347 21335
rect 1672 21097 1706 21131
rect 3801 21097 3835 21131
rect 7665 21097 7699 21131
rect 14565 21097 14599 21131
rect 19441 21097 19475 21131
rect 21465 21097 21499 21131
rect 30941 21097 30975 21131
rect 33057 21097 33091 21131
rect 38761 21097 38795 21131
rect 39865 21097 39899 21131
rect 15025 21029 15059 21063
rect 15945 21029 15979 21063
rect 17233 21029 17267 21063
rect 27077 21029 27111 21063
rect 30573 21029 30607 21063
rect 35449 21029 35483 21063
rect 1409 20961 1443 20995
rect 3157 20961 3191 20995
rect 4445 20961 4479 20995
rect 5917 20961 5951 20995
rect 6193 20961 6227 20995
rect 11897 20961 11931 20995
rect 15577 20961 15611 20995
rect 16405 20961 16439 20995
rect 19349 20961 19383 20995
rect 21373 20961 21407 20995
rect 22753 20961 22787 20995
rect 27261 20961 27295 20995
rect 29929 20961 29963 20995
rect 38945 20961 38979 20995
rect 40049 20961 40083 20995
rect 4261 20893 4295 20927
rect 5273 20893 5307 20927
rect 5457 20893 5491 20927
rect 5549 20893 5583 20927
rect 5641 20893 5675 20927
rect 11621 20893 11655 20927
rect 14473 20893 14507 20927
rect 15761 20893 15795 20927
rect 16497 20893 16531 20927
rect 16773 20893 16807 20927
rect 16957 20893 16991 20927
rect 17325 20893 17359 20927
rect 19257 20893 19291 20927
rect 21189 20893 21223 20927
rect 21465 20893 21499 20927
rect 22477 20893 22511 20927
rect 22937 20893 22971 20927
rect 23305 20893 23339 20927
rect 23489 20893 23523 20927
rect 26985 20893 27019 20927
rect 29837 20893 29871 20927
rect 30021 20893 30055 20927
rect 30113 20893 30147 20927
rect 30849 20893 30883 20927
rect 31033 20893 31067 20927
rect 31125 20893 31159 20927
rect 31309 20893 31343 20927
rect 31401 20893 31435 20927
rect 32505 20893 32539 20927
rect 32781 20893 32815 20927
rect 32873 20893 32907 20927
rect 34897 20893 34931 20927
rect 35173 20893 35207 20927
rect 35265 20893 35299 20927
rect 35541 20893 35575 20927
rect 35634 20893 35668 20927
rect 35909 20893 35943 20927
rect 36006 20893 36040 20927
rect 37381 20893 37415 20927
rect 37474 20893 37508 20927
rect 37749 20893 37783 20927
rect 37887 20893 37921 20927
rect 39037 20893 39071 20927
rect 39865 20893 39899 20927
rect 40141 20893 40175 20927
rect 40601 20893 40635 20927
rect 15025 20825 15059 20859
rect 15485 20825 15519 20859
rect 15945 20825 15979 20859
rect 16681 20825 16715 20859
rect 31585 20825 31619 20859
rect 32689 20825 32723 20859
rect 35081 20825 35115 20859
rect 35817 20825 35851 20859
rect 37657 20825 37691 20859
rect 38761 20825 38795 20859
rect 40417 20825 40451 20859
rect 4169 20757 4203 20791
rect 5825 20757 5859 20791
rect 11253 20757 11287 20791
rect 11713 20757 11747 20791
rect 19625 20757 19659 20791
rect 21649 20757 21683 20791
rect 22569 20757 22603 20791
rect 27261 20757 27295 20791
rect 29653 20757 29687 20791
rect 31769 20757 31803 20791
rect 36185 20757 36219 20791
rect 38025 20757 38059 20791
rect 39221 20757 39255 20791
rect 40325 20757 40359 20791
rect 40785 20757 40819 20791
rect 5825 20553 5859 20587
rect 8861 20553 8895 20587
rect 9873 20553 9907 20587
rect 11713 20553 11747 20587
rect 14841 20553 14875 20587
rect 16313 20553 16347 20587
rect 19901 20553 19935 20587
rect 23305 20553 23339 20587
rect 28549 20553 28583 20587
rect 37749 20553 37783 20587
rect 40325 20553 40359 20587
rect 2697 20485 2731 20519
rect 7941 20485 7975 20519
rect 9321 20485 9355 20519
rect 15669 20485 15703 20519
rect 16773 20485 16807 20519
rect 20177 20485 20211 20519
rect 20821 20485 20855 20519
rect 21051 20485 21085 20519
rect 22845 20485 22879 20519
rect 25605 20485 25639 20519
rect 28181 20485 28215 20519
rect 28381 20485 28415 20519
rect 4353 20417 4387 20451
rect 5273 20417 5307 20451
rect 5457 20417 5491 20451
rect 5549 20417 5583 20451
rect 5641 20417 5675 20451
rect 7665 20417 7699 20451
rect 7849 20417 7883 20451
rect 8033 20417 8067 20451
rect 8769 20417 8803 20451
rect 9229 20417 9263 20451
rect 9689 20417 9723 20451
rect 10793 20417 10827 20451
rect 10977 20417 11011 20451
rect 11529 20417 11563 20451
rect 11897 20417 11931 20451
rect 12081 20417 12115 20451
rect 12173 20417 12207 20451
rect 12265 20417 12299 20451
rect 12725 20417 12759 20451
rect 15025 20417 15059 20451
rect 15209 20417 15243 20451
rect 15301 20417 15335 20451
rect 15485 20417 15519 20451
rect 15577 20417 15611 20451
rect 16129 20417 16163 20451
rect 17417 20417 17451 20451
rect 19901 20417 19935 20451
rect 20729 20417 20763 20451
rect 20913 20417 20947 20451
rect 23121 20417 23155 20451
rect 25973 20417 26007 20451
rect 27445 20417 27479 20451
rect 27629 20417 27663 20451
rect 31585 20417 31619 20451
rect 37289 20417 37323 20451
rect 37473 20417 37507 20451
rect 37565 20417 37599 20451
rect 39405 20417 39439 20451
rect 39589 20417 39623 20451
rect 39957 20417 39991 20451
rect 40141 20417 40175 20451
rect 3433 20349 3467 20383
rect 3709 20349 3743 20383
rect 9505 20349 9539 20383
rect 13093 20349 13127 20383
rect 13369 20349 13403 20383
rect 16037 20349 16071 20383
rect 21189 20349 21223 20383
rect 23029 20349 23063 20383
rect 31401 20349 31435 20383
rect 19993 20281 20027 20315
rect 8217 20213 8251 20247
rect 8585 20213 8619 20247
rect 10609 20213 10643 20247
rect 11253 20213 11287 20247
rect 12449 20213 12483 20247
rect 12541 20213 12575 20247
rect 15117 20213 15151 20247
rect 16865 20213 16899 20247
rect 17233 20213 17267 20247
rect 20545 20213 20579 20247
rect 22845 20213 22879 20247
rect 27813 20213 27847 20247
rect 28365 20213 28399 20247
rect 31769 20213 31803 20247
rect 37289 20213 37323 20247
rect 39405 20213 39439 20247
rect 39773 20213 39807 20247
rect 40141 20213 40175 20247
rect 3157 20009 3191 20043
rect 4905 20009 4939 20043
rect 8401 20009 8435 20043
rect 13553 20009 13587 20043
rect 17220 20009 17254 20043
rect 23765 20009 23799 20043
rect 25605 20009 25639 20043
rect 27721 20009 27755 20043
rect 28181 20009 28215 20043
rect 30113 20009 30147 20043
rect 31309 20009 31343 20043
rect 5641 19941 5675 19975
rect 9965 19941 9999 19975
rect 14105 19941 14139 19975
rect 19717 19941 19751 19975
rect 19809 19941 19843 19975
rect 29561 19941 29595 19975
rect 1409 19873 1443 19907
rect 10425 19873 10459 19907
rect 11621 19873 11655 19907
rect 11897 19873 11931 19907
rect 14749 19873 14783 19907
rect 16957 19873 16991 19907
rect 18981 19873 19015 19907
rect 20085 19873 20119 19907
rect 20269 19873 20303 19907
rect 20729 19873 20763 19907
rect 34069 19873 34103 19907
rect 34161 19873 34195 19907
rect 3985 19805 4019 19839
rect 4261 19805 4295 19839
rect 4354 19805 4388 19839
rect 4629 19805 4663 19839
rect 4767 19805 4801 19839
rect 4997 19805 5031 19839
rect 5090 19805 5124 19839
rect 5503 19805 5537 19839
rect 7757 19805 7791 19839
rect 7850 19805 7884 19839
rect 8222 19805 8256 19839
rect 9045 19805 9079 19839
rect 9229 19805 9263 19839
rect 9413 19805 9447 19839
rect 9689 19805 9723 19839
rect 10609 19805 10643 19839
rect 10977 19805 11011 19839
rect 11529 19805 11563 19839
rect 13737 19805 13771 19839
rect 14565 19805 14599 19839
rect 15209 19805 15243 19839
rect 15301 19805 15335 19839
rect 19625 19805 19659 19839
rect 19901 19805 19935 19839
rect 20361 19805 20395 19839
rect 23581 19805 23615 19839
rect 23857 19805 23891 19839
rect 24961 19805 24995 19839
rect 25109 19805 25143 19839
rect 25467 19805 25501 19839
rect 27445 19805 27479 19839
rect 28365 19805 28399 19839
rect 28549 19805 28583 19839
rect 28641 19805 28675 19839
rect 28989 19805 29023 19839
rect 29101 19805 29135 19839
rect 29193 19805 29227 19839
rect 29389 19805 29423 19839
rect 29837 19805 29871 19839
rect 29929 19805 29963 19839
rect 30021 19805 30055 19839
rect 30297 19805 30331 19839
rect 31493 19805 31527 19839
rect 31953 19805 31987 19839
rect 33333 19805 33367 19839
rect 33793 19805 33827 19839
rect 34253 19805 34287 19839
rect 34345 19805 34379 19839
rect 34713 19805 34747 19839
rect 34989 19805 35023 19839
rect 35081 19805 35115 19839
rect 1685 19737 1719 19771
rect 4537 19737 4571 19771
rect 5273 19737 5307 19771
rect 5365 19737 5399 19771
rect 8033 19737 8067 19771
rect 8125 19737 8159 19771
rect 8585 19737 8619 19771
rect 9321 19737 9355 19771
rect 25237 19737 25271 19771
rect 25329 19737 25363 19771
rect 27629 19737 27663 19771
rect 31585 19737 31619 19771
rect 31677 19737 31711 19771
rect 31815 19737 31849 19771
rect 33425 19737 33459 19771
rect 33517 19737 33551 19771
rect 33635 19737 33669 19771
rect 34897 19737 34931 19771
rect 3801 19669 3835 19703
rect 8677 19669 8711 19703
rect 9597 19669 9631 19703
rect 13369 19669 13403 19703
rect 14473 19669 14507 19703
rect 15485 19669 15519 19703
rect 19441 19669 19475 19703
rect 20453 19669 20487 19703
rect 20637 19669 20671 19703
rect 23397 19669 23431 19703
rect 28733 19669 28767 19703
rect 33149 19669 33183 19703
rect 33885 19669 33919 19703
rect 35265 19669 35299 19703
rect 1869 19465 1903 19499
rect 2237 19465 2271 19499
rect 2605 19465 2639 19499
rect 4813 19465 4847 19499
rect 5549 19465 5583 19499
rect 9873 19465 9907 19499
rect 12173 19465 12207 19499
rect 16957 19465 16991 19499
rect 25421 19465 25455 19499
rect 31401 19465 31435 19499
rect 3341 19397 3375 19431
rect 7297 19397 7331 19431
rect 8401 19397 8435 19431
rect 10057 19397 10091 19431
rect 18245 19397 18279 19431
rect 24685 19397 24719 19431
rect 25237 19397 25271 19431
rect 25789 19397 25823 19431
rect 27353 19397 27387 19431
rect 27445 19397 27479 19431
rect 27997 19397 28031 19431
rect 28181 19397 28215 19431
rect 30573 19397 30607 19431
rect 39405 19397 39439 19431
rect 2053 19329 2087 19363
rect 2697 19329 2731 19363
rect 3065 19329 3099 19363
rect 4905 19329 4939 19363
rect 4998 19329 5032 19363
rect 5181 19329 5215 19363
rect 5273 19329 5307 19363
rect 5411 19329 5445 19363
rect 7389 19329 7423 19363
rect 8125 19329 8159 19363
rect 12541 19329 12575 19363
rect 12633 19329 12667 19363
rect 15117 19329 15151 19363
rect 15301 19329 15335 19363
rect 15761 19329 15795 19363
rect 16221 19329 16255 19363
rect 17325 19329 17359 19363
rect 17417 19329 17451 19363
rect 18889 19329 18923 19363
rect 22017 19329 22051 19363
rect 22293 19329 22327 19363
rect 22661 19329 22695 19363
rect 23397 19329 23431 19363
rect 23489 19329 23523 19363
rect 23673 19329 23707 19363
rect 23765 19329 23799 19363
rect 24409 19329 24443 19363
rect 25053 19329 25087 19363
rect 25329 19329 25363 19363
rect 25605 19329 25639 19363
rect 25881 19329 25915 19363
rect 26525 19329 26559 19363
rect 27077 19329 27111 19363
rect 27170 19329 27204 19363
rect 27583 19329 27617 19363
rect 28733 19329 28767 19363
rect 28917 19329 28951 19363
rect 30389 19329 30423 19363
rect 30665 19329 30699 19363
rect 30757 19329 30791 19363
rect 31033 19329 31067 19363
rect 39589 19329 39623 19363
rect 39681 19329 39715 19363
rect 2881 19261 2915 19295
rect 7481 19261 7515 19295
rect 10793 19261 10827 19295
rect 12817 19261 12851 19295
rect 17601 19261 17635 19295
rect 18981 19261 19015 19295
rect 19165 19261 19199 19295
rect 21833 19261 21867 19295
rect 22385 19261 22419 19295
rect 22569 19261 22603 19295
rect 24225 19261 24259 19295
rect 24777 19261 24811 19295
rect 24869 19261 24903 19295
rect 26801 19261 26835 19295
rect 28549 19261 28583 19295
rect 31125 19261 31159 19295
rect 14565 19193 14599 19227
rect 14933 19193 14967 19227
rect 26341 19193 26375 19227
rect 26709 19193 26743 19227
rect 28365 19193 28399 19227
rect 6929 19125 6963 19159
rect 18337 19125 18371 19159
rect 19073 19125 19107 19159
rect 23213 19125 23247 19159
rect 27721 19125 27755 19159
rect 30941 19125 30975 19159
rect 31217 19125 31251 19159
rect 39405 19125 39439 19159
rect 39865 19125 39899 19159
rect 3801 18921 3835 18955
rect 6009 18921 6043 18955
rect 7849 18921 7883 18955
rect 8585 18921 8619 18955
rect 11989 18921 12023 18955
rect 12725 18921 12759 18955
rect 21465 18921 21499 18955
rect 22937 18921 22971 18955
rect 25513 18921 25547 18955
rect 26525 18921 26559 18955
rect 31309 18921 31343 18955
rect 36001 18921 36035 18955
rect 36461 18921 36495 18955
rect 37841 18921 37875 18955
rect 38485 18921 38519 18955
rect 40049 18921 40083 18955
rect 40233 18921 40267 18955
rect 23121 18853 23155 18887
rect 26709 18853 26743 18887
rect 33425 18853 33459 18887
rect 36645 18853 36679 18887
rect 4353 18785 4387 18819
rect 4721 18785 4755 18819
rect 7941 18785 7975 18819
rect 10517 18785 10551 18819
rect 16957 18785 16991 18819
rect 21189 18785 21223 18819
rect 22017 18785 22051 18819
rect 22845 18785 22879 18819
rect 23857 18785 23891 18819
rect 31953 18785 31987 18819
rect 36277 18785 36311 18819
rect 37105 18785 37139 18819
rect 5457 18717 5491 18751
rect 5641 18717 5675 18751
rect 5825 18717 5859 18751
rect 6101 18717 6135 18751
rect 10241 18717 10275 18751
rect 12081 18717 12115 18751
rect 12174 18717 12208 18751
rect 12357 18717 12391 18751
rect 12587 18717 12621 18751
rect 17141 18717 17175 18751
rect 20453 18717 20487 18751
rect 20729 18717 20763 18751
rect 21281 18717 21315 18751
rect 21741 18717 21775 18751
rect 21925 18717 21959 18751
rect 22937 18717 22971 18751
rect 23581 18717 23615 18751
rect 23673 18717 23707 18751
rect 23949 18717 23983 18751
rect 25145 18717 25179 18751
rect 25605 18717 25639 18751
rect 25698 18717 25732 18751
rect 26070 18717 26104 18751
rect 31493 18717 31527 18751
rect 31677 18717 31711 18751
rect 31795 18717 31829 18751
rect 32873 18717 32907 18751
rect 33057 18717 33091 18751
rect 33149 18717 33183 18751
rect 33241 18717 33275 18751
rect 33517 18717 33551 18751
rect 33793 18717 33827 18751
rect 33885 18717 33919 18751
rect 35449 18717 35483 18751
rect 35725 18717 35759 18751
rect 35817 18717 35851 18751
rect 36461 18717 36495 18751
rect 36737 18717 36771 18751
rect 36921 18717 36955 18751
rect 37841 18717 37875 18751
rect 38025 18717 38059 18751
rect 38485 18717 38519 18751
rect 38669 18717 38703 18751
rect 38761 18717 38795 18751
rect 39870 18717 39904 18751
rect 39957 18717 39991 18751
rect 4169 18649 4203 18683
rect 5273 18649 5307 18683
rect 5733 18649 5767 18683
rect 6377 18649 6411 18683
rect 12449 18649 12483 18683
rect 16497 18649 16531 18683
rect 17325 18649 17359 18683
rect 18613 18649 18647 18683
rect 20821 18649 20855 18683
rect 22661 18649 22695 18683
rect 25329 18649 25363 18683
rect 25881 18649 25915 18683
rect 25973 18649 26007 18683
rect 26341 18649 26375 18683
rect 31585 18649 31619 18683
rect 33701 18649 33735 18683
rect 35633 18649 35667 18683
rect 36185 18649 36219 18683
rect 37565 18649 37599 18683
rect 4261 18581 4295 18615
rect 16589 18581 16623 18615
rect 18705 18581 18739 18615
rect 20551 18581 20585 18615
rect 20637 18581 20671 18615
rect 21557 18581 21591 18615
rect 23397 18581 23431 18615
rect 26249 18581 26283 18615
rect 26541 18581 26575 18615
rect 34069 18581 34103 18615
rect 38209 18581 38243 18615
rect 38945 18581 38979 18615
rect 4997 18377 5031 18411
rect 7113 18377 7147 18411
rect 9137 18377 9171 18411
rect 14473 18377 14507 18411
rect 18705 18377 18739 18411
rect 35541 18377 35575 18411
rect 39957 18377 39991 18411
rect 40877 18377 40911 18411
rect 14565 18309 14599 18343
rect 37657 18309 37691 18343
rect 2881 18241 2915 18275
rect 3985 18241 4019 18275
rect 4905 18241 4939 18275
rect 5365 18241 5399 18275
rect 7297 18241 7331 18275
rect 15761 18241 15795 18275
rect 16037 18241 16071 18275
rect 16313 18241 16347 18275
rect 16497 18241 16531 18275
rect 16957 18241 16991 18275
rect 17049 18241 17083 18275
rect 18061 18241 18095 18275
rect 18245 18241 18279 18275
rect 18521 18241 18555 18275
rect 19349 18241 19383 18275
rect 29837 18241 29871 18275
rect 30389 18241 30423 18275
rect 30665 18241 30699 18275
rect 31401 18241 31435 18275
rect 34897 18241 34931 18275
rect 34990 18241 35024 18275
rect 35173 18241 35207 18275
rect 35265 18241 35299 18275
rect 35362 18241 35396 18275
rect 36461 18241 36495 18275
rect 36737 18241 36771 18275
rect 37841 18241 37875 18275
rect 37933 18241 37967 18275
rect 39497 18241 39531 18275
rect 39681 18241 39715 18275
rect 39773 18241 39807 18275
rect 40049 18241 40083 18275
rect 40509 18241 40543 18275
rect 40693 18241 40727 18275
rect 2973 18173 3007 18207
rect 3157 18173 3191 18207
rect 3433 18173 3467 18207
rect 5457 18173 5491 18207
rect 5549 18173 5583 18207
rect 6377 18173 6411 18207
rect 7021 18173 7055 18207
rect 9229 18173 9263 18207
rect 9413 18173 9447 18207
rect 14749 18173 14783 18207
rect 15853 18173 15887 18207
rect 16865 18173 16899 18207
rect 17141 18173 17175 18207
rect 18337 18173 18371 18207
rect 19441 18173 19475 18207
rect 19625 18173 19659 18207
rect 30021 18173 30055 18207
rect 30113 18173 30147 18207
rect 31493 18173 31527 18207
rect 36645 18173 36679 18207
rect 40141 18173 40175 18207
rect 16221 18105 16255 18139
rect 29653 18105 29687 18139
rect 30573 18105 30607 18139
rect 36921 18105 36955 18139
rect 40417 18105 40451 18139
rect 2513 18037 2547 18071
rect 4721 18037 4755 18071
rect 8769 18037 8803 18071
rect 14105 18037 14139 18071
rect 15761 18037 15795 18071
rect 16313 18037 16347 18071
rect 16681 18037 16715 18071
rect 18153 18037 18187 18071
rect 18981 18037 19015 18071
rect 30205 18037 30239 18071
rect 36553 18037 36587 18071
rect 37657 18037 37691 18071
rect 38117 18037 38151 18071
rect 39773 18037 39807 18071
rect 40049 18037 40083 18071
rect 13737 17833 13771 17867
rect 15656 17833 15690 17867
rect 19625 17833 19659 17867
rect 21281 17833 21315 17867
rect 24409 17833 24443 17867
rect 27813 17833 27847 17867
rect 28089 17833 28123 17867
rect 28457 17833 28491 17867
rect 35265 17833 35299 17867
rect 37473 17833 37507 17867
rect 37933 17833 37967 17867
rect 38853 17833 38887 17867
rect 39313 17833 39347 17867
rect 39681 17833 39715 17867
rect 3157 17765 3191 17799
rect 11713 17765 11747 17799
rect 13369 17765 13403 17799
rect 19533 17765 19567 17799
rect 31585 17765 31619 17799
rect 34345 17765 34379 17799
rect 39129 17765 39163 17799
rect 1409 17697 1443 17731
rect 4261 17697 4295 17731
rect 6009 17697 6043 17731
rect 9965 17697 9999 17731
rect 12449 17697 12483 17731
rect 12633 17697 12667 17731
rect 13277 17697 13311 17731
rect 13829 17697 13863 17731
rect 15393 17697 15427 17731
rect 18337 17697 18371 17731
rect 19625 17697 19659 17731
rect 25053 17697 25087 17731
rect 27721 17697 27755 17731
rect 29561 17697 29595 17731
rect 37565 17697 37599 17731
rect 38761 17697 38795 17731
rect 7941 17629 7975 17663
rect 8769 17629 8803 17663
rect 12265 17629 12299 17663
rect 13553 17629 13587 17663
rect 14289 17629 14323 17663
rect 17417 17629 17451 17663
rect 17785 17629 17819 17663
rect 18061 17629 18095 17663
rect 18429 17629 18463 17663
rect 18521 17629 18555 17663
rect 18613 17629 18647 17663
rect 19349 17629 19383 17663
rect 19809 17629 19843 17663
rect 20085 17629 20119 17663
rect 21097 17629 21131 17663
rect 21281 17629 21315 17663
rect 24593 17629 24627 17663
rect 24685 17629 24719 17663
rect 24915 17629 24949 17663
rect 27813 17629 27847 17663
rect 28273 17629 28307 17663
rect 28549 17629 28583 17663
rect 28733 17629 28767 17663
rect 30113 17629 30147 17663
rect 30389 17629 30423 17663
rect 30573 17629 30607 17663
rect 31401 17629 31435 17663
rect 33701 17629 33735 17663
rect 33794 17629 33828 17663
rect 34066 17629 34100 17663
rect 34166 17629 34200 17663
rect 35449 17629 35483 17663
rect 35541 17629 35575 17663
rect 35817 17629 35851 17663
rect 35909 17629 35943 17663
rect 37749 17629 37783 17663
rect 38945 17629 38979 17663
rect 39313 17629 39347 17663
rect 39497 17629 39531 17663
rect 1685 17561 1719 17595
rect 4537 17561 4571 17595
rect 10241 17561 10275 17595
rect 12173 17561 12207 17595
rect 17601 17561 17635 17595
rect 19257 17561 19291 17595
rect 24777 17561 24811 17595
rect 27537 17561 27571 17595
rect 29101 17561 29135 17595
rect 33977 17561 34011 17595
rect 35633 17561 35667 17595
rect 37473 17561 37507 17595
rect 38669 17561 38703 17595
rect 8493 17493 8527 17527
rect 8585 17493 8619 17527
rect 11805 17493 11839 17527
rect 14105 17493 14139 17527
rect 17969 17493 18003 17527
rect 18153 17493 18187 17527
rect 21465 17493 21499 17527
rect 27997 17493 28031 17527
rect 1869 17289 1903 17323
rect 7481 17289 7515 17323
rect 9781 17289 9815 17323
rect 10517 17289 10551 17323
rect 11529 17289 11563 17323
rect 11989 17289 12023 17323
rect 14933 17289 14967 17323
rect 16313 17289 16347 17323
rect 17049 17289 17083 17323
rect 21649 17289 21683 17323
rect 23673 17289 23707 17323
rect 26709 17289 26743 17323
rect 27169 17289 27203 17323
rect 27997 17289 28031 17323
rect 30021 17289 30055 17323
rect 40049 17289 40083 17323
rect 3249 17221 3283 17255
rect 8309 17221 8343 17255
rect 13461 17221 13495 17255
rect 15853 17221 15887 17255
rect 19625 17221 19659 17255
rect 20637 17221 20671 17255
rect 23121 17221 23155 17255
rect 24041 17221 24075 17255
rect 34253 17221 34287 17255
rect 39589 17221 39623 17255
rect 2053 17153 2087 17187
rect 2421 17153 2455 17187
rect 3157 17153 3191 17187
rect 4261 17153 4295 17187
rect 6929 17153 6963 17187
rect 8033 17153 8067 17187
rect 10701 17153 10735 17187
rect 11161 17153 11195 17187
rect 11897 17153 11931 17187
rect 13001 17153 13035 17187
rect 16129 17153 16163 17187
rect 17601 17153 17635 17187
rect 20085 17153 20119 17187
rect 20269 17153 20303 17187
rect 21281 17153 21315 17187
rect 21833 17153 21867 17187
rect 22109 17153 22143 17187
rect 22753 17153 22787 17187
rect 23029 17153 23063 17187
rect 23305 17153 23339 17187
rect 23790 17153 23824 17187
rect 24317 17153 24351 17187
rect 24409 17153 24443 17187
rect 24501 17153 24535 17187
rect 24685 17153 24719 17187
rect 26433 17153 26467 17187
rect 26525 17153 26559 17187
rect 26985 17153 27019 17187
rect 27353 17153 27387 17187
rect 27629 17153 27663 17187
rect 28273 17153 28307 17187
rect 28641 17153 28675 17187
rect 28825 17153 28859 17187
rect 29101 17153 29135 17187
rect 29377 17153 29411 17187
rect 29929 17153 29963 17187
rect 33517 17153 33551 17187
rect 33977 17153 34011 17187
rect 34161 17153 34195 17187
rect 34345 17153 34379 17187
rect 39865 17153 39899 17187
rect 40141 17153 40175 17187
rect 40325 17153 40359 17187
rect 40509 17153 40543 17187
rect 3341 17085 3375 17119
rect 3709 17085 3743 17119
rect 7573 17085 7607 17119
rect 7757 17085 7791 17119
rect 12081 17085 12115 17119
rect 12357 17085 12391 17119
rect 13185 17085 13219 17119
rect 15945 17085 15979 17119
rect 17141 17085 17175 17119
rect 17233 17085 17267 17119
rect 17877 17085 17911 17119
rect 21373 17085 21407 17119
rect 21925 17085 21959 17119
rect 23581 17085 23615 17119
rect 27721 17085 27755 17119
rect 28549 17085 28583 17119
rect 33425 17085 33459 17119
rect 33793 17085 33827 17119
rect 33885 17085 33919 17119
rect 39773 17085 39807 17119
rect 2789 17017 2823 17051
rect 7113 17017 7147 17051
rect 20453 17017 20487 17051
rect 22293 17017 22327 17051
rect 22937 17017 22971 17051
rect 28089 17017 28123 17051
rect 28457 17017 28491 17051
rect 28917 17017 28951 17051
rect 29009 17017 29043 17051
rect 2237 16949 2271 16983
rect 6745 16949 6779 16983
rect 10977 16949 11011 16983
rect 15853 16949 15887 16983
rect 16681 16949 16715 16983
rect 20085 16949 20119 16983
rect 20729 16949 20763 16983
rect 21465 16949 21499 16983
rect 22017 16949 22051 16983
rect 22569 16949 22603 16983
rect 22845 16949 22879 16983
rect 23949 16949 23983 16983
rect 27537 16949 27571 16983
rect 27629 16949 27663 16983
rect 29469 16949 29503 16983
rect 33241 16949 33275 16983
rect 34529 16949 34563 16983
rect 39681 16949 39715 16983
rect 8033 16745 8067 16779
rect 12173 16745 12207 16779
rect 22017 16745 22051 16779
rect 23673 16745 23707 16779
rect 25697 16745 25731 16779
rect 26433 16745 26467 16779
rect 28733 16745 28767 16779
rect 32045 16745 32079 16779
rect 34345 16745 34379 16779
rect 34529 16745 34563 16779
rect 34897 16745 34931 16779
rect 37473 16745 37507 16779
rect 37657 16745 37691 16779
rect 39865 16745 39899 16779
rect 40325 16745 40359 16779
rect 21189 16677 21223 16711
rect 1777 16609 1811 16643
rect 2053 16609 2087 16643
rect 3525 16609 3559 16643
rect 4813 16609 4847 16643
rect 4905 16609 4939 16643
rect 5273 16609 5307 16643
rect 6285 16609 6319 16643
rect 6561 16609 6595 16643
rect 9597 16609 9631 16643
rect 10425 16609 10459 16643
rect 10701 16609 10735 16643
rect 14105 16609 14139 16643
rect 20177 16609 20211 16643
rect 21649 16609 21683 16643
rect 21925 16609 21959 16643
rect 28365 16609 28399 16643
rect 28825 16609 28859 16643
rect 30665 16609 30699 16643
rect 32689 16609 32723 16643
rect 33425 16609 33459 16643
rect 35541 16609 35575 16643
rect 40049 16609 40083 16643
rect 6101 16541 6135 16575
rect 13921 16541 13955 16575
rect 19901 16541 19935 16575
rect 19993 16541 20027 16575
rect 21373 16541 21407 16575
rect 21557 16541 21591 16575
rect 22017 16541 22051 16575
rect 23305 16541 23339 16575
rect 23489 16541 23523 16575
rect 25053 16541 25087 16575
rect 25201 16541 25235 16575
rect 25518 16541 25552 16575
rect 25789 16541 25823 16575
rect 25882 16541 25916 16575
rect 26157 16541 26191 16575
rect 26254 16541 26288 16575
rect 28549 16541 28583 16575
rect 30297 16541 30331 16575
rect 31309 16541 31343 16575
rect 31611 16541 31645 16575
rect 31769 16541 31803 16575
rect 32229 16541 32263 16575
rect 32413 16541 32447 16575
rect 33609 16541 33643 16575
rect 33885 16541 33919 16575
rect 35081 16541 35115 16575
rect 37289 16541 37323 16575
rect 37473 16541 37507 16575
rect 40141 16541 40175 16575
rect 4721 16473 4755 16507
rect 5825 16473 5859 16507
rect 9413 16473 9447 16507
rect 14381 16473 14415 16507
rect 21741 16473 21775 16507
rect 25329 16473 25363 16507
rect 25421 16473 25455 16507
rect 26065 16473 26099 16507
rect 30481 16473 30515 16507
rect 31401 16473 31435 16507
rect 31493 16473 31527 16507
rect 32321 16473 32355 16507
rect 32551 16473 32585 16507
rect 34161 16473 34195 16507
rect 34377 16473 34411 16507
rect 35173 16473 35207 16507
rect 35265 16473 35299 16507
rect 35383 16473 35417 16507
rect 39865 16473 39899 16507
rect 4353 16405 4387 16439
rect 5917 16405 5951 16439
rect 8953 16405 8987 16439
rect 9321 16405 9355 16439
rect 13737 16405 13771 16439
rect 15853 16405 15887 16439
rect 22201 16405 22235 16439
rect 31125 16405 31159 16439
rect 33793 16405 33827 16439
rect 5273 16201 5307 16235
rect 5457 16201 5491 16235
rect 10517 16201 10551 16235
rect 14105 16201 14139 16235
rect 14473 16201 14507 16235
rect 18067 16201 18101 16235
rect 18153 16201 18187 16235
rect 25513 16201 25547 16235
rect 35173 16201 35207 16235
rect 23581 16133 23615 16167
rect 26157 16133 26191 16167
rect 31217 16133 31251 16167
rect 35541 16133 35575 16167
rect 35659 16133 35693 16167
rect 39221 16133 39255 16167
rect 3525 16065 3559 16099
rect 5825 16065 5859 16099
rect 7021 16065 7055 16099
rect 8033 16065 8067 16099
rect 9965 16065 9999 16099
rect 12541 16065 12575 16099
rect 12633 16065 12667 16099
rect 13185 16065 13219 16099
rect 13277 16065 13311 16099
rect 13369 16065 13403 16099
rect 13553 16065 13587 16099
rect 16037 16065 16071 16099
rect 17049 16065 17083 16099
rect 17969 16065 18003 16099
rect 18245 16065 18279 16099
rect 18889 16065 18923 16099
rect 19165 16065 19199 16099
rect 25789 16065 25823 16099
rect 31401 16065 31435 16099
rect 35357 16065 35391 16099
rect 35449 16065 35483 16099
rect 37289 16065 37323 16099
rect 37565 16065 37599 16099
rect 39497 16065 39531 16099
rect 3801 15997 3835 16031
rect 5917 15997 5951 16031
rect 6101 15997 6135 16031
rect 6377 15997 6411 16031
rect 8309 15997 8343 16031
rect 12817 15997 12851 16031
rect 14565 15997 14599 16031
rect 14749 15997 14783 16031
rect 16865 15997 16899 16031
rect 18521 15997 18555 16031
rect 23949 15997 23983 16031
rect 24041 15997 24075 16031
rect 25697 15997 25731 16031
rect 26065 15997 26099 16031
rect 31585 15997 31619 16031
rect 35817 15997 35851 16031
rect 37381 15997 37415 16031
rect 39313 15997 39347 16031
rect 9781 15929 9815 15963
rect 19165 15929 19199 15963
rect 37749 15929 37783 15963
rect 12725 15861 12759 15895
rect 12909 15861 12943 15895
rect 16221 15861 16255 15895
rect 17233 15861 17267 15895
rect 24225 15861 24259 15895
rect 37565 15861 37599 15895
rect 39221 15861 39255 15895
rect 39681 15861 39715 15895
rect 3985 15657 4019 15691
rect 4892 15657 4926 15691
rect 6377 15657 6411 15691
rect 8493 15657 8527 15691
rect 25605 15657 25639 15691
rect 26893 15657 26927 15691
rect 30297 15657 30331 15691
rect 32873 15657 32907 15691
rect 35449 15657 35483 15691
rect 37933 15657 37967 15691
rect 39865 15657 39899 15691
rect 40325 15657 40359 15691
rect 2697 15589 2731 15623
rect 17693 15589 17727 15623
rect 30205 15589 30239 15623
rect 30389 15589 30423 15623
rect 3341 15521 3375 15555
rect 4629 15521 4663 15555
rect 11437 15521 11471 15555
rect 26157 15521 26191 15555
rect 26985 15521 27019 15555
rect 36093 15521 36127 15555
rect 39957 15521 39991 15555
rect 2237 15453 2271 15487
rect 3065 15453 3099 15487
rect 4169 15453 4203 15487
rect 7849 15453 7883 15487
rect 8033 15453 8067 15487
rect 8125 15453 8159 15487
rect 8309 15453 8343 15487
rect 8677 15453 8711 15487
rect 13369 15453 13403 15487
rect 13461 15453 13495 15487
rect 13645 15453 13679 15487
rect 13737 15453 13771 15487
rect 17049 15453 17083 15487
rect 17325 15453 17359 15487
rect 18153 15453 18187 15487
rect 18455 15453 18489 15487
rect 18613 15453 18647 15487
rect 21281 15453 21315 15487
rect 21465 15453 21499 15487
rect 21833 15453 21867 15487
rect 21925 15453 21959 15487
rect 22017 15453 22051 15487
rect 22201 15453 22235 15487
rect 23857 15453 23891 15487
rect 23949 15453 23983 15487
rect 24133 15453 24167 15487
rect 24225 15453 24259 15487
rect 25513 15453 25547 15487
rect 25881 15453 25915 15487
rect 26065 15453 26099 15487
rect 26341 15453 26375 15487
rect 26525 15453 26559 15487
rect 26709 15453 26743 15487
rect 26801 15453 26835 15487
rect 30113 15453 30147 15487
rect 30573 15453 30607 15487
rect 32597 15453 32631 15487
rect 32689 15453 32723 15487
rect 35633 15453 35667 15487
rect 37289 15453 37323 15487
rect 37437 15453 37471 15487
rect 37657 15453 37691 15487
rect 37795 15453 37829 15487
rect 39865 15453 39899 15487
rect 40141 15453 40175 15487
rect 1501 15385 1535 15419
rect 11161 15385 11195 15419
rect 17509 15385 17543 15419
rect 18245 15385 18279 15419
rect 18337 15385 18371 15419
rect 29837 15385 29871 15419
rect 35725 15385 35759 15419
rect 35817 15385 35851 15419
rect 35955 15385 35989 15419
rect 37565 15385 37599 15419
rect 1593 15317 1627 15351
rect 2053 15317 2087 15351
rect 3157 15317 3191 15351
rect 8033 15317 8067 15351
rect 8309 15317 8343 15351
rect 10793 15317 10827 15351
rect 11253 15317 11287 15351
rect 13185 15317 13219 15351
rect 16865 15317 16899 15351
rect 17233 15317 17267 15351
rect 17969 15317 18003 15351
rect 21373 15317 21407 15351
rect 21557 15317 21591 15351
rect 23673 15317 23707 15351
rect 3341 15113 3375 15147
rect 8125 15113 8159 15147
rect 10149 15113 10183 15147
rect 10977 15113 11011 15147
rect 12081 15113 12115 15147
rect 12541 15113 12575 15147
rect 12909 15113 12943 15147
rect 15301 15113 15335 15147
rect 21189 15113 21223 15147
rect 22661 15113 22695 15147
rect 23857 15113 23891 15147
rect 26985 15113 27019 15147
rect 28457 15113 28491 15147
rect 34069 15113 34103 15147
rect 38853 15113 38887 15147
rect 1869 15045 1903 15079
rect 10241 15045 10275 15079
rect 12173 15045 12207 15079
rect 14657 15045 14691 15079
rect 14749 15045 14783 15079
rect 16129 15045 16163 15079
rect 16957 15045 16991 15079
rect 19718 15045 19752 15079
rect 19855 15045 19889 15079
rect 28273 15045 28307 15079
rect 33793 15045 33827 15079
rect 34437 15045 34471 15079
rect 38485 15045 38519 15079
rect 38577 15045 38611 15079
rect 8217 14977 8251 15011
rect 8401 14977 8435 15011
rect 8493 14977 8527 15011
rect 8677 14977 8711 15011
rect 11069 14977 11103 15011
rect 16681 14977 16715 15011
rect 19533 14977 19567 15011
rect 19626 14977 19660 15011
rect 19993 14977 20027 15011
rect 21097 14977 21131 15011
rect 21281 14977 21315 15011
rect 21649 14977 21683 15011
rect 22017 14977 22051 15011
rect 22385 14977 22419 15011
rect 22845 14977 22879 15011
rect 23765 14977 23799 15011
rect 24041 14977 24075 15011
rect 24225 14977 24259 15011
rect 24501 14977 24535 15011
rect 27169 14977 27203 15011
rect 27445 14977 27479 15011
rect 27629 14977 27663 15011
rect 27905 14977 27939 15011
rect 29009 14977 29043 15011
rect 29561 14977 29595 15011
rect 29745 14977 29779 15011
rect 32321 14977 32355 15011
rect 32413 14977 32447 15011
rect 32505 14977 32539 15011
rect 32623 14977 32657 15011
rect 33425 14977 33459 15011
rect 33518 14977 33552 15011
rect 33701 14977 33735 15011
rect 33890 14977 33924 15011
rect 34161 14977 34195 15011
rect 34345 14977 34379 15011
rect 34529 14977 34563 15011
rect 38209 14977 38243 15011
rect 38302 14977 38336 15011
rect 38715 14977 38749 15011
rect 1593 14909 1627 14943
rect 6377 14909 6411 14943
rect 6653 14909 6687 14943
rect 10425 14909 10459 14943
rect 11161 14909 11195 14943
rect 12357 14909 12391 14943
rect 13001 14909 13035 14943
rect 13185 14909 13219 14943
rect 14179 14909 14213 14943
rect 14657 14909 14691 14943
rect 15393 14909 15427 14943
rect 15577 14909 15611 14943
rect 16405 14909 16439 14943
rect 21925 14909 21959 14943
rect 24593 14909 24627 14943
rect 28825 14909 28859 14943
rect 29285 14909 29319 14943
rect 29837 14909 29871 14943
rect 32781 14909 32815 14943
rect 8309 14841 8343 14875
rect 14933 14841 14967 14875
rect 18429 14841 18463 14875
rect 21465 14841 21499 14875
rect 23489 14841 23523 14875
rect 24409 14841 24443 14875
rect 27261 14841 27295 14875
rect 27353 14841 27387 14875
rect 29193 14841 29227 14875
rect 8585 14773 8619 14807
rect 9781 14773 9815 14807
rect 10609 14773 10643 14807
rect 11713 14773 11747 14807
rect 19349 14773 19383 14807
rect 22293 14773 22327 14807
rect 22569 14773 22603 14807
rect 23305 14773 23339 14807
rect 23581 14773 23615 14807
rect 23673 14773 23707 14807
rect 24133 14773 24167 14807
rect 28273 14773 28307 14807
rect 29377 14773 29411 14807
rect 32137 14773 32171 14807
rect 34713 14773 34747 14807
rect 14841 14569 14875 14603
rect 17785 14569 17819 14603
rect 18521 14569 18555 14603
rect 19625 14569 19659 14603
rect 25329 14569 25363 14603
rect 25789 14569 25823 14603
rect 26709 14569 26743 14603
rect 26985 14569 27019 14603
rect 27445 14569 27479 14603
rect 27629 14569 27663 14603
rect 33425 14569 33459 14603
rect 36645 14569 36679 14603
rect 38669 14569 38703 14603
rect 39037 14569 39071 14603
rect 39865 14569 39899 14603
rect 40325 14569 40359 14603
rect 14197 14501 14231 14535
rect 19257 14501 19291 14535
rect 19901 14501 19935 14535
rect 20453 14501 20487 14535
rect 21741 14501 21775 14535
rect 24409 14501 24443 14535
rect 26249 14501 26283 14535
rect 26617 14501 26651 14535
rect 31953 14501 31987 14535
rect 3341 14433 3375 14467
rect 3525 14433 3559 14467
rect 7113 14433 7147 14467
rect 10977 14433 11011 14467
rect 18981 14433 19015 14467
rect 26433 14433 26467 14467
rect 26801 14433 26835 14467
rect 27169 14433 27203 14467
rect 28825 14433 28859 14467
rect 34069 14433 34103 14467
rect 38761 14433 38795 14467
rect 39957 14433 39991 14467
rect 3801 14365 3835 14399
rect 10701 14365 10735 14399
rect 11805 14365 11839 14399
rect 11989 14365 12023 14399
rect 14473 14365 14507 14399
rect 14565 14365 14599 14399
rect 15301 14365 15335 14399
rect 15393 14365 15427 14399
rect 17325 14365 17359 14399
rect 17509 14365 17543 14399
rect 18337 14365 18371 14399
rect 18797 14365 18831 14399
rect 19073 14365 19107 14399
rect 20054 14365 20088 14399
rect 20545 14365 20579 14399
rect 21741 14365 21775 14399
rect 21833 14365 21867 14399
rect 23213 14365 23247 14399
rect 24685 14365 24719 14399
rect 25513 14365 25547 14399
rect 25605 14365 25639 14399
rect 25973 14365 26007 14399
rect 26525 14365 26559 14399
rect 26893 14365 26927 14399
rect 29009 14365 29043 14399
rect 30665 14365 30699 14399
rect 30849 14365 30883 14399
rect 30941 14365 30975 14399
rect 31033 14365 31067 14399
rect 31309 14365 31343 14399
rect 31457 14365 31491 14399
rect 31585 14365 31619 14399
rect 31677 14365 31711 14399
rect 31815 14365 31849 14399
rect 33609 14365 33643 14399
rect 33931 14365 33965 14399
rect 34897 14365 34931 14399
rect 35357 14365 35391 14399
rect 36829 14365 36863 14399
rect 36921 14365 36955 14399
rect 37105 14365 37139 14399
rect 37197 14365 37231 14399
rect 38577 14365 38611 14399
rect 38853 14365 38887 14399
rect 40141 14365 40175 14399
rect 3249 14297 3283 14331
rect 4445 14297 4479 14331
rect 14197 14297 14231 14331
rect 15117 14297 15151 14331
rect 17601 14297 17635 14331
rect 17817 14297 17851 14331
rect 18153 14297 18187 14331
rect 20151 14297 20185 14331
rect 22017 14297 22051 14331
rect 24409 14297 24443 14331
rect 25329 14297 25363 14331
rect 27292 14297 27326 14331
rect 29193 14297 29227 14331
rect 33701 14297 33735 14331
rect 33793 14297 33827 14331
rect 34989 14297 35023 14331
rect 35081 14297 35115 14331
rect 35199 14297 35233 14331
rect 39865 14297 39899 14331
rect 2881 14229 2915 14263
rect 7665 14229 7699 14263
rect 10333 14229 10367 14263
rect 10793 14229 10827 14263
rect 11989 14229 12023 14263
rect 14381 14229 14415 14263
rect 15025 14229 15059 14263
rect 15301 14229 15335 14263
rect 17417 14229 17451 14263
rect 17969 14229 18003 14263
rect 18613 14229 18647 14263
rect 19625 14229 19659 14263
rect 19809 14229 19843 14263
rect 23029 14229 23063 14263
rect 24593 14229 24627 14263
rect 27169 14229 27203 14263
rect 27445 14229 27479 14263
rect 31217 14229 31251 14263
rect 34713 14229 34747 14263
rect 6929 14025 6963 14059
rect 9505 14025 9539 14059
rect 12265 14025 12299 14059
rect 20453 14025 20487 14059
rect 25789 14025 25823 14059
rect 27721 14025 27755 14059
rect 28365 14025 28399 14059
rect 28641 14025 28675 14059
rect 29561 14025 29595 14059
rect 29929 14025 29963 14059
rect 31585 14025 31619 14059
rect 32597 14025 32631 14059
rect 37841 14025 37875 14059
rect 6653 13957 6687 13991
rect 8033 13957 8067 13991
rect 8861 13957 8895 13991
rect 10057 13957 10091 13991
rect 17417 13957 17451 13991
rect 26801 13957 26835 13991
rect 27997 13957 28031 13991
rect 31217 13957 31251 13991
rect 31309 13957 31343 13991
rect 32137 13957 32171 13991
rect 34253 13957 34287 13991
rect 37565 13957 37599 13991
rect 1501 13889 1535 13923
rect 3433 13889 3467 13923
rect 5365 13889 5399 13923
rect 6377 13889 6411 13923
rect 6561 13889 6595 13923
rect 6745 13889 6779 13923
rect 7757 13889 7791 13923
rect 7941 13889 7975 13923
rect 8217 13889 8251 13923
rect 8677 13889 8711 13923
rect 9321 13889 9355 13923
rect 9413 13889 9447 13923
rect 9873 13889 9907 13923
rect 12817 13889 12851 13923
rect 13001 13889 13035 13923
rect 16681 13889 16715 13923
rect 17693 13889 17727 13923
rect 18245 13889 18279 13923
rect 18429 13889 18463 13923
rect 18521 13889 18555 13923
rect 18889 13889 18923 13923
rect 19441 13889 19475 13923
rect 19809 13889 19843 13923
rect 20637 13889 20671 13923
rect 20821 13889 20855 13923
rect 25697 13889 25731 13923
rect 25881 13889 25915 13923
rect 26433 13889 26467 13923
rect 26985 13889 27019 13923
rect 27169 13889 27203 13923
rect 27270 13889 27304 13923
rect 27537 13889 27571 13923
rect 27813 13889 27847 13923
rect 28081 13889 28115 13923
rect 28181 13889 28215 13923
rect 28825 13889 28859 13923
rect 29009 13889 29043 13923
rect 29101 13889 29135 13923
rect 31033 13889 31067 13923
rect 31401 13889 31435 13923
rect 32413 13889 32447 13923
rect 34437 13889 34471 13923
rect 34529 13889 34563 13923
rect 35817 13889 35851 13923
rect 35909 13889 35943 13923
rect 36001 13889 36035 13923
rect 36119 13889 36153 13923
rect 36277 13889 36311 13923
rect 37289 13889 37323 13923
rect 37473 13889 37507 13923
rect 37657 13889 37691 13923
rect 1777 13821 1811 13855
rect 3249 13821 3283 13855
rect 3709 13821 3743 13855
rect 5181 13821 5215 13855
rect 8493 13821 8527 13855
rect 9689 13821 9723 13855
rect 12725 13821 12759 13855
rect 17877 13821 17911 13855
rect 18337 13821 18371 13855
rect 19533 13821 19567 13855
rect 26341 13821 26375 13855
rect 27353 13821 27387 13855
rect 30021 13821 30055 13855
rect 30205 13821 30239 13855
rect 32229 13821 32263 13855
rect 7757 13753 7791 13787
rect 12541 13753 12575 13787
rect 26433 13753 26467 13787
rect 34713 13753 34747 13787
rect 6009 13685 6043 13719
rect 8309 13685 8343 13719
rect 12633 13685 12667 13719
rect 18889 13685 18923 13719
rect 19073 13685 19107 13719
rect 32137 13685 32171 13719
rect 34529 13685 34563 13719
rect 35633 13685 35667 13719
rect 2237 13481 2271 13515
rect 4721 13481 4755 13515
rect 5549 13481 5583 13515
rect 7389 13481 7423 13515
rect 14841 13481 14875 13515
rect 15669 13481 15703 13515
rect 16405 13481 16439 13515
rect 29745 13481 29779 13515
rect 35817 13481 35851 13515
rect 37841 13481 37875 13515
rect 39865 13481 39899 13515
rect 40233 13481 40267 13515
rect 9689 13413 9723 13447
rect 11253 13413 11287 13447
rect 12449 13413 12483 13447
rect 12817 13413 12851 13447
rect 16589 13413 16623 13447
rect 26893 13413 26927 13447
rect 9321 13345 9355 13379
rect 10609 13345 10643 13379
rect 13093 13345 13127 13379
rect 17969 13345 18003 13379
rect 18061 13345 18095 13379
rect 27077 13345 27111 13379
rect 27261 13345 27295 13379
rect 30481 13345 30515 13379
rect 36185 13345 36219 13379
rect 36277 13345 36311 13379
rect 39957 13345 39991 13379
rect 2421 13277 2455 13311
rect 4905 13277 4939 13311
rect 4997 13277 5031 13311
rect 5181 13277 5215 13311
rect 5273 13277 5307 13311
rect 5457 13277 5491 13311
rect 5641 13277 5675 13311
rect 6561 13277 6595 13311
rect 6745 13277 6779 13311
rect 7113 13277 7147 13311
rect 7665 13277 7699 13311
rect 7941 13277 7975 13311
rect 8217 13277 8251 13311
rect 8585 13277 8619 13311
rect 8953 13277 8987 13311
rect 9137 13277 9171 13311
rect 9229 13277 9263 13311
rect 9516 13277 9550 13311
rect 10425 13277 10459 13311
rect 11069 13277 11103 13311
rect 11345 13277 11379 13311
rect 11805 13277 11839 13311
rect 11989 13277 12023 13311
rect 12265 13277 12299 13311
rect 12357 13277 12391 13311
rect 12541 13277 12575 13311
rect 12717 13287 12751 13321
rect 13001 13277 13035 13311
rect 13185 13277 13219 13311
rect 14749 13277 14783 13311
rect 15301 13277 15335 13311
rect 15485 13277 15519 13311
rect 15669 13277 15703 13311
rect 15853 13277 15887 13311
rect 16129 13277 16163 13311
rect 16221 13277 16255 13311
rect 16773 13277 16807 13311
rect 17233 13277 17267 13311
rect 17509 13277 17543 13311
rect 21005 13277 21039 13311
rect 21465 13277 21499 13311
rect 21725 13277 21759 13311
rect 21833 13277 21867 13311
rect 22661 13277 22695 13311
rect 22937 13277 22971 13311
rect 26801 13277 26835 13311
rect 27169 13277 27203 13311
rect 27353 13277 27387 13311
rect 29653 13277 29687 13311
rect 30389 13277 30423 13311
rect 33977 13277 34011 13311
rect 34253 13277 34287 13311
rect 34345 13277 34379 13311
rect 36001 13277 36035 13311
rect 36093 13277 36127 13311
rect 37289 13277 37323 13311
rect 37565 13277 37599 13311
rect 37657 13277 37691 13311
rect 38761 13277 38795 13311
rect 39037 13277 39071 13311
rect 39129 13277 39163 13311
rect 39865 13277 39899 13311
rect 7389 13209 7423 13243
rect 7573 13209 7607 13243
rect 8401 13209 8435 13243
rect 8493 13209 8527 13243
rect 20821 13209 20855 13243
rect 21373 13209 21407 13243
rect 22201 13209 22235 13243
rect 27077 13209 27111 13243
rect 32321 13209 32355 13243
rect 34161 13209 34195 13243
rect 36553 13209 36587 13243
rect 37473 13209 37507 13243
rect 38945 13209 38979 13243
rect 6745 13141 6779 13175
rect 7205 13141 7239 13175
rect 8033 13141 8067 13175
rect 8769 13141 8803 13175
rect 10057 13141 10091 13175
rect 10517 13141 10551 13175
rect 10885 13141 10919 13175
rect 11897 13141 11931 13175
rect 12081 13141 12115 13175
rect 15209 13141 15243 13175
rect 15393 13141 15427 13175
rect 17693 13141 17727 13175
rect 21097 13141 21131 13175
rect 21189 13141 21223 13175
rect 22753 13141 22787 13175
rect 32413 13141 32447 13175
rect 34529 13141 34563 13175
rect 36645 13141 36679 13175
rect 39313 13141 39347 13175
rect 6561 12937 6595 12971
rect 7757 12937 7791 12971
rect 8769 12937 8803 12971
rect 10241 12937 10275 12971
rect 10425 12937 10459 12971
rect 10609 12937 10643 12971
rect 11069 12937 11103 12971
rect 12357 12937 12391 12971
rect 16957 12937 16991 12971
rect 17785 12937 17819 12971
rect 22293 12937 22327 12971
rect 24317 12937 24351 12971
rect 26433 12937 26467 12971
rect 29653 12937 29687 12971
rect 29837 12937 29871 12971
rect 32413 12937 32447 12971
rect 32781 12937 32815 12971
rect 34897 12937 34931 12971
rect 36737 12937 36771 12971
rect 39405 12937 39439 12971
rect 15301 12869 15335 12903
rect 15853 12869 15887 12903
rect 22385 12869 22419 12903
rect 23949 12869 23983 12903
rect 24149 12869 24183 12903
rect 24593 12869 24627 12903
rect 24685 12869 24719 12903
rect 25881 12869 25915 12903
rect 28917 12869 28951 12903
rect 29285 12869 29319 12903
rect 32229 12869 32263 12903
rect 39037 12869 39071 12903
rect 39129 12869 39163 12903
rect 6377 12801 6411 12835
rect 6653 12801 6687 12835
rect 6745 12801 6779 12835
rect 6929 12801 6963 12835
rect 7297 12801 7331 12835
rect 7573 12801 7607 12835
rect 7849 12801 7883 12835
rect 8401 12801 8435 12835
rect 8593 12801 8627 12835
rect 8861 12801 8895 12835
rect 9045 12801 9079 12835
rect 9873 12801 9907 12835
rect 10057 12801 10091 12835
rect 10333 12801 10367 12835
rect 10977 12801 11011 12835
rect 11805 12801 11839 12835
rect 12265 12801 12299 12835
rect 12541 12801 12575 12835
rect 12633 12801 12667 12835
rect 14289 12801 14323 12835
rect 15117 12801 15151 12835
rect 15393 12801 15427 12835
rect 15669 12801 15703 12835
rect 15761 12801 15795 12835
rect 15971 12801 16005 12835
rect 16129 12801 16163 12835
rect 16773 12801 16807 12835
rect 17417 12801 17451 12835
rect 17601 12801 17635 12835
rect 17877 12801 17911 12835
rect 18613 12801 18647 12835
rect 18705 12801 18739 12835
rect 22109 12801 22143 12835
rect 24409 12801 24443 12835
rect 24777 12801 24811 12835
rect 26065 12801 26099 12835
rect 26341 12801 26375 12835
rect 26525 12801 26559 12835
rect 29834 12801 29868 12835
rect 32965 12801 32999 12835
rect 33057 12801 33091 12835
rect 33241 12801 33275 12835
rect 33333 12801 33367 12835
rect 33793 12801 33827 12835
rect 33941 12801 33975 12835
rect 34069 12801 34103 12835
rect 34161 12801 34195 12835
rect 34258 12801 34292 12835
rect 34713 12801 34747 12835
rect 36369 12801 36403 12835
rect 36553 12801 36587 12835
rect 38853 12801 38887 12835
rect 39221 12801 39255 12835
rect 8953 12733 8987 12767
rect 11253 12733 11287 12767
rect 11897 12733 11931 12767
rect 11989 12733 12023 12767
rect 12081 12733 12115 12767
rect 12909 12733 12943 12767
rect 13001 12733 13035 12767
rect 14381 12733 14415 12767
rect 18337 12733 18371 12767
rect 18521 12733 18555 12767
rect 18797 12733 18831 12767
rect 30205 12733 30239 12767
rect 30297 12733 30331 12767
rect 34529 12733 34563 12767
rect 7205 12665 7239 12699
rect 7389 12665 7423 12699
rect 11621 12665 11655 12699
rect 32597 12665 32631 12699
rect 34437 12665 34471 12699
rect 6377 12597 6411 12631
rect 10057 12597 10091 12631
rect 14657 12597 14691 12631
rect 14933 12597 14967 12631
rect 15485 12597 15519 12631
rect 21925 12597 21959 12631
rect 24133 12597 24167 12631
rect 24961 12597 24995 12631
rect 26157 12597 26191 12631
rect 32413 12597 32447 12631
rect 36369 12597 36403 12631
rect 4353 12393 4387 12427
rect 5273 12393 5307 12427
rect 7113 12393 7147 12427
rect 10425 12393 10459 12427
rect 14933 12393 14967 12427
rect 18981 12393 19015 12427
rect 19441 12393 19475 12427
rect 19625 12393 19659 12427
rect 23489 12393 23523 12427
rect 24961 12393 24995 12427
rect 25881 12393 25915 12427
rect 26065 12393 26099 12427
rect 26157 12393 26191 12427
rect 26617 12393 26651 12427
rect 26709 12393 26743 12427
rect 32229 12393 32263 12427
rect 33425 12393 33459 12427
rect 33609 12393 33643 12427
rect 34253 12393 34287 12427
rect 5641 12325 5675 12359
rect 14381 12325 14415 12359
rect 15025 12325 15059 12359
rect 23305 12325 23339 12359
rect 31033 12325 31067 12359
rect 12173 12257 12207 12291
rect 21373 12257 21407 12291
rect 21557 12257 21591 12291
rect 21925 12257 21959 12291
rect 23765 12257 23799 12291
rect 23857 12257 23891 12291
rect 25789 12257 25823 12291
rect 30389 12257 30423 12291
rect 31309 12257 31343 12291
rect 32321 12257 32355 12291
rect 3985 12189 4019 12223
rect 4077 12189 4111 12223
rect 4445 12189 4479 12223
rect 4813 12189 4847 12223
rect 4905 12189 4939 12223
rect 4997 12189 5031 12223
rect 5089 12189 5123 12223
rect 5457 12189 5491 12223
rect 5549 12189 5583 12223
rect 5733 12189 5767 12223
rect 5917 12189 5951 12223
rect 9045 12189 9079 12223
rect 9137 12189 9171 12223
rect 9321 12189 9355 12223
rect 10609 12189 10643 12223
rect 10701 12189 10735 12223
rect 14289 12189 14323 12223
rect 14473 12189 14507 12223
rect 14841 12189 14875 12223
rect 15117 12189 15151 12223
rect 15301 12189 15335 12223
rect 17325 12189 17359 12223
rect 17509 12189 17543 12223
rect 18797 12189 18831 12223
rect 18889 12189 18923 12223
rect 19073 12189 19107 12223
rect 19717 12189 19751 12223
rect 19855 12189 19889 12223
rect 21741 12189 21775 12223
rect 23213 12189 23247 12223
rect 23397 12189 23431 12223
rect 23673 12189 23707 12223
rect 23949 12189 23983 12223
rect 24777 12189 24811 12223
rect 25605 12189 25639 12223
rect 25881 12189 25915 12223
rect 26341 12189 26375 12223
rect 26433 12189 26467 12223
rect 26893 12189 26927 12223
rect 26985 12189 27019 12223
rect 27169 12189 27203 12223
rect 27261 12189 27295 12223
rect 27537 12189 27571 12223
rect 27629 12189 27663 12223
rect 27813 12189 27847 12223
rect 27905 12189 27939 12223
rect 29561 12189 29595 12223
rect 29837 12189 29871 12223
rect 30021 12189 30055 12223
rect 30205 12189 30239 12223
rect 30481 12189 30515 12223
rect 30665 12189 30699 12223
rect 31585 12189 31619 12223
rect 32045 12189 32079 12223
rect 32137 12189 32171 12223
rect 34069 12189 34103 12223
rect 6653 12121 6687 12155
rect 6929 12121 6963 12155
rect 7145 12121 7179 12155
rect 10425 12121 10459 12155
rect 12449 12121 12483 12155
rect 14565 12121 14599 12155
rect 19257 12121 19291 12155
rect 19473 12121 19507 12155
rect 24593 12121 24627 12155
rect 26157 12121 26191 12155
rect 27353 12121 27387 12155
rect 30849 12121 30883 12155
rect 31677 12121 31711 12155
rect 31794 12121 31828 12155
rect 32781 12121 32815 12155
rect 33149 12121 33183 12155
rect 33241 12121 33275 12155
rect 33441 12121 33475 12155
rect 4169 12053 4203 12087
rect 4445 12053 4479 12087
rect 4629 12053 4663 12087
rect 7297 12053 7331 12087
rect 13921 12053 13955 12087
rect 17417 12053 17451 12087
rect 18613 12053 18647 12087
rect 20085 12053 20119 12087
rect 20913 12053 20947 12087
rect 21281 12053 21315 12087
rect 30665 12053 30699 12087
rect 31953 12053 31987 12087
rect 4077 11849 4111 11883
rect 4905 11849 4939 11883
rect 5825 11849 5859 11883
rect 8125 11849 8159 11883
rect 14565 11849 14599 11883
rect 23765 11849 23799 11883
rect 26709 11849 26743 11883
rect 27445 11849 27479 11883
rect 29653 11849 29687 11883
rect 31309 11849 31343 11883
rect 36277 11849 36311 11883
rect 40325 11849 40359 11883
rect 14197 11781 14231 11815
rect 18705 11781 18739 11815
rect 20453 11781 20487 11815
rect 24133 11781 24167 11815
rect 25973 11781 26007 11815
rect 26985 11781 27019 11815
rect 30205 11781 30239 11815
rect 30389 11781 30423 11815
rect 34989 11781 35023 11815
rect 35081 11781 35115 11815
rect 35909 11781 35943 11815
rect 36001 11781 36035 11815
rect 1409 11713 1443 11747
rect 3065 11713 3099 11747
rect 3709 11713 3743 11747
rect 4353 11713 4387 11747
rect 4721 11713 4755 11747
rect 5733 11713 5767 11747
rect 5917 11713 5951 11747
rect 6561 11713 6595 11747
rect 6745 11713 6779 11747
rect 8033 11713 8067 11747
rect 8217 11713 8251 11747
rect 10885 11713 10919 11747
rect 11069 11713 11103 11747
rect 13369 11713 13403 11747
rect 14013 11713 14047 11747
rect 14289 11713 14323 11747
rect 14381 11713 14415 11747
rect 18429 11713 18463 11747
rect 20913 11713 20947 11747
rect 23673 11713 23707 11747
rect 23857 11713 23891 11747
rect 23949 11713 23983 11747
rect 24225 11713 24259 11747
rect 25789 11713 25823 11747
rect 26157 11713 26191 11747
rect 26249 11713 26283 11747
rect 26709 11713 26743 11747
rect 27261 11713 27295 11747
rect 29009 11713 29043 11747
rect 29377 11713 29411 11747
rect 29561 11713 29595 11747
rect 30021 11713 30055 11747
rect 30481 11713 30515 11747
rect 30665 11713 30699 11747
rect 30941 11713 30975 11747
rect 34069 11713 34103 11747
rect 34805 11713 34839 11747
rect 35173 11713 35207 11747
rect 35633 11713 35667 11747
rect 35726 11713 35760 11747
rect 36098 11713 36132 11747
rect 39397 11735 39431 11769
rect 39497 11713 39531 11747
rect 39681 11713 39715 11747
rect 39773 11713 39807 11747
rect 39865 11713 39899 11747
rect 40141 11713 40175 11747
rect 1685 11645 1719 11679
rect 3157 11645 3191 11679
rect 3617 11645 3651 11679
rect 6837 11645 6871 11679
rect 13921 11645 13955 11679
rect 27077 11645 27111 11679
rect 29285 11645 29319 11679
rect 31033 11645 31067 11679
rect 39221 11645 39255 11679
rect 40049 11645 40083 11679
rect 3433 11577 3467 11611
rect 23949 11577 23983 11611
rect 26387 11577 26421 11611
rect 30757 11577 30791 11611
rect 35357 11577 35391 11611
rect 4721 11509 4755 11543
rect 6377 11509 6411 11543
rect 11253 11509 11287 11543
rect 20729 11509 20763 11543
rect 26525 11509 26559 11543
rect 27169 11509 27203 11543
rect 30941 11509 30975 11543
rect 34161 11509 34195 11543
rect 39865 11509 39899 11543
rect 6193 11305 6227 11339
rect 6377 11305 6411 11339
rect 7573 11305 7607 11339
rect 8217 11305 8251 11339
rect 15853 11305 15887 11339
rect 21373 11305 21407 11339
rect 26709 11305 26743 11339
rect 31033 11305 31067 11339
rect 38485 11305 38519 11339
rect 39313 11305 39347 11339
rect 22385 11237 22419 11271
rect 30849 11237 30883 11271
rect 32137 11237 32171 11271
rect 33793 11237 33827 11271
rect 36369 11237 36403 11271
rect 38025 11237 38059 11271
rect 5917 11169 5951 11203
rect 7849 11169 7883 11203
rect 8033 11169 8067 11203
rect 9597 11169 9631 11203
rect 10977 11169 11011 11203
rect 11713 11169 11747 11203
rect 11897 11169 11931 11203
rect 12265 11169 12299 11203
rect 15485 11169 15519 11203
rect 17509 11169 17543 11203
rect 17693 11169 17727 11203
rect 19901 11169 19935 11203
rect 21925 11169 21959 11203
rect 32965 11169 32999 11203
rect 6009 11101 6043 11135
rect 6285 11101 6319 11135
rect 6469 11101 6503 11135
rect 7757 11101 7791 11135
rect 7941 11101 7975 11135
rect 8401 11101 8435 11135
rect 8677 11101 8711 11135
rect 9505 11101 9539 11135
rect 9781 11101 9815 11135
rect 10885 11101 10919 11135
rect 12449 11101 12483 11135
rect 12909 11101 12943 11135
rect 13093 11101 13127 11135
rect 15669 11101 15703 11135
rect 16221 11101 16255 11135
rect 16405 11101 16439 11135
rect 16497 11101 16531 11135
rect 19625 11101 19659 11135
rect 22017 11101 22051 11135
rect 22661 11101 22695 11135
rect 23121 11101 23155 11135
rect 29101 11101 29135 11135
rect 31861 11101 31895 11135
rect 33149 11101 33183 11135
rect 33609 11101 33643 11135
rect 33701 11103 33735 11137
rect 35817 11101 35851 11135
rect 36093 11101 36127 11135
rect 36185 11101 36219 11135
rect 36461 11101 36495 11135
rect 36645 11101 36679 11135
rect 37473 11101 37507 11135
rect 37657 11101 37691 11135
rect 37841 11101 37875 11135
rect 38669 11101 38703 11135
rect 38762 11101 38796 11135
rect 39037 11101 39071 11135
rect 39134 11101 39168 11135
rect 5549 11033 5583 11067
rect 10793 11033 10827 11067
rect 11621 11033 11655 11067
rect 13277 11033 13311 11067
rect 16589 11033 16623 11067
rect 26617 11033 26651 11067
rect 30573 11033 30607 11067
rect 31585 11033 31619 11067
rect 31953 11033 31987 11067
rect 33241 11033 33275 11067
rect 33333 11033 33367 11067
rect 33451 11033 33485 11067
rect 36001 11033 36035 11067
rect 37749 11033 37783 11067
rect 38209 11033 38243 11067
rect 38945 11033 38979 11067
rect 8585 10965 8619 10999
rect 9965 10965 9999 10999
rect 10425 10965 10459 10999
rect 11253 10965 11287 10999
rect 12633 10965 12667 10999
rect 16313 10965 16347 10999
rect 17049 10965 17083 10999
rect 17417 10965 17451 10999
rect 29285 10965 29319 10999
rect 31769 10965 31803 10999
rect 36829 10965 36863 10999
rect 6469 10761 6503 10795
rect 7113 10761 7147 10795
rect 11897 10761 11931 10795
rect 11989 10761 12023 10795
rect 20269 10761 20303 10795
rect 30113 10761 30147 10795
rect 30573 10761 30607 10795
rect 31769 10761 31803 10795
rect 32965 10761 32999 10795
rect 33149 10761 33183 10795
rect 9689 10693 9723 10727
rect 10517 10693 10551 10727
rect 16313 10693 16347 10727
rect 17693 10693 17727 10727
rect 20177 10693 20211 10727
rect 25513 10693 25547 10727
rect 27721 10693 27755 10727
rect 32597 10693 32631 10727
rect 32797 10693 32831 10727
rect 37565 10693 37599 10727
rect 6653 10625 6687 10659
rect 6837 10625 6871 10659
rect 6929 10625 6963 10659
rect 7021 10625 7055 10659
rect 7205 10625 7239 10659
rect 7297 10625 7331 10659
rect 7941 10625 7975 10659
rect 8125 10625 8159 10659
rect 8585 10625 8619 10659
rect 8769 10625 8803 10659
rect 8953 10625 8987 10659
rect 9137 10625 9171 10659
rect 9321 10625 9355 10659
rect 9505 10625 9539 10659
rect 9965 10625 9999 10659
rect 10241 10625 10275 10659
rect 12817 10625 12851 10659
rect 13001 10625 13035 10659
rect 16129 10625 16163 10659
rect 17417 10625 17451 10659
rect 19809 10625 19843 10659
rect 26065 10625 26099 10659
rect 27445 10625 27479 10659
rect 29469 10625 29503 10659
rect 29561 10625 29595 10659
rect 29745 10625 29779 10659
rect 29837 10625 29871 10659
rect 29929 10625 29963 10659
rect 30205 10625 30239 10659
rect 30389 10625 30423 10659
rect 31677 10625 31711 10659
rect 31861 10625 31895 10659
rect 33241 10625 33275 10659
rect 33793 10625 33827 10659
rect 37289 10625 37323 10659
rect 37473 10625 37507 10659
rect 37657 10625 37691 10659
rect 8309 10557 8343 10591
rect 8861 10557 8895 10591
rect 9229 10557 9263 10591
rect 10977 10557 11011 10591
rect 12081 10557 12115 10591
rect 16405 10557 16439 10591
rect 19165 10557 19199 10591
rect 19349 10557 19383 10591
rect 19717 10557 19751 10591
rect 23305 10557 23339 10591
rect 31125 10557 31159 10591
rect 31309 10557 31343 10591
rect 33885 10557 33919 10591
rect 9781 10489 9815 10523
rect 10149 10489 10183 10523
rect 10793 10489 10827 10523
rect 8401 10421 8435 10455
rect 11529 10421 11563 10455
rect 12909 10421 12943 10455
rect 15853 10421 15887 10455
rect 19993 10421 20027 10455
rect 23857 10421 23891 10455
rect 25605 10421 25639 10455
rect 26341 10421 26375 10455
rect 32781 10421 32815 10455
rect 37841 10421 37875 10455
rect 4905 10217 4939 10251
rect 5181 10217 5215 10251
rect 5825 10217 5859 10251
rect 9781 10217 9815 10251
rect 20085 10217 20119 10251
rect 20453 10217 20487 10251
rect 21465 10217 21499 10251
rect 22385 10217 22419 10251
rect 26157 10217 26191 10251
rect 28825 10217 28859 10251
rect 38117 10217 38151 10251
rect 38577 10217 38611 10251
rect 5089 10149 5123 10183
rect 7941 10149 7975 10183
rect 16037 10149 16071 10183
rect 22109 10149 22143 10183
rect 23397 10149 23431 10183
rect 30113 10149 30147 10183
rect 5917 10081 5951 10115
rect 24409 10081 24443 10115
rect 26893 10081 26927 10115
rect 27077 10081 27111 10115
rect 31677 10081 31711 10115
rect 38209 10081 38243 10115
rect 5457 10013 5491 10047
rect 5825 10013 5859 10047
rect 7941 10013 7975 10047
rect 8125 10013 8159 10047
rect 8217 10013 8251 10047
rect 9229 10013 9263 10047
rect 9413 10013 9447 10047
rect 9689 10013 9723 10047
rect 12081 10013 12115 10047
rect 13645 10013 13679 10047
rect 13737 10013 13771 10047
rect 14105 10013 14139 10047
rect 15761 10013 15795 10047
rect 16129 10013 16163 10047
rect 16773 10013 16807 10047
rect 16957 10013 16991 10047
rect 20269 10013 20303 10047
rect 20453 10013 20487 10047
rect 20821 10013 20855 10047
rect 21557 10013 21591 10047
rect 21925 10013 21959 10047
rect 22293 10013 22327 10047
rect 22569 10013 22603 10047
rect 23397 10013 23431 10047
rect 23581 10013 23615 10047
rect 26801 10013 26835 10047
rect 28089 10013 28123 10047
rect 28249 10013 28283 10047
rect 30297 10013 30331 10047
rect 30389 10013 30423 10047
rect 31585 10013 31619 10047
rect 31769 10013 31803 10047
rect 32781 10013 32815 10047
rect 32965 10013 32999 10047
rect 33149 10013 33183 10047
rect 33517 10013 33551 10047
rect 38117 10013 38151 10047
rect 38393 10013 38427 10047
rect 4721 9945 4755 9979
rect 4926 9945 4960 9979
rect 5181 9945 5215 9979
rect 5365 9945 5399 9979
rect 14289 9945 14323 9979
rect 19809 9945 19843 9979
rect 20729 9945 20763 9979
rect 21741 9945 21775 9979
rect 21833 9945 21867 9979
rect 24685 9945 24719 9979
rect 28733 9945 28767 9979
rect 30113 9945 30147 9979
rect 32873 9945 32907 9979
rect 33333 9945 33367 9979
rect 33425 9945 33459 9979
rect 6193 9877 6227 9911
rect 9597 9877 9631 9911
rect 12173 9877 12207 9911
rect 13921 9877 13955 9911
rect 14473 9877 14507 9911
rect 17141 9877 17175 9911
rect 26433 9877 26467 9911
rect 28181 9877 28215 9911
rect 33701 9877 33735 9911
rect 7205 9673 7239 9707
rect 25973 9673 26007 9707
rect 35173 9673 35207 9707
rect 5549 9605 5583 9639
rect 5917 9605 5951 9639
rect 7481 9605 7515 9639
rect 9689 9605 9723 9639
rect 9873 9605 9907 9639
rect 11345 9605 11379 9639
rect 19349 9605 19383 9639
rect 19901 9605 19935 9639
rect 21649 9605 21683 9639
rect 22109 9605 22143 9639
rect 26249 9605 26283 9639
rect 26341 9605 26375 9639
rect 27353 9605 27387 9639
rect 28365 9605 28399 9639
rect 31401 9605 31435 9639
rect 32505 9605 32539 9639
rect 33977 9605 34011 9639
rect 35633 9605 35667 9639
rect 39037 9605 39071 9639
rect 39405 9605 39439 9639
rect 4997 9537 5031 9571
rect 5641 9537 5675 9571
rect 5825 9537 5859 9571
rect 6009 9537 6043 9571
rect 6561 9537 6595 9571
rect 6745 9537 6779 9571
rect 7389 9537 7423 9571
rect 7573 9537 7607 9571
rect 7757 9537 7791 9571
rect 7847 9559 7881 9593
rect 8861 9537 8895 9571
rect 9045 9537 9079 9571
rect 9413 9537 9447 9571
rect 11161 9537 11195 9571
rect 11529 9537 11563 9571
rect 11713 9537 11747 9571
rect 12081 9537 12115 9571
rect 12449 9537 12483 9571
rect 12633 9537 12667 9571
rect 12725 9537 12759 9571
rect 13001 9537 13035 9571
rect 13829 9537 13863 9571
rect 14381 9537 14415 9571
rect 15301 9537 15335 9571
rect 15485 9537 15519 9571
rect 16037 9537 16071 9571
rect 16129 9537 16163 9571
rect 16221 9537 16255 9571
rect 16405 9537 16439 9571
rect 16865 9537 16899 9571
rect 16957 9537 16991 9571
rect 17141 9537 17175 9571
rect 17325 9537 17359 9571
rect 19165 9537 19199 9571
rect 22017 9537 22051 9571
rect 22201 9537 22235 9571
rect 22661 9537 22695 9571
rect 26065 9537 26099 9571
rect 26433 9537 26467 9571
rect 27077 9537 27111 9571
rect 27261 9537 27295 9571
rect 27445 9537 27479 9571
rect 31309 9537 31343 9571
rect 31493 9537 31527 9571
rect 32137 9537 32171 9571
rect 32321 9537 32355 9571
rect 33609 9537 33643 9571
rect 33793 9537 33827 9571
rect 33885 9537 33919 9571
rect 34161 9537 34195 9571
rect 34437 9537 34471 9571
rect 34621 9537 34655 9571
rect 35081 9537 35115 9571
rect 35541 9537 35575 9571
rect 9137 9469 9171 9503
rect 9229 9469 9263 9503
rect 10977 9469 11011 9503
rect 11805 9469 11839 9503
rect 11897 9469 11931 9503
rect 12817 9469 12851 9503
rect 16681 9469 16715 9503
rect 17049 9469 17083 9503
rect 19625 9469 19659 9503
rect 22293 9469 22327 9503
rect 24087 9469 24121 9503
rect 24225 9469 24259 9503
rect 24501 9469 24535 9503
rect 27813 9469 27847 9503
rect 34345 9469 34379 9503
rect 35265 9469 35299 9503
rect 35449 9469 35483 9503
rect 6561 9401 6595 9435
rect 9597 9401 9631 9435
rect 10057 9401 10091 9435
rect 14565 9401 14599 9435
rect 15301 9401 15335 9435
rect 26617 9401 26651 9435
rect 33609 9401 33643 9435
rect 34253 9401 34287 9435
rect 6193 9333 6227 9367
rect 12265 9333 12299 9367
rect 13185 9333 13219 9367
rect 15761 9333 15795 9367
rect 19533 9333 19567 9367
rect 27629 9333 27663 9367
rect 35357 9333 35391 9367
rect 4432 9129 4466 9163
rect 6561 9129 6595 9163
rect 6837 9129 6871 9163
rect 7389 9129 7423 9163
rect 8033 9129 8067 9163
rect 9505 9129 9539 9163
rect 11713 9129 11747 9163
rect 20821 9129 20855 9163
rect 24869 9129 24903 9163
rect 27813 9129 27847 9163
rect 30573 9129 30607 9163
rect 30665 9129 30699 9163
rect 33517 9129 33551 9163
rect 33977 9129 34011 9163
rect 36001 9129 36035 9163
rect 37473 9129 37507 9163
rect 5917 9061 5951 9095
rect 11529 9061 11563 9095
rect 14933 9061 14967 9095
rect 21189 9061 21223 9095
rect 28089 9061 28123 9095
rect 31861 9061 31895 9095
rect 33885 9061 33919 9095
rect 9965 8993 9999 9027
rect 11253 8993 11287 9027
rect 11897 8993 11931 9027
rect 15853 8993 15887 9027
rect 17325 8993 17359 9027
rect 20913 8993 20947 9027
rect 21741 8993 21775 9027
rect 22017 8993 22051 9027
rect 23765 8993 23799 9027
rect 26065 8993 26099 9027
rect 26341 8993 26375 9027
rect 28641 8993 28675 9027
rect 30113 8993 30147 9027
rect 31493 8993 31527 9027
rect 4169 8925 4203 8959
rect 6745 8925 6779 8959
rect 7021 8925 7055 8959
rect 7297 8925 7331 8959
rect 7573 8925 7607 8959
rect 7849 8925 7883 8959
rect 8217 8925 8251 8959
rect 8953 8925 8987 8959
rect 9137 8925 9171 8959
rect 9229 8925 9263 8959
rect 9321 8925 9355 8959
rect 9781 8925 9815 8959
rect 11161 8925 11195 8959
rect 11621 8925 11655 8959
rect 11989 8925 12023 8959
rect 12081 8925 12115 8959
rect 12173 8925 12207 8959
rect 14381 8925 14415 8959
rect 14473 8925 14507 8959
rect 14565 8925 14599 8959
rect 14749 8925 14783 8959
rect 15025 8925 15059 8959
rect 15393 8925 15427 8959
rect 16129 8925 16163 8959
rect 16221 8925 16255 8959
rect 16313 8925 16347 8959
rect 19441 8925 19475 8959
rect 20821 8925 20855 8959
rect 25053 8925 25087 8959
rect 28825 8925 28859 8959
rect 29561 8925 29595 8959
rect 29653 8925 29687 8959
rect 29929 8925 29963 8959
rect 30021 8925 30055 8959
rect 30665 8925 30699 8959
rect 30849 8925 30883 8959
rect 32137 8925 32171 8959
rect 32321 8925 32355 8959
rect 33517 8925 33551 8959
rect 33609 8925 33643 8959
rect 34161 8925 34195 8959
rect 34437 8925 34471 8959
rect 35817 8925 35851 8959
rect 37657 8925 37691 8959
rect 37749 8925 37783 8959
rect 37933 8925 37967 8959
rect 38025 8925 38059 8959
rect 6469 8857 6503 8891
rect 6653 8857 6687 8891
rect 7205 8857 7239 8891
rect 7941 8857 7975 8891
rect 8125 8857 8159 8891
rect 9597 8857 9631 8891
rect 11897 8857 11931 8891
rect 17601 8857 17635 8891
rect 28089 8857 28123 8891
rect 28549 8857 28583 8891
rect 29837 8857 29871 8891
rect 30205 8857 30239 8891
rect 30389 8857 30423 8891
rect 35633 8857 35667 8891
rect 7757 8789 7791 8823
rect 14105 8789 14139 8823
rect 19073 8789 19107 8823
rect 20085 8789 20119 8823
rect 31953 8789 31987 8823
rect 32229 8789 32263 8823
rect 34345 8789 34379 8823
rect 28549 8585 28583 8619
rect 28917 8585 28951 8619
rect 33425 8585 33459 8619
rect 33701 8585 33735 8619
rect 37657 8585 37691 8619
rect 37841 8585 37875 8619
rect 17325 8517 17359 8551
rect 27998 8517 28032 8551
rect 28227 8517 28261 8551
rect 32505 8517 32539 8551
rect 37289 8517 37323 8551
rect 38301 8517 38335 8551
rect 8861 8449 8895 8483
rect 9045 8449 9079 8483
rect 9137 8449 9171 8483
rect 11805 8449 11839 8483
rect 11897 8449 11931 8483
rect 11989 8449 12023 8483
rect 12173 8449 12207 8483
rect 12265 8449 12299 8483
rect 13553 8449 13587 8483
rect 13829 8449 13863 8483
rect 15577 8449 15611 8483
rect 16037 8449 16071 8483
rect 16957 8449 16991 8483
rect 19257 8449 19291 8483
rect 19441 8449 19475 8483
rect 19533 8449 19567 8483
rect 19625 8449 19659 8483
rect 27905 8449 27939 8483
rect 28089 8449 28123 8483
rect 28457 8449 28491 8483
rect 28641 8449 28675 8483
rect 28733 8449 28767 8483
rect 29837 8449 29871 8483
rect 30113 8449 30147 8483
rect 31401 8449 31435 8483
rect 31677 8449 31711 8483
rect 31769 8449 31803 8483
rect 32321 8449 32355 8483
rect 34253 8449 34287 8483
rect 37473 8449 37507 8483
rect 37565 8449 37599 8483
rect 38117 8449 38151 8483
rect 38393 8449 38427 8483
rect 9229 8381 9263 8415
rect 16313 8381 16347 8415
rect 16865 8381 16899 8415
rect 17233 8381 17267 8415
rect 26985 8381 27019 8415
rect 28365 8381 28399 8415
rect 32137 8381 32171 8415
rect 33057 8381 33091 8415
rect 33333 8381 33367 8415
rect 33517 8381 33551 8415
rect 37933 8381 37967 8415
rect 11529 8313 11563 8347
rect 19809 8313 19843 8347
rect 8953 8245 8987 8279
rect 12357 8245 12391 8279
rect 16681 8245 16715 8279
rect 27629 8245 27663 8279
rect 27721 8245 27755 8279
rect 29929 8245 29963 8279
rect 34345 8245 34379 8279
rect 1777 8041 1811 8075
rect 18705 8041 18739 8075
rect 21741 8041 21775 8075
rect 26157 8041 26191 8075
rect 35357 8041 35391 8075
rect 36645 8041 36679 8075
rect 11069 7973 11103 8007
rect 8585 7905 8619 7939
rect 12449 7905 12483 7939
rect 13185 7905 13219 7939
rect 18613 7905 18647 7939
rect 19625 7905 19659 7939
rect 19717 7905 19751 7939
rect 19993 7905 20027 7939
rect 22753 7905 22787 7939
rect 24409 7905 24443 7939
rect 24685 7905 24719 7939
rect 34713 7905 34747 7939
rect 37105 7905 37139 7939
rect 7947 7837 7981 7871
rect 8125 7837 8159 7871
rect 8217 7837 8251 7871
rect 11069 7837 11103 7871
rect 11253 7837 11287 7871
rect 11345 7837 11379 7871
rect 11621 7837 11655 7871
rect 11713 7837 11747 7871
rect 11897 7837 11931 7871
rect 11989 7837 12023 7871
rect 12817 7837 12851 7871
rect 13093 7837 13127 7871
rect 18337 7837 18371 7871
rect 23489 7837 23523 7871
rect 29837 7837 29871 7871
rect 35173 7837 35207 7871
rect 35449 7837 35483 7871
rect 36829 7837 36863 7871
rect 36921 7837 36955 7871
rect 37013 7837 37047 7871
rect 1501 7769 1535 7803
rect 8401 7769 8435 7803
rect 19901 7769 19935 7803
rect 20269 7769 20303 7803
rect 21925 7769 21959 7803
rect 29561 7769 29595 7803
rect 29745 7769 29779 7803
rect 35081 7769 35115 7803
rect 35541 7769 35575 7803
rect 35725 7769 35759 7803
rect 35909 7769 35943 7803
rect 8125 7701 8159 7735
rect 11437 7701 11471 7735
rect 18889 7701 18923 7735
rect 19257 7701 19291 7735
rect 23581 7701 23615 7735
rect 29653 7701 29687 7735
rect 34995 7701 35029 7735
rect 8585 7497 8619 7531
rect 10885 7497 10919 7531
rect 16497 7497 16531 7531
rect 21097 7497 21131 7531
rect 36185 7497 36219 7531
rect 7113 7429 7147 7463
rect 9137 7429 9171 7463
rect 12725 7429 12759 7463
rect 14013 7429 14047 7463
rect 15393 7429 15427 7463
rect 18429 7429 18463 7463
rect 25513 7429 25547 7463
rect 26249 7429 26283 7463
rect 26341 7429 26375 7463
rect 27169 7429 27203 7463
rect 27261 7429 27295 7463
rect 28273 7429 28307 7463
rect 31585 7429 31619 7463
rect 32413 7429 32447 7463
rect 32505 7429 32539 7463
rect 32623 7429 32657 7463
rect 33517 7429 33551 7463
rect 35357 7429 35391 7463
rect 35817 7429 35851 7463
rect 36001 7429 36035 7463
rect 31815 7395 31849 7429
rect 35587 7395 35621 7429
rect 7297 7361 7331 7395
rect 7389 7361 7423 7395
rect 7665 7361 7699 7395
rect 7757 7361 7791 7395
rect 7849 7361 7883 7395
rect 7987 7361 8021 7395
rect 8401 7361 8435 7395
rect 8677 7361 8711 7395
rect 8953 7361 8987 7395
rect 9229 7361 9263 7395
rect 10885 7361 10919 7395
rect 11253 7361 11287 7395
rect 11805 7361 11839 7395
rect 11989 7361 12023 7395
rect 12265 7361 12299 7395
rect 12449 7361 12483 7395
rect 12633 7361 12667 7395
rect 14197 7361 14231 7395
rect 14473 7361 14507 7395
rect 14657 7361 14691 7395
rect 15117 7361 15151 7395
rect 15669 7361 15703 7395
rect 15762 7361 15796 7395
rect 15945 7361 15979 7395
rect 16129 7361 16163 7395
rect 16221 7361 16255 7395
rect 18153 7361 18187 7395
rect 20453 7361 20487 7395
rect 21281 7361 21315 7395
rect 21925 7361 21959 7395
rect 22109 7361 22143 7395
rect 23489 7361 23523 7395
rect 26065 7361 26099 7395
rect 26479 7361 26513 7395
rect 26985 7361 27019 7395
rect 27353 7361 27387 7395
rect 27629 7361 27663 7395
rect 28549 7361 28583 7395
rect 28733 7361 28767 7395
rect 28825 7361 28859 7395
rect 28917 7361 28951 7395
rect 29193 7361 29227 7395
rect 29377 7361 29411 7395
rect 29653 7361 29687 7395
rect 29929 7361 29963 7395
rect 30205 7361 30239 7395
rect 30389 7361 30423 7395
rect 30573 7361 30607 7395
rect 30757 7361 30791 7395
rect 30849 7361 30883 7395
rect 31033 7361 31067 7395
rect 31309 7361 31343 7395
rect 31493 7361 31527 7395
rect 32321 7361 32355 7395
rect 32781 7361 32815 7395
rect 33057 7361 33091 7395
rect 33425 7361 33459 7395
rect 33609 7361 33643 7395
rect 34529 7361 34563 7395
rect 34713 7361 34747 7395
rect 34805 7361 34839 7395
rect 35081 7361 35115 7395
rect 36461 7361 36495 7395
rect 8125 7293 8159 7327
rect 10701 7293 10735 7327
rect 12081 7293 12115 7327
rect 15209 7293 15243 7327
rect 15393 7293 15427 7327
rect 15854 7293 15888 7327
rect 20177 7293 20211 7327
rect 21005 7293 21039 7327
rect 21557 7293 21591 7327
rect 23765 7293 23799 7327
rect 29101 7293 29135 7327
rect 30021 7293 30055 7327
rect 33333 7293 33367 7327
rect 8769 7225 8803 7259
rect 26617 7225 26651 7259
rect 29561 7225 29595 7259
rect 30389 7225 30423 7259
rect 30849 7225 30883 7259
rect 31953 7225 31987 7259
rect 35725 7225 35759 7259
rect 7113 7157 7147 7191
rect 7481 7157 7515 7191
rect 8217 7157 8251 7191
rect 15485 7157 15519 7191
rect 16313 7157 16347 7191
rect 21465 7157 21499 7191
rect 21925 7157 21959 7191
rect 27537 7157 27571 7191
rect 28641 7157 28675 7191
rect 29009 7157 29043 7191
rect 30573 7157 30607 7191
rect 31309 7157 31343 7191
rect 31769 7157 31803 7191
rect 32137 7157 32171 7191
rect 32873 7157 32907 7191
rect 33241 7157 33275 7191
rect 34529 7157 34563 7191
rect 35501 7157 35535 7191
rect 36001 7157 36035 7191
rect 36553 7157 36587 7191
rect 8585 6953 8619 6987
rect 12173 6953 12207 6987
rect 13001 6953 13035 6987
rect 14933 6953 14967 6987
rect 15926 6953 15960 6987
rect 26328 6953 26362 6987
rect 27813 6953 27847 6987
rect 28825 6953 28859 6987
rect 29745 6953 29779 6987
rect 32229 6953 32263 6987
rect 35173 6953 35207 6987
rect 36277 6953 36311 6987
rect 12725 6885 12759 6919
rect 13185 6885 13219 6919
rect 29285 6885 29319 6919
rect 33149 6885 33183 6919
rect 6929 6817 6963 6851
rect 12449 6817 12483 6851
rect 13369 6817 13403 6851
rect 14657 6817 14691 6851
rect 15025 6817 15059 6851
rect 15669 6817 15703 6851
rect 17417 6817 17451 6851
rect 18429 6817 18463 6851
rect 21833 6817 21867 6851
rect 26065 6817 26099 6851
rect 30389 6817 30423 6851
rect 31861 6817 31895 6851
rect 32045 6817 32079 6851
rect 32321 6817 32355 6851
rect 5181 6749 5215 6783
rect 7113 6749 7147 6783
rect 8033 6749 8067 6783
rect 8493 6749 8527 6783
rect 8677 6749 8711 6783
rect 8769 6749 8803 6783
rect 11345 6749 11379 6783
rect 11493 6749 11527 6783
rect 11621 6749 11655 6783
rect 11810 6749 11844 6783
rect 12541 6749 12575 6783
rect 13277 6749 13311 6783
rect 13461 6749 13495 6783
rect 13645 6749 13679 6783
rect 13737 6749 13771 6783
rect 14473 6749 14507 6783
rect 14933 6749 14967 6783
rect 18245 6749 18279 6783
rect 19441 6749 19475 6783
rect 20085 6749 20119 6783
rect 21557 6739 21591 6773
rect 21741 6749 21775 6783
rect 25421 6749 25455 6783
rect 29193 6749 29227 6783
rect 29377 6749 29411 6783
rect 31769 6749 31803 6783
rect 31953 6749 31987 6783
rect 32229 6749 32263 6783
rect 32505 6749 32539 6783
rect 33333 6749 33367 6783
rect 33425 6749 33459 6783
rect 33609 6749 33643 6783
rect 33701 6749 33735 6783
rect 33793 6749 33827 6783
rect 33977 6749 34011 6783
rect 34161 6749 34195 6783
rect 34437 6749 34471 6783
rect 35081 6749 35115 6783
rect 35449 6749 35483 6783
rect 35725 6749 35759 6783
rect 35909 6749 35943 6783
rect 36093 6749 36127 6783
rect 29791 6715 29825 6749
rect 5457 6681 5491 6715
rect 8217 6681 8251 6715
rect 11713 6681 11747 6715
rect 12081 6681 12115 6715
rect 12817 6681 12851 6715
rect 13022 6681 13056 6715
rect 13921 6681 13955 6715
rect 21649 6681 21683 6715
rect 22109 6681 22143 6715
rect 23857 6681 23891 6715
rect 28641 6681 28675 6715
rect 29561 6681 29595 6715
rect 30113 6681 30147 6715
rect 34069 6681 34103 6715
rect 34299 6681 34333 6715
rect 34897 6681 34931 6715
rect 7665 6613 7699 6647
rect 8401 6613 8435 6647
rect 11989 6613 12023 6647
rect 14105 6613 14139 6647
rect 14565 6613 14599 6647
rect 15301 6613 15335 6647
rect 19257 6613 19291 6647
rect 20637 6613 20671 6647
rect 25973 6613 26007 6647
rect 28846 6613 28880 6647
rect 29009 6613 29043 6647
rect 29929 6613 29963 6647
rect 31585 6613 31619 6647
rect 32689 6613 32723 6647
rect 35541 6613 35575 6647
rect 5549 6409 5583 6443
rect 6377 6409 6411 6443
rect 6745 6409 6779 6443
rect 10885 6409 10919 6443
rect 11529 6409 11563 6443
rect 12449 6409 12483 6443
rect 13277 6409 13311 6443
rect 14473 6409 14507 6443
rect 18337 6409 18371 6443
rect 20545 6409 20579 6443
rect 20637 6409 20671 6443
rect 26249 6409 26283 6443
rect 26709 6409 26743 6443
rect 35449 6409 35483 6443
rect 6837 6341 6871 6375
rect 10333 6341 10367 6375
rect 18797 6341 18831 6375
rect 19165 6341 19199 6375
rect 19901 6341 19935 6375
rect 22385 6341 22419 6375
rect 29561 6341 29595 6375
rect 33701 6341 33735 6375
rect 5733 6273 5767 6307
rect 8033 6273 8067 6307
rect 8309 6273 8343 6307
rect 10793 6273 10827 6307
rect 11713 6273 11747 6307
rect 11989 6273 12023 6307
rect 12081 6273 12115 6307
rect 13185 6273 13219 6307
rect 14105 6273 14139 6307
rect 18705 6273 18739 6307
rect 21189 6273 21223 6307
rect 22293 6273 22327 6307
rect 22477 6273 22511 6307
rect 24501 6273 24535 6307
rect 26525 6273 26559 6307
rect 26801 6273 26835 6307
rect 29469 6273 29503 6307
rect 29653 6271 29687 6305
rect 31217 6273 31251 6307
rect 31401 6273 31435 6307
rect 35633 6273 35667 6307
rect 6929 6205 6963 6239
rect 8585 6205 8619 6239
rect 10977 6205 11011 6239
rect 12173 6205 12207 6239
rect 14197 6205 14231 6239
rect 18981 6205 19015 6239
rect 20821 6205 20855 6239
rect 24777 6205 24811 6239
rect 26341 6205 26375 6239
rect 34069 6205 34103 6239
rect 34805 6205 34839 6239
rect 20177 6137 20211 6171
rect 33701 6137 33735 6171
rect 33977 6137 34011 6171
rect 7849 6069 7883 6103
rect 10425 6069 10459 6103
rect 11897 6069 11931 6103
rect 12265 6069 12299 6103
rect 21005 6069 21039 6103
rect 31217 6069 31251 6103
rect 33885 6069 33919 6103
rect 35725 6069 35759 6103
rect 10885 5865 10919 5899
rect 21097 5865 21131 5899
rect 28641 5865 28675 5899
rect 33885 5865 33919 5899
rect 40969 5865 41003 5899
rect 9137 5729 9171 5763
rect 19349 5729 19383 5763
rect 19625 5729 19659 5763
rect 21189 5729 21223 5763
rect 34069 5729 34103 5763
rect 16129 5661 16163 5695
rect 27721 5661 27755 5695
rect 27813 5661 27847 5695
rect 28181 5661 28215 5695
rect 28273 5661 28307 5695
rect 28457 5661 28491 5695
rect 28733 5661 28767 5695
rect 29561 5661 29595 5695
rect 30573 5661 30607 5695
rect 30757 5661 30791 5695
rect 30941 5661 30975 5695
rect 33241 5661 33275 5695
rect 33885 5661 33919 5695
rect 34161 5661 34195 5695
rect 35357 5661 35391 5695
rect 35633 5661 35667 5695
rect 36277 5661 36311 5695
rect 40785 5661 40819 5695
rect 9413 5593 9447 5627
rect 16405 5593 16439 5627
rect 18153 5593 18187 5627
rect 21465 5593 21499 5627
rect 23213 5593 23247 5627
rect 30297 5593 30331 5627
rect 30849 5593 30883 5627
rect 28917 5525 28951 5559
rect 31125 5525 31159 5559
rect 33793 5525 33827 5559
rect 34345 5525 34379 5559
rect 35173 5525 35207 5559
rect 35541 5525 35575 5559
rect 36829 5525 36863 5559
rect 9597 5321 9631 5355
rect 13277 5321 13311 5355
rect 21833 5321 21867 5355
rect 22477 5321 22511 5355
rect 31401 5321 31435 5355
rect 32321 5321 32355 5355
rect 36921 5321 36955 5355
rect 11805 5253 11839 5287
rect 16681 5253 16715 5287
rect 17049 5253 17083 5287
rect 18429 5253 18463 5287
rect 33609 5253 33643 5287
rect 35449 5253 35483 5287
rect 9781 5185 9815 5219
rect 16865 5185 16899 5219
rect 17141 5185 17175 5219
rect 18153 5185 18187 5219
rect 22293 5185 22327 5219
rect 27169 5185 27203 5219
rect 27261 5185 27295 5219
rect 27537 5185 27571 5219
rect 27629 5191 27663 5225
rect 28365 5185 28399 5219
rect 31309 5185 31343 5219
rect 32689 5185 32723 5219
rect 33333 5185 33367 5219
rect 35173 5185 35207 5219
rect 9965 5117 9999 5151
rect 11529 5117 11563 5151
rect 22201 5117 22235 5151
rect 27905 5117 27939 5151
rect 28641 5117 28675 5151
rect 30389 5117 30423 5151
rect 31493 5117 31527 5151
rect 32781 5117 32815 5151
rect 35081 5117 35115 5151
rect 10609 4981 10643 5015
rect 19901 4981 19935 5015
rect 26985 4981 27019 5015
rect 27445 4981 27479 5015
rect 27721 4981 27755 5015
rect 27813 4981 27847 5015
rect 30941 4981 30975 5015
rect 32965 4981 32999 5015
rect 3617 4777 3651 4811
rect 16294 4777 16328 4811
rect 17785 4777 17819 4811
rect 27951 4777 27985 4811
rect 31769 4777 31803 4811
rect 33655 4777 33689 4811
rect 1869 4641 1903 4675
rect 16037 4641 16071 4675
rect 26157 4641 26191 4675
rect 26525 4641 26559 4675
rect 30021 4641 30055 4675
rect 31861 4641 31895 4675
rect 32229 4641 32263 4675
rect 36001 4573 36035 4607
rect 2145 4505 2179 4539
rect 30297 4505 30331 4539
rect 36185 4437 36219 4471
rect 1961 4233 1995 4267
rect 30573 4233 30607 4267
rect 1869 4097 1903 4131
rect 10793 4097 10827 4131
rect 30757 4097 30791 4131
rect 10977 3893 11011 3927
rect 15025 3553 15059 3587
rect 14749 3485 14783 3519
rect 14841 3485 14875 3519
rect 14105 3009 14139 3043
rect 14197 2805 14231 2839
rect 40785 2601 40819 2635
rect 29837 2465 29871 2499
rect 7297 2397 7331 2431
rect 22109 2397 22143 2431
rect 29561 2397 29595 2431
rect 33057 2397 33091 2431
rect 40693 2329 40727 2363
rect 7389 2261 7423 2295
rect 22201 2261 22235 2295
rect 33149 2261 33183 2295
<< metal1 >>
rect 1104 42458 41400 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 41400 42458
rect 1104 42384 41400 42406
rect 1302 42304 1308 42356
rect 1360 42344 1366 42356
rect 1581 42347 1639 42353
rect 1581 42344 1593 42347
rect 1360 42316 1593 42344
rect 1360 42304 1366 42316
rect 1581 42313 1593 42316
rect 1627 42313 1639 42347
rect 1581 42307 1639 42313
rect 35066 42304 35072 42356
rect 35124 42304 35130 42356
rect 9030 42236 9036 42288
rect 9088 42276 9094 42288
rect 9217 42279 9275 42285
rect 9217 42276 9229 42279
rect 9088 42248 9229 42276
rect 9088 42236 9094 42248
rect 9217 42245 9229 42248
rect 9263 42245 9275 42279
rect 9217 42239 9275 42245
rect 1486 42168 1492 42220
rect 1544 42168 1550 42220
rect 17494 42168 17500 42220
rect 17552 42168 17558 42220
rect 19426 42168 19432 42220
rect 19484 42208 19490 42220
rect 19705 42211 19763 42217
rect 19705 42208 19717 42211
rect 19484 42180 19717 42208
rect 19484 42168 19490 42180
rect 19705 42177 19717 42180
rect 19751 42177 19763 42211
rect 19705 42171 19763 42177
rect 30926 42168 30932 42220
rect 30984 42208 30990 42220
rect 31021 42211 31079 42217
rect 31021 42208 31033 42211
rect 30984 42180 31033 42208
rect 30984 42168 30990 42180
rect 31021 42177 31033 42180
rect 31067 42177 31079 42211
rect 31021 42171 31079 42177
rect 34514 42168 34520 42220
rect 34572 42208 34578 42220
rect 34977 42211 35035 42217
rect 34977 42208 34989 42211
rect 34572 42180 34989 42208
rect 34572 42168 34578 42180
rect 34977 42177 34989 42180
rect 35023 42208 35035 42211
rect 35621 42211 35679 42217
rect 35621 42208 35633 42211
rect 35023 42180 35633 42208
rect 35023 42177 35035 42180
rect 34977 42171 35035 42177
rect 35621 42177 35633 42180
rect 35667 42177 35679 42211
rect 35621 42171 35679 42177
rect 38654 42168 38660 42220
rect 38712 42208 38718 42220
rect 38749 42211 38807 42217
rect 38749 42208 38761 42211
rect 38712 42180 38761 42208
rect 38712 42168 38718 42180
rect 38749 42177 38761 42180
rect 38795 42177 38807 42211
rect 38749 42171 38807 42177
rect 31294 42100 31300 42152
rect 31352 42100 31358 42152
rect 37182 42100 37188 42152
rect 37240 42140 37246 42152
rect 38933 42143 38991 42149
rect 38933 42140 38945 42143
rect 37240 42112 38945 42140
rect 37240 42100 37246 42112
rect 38933 42109 38945 42112
rect 38979 42109 38991 42143
rect 38933 42103 38991 42109
rect 9306 41964 9312 42016
rect 9364 41964 9370 42016
rect 17310 41964 17316 42016
rect 17368 41964 17374 42016
rect 19521 42007 19579 42013
rect 19521 41973 19533 42007
rect 19567 42004 19579 42007
rect 19610 42004 19616 42016
rect 19567 41976 19616 42004
rect 19567 41973 19579 41976
rect 19521 41967 19579 41973
rect 19610 41964 19616 41976
rect 19668 41964 19674 42016
rect 1104 41914 41400 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 41400 41914
rect 1104 41840 41400 41862
rect 17116 41803 17174 41809
rect 17116 41769 17128 41803
rect 17162 41800 17174 41803
rect 17310 41800 17316 41812
rect 17162 41772 17316 41800
rect 17162 41769 17174 41772
rect 17116 41763 17174 41769
rect 17310 41760 17316 41772
rect 17368 41760 17374 41812
rect 10137 41667 10195 41673
rect 10137 41633 10149 41667
rect 10183 41664 10195 41667
rect 11146 41664 11152 41676
rect 10183 41636 11152 41664
rect 10183 41633 10195 41636
rect 10137 41627 10195 41633
rect 11146 41624 11152 41636
rect 11204 41624 11210 41676
rect 14093 41667 14151 41673
rect 14093 41633 14105 41667
rect 14139 41664 14151 41667
rect 16853 41667 16911 41673
rect 16853 41664 16865 41667
rect 14139 41636 16865 41664
rect 14139 41633 14151 41636
rect 14093 41627 14151 41633
rect 16853 41633 16865 41636
rect 16899 41664 16911 41667
rect 19334 41664 19340 41676
rect 16899 41636 19340 41664
rect 16899 41633 16911 41636
rect 16853 41627 16911 41633
rect 19334 41624 19340 41636
rect 19392 41624 19398 41676
rect 19610 41624 19616 41676
rect 19668 41624 19674 41676
rect 19978 41624 19984 41676
rect 20036 41664 20042 41676
rect 21361 41667 21419 41673
rect 21361 41664 21373 41667
rect 20036 41636 21373 41664
rect 20036 41624 20042 41636
rect 21361 41633 21373 41636
rect 21407 41633 21419 41667
rect 21361 41627 21419 41633
rect 9861 41599 9919 41605
rect 9861 41565 9873 41599
rect 9907 41565 9919 41599
rect 11793 41599 11851 41605
rect 11793 41596 11805 41599
rect 9861 41559 9919 41565
rect 11440 41568 11805 41596
rect 9876 41460 9904 41559
rect 10594 41488 10600 41540
rect 10652 41488 10658 41540
rect 10962 41460 10968 41472
rect 9876 41432 10968 41460
rect 10962 41420 10968 41432
rect 11020 41460 11026 41472
rect 11440 41460 11468 41568
rect 11793 41565 11805 41568
rect 11839 41565 11851 41599
rect 13202 41568 14044 41596
rect 11793 41559 11851 41565
rect 14016 41540 14044 41568
rect 16114 41556 16120 41608
rect 16172 41556 16178 41608
rect 18782 41596 18788 41608
rect 18262 41568 18788 41596
rect 18782 41556 18788 41568
rect 18840 41556 18846 41608
rect 18877 41599 18935 41605
rect 18877 41565 18889 41599
rect 18923 41596 18935 41599
rect 18923 41568 19012 41596
rect 18923 41565 18935 41568
rect 18877 41559 18935 41565
rect 12066 41488 12072 41540
rect 12124 41488 12130 41540
rect 13817 41531 13875 41537
rect 13817 41528 13829 41531
rect 13372 41500 13829 41528
rect 11020 41432 11468 41460
rect 11020 41420 11026 41432
rect 11514 41420 11520 41472
rect 11572 41460 11578 41472
rect 11609 41463 11667 41469
rect 11609 41460 11621 41463
rect 11572 41432 11621 41460
rect 11572 41420 11578 41432
rect 11609 41429 11621 41432
rect 11655 41429 11667 41463
rect 11609 41423 11667 41429
rect 12894 41420 12900 41472
rect 12952 41460 12958 41472
rect 13372 41460 13400 41500
rect 13817 41497 13829 41500
rect 13863 41497 13875 41531
rect 13817 41491 13875 41497
rect 13998 41488 14004 41540
rect 14056 41488 14062 41540
rect 14366 41488 14372 41540
rect 14424 41488 14430 41540
rect 14476 41500 14858 41528
rect 12952 41432 13400 41460
rect 14016 41460 14044 41488
rect 14476 41460 14504 41500
rect 17402 41488 17408 41540
rect 17460 41488 17466 41540
rect 14016 41432 14504 41460
rect 17420 41460 17448 41488
rect 18984 41460 19012 41568
rect 22094 41556 22100 41608
rect 22152 41596 22158 41608
rect 22189 41599 22247 41605
rect 22189 41596 22201 41599
rect 22152 41568 22201 41596
rect 22152 41556 22158 41568
rect 22189 41565 22201 41568
rect 22235 41565 22247 41599
rect 22189 41559 22247 41565
rect 20898 41528 20904 41540
rect 20838 41500 20904 41528
rect 20898 41488 20904 41500
rect 20956 41488 20962 41540
rect 22462 41488 22468 41540
rect 22520 41488 22526 41540
rect 23934 41528 23940 41540
rect 23690 41500 23940 41528
rect 23934 41488 23940 41500
rect 23992 41488 23998 41540
rect 24210 41488 24216 41540
rect 24268 41488 24274 41540
rect 17420 41432 19012 41460
rect 12952 41420 12958 41432
rect 1104 41370 41400 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 41400 41370
rect 1104 41296 41400 41318
rect 12066 41216 12072 41268
rect 12124 41256 12130 41268
rect 12345 41259 12403 41265
rect 12345 41256 12357 41259
rect 12124 41228 12357 41256
rect 12124 41216 12130 41228
rect 12345 41225 12357 41228
rect 12391 41225 12403 41259
rect 12345 41219 12403 41225
rect 14277 41259 14335 41265
rect 14277 41225 14289 41259
rect 14323 41256 14335 41259
rect 14366 41256 14372 41268
rect 14323 41228 14372 41256
rect 14323 41225 14335 41228
rect 14277 41219 14335 41225
rect 14366 41216 14372 41228
rect 14424 41216 14430 41268
rect 16853 41259 16911 41265
rect 16853 41225 16865 41259
rect 16899 41256 16911 41259
rect 17494 41256 17500 41268
rect 16899 41228 17500 41256
rect 16899 41225 16911 41228
rect 16853 41219 16911 41225
rect 17494 41216 17500 41228
rect 17552 41216 17558 41268
rect 19426 41216 19432 41268
rect 19484 41216 19490 41268
rect 19797 41259 19855 41265
rect 19797 41225 19809 41259
rect 19843 41256 19855 41259
rect 19978 41256 19984 41268
rect 19843 41228 19984 41256
rect 19843 41225 19855 41228
rect 19797 41219 19855 41225
rect 19978 41216 19984 41228
rect 20036 41216 20042 41268
rect 21545 41259 21603 41265
rect 21545 41225 21557 41259
rect 21591 41256 21603 41259
rect 23842 41256 23848 41268
rect 21591 41228 23848 41256
rect 21591 41225 21603 41228
rect 21545 41219 21603 41225
rect 23842 41216 23848 41228
rect 23900 41216 23906 41268
rect 24210 41216 24216 41268
rect 24268 41256 24274 41268
rect 41874 41256 41880 41268
rect 24268 41228 41880 41256
rect 24268 41216 24274 41228
rect 41874 41216 41880 41228
rect 41932 41216 41938 41268
rect 1670 41148 1676 41200
rect 1728 41148 1734 41200
rect 12713 41191 12771 41197
rect 12713 41188 12725 41191
rect 12268 41160 12725 41188
rect 3602 41120 3608 41132
rect 2806 41092 3608 41120
rect 3602 41080 3608 41092
rect 3660 41080 3666 41132
rect 12268 41129 12296 41160
rect 12713 41157 12725 41160
rect 12759 41157 12771 41191
rect 14921 41191 14979 41197
rect 14921 41188 14933 41191
rect 12713 41151 12771 41157
rect 14108 41160 14933 41188
rect 12253 41123 12311 41129
rect 5198 41092 5304 41120
rect 1397 41055 1455 41061
rect 1397 41021 1409 41055
rect 1443 41052 1455 41055
rect 2682 41052 2688 41064
rect 1443 41024 2688 41052
rect 1443 41021 1455 41024
rect 1397 41015 1455 41021
rect 2682 41012 2688 41024
rect 2740 41052 2746 41064
rect 2740 41024 2820 41052
rect 2740 41012 2746 41024
rect 2792 40984 2820 41024
rect 2866 41012 2872 41064
rect 2924 41052 2930 41064
rect 3418 41052 3424 41064
rect 2924 41024 3424 41052
rect 2924 41012 2930 41024
rect 3418 41012 3424 41024
rect 3476 41012 3482 41064
rect 3789 41055 3847 41061
rect 3789 41021 3801 41055
rect 3835 41021 3847 41055
rect 3789 41015 3847 41021
rect 3804 40984 3832 41015
rect 4062 41012 4068 41064
rect 4120 41012 4126 41064
rect 2792 40956 3832 40984
rect 5276 40928 5304 41092
rect 12253 41089 12265 41123
rect 12299 41089 12311 41123
rect 12253 41083 12311 41089
rect 12437 41123 12495 41129
rect 12437 41089 12449 41123
rect 12483 41120 12495 41123
rect 12526 41120 12532 41132
rect 12483 41092 12532 41120
rect 12483 41089 12495 41092
rect 12437 41083 12495 41089
rect 12526 41080 12532 41092
rect 12584 41080 12590 41132
rect 12621 41123 12679 41129
rect 12621 41089 12633 41123
rect 12667 41089 12679 41123
rect 12621 41083 12679 41089
rect 5350 41012 5356 41064
rect 5408 41052 5414 41064
rect 5813 41055 5871 41061
rect 5813 41052 5825 41055
rect 5408 41024 5825 41052
rect 5408 41012 5414 41024
rect 5813 41021 5825 41024
rect 5859 41021 5871 41055
rect 5813 41015 5871 41021
rect 10505 41055 10563 41061
rect 10505 41021 10517 41055
rect 10551 41052 10563 41055
rect 11514 41052 11520 41064
rect 10551 41024 11520 41052
rect 10551 41021 10563 41024
rect 10505 41015 10563 41021
rect 11514 41012 11520 41024
rect 11572 41012 11578 41064
rect 12636 40984 12664 41083
rect 12802 41080 12808 41132
rect 12860 41080 12866 41132
rect 14108 41129 14136 41160
rect 14921 41157 14933 41160
rect 14967 41157 14979 41191
rect 22094 41188 22100 41200
rect 14921 41151 14979 41157
rect 16224 41160 21680 41188
rect 14093 41123 14151 41129
rect 14093 41089 14105 41123
rect 14139 41089 14151 41123
rect 14093 41083 14151 41089
rect 14274 41080 14280 41132
rect 14332 41080 14338 41132
rect 14829 41123 14887 41129
rect 14829 41089 14841 41123
rect 14875 41089 14887 41123
rect 14829 41083 14887 41089
rect 15013 41123 15071 41129
rect 15013 41089 15025 41123
rect 15059 41120 15071 41123
rect 16114 41120 16120 41132
rect 15059 41092 16120 41120
rect 15059 41089 15071 41092
rect 15013 41083 15071 41089
rect 14844 41052 14872 41083
rect 16114 41080 16120 41092
rect 16172 41080 16178 41132
rect 16224 41052 16252 41160
rect 21652 41132 21680 41160
rect 21836 41160 22100 41188
rect 17218 41080 17224 41132
rect 17276 41080 17282 41132
rect 17420 41092 20116 41120
rect 14844 41024 16252 41052
rect 14844 40984 14872 41024
rect 17310 41012 17316 41064
rect 17368 41012 17374 41064
rect 12636 40956 14872 40984
rect 15378 40944 15384 40996
rect 15436 40984 15442 40996
rect 17420 40984 17448 41092
rect 17497 41055 17555 41061
rect 17497 41021 17509 41055
rect 17543 41052 17555 41055
rect 17586 41052 17592 41064
rect 17543 41024 17592 41052
rect 17543 41021 17555 41024
rect 17497 41015 17555 41021
rect 17586 41012 17592 41024
rect 17644 41012 17650 41064
rect 20088 41061 20116 41092
rect 21358 41080 21364 41132
rect 21416 41080 21422 41132
rect 21634 41080 21640 41132
rect 21692 41080 21698 41132
rect 21836 41064 21864 41160
rect 22094 41148 22100 41160
rect 22152 41148 22158 41200
rect 23382 41120 23388 41132
rect 23230 41092 23388 41120
rect 23382 41080 23388 41092
rect 23440 41120 23446 41132
rect 23934 41120 23940 41132
rect 23440 41092 23940 41120
rect 23440 41080 23446 41092
rect 23934 41080 23940 41092
rect 23992 41080 23998 41132
rect 40770 41080 40776 41132
rect 40828 41080 40834 41132
rect 19889 41055 19947 41061
rect 19889 41021 19901 41055
rect 19935 41021 19947 41055
rect 19889 41015 19947 41021
rect 20073 41055 20131 41061
rect 20073 41021 20085 41055
rect 20119 41052 20131 41055
rect 21082 41052 21088 41064
rect 20119 41024 21088 41052
rect 20119 41021 20131 41024
rect 20073 41015 20131 41021
rect 15436 40956 17448 40984
rect 15436 40944 15442 40956
rect 5258 40876 5264 40928
rect 5316 40876 5322 40928
rect 11054 40876 11060 40928
rect 11112 40876 11118 40928
rect 16022 40876 16028 40928
rect 16080 40916 16086 40928
rect 19904 40916 19932 41015
rect 21082 41012 21088 41024
rect 21140 41012 21146 41064
rect 21818 41012 21824 41064
rect 21876 41012 21882 41064
rect 22097 41055 22155 41061
rect 22097 41052 22109 41055
rect 21928 41024 22109 41052
rect 21177 40987 21235 40993
rect 21177 40953 21189 40987
rect 21223 40984 21235 40987
rect 21928 40984 21956 41024
rect 22097 41021 22109 41024
rect 22143 41021 22155 41055
rect 22097 41015 22155 41021
rect 23842 41012 23848 41064
rect 23900 41012 23906 41064
rect 21223 40956 21956 40984
rect 21223 40953 21235 40956
rect 21177 40947 21235 40953
rect 16080 40888 19932 40916
rect 16080 40876 16086 40888
rect 40954 40876 40960 40928
rect 41012 40876 41018 40928
rect 1104 40826 41400 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 41400 40826
rect 1104 40752 41400 40774
rect 1670 40672 1676 40724
rect 1728 40712 1734 40724
rect 2041 40715 2099 40721
rect 2041 40712 2053 40715
rect 1728 40684 2053 40712
rect 1728 40672 1734 40684
rect 2041 40681 2053 40684
rect 2087 40681 2099 40715
rect 2041 40675 2099 40681
rect 4062 40672 4068 40724
rect 4120 40712 4126 40724
rect 4249 40715 4307 40721
rect 4249 40712 4261 40715
rect 4120 40684 4261 40712
rect 4120 40672 4126 40684
rect 4249 40681 4261 40684
rect 4295 40681 4307 40715
rect 11057 40715 11115 40721
rect 4249 40675 4307 40681
rect 5368 40684 9904 40712
rect 2501 40647 2559 40653
rect 2501 40613 2513 40647
rect 2547 40613 2559 40647
rect 2501 40607 2559 40613
rect 2225 40511 2283 40517
rect 2225 40477 2237 40511
rect 2271 40508 2283 40511
rect 2516 40508 2544 40607
rect 3145 40579 3203 40585
rect 3145 40545 3157 40579
rect 3191 40576 3203 40579
rect 3418 40576 3424 40588
rect 3191 40548 3424 40576
rect 3191 40545 3203 40548
rect 3145 40539 3203 40545
rect 3418 40536 3424 40548
rect 3476 40576 3482 40588
rect 5261 40579 5319 40585
rect 5261 40576 5273 40579
rect 3476 40548 5273 40576
rect 3476 40536 3482 40548
rect 5261 40545 5273 40548
rect 5307 40576 5319 40579
rect 5368 40576 5396 40684
rect 9766 40644 9772 40656
rect 5307 40548 5396 40576
rect 6288 40616 9772 40644
rect 5307 40545 5319 40548
rect 5261 40539 5319 40545
rect 2271 40480 2544 40508
rect 2271 40477 2283 40480
rect 2225 40471 2283 40477
rect 2866 40468 2872 40520
rect 2924 40468 2930 40520
rect 4433 40511 4491 40517
rect 4433 40477 4445 40511
rect 4479 40508 4491 40511
rect 4614 40508 4620 40520
rect 4479 40480 4620 40508
rect 4479 40477 4491 40480
rect 4433 40471 4491 40477
rect 4614 40468 4620 40480
rect 4672 40468 4678 40520
rect 4985 40511 5043 40517
rect 4985 40477 4997 40511
rect 5031 40508 5043 40511
rect 5350 40508 5356 40520
rect 5031 40480 5356 40508
rect 5031 40477 5043 40480
rect 4985 40471 5043 40477
rect 5350 40468 5356 40480
rect 5408 40468 5414 40520
rect 2961 40443 3019 40449
rect 2961 40409 2973 40443
rect 3007 40440 3019 40443
rect 6288 40440 6316 40616
rect 9766 40604 9772 40616
rect 9824 40604 9830 40656
rect 9876 40644 9904 40684
rect 11057 40681 11069 40715
rect 11103 40712 11115 40715
rect 11146 40712 11152 40724
rect 11103 40684 11152 40712
rect 11103 40681 11115 40684
rect 11057 40675 11115 40681
rect 11146 40672 11152 40684
rect 11204 40672 11210 40724
rect 15378 40712 15384 40724
rect 12406 40684 15384 40712
rect 12406 40644 12434 40684
rect 15378 40672 15384 40684
rect 15436 40672 15442 40724
rect 15470 40672 15476 40724
rect 15528 40712 15534 40724
rect 17037 40715 17095 40721
rect 15528 40684 16068 40712
rect 15528 40672 15534 40684
rect 15654 40644 15660 40656
rect 9876 40616 12434 40644
rect 14844 40616 15660 40644
rect 13262 40576 13268 40588
rect 8864 40548 13268 40576
rect 3007 40412 6316 40440
rect 3007 40409 3019 40412
rect 2961 40403 3019 40409
rect 8018 40400 8024 40452
rect 8076 40400 8082 40452
rect 8864 40384 8892 40548
rect 10410 40468 10416 40520
rect 10468 40468 10474 40520
rect 10561 40511 10619 40517
rect 10561 40477 10573 40511
rect 10607 40477 10619 40511
rect 10704 40508 10732 40548
rect 13262 40536 13268 40548
rect 13320 40536 13326 40588
rect 14369 40579 14427 40585
rect 14369 40545 14381 40579
rect 14415 40576 14427 40579
rect 14415 40548 14596 40576
rect 14415 40545 14427 40548
rect 14369 40539 14427 40545
rect 10878 40511 10936 40517
rect 10878 40508 10890 40511
rect 10704 40480 10890 40508
rect 10561 40471 10619 40477
rect 10878 40477 10890 40480
rect 10924 40477 10936 40511
rect 10878 40471 10936 40477
rect 4614 40332 4620 40384
rect 4672 40332 4678 40384
rect 4798 40332 4804 40384
rect 4856 40372 4862 40384
rect 5077 40375 5135 40381
rect 5077 40372 5089 40375
rect 4856 40344 5089 40372
rect 4856 40332 4862 40344
rect 5077 40341 5089 40344
rect 5123 40341 5135 40375
rect 5077 40335 5135 40341
rect 8297 40375 8355 40381
rect 8297 40341 8309 40375
rect 8343 40372 8355 40375
rect 8846 40372 8852 40384
rect 8343 40344 8852 40372
rect 8343 40341 8355 40344
rect 8297 40335 8355 40341
rect 8846 40332 8852 40344
rect 8904 40332 8910 40384
rect 9950 40332 9956 40384
rect 10008 40372 10014 40384
rect 10576 40372 10604 40471
rect 11054 40468 11060 40520
rect 11112 40468 11118 40520
rect 11241 40511 11299 40517
rect 11241 40477 11253 40511
rect 11287 40477 11299 40511
rect 11241 40471 11299 40477
rect 11425 40511 11483 40517
rect 11425 40477 11437 40511
rect 11471 40508 11483 40511
rect 11514 40508 11520 40520
rect 11471 40480 11520 40508
rect 11471 40477 11483 40480
rect 11425 40471 11483 40477
rect 10686 40400 10692 40452
rect 10744 40400 10750 40452
rect 10781 40443 10839 40449
rect 10781 40409 10793 40443
rect 10827 40440 10839 40443
rect 11072 40440 11100 40468
rect 10827 40412 11100 40440
rect 11256 40440 11284 40471
rect 11514 40468 11520 40480
rect 11572 40468 11578 40520
rect 14182 40468 14188 40520
rect 14240 40508 14246 40520
rect 14568 40517 14596 40548
rect 14277 40511 14335 40517
rect 14277 40508 14289 40511
rect 14240 40480 14289 40508
rect 14240 40468 14246 40480
rect 14277 40477 14289 40480
rect 14323 40477 14335 40511
rect 14277 40471 14335 40477
rect 14461 40511 14519 40517
rect 14461 40477 14473 40511
rect 14507 40477 14519 40511
rect 14461 40471 14519 40477
rect 14553 40511 14611 40517
rect 14553 40477 14565 40511
rect 14599 40477 14611 40511
rect 14553 40471 14611 40477
rect 11256 40412 11468 40440
rect 10827 40409 10839 40412
rect 10781 40403 10839 40409
rect 11440 40384 11468 40412
rect 11238 40372 11244 40384
rect 10008 40344 11244 40372
rect 10008 40332 10014 40344
rect 11238 40332 11244 40344
rect 11296 40332 11302 40384
rect 11330 40332 11336 40384
rect 11388 40332 11394 40384
rect 11422 40332 11428 40384
rect 11480 40332 11486 40384
rect 12342 40332 12348 40384
rect 12400 40372 12406 40384
rect 14274 40372 14280 40384
rect 12400 40344 14280 40372
rect 12400 40332 12406 40344
rect 14274 40332 14280 40344
rect 14332 40332 14338 40384
rect 14476 40372 14504 40471
rect 14734 40468 14740 40520
rect 14792 40468 14798 40520
rect 14844 40517 14872 40616
rect 15654 40604 15660 40616
rect 15712 40604 15718 40656
rect 16040 40653 16068 40684
rect 17037 40681 17049 40715
rect 17083 40712 17095 40715
rect 17218 40712 17224 40724
rect 17083 40684 17224 40712
rect 17083 40681 17095 40684
rect 17037 40675 17095 40681
rect 17218 40672 17224 40684
rect 17276 40672 17282 40724
rect 21358 40712 21364 40724
rect 18800 40684 21364 40712
rect 16025 40647 16083 40653
rect 16025 40613 16037 40647
rect 16071 40613 16083 40647
rect 16025 40607 16083 40613
rect 17957 40647 18015 40653
rect 17957 40613 17969 40647
rect 18003 40644 18015 40647
rect 18800 40644 18828 40684
rect 21358 40672 21364 40684
rect 21416 40672 21422 40724
rect 22462 40672 22468 40724
rect 22520 40672 22526 40724
rect 18003 40616 18828 40644
rect 18003 40613 18015 40616
rect 17957 40607 18015 40613
rect 14921 40579 14979 40585
rect 14921 40545 14933 40579
rect 14967 40576 14979 40579
rect 16209 40579 16267 40585
rect 14967 40548 15792 40576
rect 14967 40545 14979 40548
rect 14921 40539 14979 40545
rect 14829 40511 14887 40517
rect 14829 40477 14841 40511
rect 14875 40477 14887 40511
rect 14829 40471 14887 40477
rect 15010 40468 15016 40520
rect 15068 40468 15074 40520
rect 15289 40511 15347 40517
rect 15289 40508 15301 40511
rect 15212 40480 15301 40508
rect 14645 40443 14703 40449
rect 14645 40409 14657 40443
rect 14691 40440 14703 40443
rect 15212 40440 15240 40480
rect 15289 40477 15301 40480
rect 15335 40508 15347 40511
rect 15378 40508 15384 40520
rect 15335 40480 15384 40508
rect 15335 40477 15347 40480
rect 15289 40471 15347 40477
rect 15378 40468 15384 40480
rect 15436 40468 15442 40520
rect 15473 40511 15531 40517
rect 15473 40477 15485 40511
rect 15519 40477 15531 40511
rect 15764 40508 15792 40548
rect 16209 40545 16221 40579
rect 16255 40576 16267 40579
rect 16393 40579 16451 40585
rect 16393 40576 16405 40579
rect 16255 40548 16405 40576
rect 16255 40545 16267 40548
rect 16209 40539 16267 40545
rect 16393 40545 16405 40548
rect 16439 40545 16451 40579
rect 16393 40539 16451 40545
rect 16574 40536 16580 40588
rect 16632 40576 16638 40588
rect 18800 40585 18828 40616
rect 17681 40579 17739 40585
rect 17681 40576 17693 40579
rect 16632 40548 17693 40576
rect 16632 40536 16638 40548
rect 17681 40545 17693 40548
rect 17727 40576 17739 40579
rect 18785 40579 18843 40585
rect 17727 40548 18000 40576
rect 17727 40545 17739 40548
rect 17681 40539 17739 40545
rect 16485 40511 16543 40517
rect 16485 40508 16497 40511
rect 15764 40480 16497 40508
rect 15473 40471 15531 40477
rect 16485 40477 16497 40480
rect 16531 40477 16543 40511
rect 16485 40471 16543 40477
rect 15488 40440 15516 40471
rect 16942 40468 16948 40520
rect 17000 40508 17006 40520
rect 17865 40511 17923 40517
rect 17865 40508 17877 40511
rect 17000 40480 17877 40508
rect 17000 40468 17006 40480
rect 17865 40477 17877 40480
rect 17911 40477 17923 40511
rect 17972 40508 18000 40548
rect 18785 40545 18797 40579
rect 18831 40545 18843 40579
rect 18785 40539 18843 40545
rect 18877 40579 18935 40585
rect 18877 40545 18889 40579
rect 18923 40545 18935 40579
rect 18877 40539 18935 40545
rect 18892 40508 18920 40539
rect 19426 40536 19432 40588
rect 19484 40576 19490 40588
rect 19484 40548 20760 40576
rect 19484 40536 19490 40548
rect 20732 40520 20760 40548
rect 21634 40536 21640 40588
rect 21692 40576 21698 40588
rect 22278 40576 22284 40588
rect 21692 40548 22284 40576
rect 21692 40536 21698 40548
rect 22278 40536 22284 40548
rect 22336 40576 22342 40588
rect 22336 40548 22692 40576
rect 22336 40536 22342 40548
rect 17972 40480 18920 40508
rect 17865 40471 17923 40477
rect 20714 40468 20720 40520
rect 20772 40468 20778 40520
rect 22373 40511 22431 40517
rect 22373 40477 22385 40511
rect 22419 40477 22431 40511
rect 22373 40471 22431 40477
rect 14691 40412 15240 40440
rect 15304 40412 15516 40440
rect 15749 40443 15807 40449
rect 14691 40409 14703 40412
rect 14645 40403 14703 40409
rect 15304 40384 15332 40412
rect 15749 40409 15761 40443
rect 15795 40409 15807 40443
rect 15749 40403 15807 40409
rect 14734 40372 14740 40384
rect 14476 40344 14740 40372
rect 14734 40332 14740 40344
rect 14792 40332 14798 40384
rect 15286 40332 15292 40384
rect 15344 40332 15350 40384
rect 15764 40372 15792 40403
rect 19426 40400 19432 40452
rect 19484 40440 19490 40452
rect 19705 40443 19763 40449
rect 19705 40440 19717 40443
rect 19484 40412 19717 40440
rect 19484 40400 19490 40412
rect 19705 40409 19717 40412
rect 19751 40409 19763 40443
rect 21174 40440 21180 40452
rect 20930 40412 21180 40440
rect 19705 40403 19763 40409
rect 21174 40400 21180 40412
rect 21232 40400 21238 40452
rect 21453 40443 21511 40449
rect 21453 40409 21465 40443
rect 21499 40409 21511 40443
rect 22388 40440 22416 40471
rect 22462 40468 22468 40520
rect 22520 40508 22526 40520
rect 22664 40517 22692 40548
rect 22557 40511 22615 40517
rect 22557 40508 22569 40511
rect 22520 40480 22569 40508
rect 22520 40468 22526 40480
rect 22557 40477 22569 40480
rect 22603 40477 22615 40511
rect 22557 40471 22615 40477
rect 22649 40511 22707 40517
rect 22649 40477 22661 40511
rect 22695 40477 22707 40511
rect 22649 40471 22707 40477
rect 22833 40511 22891 40517
rect 22833 40477 22845 40511
rect 22879 40508 22891 40511
rect 24210 40508 24216 40520
rect 22879 40480 24216 40508
rect 22879 40477 22891 40480
rect 22833 40471 22891 40477
rect 24210 40468 24216 40480
rect 24268 40468 24274 40520
rect 22741 40443 22799 40449
rect 22741 40440 22753 40443
rect 22388 40412 22753 40440
rect 21453 40403 21511 40409
rect 22741 40409 22753 40412
rect 22787 40409 22799 40443
rect 22741 40403 22799 40409
rect 15838 40372 15844 40384
rect 15764 40344 15844 40372
rect 15838 40332 15844 40344
rect 15896 40332 15902 40384
rect 16853 40375 16911 40381
rect 16853 40341 16865 40375
rect 16899 40372 16911 40375
rect 17405 40375 17463 40381
rect 17405 40372 17417 40375
rect 16899 40344 17417 40372
rect 16899 40341 16911 40344
rect 16853 40335 16911 40341
rect 17405 40341 17417 40344
rect 17451 40341 17463 40375
rect 17405 40335 17463 40341
rect 17494 40332 17500 40384
rect 17552 40332 17558 40384
rect 18322 40332 18328 40384
rect 18380 40332 18386 40384
rect 18693 40375 18751 40381
rect 18693 40341 18705 40375
rect 18739 40372 18751 40375
rect 20070 40372 20076 40384
rect 18739 40344 20076 40372
rect 18739 40341 18751 40344
rect 18693 40335 18751 40341
rect 20070 40332 20076 40344
rect 20128 40372 20134 40384
rect 21468 40372 21496 40403
rect 20128 40344 21496 40372
rect 20128 40332 20134 40344
rect 1104 40282 41400 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 41400 40282
rect 1104 40208 41400 40230
rect 9858 40168 9864 40180
rect 8220 40140 9864 40168
rect 8220 40112 8248 40140
rect 9858 40128 9864 40140
rect 9916 40128 9922 40180
rect 10342 40171 10400 40177
rect 10342 40137 10354 40171
rect 10388 40168 10400 40171
rect 10388 40140 10456 40168
rect 10388 40137 10400 40140
rect 10342 40131 10400 40137
rect 7466 40060 7472 40112
rect 7524 40060 7530 40112
rect 8202 40060 8208 40112
rect 8260 40060 8266 40112
rect 8665 40103 8723 40109
rect 8665 40100 8677 40103
rect 8312 40072 8677 40100
rect 7282 39992 7288 40044
rect 7340 40032 7346 40044
rect 8312 40032 8340 40072
rect 8665 40069 8677 40072
rect 8711 40069 8723 40103
rect 8665 40063 8723 40069
rect 10134 40060 10140 40112
rect 10192 40109 10198 40112
rect 10192 40103 10221 40109
rect 10209 40069 10221 40103
rect 10428 40100 10456 40140
rect 10502 40128 10508 40180
rect 10560 40128 10566 40180
rect 10594 40128 10600 40180
rect 10652 40168 10658 40180
rect 11146 40168 11152 40180
rect 10652 40140 11152 40168
rect 10652 40128 10658 40140
rect 11146 40128 11152 40140
rect 11204 40128 11210 40180
rect 11330 40128 11336 40180
rect 11388 40128 11394 40180
rect 14182 40168 14188 40180
rect 12912 40140 14188 40168
rect 10612 40100 10640 40128
rect 11054 40100 11060 40112
rect 10428 40072 10640 40100
rect 10704 40072 11060 40100
rect 10192 40063 10221 40069
rect 10192 40060 10198 40063
rect 7340 40004 8340 40032
rect 7340 39992 7346 40004
rect 8478 39992 8484 40044
rect 8536 39992 8542 40044
rect 9861 40035 9919 40041
rect 9861 40001 9873 40035
rect 9907 40001 9919 40035
rect 9861 39995 9919 40001
rect 2682 39924 2688 39976
rect 2740 39964 2746 39976
rect 8205 39967 8263 39973
rect 8205 39964 8217 39967
rect 2740 39936 8217 39964
rect 2740 39924 2746 39936
rect 8205 39933 8217 39936
rect 8251 39964 8263 39967
rect 8570 39964 8576 39976
rect 8251 39936 8576 39964
rect 8251 39933 8263 39936
rect 8205 39927 8263 39933
rect 8570 39924 8576 39936
rect 8628 39924 8634 39976
rect 9876 39964 9904 39995
rect 10042 39992 10048 40044
rect 10100 39992 10106 40044
rect 10597 40035 10655 40041
rect 10597 40001 10609 40035
rect 10643 40032 10655 40035
rect 10704 40032 10732 40072
rect 11054 40060 11060 40072
rect 11112 40060 11118 40112
rect 11348 40100 11376 40128
rect 11164 40072 11376 40100
rect 10643 40004 10732 40032
rect 10643 40001 10655 40004
rect 10597 39995 10655 40001
rect 10778 39992 10784 40044
rect 10836 40032 10842 40044
rect 11164 40041 11192 40072
rect 11422 40060 11428 40112
rect 11480 40100 11486 40112
rect 11480 40072 11744 40100
rect 11480 40060 11486 40072
rect 11716 40041 11744 40072
rect 11149 40035 11207 40041
rect 10836 40004 11100 40032
rect 10836 39992 10842 40004
rect 10134 39964 10140 39976
rect 9876 39936 10140 39964
rect 10134 39924 10140 39936
rect 10192 39924 10198 39976
rect 10410 39924 10416 39976
rect 10468 39964 10474 39976
rect 10965 39967 11023 39973
rect 10965 39964 10977 39967
rect 10468 39936 10977 39964
rect 10468 39924 10474 39936
rect 10965 39933 10977 39936
rect 11011 39933 11023 39967
rect 11072 39964 11100 40004
rect 11149 40001 11161 40035
rect 11195 40001 11207 40035
rect 11149 39995 11207 40001
rect 11333 40035 11391 40041
rect 11333 40001 11345 40035
rect 11379 40032 11391 40035
rect 11701 40035 11759 40041
rect 11379 40004 11652 40032
rect 11379 40001 11391 40004
rect 11333 39995 11391 40001
rect 11241 39967 11299 39973
rect 11241 39964 11253 39967
rect 11072 39936 11253 39964
rect 10965 39927 11023 39933
rect 11241 39933 11253 39936
rect 11287 39933 11299 39967
rect 11241 39927 11299 39933
rect 11514 39924 11520 39976
rect 11572 39924 11578 39976
rect 11624 39964 11652 40004
rect 11701 40001 11713 40035
rect 11747 40032 11759 40035
rect 12912 40032 12940 40140
rect 14182 40128 14188 40140
rect 14240 40128 14246 40180
rect 15838 40128 15844 40180
rect 15896 40168 15902 40180
rect 17037 40171 17095 40177
rect 17037 40168 17049 40171
rect 15896 40140 17049 40168
rect 15896 40128 15902 40140
rect 17037 40137 17049 40140
rect 17083 40137 17095 40171
rect 17037 40131 17095 40137
rect 19245 40171 19303 40177
rect 19245 40137 19257 40171
rect 19291 40168 19303 40171
rect 19426 40168 19432 40180
rect 19291 40140 19432 40168
rect 19291 40137 19303 40140
rect 19245 40131 19303 40137
rect 19426 40128 19432 40140
rect 19484 40128 19490 40180
rect 22925 40171 22983 40177
rect 22925 40137 22937 40171
rect 22971 40168 22983 40171
rect 22971 40140 23520 40168
rect 22971 40137 22983 40140
rect 22925 40131 22983 40137
rect 13906 40060 13912 40112
rect 13964 40060 13970 40112
rect 15378 40060 15384 40112
rect 15436 40100 15442 40112
rect 15562 40100 15568 40112
rect 15436 40072 15568 40100
rect 15436 40060 15442 40072
rect 15562 40060 15568 40072
rect 15620 40060 15626 40112
rect 15856 40100 15884 40128
rect 15764 40072 15884 40100
rect 11747 40004 12940 40032
rect 11747 40001 11759 40004
rect 11701 39995 11759 40001
rect 15010 39992 15016 40044
rect 15068 39992 15074 40044
rect 15286 39992 15292 40044
rect 15344 39992 15350 40044
rect 15470 39992 15476 40044
rect 15528 39992 15534 40044
rect 15764 40041 15792 40072
rect 16206 40060 16212 40112
rect 16264 40060 16270 40112
rect 19334 40060 19340 40112
rect 19392 40100 19398 40112
rect 23492 40109 23520 40140
rect 24946 40128 24952 40180
rect 25004 40168 25010 40180
rect 40770 40168 40776 40180
rect 25004 40140 40776 40168
rect 25004 40128 25010 40140
rect 40770 40128 40776 40140
rect 40828 40128 40834 40180
rect 19981 40103 20039 40109
rect 19981 40100 19993 40103
rect 19392 40072 19993 40100
rect 19392 40060 19398 40072
rect 19981 40069 19993 40072
rect 20027 40069 20039 40103
rect 19981 40063 20039 40069
rect 23477 40103 23535 40109
rect 23477 40069 23489 40103
rect 23523 40069 23535 40103
rect 23477 40063 23535 40069
rect 23566 40060 23572 40112
rect 23624 40100 23630 40112
rect 23624 40072 23966 40100
rect 23624 40060 23630 40072
rect 15657 40035 15715 40041
rect 15657 40001 15669 40035
rect 15703 40001 15715 40035
rect 15657 39995 15715 40001
rect 15749 40035 15807 40041
rect 15749 40001 15761 40035
rect 15795 40001 15807 40035
rect 15749 39995 15807 40001
rect 11882 39964 11888 39976
rect 11624 39936 11888 39964
rect 11882 39924 11888 39936
rect 11940 39924 11946 39976
rect 12897 39967 12955 39973
rect 12897 39964 12909 39967
rect 12636 39936 12909 39964
rect 8588 39896 8616 39924
rect 10870 39896 10876 39908
rect 8588 39868 10876 39896
rect 10870 39856 10876 39868
rect 10928 39896 10934 39908
rect 12636 39896 12664 39936
rect 12897 39933 12909 39936
rect 12943 39933 12955 39967
rect 12897 39927 12955 39933
rect 13170 39924 13176 39976
rect 13228 39924 13234 39976
rect 14734 39924 14740 39976
rect 14792 39964 14798 39976
rect 14921 39967 14979 39973
rect 14921 39964 14933 39967
rect 14792 39936 14933 39964
rect 14792 39924 14798 39936
rect 14921 39933 14933 39936
rect 14967 39933 14979 39967
rect 15028 39964 15056 39992
rect 15672 39964 15700 39995
rect 15838 39992 15844 40044
rect 15896 40032 15902 40044
rect 16853 40035 16911 40041
rect 16853 40032 16865 40035
rect 15896 40004 16865 40032
rect 15896 39992 15902 40004
rect 16853 40001 16865 40004
rect 16899 40001 16911 40035
rect 16853 39995 16911 40001
rect 18874 39992 18880 40044
rect 18932 39992 18938 40044
rect 22002 39992 22008 40044
rect 22060 39992 22066 40044
rect 23106 39992 23112 40044
rect 23164 39992 23170 40044
rect 15028 39936 15700 39964
rect 14921 39927 14979 39933
rect 16666 39924 16672 39976
rect 16724 39964 16730 39976
rect 17402 39964 17408 39976
rect 16724 39936 17408 39964
rect 16724 39924 16730 39936
rect 17402 39924 17408 39936
rect 17460 39964 17466 39976
rect 18046 39964 18052 39976
rect 17460 39936 18052 39964
rect 17460 39924 17466 39936
rect 18046 39924 18052 39936
rect 18104 39924 18110 39976
rect 18322 39924 18328 39976
rect 18380 39964 18386 39976
rect 18785 39967 18843 39973
rect 18785 39964 18797 39967
rect 18380 39936 18797 39964
rect 18380 39924 18386 39936
rect 18785 39933 18797 39936
rect 18831 39933 18843 39967
rect 18785 39927 18843 39933
rect 20714 39924 20720 39976
rect 20772 39964 20778 39976
rect 21818 39964 21824 39976
rect 20772 39936 21824 39964
rect 20772 39924 20778 39936
rect 21818 39924 21824 39936
rect 21876 39964 21882 39976
rect 23201 39967 23259 39973
rect 23201 39964 23213 39967
rect 21876 39936 23213 39964
rect 21876 39924 21882 39936
rect 23201 39933 23213 39936
rect 23247 39933 23259 39967
rect 23201 39927 23259 39933
rect 10928 39868 12664 39896
rect 10928 39856 10934 39868
rect 12636 39840 12664 39868
rect 15654 39856 15660 39908
rect 15712 39896 15718 39908
rect 15841 39899 15899 39905
rect 15841 39896 15853 39899
rect 15712 39868 15853 39896
rect 15712 39856 15718 39868
rect 15841 39865 15853 39868
rect 15887 39865 15899 39899
rect 15841 39859 15899 39865
rect 8110 39788 8116 39840
rect 8168 39828 8174 39840
rect 8849 39831 8907 39837
rect 8849 39828 8861 39831
rect 8168 39800 8861 39828
rect 8168 39788 8174 39800
rect 8849 39797 8861 39800
rect 8895 39797 8907 39831
rect 8849 39791 8907 39797
rect 9953 39831 10011 39837
rect 9953 39797 9965 39831
rect 9999 39828 10011 39831
rect 10321 39831 10379 39837
rect 10321 39828 10333 39831
rect 9999 39800 10333 39828
rect 9999 39797 10011 39800
rect 9953 39791 10011 39797
rect 10321 39797 10333 39800
rect 10367 39797 10379 39831
rect 10321 39791 10379 39797
rect 12618 39788 12624 39840
rect 12676 39788 12682 39840
rect 12710 39788 12716 39840
rect 12768 39828 12774 39840
rect 15105 39831 15163 39837
rect 15105 39828 15117 39831
rect 12768 39800 15117 39828
rect 12768 39788 12774 39800
rect 15105 39797 15117 39800
rect 15151 39797 15163 39831
rect 15105 39791 15163 39797
rect 15930 39788 15936 39840
rect 15988 39828 15994 39840
rect 16209 39831 16267 39837
rect 16209 39828 16221 39831
rect 15988 39800 16221 39828
rect 15988 39788 15994 39800
rect 16209 39797 16221 39800
rect 16255 39797 16267 39831
rect 16209 39791 16267 39797
rect 16390 39788 16396 39840
rect 16448 39788 16454 39840
rect 21818 39788 21824 39840
rect 21876 39788 21882 39840
rect 1104 39738 41400 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 41400 39738
rect 1104 39664 41400 39686
rect 7374 39584 7380 39636
rect 7432 39624 7438 39636
rect 8202 39624 8208 39636
rect 7432 39596 8208 39624
rect 7432 39584 7438 39596
rect 8202 39584 8208 39596
rect 8260 39584 8266 39636
rect 8570 39584 8576 39636
rect 8628 39584 8634 39636
rect 8662 39584 8668 39636
rect 8720 39624 8726 39636
rect 11057 39627 11115 39633
rect 11057 39624 11069 39627
rect 8720 39596 11069 39624
rect 8720 39584 8726 39596
rect 11057 39593 11069 39596
rect 11103 39593 11115 39627
rect 11057 39587 11115 39593
rect 11238 39584 11244 39636
rect 11296 39624 11302 39636
rect 12894 39624 12900 39636
rect 11296 39596 12900 39624
rect 11296 39584 11302 39596
rect 12894 39584 12900 39596
rect 12952 39584 12958 39636
rect 13170 39584 13176 39636
rect 13228 39624 13234 39636
rect 13449 39627 13507 39633
rect 13449 39624 13461 39627
rect 13228 39596 13461 39624
rect 13228 39584 13234 39596
rect 13449 39593 13461 39596
rect 13495 39593 13507 39627
rect 13449 39587 13507 39593
rect 15010 39584 15016 39636
rect 15068 39624 15074 39636
rect 15105 39627 15163 39633
rect 15105 39624 15117 39627
rect 15068 39596 15117 39624
rect 15068 39584 15074 39596
rect 15105 39593 15117 39596
rect 15151 39593 15163 39627
rect 15105 39587 15163 39593
rect 15749 39627 15807 39633
rect 15749 39593 15761 39627
rect 15795 39624 15807 39627
rect 16206 39624 16212 39636
rect 15795 39596 16212 39624
rect 15795 39593 15807 39596
rect 15749 39587 15807 39593
rect 16206 39584 16212 39596
rect 16264 39584 16270 39636
rect 23017 39627 23075 39633
rect 16500 39596 22784 39624
rect 1486 39448 1492 39500
rect 1544 39488 1550 39500
rect 3789 39491 3847 39497
rect 3789 39488 3801 39491
rect 1544 39460 3801 39488
rect 1544 39448 1550 39460
rect 3789 39457 3801 39460
rect 3835 39488 3847 39491
rect 4062 39488 4068 39500
rect 3835 39460 4068 39488
rect 3835 39457 3847 39460
rect 3789 39451 3847 39457
rect 4062 39448 4068 39460
rect 4120 39448 4126 39500
rect 7282 39448 7288 39500
rect 7340 39488 7346 39500
rect 7377 39491 7435 39497
rect 7377 39488 7389 39491
rect 7340 39460 7389 39488
rect 7340 39448 7346 39460
rect 7377 39457 7389 39460
rect 7423 39457 7435 39491
rect 8478 39488 8484 39500
rect 7377 39451 7435 39457
rect 7668 39460 8484 39488
rect 7561 39423 7619 39429
rect 7561 39389 7573 39423
rect 7607 39422 7619 39423
rect 7668 39422 7696 39460
rect 8478 39448 8484 39460
rect 8536 39448 8542 39500
rect 8588 39488 8616 39584
rect 11790 39516 11796 39568
rect 11848 39516 11854 39568
rect 12710 39516 12716 39568
rect 12768 39516 12774 39568
rect 15194 39516 15200 39568
rect 15252 39556 15258 39568
rect 16500 39556 16528 39596
rect 15252 39528 16528 39556
rect 15252 39516 15258 39528
rect 8941 39491 8999 39497
rect 8941 39488 8953 39491
rect 8588 39460 8953 39488
rect 8941 39457 8953 39460
rect 8987 39457 8999 39491
rect 8941 39451 8999 39457
rect 9214 39448 9220 39500
rect 9272 39448 9278 39500
rect 9582 39448 9588 39500
rect 9640 39488 9646 39500
rect 9640 39460 10732 39488
rect 9640 39448 9646 39460
rect 7607 39394 7696 39422
rect 7607 39389 7619 39394
rect 7561 39383 7619 39389
rect 7834 39380 7840 39432
rect 7892 39380 7898 39432
rect 7944 39392 8340 39420
rect 5718 39312 5724 39364
rect 5776 39352 5782 39364
rect 7944 39352 7972 39392
rect 5776 39324 7972 39352
rect 5776 39312 5782 39324
rect 8110 39312 8116 39364
rect 8168 39352 8174 39364
rect 8205 39355 8263 39361
rect 8205 39352 8217 39355
rect 8168 39324 8217 39352
rect 8168 39312 8174 39324
rect 8205 39321 8217 39324
rect 8251 39321 8263 39355
rect 8312 39352 8340 39392
rect 9674 39352 9680 39364
rect 8312 39324 9680 39352
rect 8205 39315 8263 39321
rect 9674 39312 9680 39324
rect 9732 39312 9738 39364
rect 10704 39352 10732 39460
rect 10796 39460 11468 39488
rect 10796 39432 10824 39460
rect 10778 39380 10784 39432
rect 10836 39380 10842 39432
rect 11238 39380 11244 39432
rect 11296 39380 11302 39432
rect 11440 39429 11468 39460
rect 11882 39448 11888 39500
rect 11940 39448 11946 39500
rect 11425 39423 11483 39429
rect 11425 39389 11437 39423
rect 11471 39389 11483 39423
rect 11425 39383 11483 39389
rect 10965 39355 11023 39361
rect 10965 39352 10977 39355
rect 10704 39324 10977 39352
rect 10965 39321 10977 39324
rect 11011 39321 11023 39355
rect 10965 39315 11023 39321
rect 11054 39312 11060 39364
rect 11112 39352 11118 39364
rect 11333 39355 11391 39361
rect 11333 39352 11345 39355
rect 11112 39324 11345 39352
rect 11112 39312 11118 39324
rect 11333 39321 11345 39324
rect 11379 39321 11391 39355
rect 11440 39352 11468 39383
rect 11606 39380 11612 39432
rect 11664 39380 11670 39432
rect 11701 39423 11759 39429
rect 11701 39389 11713 39423
rect 11747 39420 11759 39423
rect 11793 39423 11851 39429
rect 11793 39420 11805 39423
rect 11747 39392 11805 39420
rect 11747 39389 11759 39392
rect 11701 39383 11759 39389
rect 11793 39389 11805 39392
rect 11839 39420 11851 39423
rect 11900 39420 11928 39448
rect 11839 39392 11928 39420
rect 12069 39423 12127 39429
rect 11839 39389 11851 39392
rect 11793 39383 11851 39389
rect 12069 39389 12081 39423
rect 12115 39420 12127 39423
rect 12728 39420 12756 39516
rect 16390 39488 16396 39500
rect 12820 39460 16396 39488
rect 12820 39429 12848 39460
rect 16390 39448 16396 39460
rect 16448 39448 16454 39500
rect 21453 39491 21511 39497
rect 21453 39457 21465 39491
rect 21499 39488 21511 39491
rect 21818 39488 21824 39500
rect 21499 39460 21824 39488
rect 21499 39457 21511 39460
rect 21453 39451 21511 39457
rect 21818 39448 21824 39460
rect 21876 39448 21882 39500
rect 22756 39488 22784 39596
rect 23017 39593 23029 39627
rect 23063 39624 23075 39627
rect 23106 39624 23112 39636
rect 23063 39596 23112 39624
rect 23063 39593 23075 39596
rect 23017 39587 23075 39593
rect 23106 39584 23112 39596
rect 23164 39584 23170 39636
rect 22830 39516 22836 39568
rect 22888 39556 22894 39568
rect 22888 39528 23612 39556
rect 22888 39516 22894 39528
rect 23584 39497 23612 39528
rect 23477 39491 23535 39497
rect 23477 39488 23489 39491
rect 22756 39460 23489 39488
rect 23477 39457 23489 39460
rect 23523 39457 23535 39491
rect 23477 39451 23535 39457
rect 23569 39491 23627 39497
rect 23569 39457 23581 39491
rect 23615 39457 23627 39491
rect 23569 39451 23627 39457
rect 25869 39491 25927 39497
rect 25869 39457 25881 39491
rect 25915 39488 25927 39491
rect 26142 39488 26148 39500
rect 25915 39460 26148 39488
rect 25915 39457 25927 39460
rect 25869 39451 25927 39457
rect 26142 39448 26148 39460
rect 26200 39448 26206 39500
rect 12115 39392 12756 39420
rect 12805 39423 12863 39429
rect 12115 39389 12127 39392
rect 12069 39383 12127 39389
rect 12805 39389 12817 39423
rect 12851 39389 12863 39423
rect 12805 39383 12863 39389
rect 11977 39355 12035 39361
rect 11977 39352 11989 39355
rect 11440 39324 11989 39352
rect 11333 39315 11391 39321
rect 11977 39321 11989 39324
rect 12023 39321 12035 39355
rect 11977 39315 12035 39321
rect 4433 39287 4491 39293
rect 4433 39253 4445 39287
rect 4479 39284 4491 39287
rect 4614 39284 4620 39296
rect 4479 39256 4620 39284
rect 4479 39253 4491 39256
rect 4433 39247 4491 39253
rect 4614 39244 4620 39256
rect 4672 39244 4678 39296
rect 7006 39244 7012 39296
rect 7064 39284 7070 39296
rect 7745 39287 7803 39293
rect 7745 39284 7757 39287
rect 7064 39256 7757 39284
rect 7064 39244 7070 39256
rect 7745 39253 7757 39256
rect 7791 39284 7803 39287
rect 7834 39284 7840 39296
rect 7791 39256 7840 39284
rect 7791 39253 7803 39256
rect 7745 39247 7803 39253
rect 7834 39244 7840 39256
rect 7892 39244 7898 39296
rect 8386 39244 8392 39296
rect 8444 39244 8450 39296
rect 8478 39244 8484 39296
rect 8536 39284 8542 39296
rect 9950 39284 9956 39296
rect 8536 39256 9956 39284
rect 8536 39244 8542 39256
rect 9950 39244 9956 39256
rect 10008 39244 10014 39296
rect 10134 39244 10140 39296
rect 10192 39284 10198 39296
rect 11072 39284 11100 39312
rect 10192 39256 11100 39284
rect 11348 39284 11376 39315
rect 12084 39284 12112 39383
rect 12894 39380 12900 39432
rect 12952 39420 12958 39432
rect 12952 39392 12997 39420
rect 12952 39380 12958 39392
rect 13262 39380 13268 39432
rect 13320 39429 13326 39432
rect 13320 39420 13328 39429
rect 13320 39392 13365 39420
rect 13320 39383 13328 39392
rect 13320 39380 13326 39383
rect 14734 39380 14740 39432
rect 14792 39380 14798 39432
rect 14921 39423 14979 39429
rect 14921 39389 14933 39423
rect 14967 39389 14979 39423
rect 14921 39383 14979 39389
rect 13078 39312 13084 39364
rect 13136 39312 13142 39364
rect 13173 39355 13231 39361
rect 13173 39321 13185 39355
rect 13219 39352 13231 39355
rect 14752 39352 14780 39380
rect 13219 39324 14780 39352
rect 13219 39321 13231 39324
rect 13173 39315 13231 39321
rect 11348 39256 12112 39284
rect 10192 39244 10198 39256
rect 12986 39244 12992 39296
rect 13044 39284 13050 39296
rect 13188 39284 13216 39315
rect 13044 39256 13216 39284
rect 13044 39244 13050 39256
rect 14182 39244 14188 39296
rect 14240 39284 14246 39296
rect 14936 39284 14964 39383
rect 15470 39380 15476 39432
rect 15528 39420 15534 39432
rect 16209 39423 16267 39429
rect 16209 39420 16221 39423
rect 15528 39392 16221 39420
rect 15528 39380 15534 39392
rect 16209 39389 16221 39392
rect 16255 39389 16267 39423
rect 16209 39383 16267 39389
rect 16666 39380 16672 39432
rect 16724 39380 16730 39432
rect 17218 39380 17224 39432
rect 17276 39420 17282 39432
rect 18049 39423 18107 39429
rect 18049 39420 18061 39423
rect 17276 39392 18061 39420
rect 17276 39380 17282 39392
rect 18049 39389 18061 39392
rect 18095 39389 18107 39423
rect 18049 39383 18107 39389
rect 20162 39380 20168 39432
rect 20220 39420 20226 39432
rect 20714 39420 20720 39432
rect 20220 39392 20720 39420
rect 20220 39380 20226 39392
rect 20714 39380 20720 39392
rect 20772 39420 20778 39432
rect 21177 39423 21235 39429
rect 21177 39420 21189 39423
rect 20772 39392 21189 39420
rect 20772 39380 20778 39392
rect 21177 39389 21189 39392
rect 21223 39389 21235 39423
rect 21177 39383 21235 39389
rect 23385 39423 23443 39429
rect 23385 39389 23397 39423
rect 23431 39420 23443 39423
rect 24946 39420 24952 39432
rect 23431 39392 24952 39420
rect 23431 39389 23443 39392
rect 23385 39383 23443 39389
rect 24946 39380 24952 39392
rect 25004 39380 25010 39432
rect 15286 39312 15292 39364
rect 15344 39352 15350 39364
rect 15381 39355 15439 39361
rect 15381 39352 15393 39355
rect 15344 39324 15393 39352
rect 15344 39312 15350 39324
rect 15381 39321 15393 39324
rect 15427 39321 15439 39355
rect 15381 39315 15439 39321
rect 15562 39312 15568 39364
rect 15620 39312 15626 39364
rect 15838 39312 15844 39364
rect 15896 39312 15902 39364
rect 16025 39355 16083 39361
rect 16025 39321 16037 39355
rect 16071 39352 16083 39355
rect 16684 39352 16712 39380
rect 16071 39324 16712 39352
rect 22678 39324 23428 39352
rect 16071 39321 16083 39324
rect 16025 39315 16083 39321
rect 15856 39284 15884 39312
rect 23400 39296 23428 39324
rect 26050 39312 26056 39364
rect 26108 39352 26114 39364
rect 26145 39355 26203 39361
rect 26145 39352 26157 39355
rect 26108 39324 26157 39352
rect 26108 39312 26114 39324
rect 26145 39321 26157 39324
rect 26191 39321 26203 39355
rect 27706 39352 27712 39364
rect 27370 39324 27712 39352
rect 26145 39315 26203 39321
rect 27706 39312 27712 39324
rect 27764 39312 27770 39364
rect 14240 39256 15884 39284
rect 17865 39287 17923 39293
rect 14240 39244 14246 39256
rect 17865 39253 17877 39287
rect 17911 39284 17923 39287
rect 18230 39284 18236 39296
rect 17911 39256 18236 39284
rect 17911 39253 17923 39256
rect 17865 39247 17923 39253
rect 18230 39244 18236 39256
rect 18288 39244 18294 39296
rect 18782 39244 18788 39296
rect 18840 39284 18846 39296
rect 20622 39284 20628 39296
rect 18840 39256 20628 39284
rect 18840 39244 18846 39256
rect 20622 39244 20628 39256
rect 20680 39244 20686 39296
rect 22922 39244 22928 39296
rect 22980 39244 22986 39296
rect 23382 39244 23388 39296
rect 23440 39244 23446 39296
rect 27617 39287 27675 39293
rect 27617 39253 27629 39287
rect 27663 39284 27675 39287
rect 27798 39284 27804 39296
rect 27663 39256 27804 39284
rect 27663 39253 27675 39256
rect 27617 39247 27675 39253
rect 27798 39244 27804 39256
rect 27856 39244 27862 39296
rect 1104 39194 41400 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 41400 39194
rect 1104 39120 41400 39142
rect 3602 39040 3608 39092
rect 3660 39080 3666 39092
rect 3660 39052 3924 39080
rect 3660 39040 3666 39052
rect 3896 39012 3924 39052
rect 4062 39040 4068 39092
rect 4120 39040 4126 39092
rect 4356 39052 5580 39080
rect 4356 39012 4384 39052
rect 3818 38984 4384 39012
rect 4433 39015 4491 39021
rect 4433 38981 4445 39015
rect 4479 39012 4491 39015
rect 4706 39012 4712 39024
rect 4479 38984 4712 39012
rect 4479 38981 4491 38984
rect 4433 38975 4491 38981
rect 4706 38972 4712 38984
rect 4764 38972 4770 39024
rect 5552 38944 5580 39052
rect 7282 39040 7288 39092
rect 7340 39080 7346 39092
rect 7340 39052 7972 39080
rect 7340 39040 7346 39052
rect 7193 39015 7251 39021
rect 7193 38981 7205 39015
rect 7239 39012 7251 39015
rect 7239 38984 7604 39012
rect 7239 38981 7251 38984
rect 7193 38975 7251 38981
rect 5718 38944 5724 38956
rect 5552 38930 5724 38944
rect 5566 38916 5724 38930
rect 5718 38904 5724 38916
rect 5776 38904 5782 38956
rect 7006 38904 7012 38956
rect 7064 38904 7070 38956
rect 7576 38953 7604 38984
rect 7285 38947 7343 38953
rect 7285 38913 7297 38947
rect 7331 38913 7343 38947
rect 7285 38907 7343 38913
rect 7561 38947 7619 38953
rect 7561 38913 7573 38947
rect 7607 38944 7619 38947
rect 7607 38916 7880 38944
rect 7607 38913 7619 38916
rect 7561 38907 7619 38913
rect 1762 38836 1768 38888
rect 1820 38876 1826 38888
rect 2317 38879 2375 38885
rect 2317 38876 2329 38879
rect 1820 38848 2329 38876
rect 1820 38836 1826 38848
rect 2317 38845 2329 38848
rect 2363 38845 2375 38879
rect 2317 38839 2375 38845
rect 2593 38879 2651 38885
rect 2593 38845 2605 38879
rect 2639 38876 2651 38879
rect 3050 38876 3056 38888
rect 2639 38848 3056 38876
rect 2639 38845 2651 38848
rect 2593 38839 2651 38845
rect 2332 38740 2360 38839
rect 3050 38836 3056 38848
rect 3108 38836 3114 38888
rect 4157 38879 4215 38885
rect 4157 38845 4169 38879
rect 4203 38845 4215 38879
rect 4157 38839 4215 38845
rect 6181 38879 6239 38885
rect 6181 38845 6193 38879
rect 6227 38876 6239 38879
rect 6454 38876 6460 38888
rect 6227 38848 6460 38876
rect 6227 38845 6239 38848
rect 6181 38839 6239 38845
rect 4172 38808 4200 38839
rect 6454 38836 6460 38848
rect 6512 38836 6518 38888
rect 7300 38876 7328 38907
rect 7653 38879 7711 38885
rect 7653 38876 7665 38879
rect 7300 38848 7665 38876
rect 7653 38845 7665 38848
rect 7699 38845 7711 38879
rect 7653 38839 7711 38845
rect 3620 38780 4200 38808
rect 2682 38740 2688 38752
rect 2332 38712 2688 38740
rect 2682 38700 2688 38712
rect 2740 38740 2746 38752
rect 3620 38740 3648 38780
rect 2740 38712 3648 38740
rect 2740 38700 2746 38712
rect 6730 38700 6736 38752
rect 6788 38740 6794 38752
rect 6825 38743 6883 38749
rect 6825 38740 6837 38743
rect 6788 38712 6837 38740
rect 6788 38700 6794 38712
rect 6825 38709 6837 38712
rect 6871 38709 6883 38743
rect 7668 38740 7696 38839
rect 7852 38808 7880 38916
rect 7944 38885 7972 39052
rect 8386 39040 8392 39092
rect 8444 39040 8450 39092
rect 9033 39083 9091 39089
rect 9033 39049 9045 39083
rect 9079 39080 9091 39083
rect 9214 39080 9220 39092
rect 9079 39052 9220 39080
rect 9079 39049 9091 39052
rect 9033 39043 9091 39049
rect 9214 39040 9220 39052
rect 9272 39040 9278 39092
rect 11238 39040 11244 39092
rect 11296 39040 11302 39092
rect 11790 39040 11796 39092
rect 11848 39040 11854 39092
rect 12894 39040 12900 39092
rect 12952 39080 12958 39092
rect 16574 39080 16580 39092
rect 12952 39052 16580 39080
rect 12952 39040 12958 39052
rect 16574 39040 16580 39052
rect 16632 39040 16638 39092
rect 17218 39040 17224 39092
rect 17276 39040 17282 39092
rect 17589 39083 17647 39089
rect 17589 39049 17601 39083
rect 17635 39080 17647 39083
rect 17954 39080 17960 39092
rect 17635 39052 17960 39080
rect 17635 39049 17647 39052
rect 17589 39043 17647 39049
rect 17954 39040 17960 39052
rect 18012 39040 18018 39092
rect 20162 39080 20168 39092
rect 18064 39052 20168 39080
rect 8404 38953 8432 39040
rect 8757 39015 8815 39021
rect 8757 38981 8769 39015
rect 8803 39012 8815 39015
rect 11422 39012 11428 39024
rect 8803 38984 9628 39012
rect 8803 38981 8815 38984
rect 8757 38975 8815 38981
rect 8389 38947 8447 38953
rect 8389 38913 8401 38947
rect 8435 38913 8447 38947
rect 8389 38907 8447 38913
rect 8478 38904 8484 38956
rect 8536 38944 8542 38956
rect 8536 38916 8581 38944
rect 8536 38904 8542 38916
rect 8662 38904 8668 38956
rect 8720 38904 8726 38956
rect 7929 38879 7987 38885
rect 7929 38845 7941 38879
rect 7975 38845 7987 38879
rect 7929 38839 7987 38845
rect 8772 38808 8800 38975
rect 9600 38956 9628 38984
rect 10888 38984 11428 39012
rect 8846 38904 8852 38956
rect 8904 38953 8910 38956
rect 8904 38944 8912 38953
rect 8904 38916 8949 38944
rect 8904 38907 8912 38916
rect 8904 38904 8910 38907
rect 9582 38904 9588 38956
rect 9640 38904 9646 38956
rect 10778 38904 10784 38956
rect 10836 38944 10842 38956
rect 10888 38953 10916 38984
rect 11422 38972 11428 38984
rect 11480 38972 11486 39024
rect 10873 38947 10931 38953
rect 10873 38944 10885 38947
rect 10836 38916 10885 38944
rect 10836 38904 10842 38916
rect 10873 38913 10885 38916
rect 10919 38913 10931 38947
rect 10873 38907 10931 38913
rect 11057 38947 11115 38953
rect 11057 38913 11069 38947
rect 11103 38944 11115 38947
rect 11330 38944 11336 38956
rect 11103 38916 11336 38944
rect 11103 38913 11115 38916
rect 11057 38907 11115 38913
rect 11330 38904 11336 38916
rect 11388 38904 11394 38956
rect 11698 38904 11704 38956
rect 11756 38904 11762 38956
rect 11808 38885 11836 39040
rect 12986 39012 12992 39024
rect 12406 38984 12992 39012
rect 11793 38879 11851 38885
rect 11793 38845 11805 38879
rect 11839 38845 11851 38879
rect 12406 38876 12434 38984
rect 12986 38972 12992 38984
rect 13044 38972 13050 39024
rect 17681 39015 17739 39021
rect 17681 39012 17693 39015
rect 14384 38984 17693 39012
rect 12618 38904 12624 38956
rect 12676 38904 12682 38956
rect 13906 38904 13912 38956
rect 13964 38944 13970 38956
rect 13964 38916 14030 38944
rect 13964 38904 13970 38916
rect 14384 38888 14412 38984
rect 17681 38981 17693 38984
rect 17727 39012 17739 39015
rect 17727 38984 18000 39012
rect 17727 38981 17739 38984
rect 17681 38975 17739 38981
rect 11793 38839 11851 38845
rect 11900 38848 12434 38876
rect 11900 38808 11928 38848
rect 12894 38836 12900 38888
rect 12952 38836 12958 38888
rect 14366 38836 14372 38888
rect 14424 38836 14430 38888
rect 14645 38879 14703 38885
rect 14645 38845 14657 38879
rect 14691 38876 14703 38879
rect 14829 38879 14887 38885
rect 14829 38876 14841 38879
rect 14691 38848 14841 38876
rect 14691 38845 14703 38848
rect 14645 38839 14703 38845
rect 14829 38845 14841 38848
rect 14875 38876 14887 38879
rect 15470 38876 15476 38888
rect 14875 38848 15476 38876
rect 14875 38845 14887 38848
rect 14829 38839 14887 38845
rect 7852 38780 8800 38808
rect 8864 38780 11928 38808
rect 12069 38811 12127 38817
rect 8202 38740 8208 38752
rect 7668 38712 8208 38740
rect 6825 38703 6883 38709
rect 8202 38700 8208 38712
rect 8260 38700 8266 38752
rect 8478 38700 8484 38752
rect 8536 38740 8542 38752
rect 8864 38740 8892 38780
rect 12069 38777 12081 38811
rect 12115 38808 12127 38811
rect 12250 38808 12256 38820
rect 12115 38780 12256 38808
rect 12115 38777 12127 38780
rect 12069 38771 12127 38777
rect 12250 38768 12256 38780
rect 12308 38768 12314 38820
rect 8536 38712 8892 38740
rect 8536 38700 8542 38712
rect 11330 38700 11336 38752
rect 11388 38740 11394 38752
rect 14660 38740 14688 38839
rect 15470 38836 15476 38848
rect 15528 38836 15534 38888
rect 17310 38836 17316 38888
rect 17368 38876 17374 38888
rect 17586 38876 17592 38888
rect 17368 38848 17592 38876
rect 17368 38836 17374 38848
rect 17586 38836 17592 38848
rect 17644 38876 17650 38888
rect 17773 38879 17831 38885
rect 17773 38876 17785 38879
rect 17644 38848 17785 38876
rect 17644 38836 17650 38848
rect 17773 38845 17785 38848
rect 17819 38845 17831 38879
rect 17972 38876 18000 38984
rect 18064 38953 18092 39052
rect 20162 39040 20168 39052
rect 20220 39040 20226 39092
rect 21637 39083 21695 39089
rect 21637 39049 21649 39083
rect 21683 39080 21695 39083
rect 22002 39080 22008 39092
rect 21683 39052 22008 39080
rect 21683 39049 21695 39052
rect 21637 39043 21695 39049
rect 22002 39040 22008 39052
rect 22060 39040 22066 39092
rect 22922 39040 22928 39092
rect 22980 39040 22986 39092
rect 26050 39040 26056 39092
rect 26108 39080 26114 39092
rect 26145 39083 26203 39089
rect 26145 39080 26157 39083
rect 26108 39052 26157 39080
rect 26108 39040 26114 39052
rect 26145 39049 26157 39052
rect 26191 39049 26203 39083
rect 26145 39043 26203 39049
rect 18230 38972 18236 39024
rect 18288 39012 18294 39024
rect 18325 39015 18383 39021
rect 18325 39012 18337 39015
rect 18288 38984 18337 39012
rect 18288 38972 18294 38984
rect 18325 38981 18337 38984
rect 18371 38981 18383 39015
rect 18325 38975 18383 38981
rect 18782 38972 18788 39024
rect 18840 38972 18846 39024
rect 21177 39015 21235 39021
rect 21177 38981 21189 39015
rect 21223 39012 21235 39015
rect 22940 39012 22968 39040
rect 21223 38984 22968 39012
rect 21223 38981 21235 38984
rect 21177 38975 21235 38981
rect 18049 38947 18107 38953
rect 18049 38913 18061 38947
rect 18095 38913 18107 38947
rect 18049 38907 18107 38913
rect 22002 38904 22008 38956
rect 22060 38944 22066 38956
rect 22940 38953 22968 38984
rect 25869 39015 25927 39021
rect 25869 38981 25881 39015
rect 25915 39012 25927 39015
rect 27617 39015 27675 39021
rect 27617 39012 27629 39015
rect 25915 38984 27629 39012
rect 25915 38981 25927 38984
rect 25869 38975 25927 38981
rect 27617 38981 27629 38984
rect 27663 38981 27675 39015
rect 27617 38975 27675 38981
rect 22097 38947 22155 38953
rect 22097 38944 22109 38947
rect 22060 38916 22109 38944
rect 22060 38904 22066 38916
rect 22097 38913 22109 38916
rect 22143 38944 22155 38947
rect 22741 38947 22799 38953
rect 22741 38944 22753 38947
rect 22143 38916 22753 38944
rect 22143 38913 22155 38916
rect 22097 38907 22155 38913
rect 22741 38913 22753 38916
rect 22787 38913 22799 38947
rect 22741 38907 22799 38913
rect 22925 38947 22983 38953
rect 22925 38913 22937 38947
rect 22971 38913 22983 38947
rect 22925 38907 22983 38913
rect 25590 38904 25596 38956
rect 25648 38904 25654 38956
rect 25774 38904 25780 38956
rect 25832 38904 25838 38956
rect 25961 38947 26019 38953
rect 25961 38913 25973 38947
rect 26007 38944 26019 38947
rect 26050 38944 26056 38956
rect 26007 38916 26056 38944
rect 26007 38913 26019 38916
rect 25961 38907 26019 38913
rect 26050 38904 26056 38916
rect 26108 38904 26114 38956
rect 27065 38947 27123 38953
rect 27065 38913 27077 38947
rect 27111 38944 27123 38947
rect 27798 38944 27804 38956
rect 27111 38916 27804 38944
rect 27111 38913 27123 38916
rect 27065 38907 27123 38913
rect 27798 38904 27804 38916
rect 27856 38904 27862 38956
rect 20073 38879 20131 38885
rect 20073 38876 20085 38879
rect 17972 38848 20085 38876
rect 17773 38839 17831 38845
rect 19444 38820 19472 38848
rect 20073 38845 20085 38848
rect 20119 38845 20131 38879
rect 22649 38879 22707 38885
rect 22649 38876 22661 38879
rect 20073 38839 20131 38845
rect 22388 38848 22661 38876
rect 19426 38768 19432 38820
rect 19484 38768 19490 38820
rect 21545 38811 21603 38817
rect 21545 38777 21557 38811
rect 21591 38808 21603 38811
rect 22388 38808 22416 38848
rect 22649 38845 22661 38848
rect 22695 38845 22707 38879
rect 22649 38839 22707 38845
rect 21591 38780 22416 38808
rect 22572 38780 23060 38808
rect 21591 38777 21603 38780
rect 21545 38771 21603 38777
rect 11388 38712 14688 38740
rect 11388 38700 11394 38712
rect 15378 38700 15384 38752
rect 15436 38700 15442 38752
rect 20898 38700 20904 38752
rect 20956 38740 20962 38752
rect 22572 38740 22600 38780
rect 23032 38749 23060 38780
rect 20956 38712 22600 38740
rect 23017 38743 23075 38749
rect 20956 38700 20962 38712
rect 23017 38709 23029 38743
rect 23063 38709 23075 38743
rect 23017 38703 23075 38709
rect 1104 38650 41400 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 41400 38650
rect 1104 38576 41400 38598
rect 3050 38496 3056 38548
rect 3108 38536 3114 38548
rect 3421 38539 3479 38545
rect 3421 38536 3433 38539
rect 3108 38508 3433 38536
rect 3108 38496 3114 38508
rect 3421 38505 3433 38508
rect 3467 38505 3479 38539
rect 3421 38499 3479 38505
rect 4706 38496 4712 38548
rect 4764 38496 4770 38548
rect 6546 38496 6552 38548
rect 6604 38496 6610 38548
rect 6730 38496 6736 38548
rect 6788 38536 6794 38548
rect 7561 38539 7619 38545
rect 7561 38536 7573 38539
rect 6788 38508 7573 38536
rect 6788 38496 6794 38508
rect 7561 38505 7573 38508
rect 7607 38505 7619 38539
rect 11333 38539 11391 38545
rect 7561 38499 7619 38505
rect 7668 38508 8064 38536
rect 5261 38471 5319 38477
rect 5261 38437 5273 38471
rect 5307 38437 5319 38471
rect 7668 38468 7696 38508
rect 8036 38480 8064 38508
rect 11333 38505 11345 38539
rect 11379 38536 11391 38539
rect 11698 38536 11704 38548
rect 11379 38508 11704 38536
rect 11379 38505 11391 38508
rect 11333 38499 11391 38505
rect 11698 38496 11704 38508
rect 11756 38496 11762 38548
rect 12621 38539 12679 38545
rect 12621 38505 12633 38539
rect 12667 38536 12679 38539
rect 12894 38536 12900 38548
rect 12667 38508 12900 38536
rect 12667 38505 12679 38508
rect 12621 38499 12679 38505
rect 12894 38496 12900 38508
rect 12952 38496 12958 38548
rect 17954 38496 17960 38548
rect 18012 38536 18018 38548
rect 18049 38539 18107 38545
rect 18049 38536 18061 38539
rect 18012 38508 18061 38536
rect 18012 38496 18018 38508
rect 18049 38505 18061 38508
rect 18095 38505 18107 38539
rect 18049 38499 18107 38505
rect 22002 38496 22008 38548
rect 22060 38496 22066 38548
rect 23198 38496 23204 38548
rect 23256 38536 23262 38548
rect 27614 38536 27620 38548
rect 23256 38508 27620 38536
rect 23256 38496 23262 38508
rect 27614 38496 27620 38508
rect 27672 38496 27678 38548
rect 5261 38431 5319 38437
rect 5920 38440 7696 38468
rect 7837 38471 7895 38477
rect 4433 38403 4491 38409
rect 4433 38369 4445 38403
rect 4479 38400 4491 38403
rect 4479 38372 4844 38400
rect 4479 38369 4491 38372
rect 4433 38363 4491 38369
rect 3605 38335 3663 38341
rect 3605 38301 3617 38335
rect 3651 38332 3663 38335
rect 4157 38335 4215 38341
rect 3651 38304 3832 38332
rect 3651 38301 3663 38304
rect 3605 38295 3663 38301
rect 3804 38205 3832 38304
rect 4157 38301 4169 38335
rect 4203 38332 4215 38335
rect 4614 38332 4620 38344
rect 4203 38304 4620 38332
rect 4203 38301 4215 38304
rect 4157 38295 4215 38301
rect 4614 38292 4620 38304
rect 4672 38292 4678 38344
rect 4816 38264 4844 38372
rect 4893 38335 4951 38341
rect 4893 38301 4905 38335
rect 4939 38332 4951 38335
rect 5276 38332 5304 38431
rect 5350 38360 5356 38412
rect 5408 38400 5414 38412
rect 5920 38409 5948 38440
rect 7837 38437 7849 38471
rect 7883 38437 7895 38471
rect 7837 38431 7895 38437
rect 5905 38403 5963 38409
rect 5905 38400 5917 38403
rect 5408 38372 5917 38400
rect 5408 38360 5414 38372
rect 5905 38369 5917 38372
rect 5951 38369 5963 38403
rect 6730 38400 6736 38412
rect 5905 38363 5963 38369
rect 6288 38372 6736 38400
rect 6288 38341 6316 38372
rect 6730 38360 6736 38372
rect 6788 38360 6794 38412
rect 6822 38360 6828 38412
rect 6880 38400 6886 38412
rect 7101 38403 7159 38409
rect 7101 38400 7113 38403
rect 6880 38372 7113 38400
rect 6880 38360 6886 38372
rect 7101 38369 7113 38372
rect 7147 38369 7159 38403
rect 7101 38363 7159 38369
rect 7193 38403 7251 38409
rect 7193 38369 7205 38403
rect 7239 38400 7251 38403
rect 7852 38400 7880 38431
rect 8018 38428 8024 38480
rect 8076 38428 8082 38480
rect 11241 38471 11299 38477
rect 11241 38437 11253 38471
rect 11287 38468 11299 38471
rect 11606 38468 11612 38480
rect 11287 38440 11612 38468
rect 11287 38437 11299 38440
rect 11241 38431 11299 38437
rect 9398 38400 9404 38412
rect 7239 38372 7880 38400
rect 7944 38372 9404 38400
rect 7239 38369 7251 38372
rect 7193 38363 7251 38369
rect 4939 38304 5304 38332
rect 6273 38335 6331 38341
rect 4939 38301 4951 38304
rect 4893 38295 4951 38301
rect 6273 38301 6285 38335
rect 6319 38301 6331 38335
rect 6273 38295 6331 38301
rect 6638 38292 6644 38344
rect 6696 38332 6702 38344
rect 6696 38304 7052 38332
rect 6696 38292 6702 38304
rect 5629 38267 5687 38273
rect 4816 38236 5580 38264
rect 5552 38208 5580 38236
rect 5629 38233 5641 38267
rect 5675 38264 5687 38267
rect 5675 38236 6960 38264
rect 5675 38233 5687 38236
rect 5629 38227 5687 38233
rect 3789 38199 3847 38205
rect 3789 38165 3801 38199
rect 3835 38165 3847 38199
rect 3789 38159 3847 38165
rect 4249 38199 4307 38205
rect 4249 38165 4261 38199
rect 4295 38196 4307 38199
rect 4614 38196 4620 38208
rect 4295 38168 4620 38196
rect 4295 38165 4307 38168
rect 4249 38159 4307 38165
rect 4614 38156 4620 38168
rect 4672 38156 4678 38208
rect 5534 38156 5540 38208
rect 5592 38156 5598 38208
rect 5721 38199 5779 38205
rect 5721 38165 5733 38199
rect 5767 38196 5779 38199
rect 6454 38196 6460 38208
rect 5767 38168 6460 38196
rect 5767 38165 5779 38168
rect 5721 38159 5779 38165
rect 6454 38156 6460 38168
rect 6512 38156 6518 38208
rect 6822 38156 6828 38208
rect 6880 38156 6886 38208
rect 6932 38205 6960 38236
rect 6917 38199 6975 38205
rect 6917 38165 6929 38199
rect 6963 38165 6975 38199
rect 7024 38196 7052 38304
rect 7282 38292 7288 38344
rect 7340 38292 7346 38344
rect 7377 38335 7435 38341
rect 7377 38301 7389 38335
rect 7423 38301 7435 38335
rect 7377 38295 7435 38301
rect 7392 38264 7420 38295
rect 7742 38292 7748 38344
rect 7800 38332 7806 38344
rect 7837 38335 7895 38341
rect 7837 38332 7849 38335
rect 7800 38304 7849 38332
rect 7800 38292 7806 38304
rect 7837 38301 7849 38304
rect 7883 38301 7895 38335
rect 7837 38295 7895 38301
rect 7944 38264 7972 38372
rect 9398 38360 9404 38372
rect 9456 38360 9462 38412
rect 10873 38403 10931 38409
rect 10873 38369 10885 38403
rect 10919 38400 10931 38403
rect 10919 38372 11284 38400
rect 10919 38369 10931 38372
rect 10873 38363 10931 38369
rect 11256 38344 11284 38372
rect 8021 38335 8079 38341
rect 8021 38301 8033 38335
rect 8067 38301 8079 38335
rect 8021 38295 8079 38301
rect 7392 38236 7972 38264
rect 8036 38196 8064 38295
rect 8202 38292 8208 38344
rect 8260 38332 8266 38344
rect 11054 38332 11060 38344
rect 8260 38304 11060 38332
rect 8260 38292 8266 38304
rect 11054 38292 11060 38304
rect 11112 38292 11118 38344
rect 11146 38292 11152 38344
rect 11204 38292 11210 38344
rect 11238 38292 11244 38344
rect 11296 38292 11302 38344
rect 11348 38341 11376 38440
rect 11606 38428 11612 38440
rect 11664 38428 11670 38480
rect 14826 38428 14832 38480
rect 14884 38468 14890 38480
rect 14884 38440 19334 38468
rect 14884 38428 14890 38440
rect 15930 38400 15936 38412
rect 12406 38372 15936 38400
rect 11333 38335 11391 38341
rect 11333 38301 11345 38335
rect 11379 38301 11391 38335
rect 11333 38295 11391 38301
rect 11514 38292 11520 38344
rect 11572 38292 11578 38344
rect 11974 38292 11980 38344
rect 12032 38292 12038 38344
rect 12070 38335 12128 38341
rect 12070 38301 12082 38335
rect 12116 38332 12128 38335
rect 12406 38332 12434 38372
rect 15930 38360 15936 38372
rect 15988 38360 15994 38412
rect 16574 38360 16580 38412
rect 16632 38400 16638 38412
rect 19306 38400 19334 38440
rect 22462 38400 22468 38412
rect 16632 38372 17540 38400
rect 19306 38372 22468 38400
rect 16632 38360 16638 38372
rect 12116 38304 12434 38332
rect 12483 38335 12541 38341
rect 12116 38301 12128 38304
rect 12070 38295 12128 38301
rect 12483 38301 12495 38335
rect 12529 38332 12541 38335
rect 13262 38332 13268 38344
rect 12529 38304 13268 38332
rect 12529 38301 12541 38304
rect 12483 38295 12541 38301
rect 11164 38264 11192 38292
rect 12084 38264 12112 38295
rect 13262 38292 13268 38304
rect 13320 38332 13326 38344
rect 14458 38332 14464 38344
rect 13320 38304 14464 38332
rect 13320 38292 13326 38304
rect 14458 38292 14464 38304
rect 14516 38292 14522 38344
rect 17034 38292 17040 38344
rect 17092 38292 17098 38344
rect 17512 38341 17540 38372
rect 22462 38360 22468 38372
rect 22520 38360 22526 38412
rect 24673 38403 24731 38409
rect 24673 38369 24685 38403
rect 24719 38400 24731 38403
rect 24946 38400 24952 38412
rect 24719 38372 24952 38400
rect 24719 38369 24731 38372
rect 24673 38363 24731 38369
rect 24946 38360 24952 38372
rect 25004 38400 25010 38412
rect 26142 38400 26148 38412
rect 25004 38372 26148 38400
rect 25004 38360 25010 38372
rect 26142 38360 26148 38372
rect 26200 38360 26206 38412
rect 26252 38372 29132 38400
rect 17129 38335 17187 38341
rect 17129 38301 17141 38335
rect 17175 38332 17187 38335
rect 17497 38335 17555 38341
rect 17175 38304 17448 38332
rect 17175 38301 17187 38304
rect 17129 38295 17187 38301
rect 11164 38236 12112 38264
rect 12250 38224 12256 38276
rect 12308 38224 12314 38276
rect 12345 38267 12403 38273
rect 12345 38233 12357 38267
rect 12391 38264 12403 38267
rect 15378 38264 15384 38276
rect 12391 38236 15384 38264
rect 12391 38233 12403 38236
rect 12345 38227 12403 38233
rect 15378 38224 15384 38236
rect 15436 38224 15442 38276
rect 7024 38168 8064 38196
rect 6917 38159 6975 38165
rect 14274 38156 14280 38208
rect 14332 38196 14338 38208
rect 17310 38196 17316 38208
rect 14332 38168 17316 38196
rect 14332 38156 14338 38168
rect 17310 38156 17316 38168
rect 17368 38156 17374 38208
rect 17420 38196 17448 38304
rect 17497 38301 17509 38335
rect 17543 38332 17555 38335
rect 17586 38332 17592 38344
rect 17543 38304 17592 38332
rect 17543 38301 17555 38304
rect 17497 38295 17555 38301
rect 17586 38292 17592 38304
rect 17644 38292 17650 38344
rect 17865 38335 17923 38341
rect 17865 38301 17877 38335
rect 17911 38332 17923 38335
rect 18138 38332 18144 38344
rect 17911 38304 18144 38332
rect 17911 38301 17923 38304
rect 17865 38295 17923 38301
rect 18138 38292 18144 38304
rect 18196 38292 18202 38344
rect 20162 38292 20168 38344
rect 20220 38332 20226 38344
rect 20257 38335 20315 38341
rect 20257 38332 20269 38335
rect 20220 38304 20269 38332
rect 20220 38292 20226 38304
rect 20257 38301 20269 38304
rect 20303 38301 20315 38335
rect 26252 38332 26280 38372
rect 26082 38318 26280 38332
rect 20257 38295 20315 38301
rect 26068 38304 26280 38318
rect 27617 38335 27675 38341
rect 17678 38224 17684 38276
rect 17736 38224 17742 38276
rect 17770 38224 17776 38276
rect 17828 38224 17834 38276
rect 20533 38267 20591 38273
rect 20533 38233 20545 38267
rect 20579 38233 20591 38267
rect 20533 38227 20591 38233
rect 18598 38196 18604 38208
rect 17420 38168 18604 38196
rect 18598 38156 18604 38168
rect 18656 38156 18662 38208
rect 20346 38156 20352 38208
rect 20404 38196 20410 38208
rect 20548 38196 20576 38227
rect 20622 38224 20628 38276
rect 20680 38264 20686 38276
rect 20990 38264 20996 38276
rect 20680 38236 20996 38264
rect 20680 38224 20686 38236
rect 20990 38224 20996 38236
rect 21048 38224 21054 38276
rect 24949 38267 25007 38273
rect 24949 38233 24961 38267
rect 24995 38264 25007 38267
rect 25038 38264 25044 38276
rect 24995 38236 25044 38264
rect 24995 38233 25007 38236
rect 24949 38227 25007 38233
rect 25038 38224 25044 38236
rect 25096 38224 25102 38276
rect 20404 38168 20576 38196
rect 20404 38156 20410 38168
rect 23382 38156 23388 38208
rect 23440 38196 23446 38208
rect 25314 38196 25320 38208
rect 23440 38168 25320 38196
rect 23440 38156 23446 38168
rect 25314 38156 25320 38168
rect 25372 38196 25378 38208
rect 26068 38196 26096 38304
rect 27617 38301 27629 38335
rect 27663 38301 27675 38335
rect 27617 38295 27675 38301
rect 27632 38264 27660 38295
rect 27632 38236 27844 38264
rect 27816 38208 27844 38236
rect 27890 38224 27896 38276
rect 27948 38224 27954 38276
rect 29104 38264 29132 38372
rect 31202 38264 31208 38276
rect 29104 38250 31208 38264
rect 29118 38236 31208 38250
rect 31202 38224 31208 38236
rect 31260 38224 31266 38276
rect 25372 38168 26096 38196
rect 25372 38156 25378 38168
rect 26418 38156 26424 38208
rect 26476 38156 26482 38208
rect 27798 38156 27804 38208
rect 27856 38156 27862 38208
rect 29365 38199 29423 38205
rect 29365 38165 29377 38199
rect 29411 38196 29423 38199
rect 30006 38196 30012 38208
rect 29411 38168 30012 38196
rect 29411 38165 29423 38168
rect 29365 38159 29423 38165
rect 30006 38156 30012 38168
rect 30064 38156 30070 38208
rect 1104 38106 41400 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 41400 38106
rect 1104 38032 41400 38054
rect 6457 37995 6515 38001
rect 6457 37961 6469 37995
rect 6503 37992 6515 37995
rect 6638 37992 6644 38004
rect 6503 37964 6644 37992
rect 6503 37961 6515 37964
rect 6457 37955 6515 37961
rect 6638 37952 6644 37964
rect 6696 37952 6702 38004
rect 8110 37992 8116 38004
rect 6748 37964 8116 37992
rect 6748 37924 6776 37964
rect 8110 37952 8116 37964
rect 8168 37952 8174 38004
rect 9309 37995 9367 38001
rect 9309 37992 9321 37995
rect 9232 37964 9321 37992
rect 6380 37896 6776 37924
rect 7837 37927 7895 37933
rect 6270 37816 6276 37868
rect 6328 37856 6334 37868
rect 6380 37865 6408 37896
rect 7837 37893 7849 37927
rect 7883 37924 7895 37927
rect 8202 37924 8208 37936
rect 7883 37896 8208 37924
rect 7883 37893 7895 37896
rect 7837 37887 7895 37893
rect 6365 37859 6423 37865
rect 6365 37856 6377 37859
rect 6328 37828 6377 37856
rect 6328 37816 6334 37828
rect 6365 37825 6377 37828
rect 6411 37825 6423 37859
rect 6365 37819 6423 37825
rect 6454 37816 6460 37868
rect 6512 37856 6518 37868
rect 6549 37859 6607 37865
rect 6549 37856 6561 37859
rect 6512 37828 6561 37856
rect 6512 37816 6518 37828
rect 6549 37825 6561 37828
rect 6595 37825 6607 37859
rect 6549 37819 6607 37825
rect 6564 37788 6592 37819
rect 6730 37816 6736 37868
rect 6788 37856 6794 37868
rect 6917 37859 6975 37865
rect 6917 37856 6929 37859
rect 6788 37828 6929 37856
rect 6788 37816 6794 37828
rect 6917 37825 6929 37828
rect 6963 37825 6975 37859
rect 6917 37819 6975 37825
rect 7006 37816 7012 37868
rect 7064 37856 7070 37868
rect 7101 37859 7159 37865
rect 7101 37856 7113 37859
rect 7064 37828 7113 37856
rect 7064 37816 7070 37828
rect 7101 37825 7113 37828
rect 7147 37856 7159 37859
rect 7469 37859 7527 37865
rect 7469 37856 7481 37859
rect 7147 37828 7481 37856
rect 7147 37825 7159 37828
rect 7101 37819 7159 37825
rect 7469 37825 7481 37828
rect 7515 37856 7527 37859
rect 7852 37856 7880 37887
rect 8202 37884 8208 37896
rect 8260 37884 8266 37936
rect 7515 37828 7880 37856
rect 7515 37825 7527 37828
rect 7469 37819 7527 37825
rect 8938 37816 8944 37868
rect 8996 37816 9002 37868
rect 9232 37856 9260 37964
rect 9309 37961 9321 37964
rect 9355 37961 9367 37995
rect 9309 37955 9367 37961
rect 9398 37952 9404 38004
rect 9456 37992 9462 38004
rect 9493 37995 9551 38001
rect 9493 37992 9505 37995
rect 9456 37964 9505 37992
rect 9456 37952 9462 37964
rect 9493 37961 9505 37964
rect 9539 37961 9551 37995
rect 9493 37955 9551 37961
rect 10965 37995 11023 38001
rect 10965 37961 10977 37995
rect 11011 37992 11023 37995
rect 11054 37992 11060 38004
rect 11011 37964 11060 37992
rect 11011 37961 11023 37964
rect 10965 37955 11023 37961
rect 11054 37952 11060 37964
rect 11112 37952 11118 38004
rect 11609 37995 11667 38001
rect 11609 37961 11621 37995
rect 11655 37992 11667 37995
rect 11974 37992 11980 38004
rect 11655 37964 11980 37992
rect 11655 37961 11667 37964
rect 11609 37955 11667 37961
rect 11974 37952 11980 37964
rect 12032 37952 12038 38004
rect 15838 37952 15844 38004
rect 15896 37992 15902 38004
rect 16117 37995 16175 38001
rect 16117 37992 16129 37995
rect 15896 37964 16129 37992
rect 15896 37952 15902 37964
rect 16117 37961 16129 37964
rect 16163 37961 16175 37995
rect 16117 37955 16175 37961
rect 17770 37952 17776 38004
rect 17828 37992 17834 38004
rect 18049 37995 18107 38001
rect 18049 37992 18061 37995
rect 17828 37964 18061 37992
rect 17828 37952 17834 37964
rect 18049 37961 18061 37964
rect 18095 37961 18107 37995
rect 18049 37955 18107 37961
rect 18138 37952 18144 38004
rect 18196 37952 18202 38004
rect 24946 37992 24952 38004
rect 23768 37964 24952 37992
rect 11330 37884 11336 37936
rect 11388 37924 11394 37936
rect 16022 37924 16028 37936
rect 11388 37896 16028 37924
rect 11388 37884 11394 37896
rect 16022 37884 16028 37896
rect 16080 37884 16086 37936
rect 17034 37884 17040 37936
rect 17092 37924 17098 37936
rect 17862 37924 17868 37936
rect 17092 37896 17868 37924
rect 17092 37884 17098 37896
rect 17862 37884 17868 37896
rect 17920 37924 17926 37936
rect 18877 37927 18935 37933
rect 17920 37896 18644 37924
rect 17920 37884 17926 37896
rect 9401 37859 9459 37865
rect 9401 37856 9413 37859
rect 9232 37828 9413 37856
rect 9401 37825 9413 37828
rect 9447 37825 9459 37859
rect 9401 37819 9459 37825
rect 9490 37816 9496 37868
rect 9548 37856 9554 37868
rect 9585 37859 9643 37865
rect 9585 37856 9597 37859
rect 9548 37828 9597 37856
rect 9548 37816 9554 37828
rect 9585 37825 9597 37828
rect 9631 37856 9643 37859
rect 9631 37828 9812 37856
rect 9631 37825 9643 37828
rect 9585 37819 9643 37825
rect 7193 37791 7251 37797
rect 7193 37788 7205 37791
rect 6564 37760 7205 37788
rect 7193 37757 7205 37760
rect 7239 37788 7251 37791
rect 7285 37791 7343 37797
rect 7285 37788 7297 37791
rect 7239 37760 7297 37788
rect 7239 37757 7251 37760
rect 7193 37751 7251 37757
rect 7285 37757 7297 37760
rect 7331 37788 7343 37791
rect 9033 37791 9091 37797
rect 7331 37760 8432 37788
rect 7331 37757 7343 37760
rect 7285 37751 7343 37757
rect 8404 37720 8432 37760
rect 9033 37757 9045 37791
rect 9079 37788 9091 37791
rect 9674 37788 9680 37800
rect 9079 37760 9680 37788
rect 9079 37757 9091 37760
rect 9033 37751 9091 37757
rect 9674 37748 9680 37760
rect 9732 37748 9738 37800
rect 9784 37788 9812 37828
rect 10778 37816 10784 37868
rect 10836 37816 10842 37868
rect 11054 37816 11060 37868
rect 11112 37856 11118 37868
rect 11517 37859 11575 37865
rect 11517 37856 11529 37859
rect 11112 37828 11529 37856
rect 11112 37816 11118 37828
rect 11517 37825 11529 37828
rect 11563 37825 11575 37859
rect 11517 37819 11575 37825
rect 11701 37859 11759 37865
rect 11701 37825 11713 37859
rect 11747 37856 11759 37859
rect 13722 37856 13728 37868
rect 11747 37828 13728 37856
rect 11747 37825 11759 37828
rect 11701 37819 11759 37825
rect 11716 37788 11744 37819
rect 13722 37816 13728 37828
rect 13780 37816 13786 37868
rect 14550 37816 14556 37868
rect 14608 37816 14614 37868
rect 14734 37816 14740 37868
rect 14792 37816 14798 37868
rect 15933 37859 15991 37865
rect 15933 37825 15945 37859
rect 15979 37856 15991 37859
rect 16482 37856 16488 37868
rect 15979 37828 16488 37856
rect 15979 37825 15991 37828
rect 15933 37819 15991 37825
rect 16482 37816 16488 37828
rect 16540 37816 16546 37868
rect 17773 37859 17831 37865
rect 17773 37825 17785 37859
rect 17819 37856 17831 37859
rect 18325 37859 18383 37865
rect 18325 37856 18337 37859
rect 17819 37828 18337 37856
rect 17819 37825 17831 37828
rect 17773 37819 17831 37825
rect 18325 37825 18337 37828
rect 18371 37856 18383 37859
rect 18506 37856 18512 37868
rect 18371 37828 18512 37856
rect 18371 37825 18383 37828
rect 18325 37819 18383 37825
rect 18506 37816 18512 37828
rect 18564 37816 18570 37868
rect 18616 37865 18644 37896
rect 18877 37893 18889 37927
rect 18923 37924 18935 37927
rect 19058 37924 19064 37936
rect 18923 37896 19064 37924
rect 18923 37893 18935 37896
rect 18877 37887 18935 37893
rect 19058 37884 19064 37896
rect 19116 37924 19122 37936
rect 19797 37927 19855 37933
rect 19797 37924 19809 37927
rect 19116 37896 19809 37924
rect 19116 37884 19122 37896
rect 19797 37893 19809 37896
rect 19843 37893 19855 37927
rect 19797 37887 19855 37893
rect 22020 37896 23520 37924
rect 22020 37868 22048 37896
rect 23492 37868 23520 37896
rect 18601 37859 18659 37865
rect 18601 37825 18613 37859
rect 18647 37825 18659 37859
rect 18601 37819 18659 37825
rect 19518 37816 19524 37868
rect 19576 37856 19582 37868
rect 19613 37859 19671 37865
rect 19613 37856 19625 37859
rect 19576 37828 19625 37856
rect 19576 37816 19582 37828
rect 19613 37825 19625 37828
rect 19659 37825 19671 37859
rect 19613 37819 19671 37825
rect 20809 37859 20867 37865
rect 20809 37825 20821 37859
rect 20855 37825 20867 37859
rect 20809 37819 20867 37825
rect 21913 37859 21971 37865
rect 21913 37825 21925 37859
rect 21959 37825 21971 37859
rect 21913 37819 21971 37825
rect 9784 37760 11744 37788
rect 18049 37791 18107 37797
rect 18049 37757 18061 37791
rect 18095 37788 18107 37791
rect 18095 37760 18552 37788
rect 18095 37757 18107 37760
rect 18049 37751 18107 37757
rect 12986 37720 12992 37732
rect 8404 37692 12992 37720
rect 12986 37680 12992 37692
rect 13044 37680 13050 37732
rect 17865 37723 17923 37729
rect 17865 37689 17877 37723
rect 17911 37720 17923 37723
rect 18322 37720 18328 37732
rect 17911 37692 18328 37720
rect 17911 37689 17923 37692
rect 17865 37683 17923 37689
rect 18322 37680 18328 37692
rect 18380 37720 18386 37732
rect 18524 37729 18552 37760
rect 19426 37748 19432 37800
rect 19484 37748 19490 37800
rect 20824 37788 20852 37819
rect 20898 37788 20904 37800
rect 20824 37760 20904 37788
rect 20898 37748 20904 37760
rect 20956 37748 20962 37800
rect 21928 37788 21956 37819
rect 22002 37816 22008 37868
rect 22060 37816 22066 37868
rect 22646 37816 22652 37868
rect 22704 37816 22710 37868
rect 23106 37816 23112 37868
rect 23164 37816 23170 37868
rect 23198 37816 23204 37868
rect 23256 37816 23262 37868
rect 23293 37859 23351 37865
rect 23293 37825 23305 37859
rect 23339 37825 23351 37859
rect 23293 37819 23351 37825
rect 23385 37859 23443 37865
rect 23385 37825 23397 37859
rect 23431 37825 23443 37859
rect 23385 37819 23443 37825
rect 23216 37788 23244 37816
rect 21928 37760 23244 37788
rect 18417 37723 18475 37729
rect 18417 37720 18429 37723
rect 18380 37692 18429 37720
rect 18380 37680 18386 37692
rect 18417 37689 18429 37692
rect 18463 37689 18475 37723
rect 18417 37683 18475 37689
rect 18509 37723 18567 37729
rect 18509 37689 18521 37723
rect 18555 37689 18567 37723
rect 18509 37683 18567 37689
rect 6730 37612 6736 37664
rect 6788 37612 6794 37664
rect 7098 37612 7104 37664
rect 7156 37652 7162 37664
rect 7653 37655 7711 37661
rect 7653 37652 7665 37655
rect 7156 37624 7665 37652
rect 7156 37612 7162 37624
rect 7653 37621 7665 37624
rect 7699 37652 7711 37655
rect 7742 37652 7748 37664
rect 7699 37624 7748 37652
rect 7699 37621 7711 37624
rect 7653 37615 7711 37621
rect 7742 37612 7748 37624
rect 7800 37612 7806 37664
rect 8110 37612 8116 37664
rect 8168 37652 8174 37664
rect 10410 37652 10416 37664
rect 8168 37624 10416 37652
rect 8168 37612 8174 37624
rect 10410 37612 10416 37624
rect 10468 37612 10474 37664
rect 14642 37612 14648 37664
rect 14700 37612 14706 37664
rect 16574 37612 16580 37664
rect 16632 37652 16638 37664
rect 17678 37652 17684 37664
rect 16632 37624 17684 37652
rect 16632 37612 16638 37624
rect 17678 37612 17684 37624
rect 17736 37612 17742 37664
rect 18524 37652 18552 37683
rect 19242 37680 19248 37732
rect 19300 37680 19306 37732
rect 22094 37680 22100 37732
rect 22152 37680 22158 37732
rect 19337 37655 19395 37661
rect 19337 37652 19349 37655
rect 18524 37624 19349 37652
rect 19337 37621 19349 37624
rect 19383 37621 19395 37655
rect 19337 37615 19395 37621
rect 20346 37612 20352 37664
rect 20404 37652 20410 37664
rect 20901 37655 20959 37661
rect 20901 37652 20913 37655
rect 20404 37624 20913 37652
rect 20404 37612 20410 37624
rect 20901 37621 20913 37624
rect 20947 37621 20959 37655
rect 20901 37615 20959 37621
rect 22370 37612 22376 37664
rect 22428 37652 22434 37664
rect 22465 37655 22523 37661
rect 22465 37652 22477 37655
rect 22428 37624 22477 37652
rect 22428 37612 22434 37624
rect 22465 37621 22477 37624
rect 22511 37621 22523 37655
rect 23308 37652 23336 37819
rect 23400 37788 23428 37819
rect 23474 37816 23480 37868
rect 23532 37816 23538 37868
rect 23566 37816 23572 37868
rect 23624 37816 23630 37868
rect 23768 37865 23796 37964
rect 24946 37952 24952 37964
rect 25004 37952 25010 38004
rect 25314 37952 25320 38004
rect 25372 37952 25378 38004
rect 25332 37924 25360 37952
rect 25254 37896 25360 37924
rect 25682 37884 25688 37936
rect 25740 37924 25746 37936
rect 25961 37927 26019 37933
rect 25961 37924 25973 37927
rect 25740 37896 25973 37924
rect 25740 37884 25746 37896
rect 25961 37893 25973 37896
rect 26007 37924 26019 37927
rect 26418 37924 26424 37936
rect 26007 37896 26424 37924
rect 26007 37893 26019 37896
rect 25961 37887 26019 37893
rect 26418 37884 26424 37896
rect 26476 37884 26482 37936
rect 27706 37884 27712 37936
rect 27764 37884 27770 37936
rect 23753 37859 23811 37865
rect 23753 37825 23765 37859
rect 23799 37825 23811 37859
rect 23753 37819 23811 37825
rect 23584 37788 23612 37816
rect 24029 37791 24087 37797
rect 24029 37788 24041 37791
rect 23400 37760 23612 37788
rect 23676 37760 24041 37788
rect 23676 37729 23704 37760
rect 24029 37757 24041 37760
rect 24075 37757 24087 37791
rect 24029 37751 24087 37757
rect 25498 37748 25504 37800
rect 25556 37788 25562 37800
rect 25777 37791 25835 37797
rect 25777 37788 25789 37791
rect 25556 37760 25789 37788
rect 25556 37748 25562 37760
rect 25777 37757 25789 37760
rect 25823 37757 25835 37791
rect 25777 37751 25835 37757
rect 26142 37748 26148 37800
rect 26200 37788 26206 37800
rect 26973 37791 27031 37797
rect 26973 37788 26985 37791
rect 26200 37760 26985 37788
rect 26200 37748 26206 37760
rect 26973 37757 26985 37760
rect 27019 37757 27031 37791
rect 26973 37751 27031 37757
rect 23661 37723 23719 37729
rect 23661 37689 23673 37723
rect 23707 37689 23719 37723
rect 23661 37683 23719 37689
rect 24578 37652 24584 37664
rect 23308 37624 24584 37652
rect 22465 37615 22523 37621
rect 24578 37612 24584 37624
rect 24636 37612 24642 37664
rect 24762 37612 24768 37664
rect 24820 37652 24826 37664
rect 25590 37652 25596 37664
rect 24820 37624 25596 37652
rect 24820 37612 24826 37624
rect 25590 37612 25596 37624
rect 25648 37652 25654 37664
rect 26053 37655 26111 37661
rect 26053 37652 26065 37655
rect 25648 37624 26065 37652
rect 25648 37612 25654 37624
rect 26053 37621 26065 37624
rect 26099 37621 26111 37655
rect 26988 37652 27016 37751
rect 27246 37748 27252 37800
rect 27304 37748 27310 37800
rect 27798 37652 27804 37664
rect 26988 37624 27804 37652
rect 26053 37615 26111 37621
rect 27798 37612 27804 37624
rect 27856 37612 27862 37664
rect 28721 37655 28779 37661
rect 28721 37621 28733 37655
rect 28767 37652 28779 37655
rect 29362 37652 29368 37664
rect 28767 37624 29368 37652
rect 28767 37621 28779 37624
rect 28721 37615 28779 37621
rect 29362 37612 29368 37624
rect 29420 37612 29426 37664
rect 1104 37562 41400 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 41400 37562
rect 1104 37488 41400 37510
rect 6546 37408 6552 37460
rect 6604 37408 6610 37460
rect 6730 37408 6736 37460
rect 6788 37448 6794 37460
rect 6825 37451 6883 37457
rect 6825 37448 6837 37451
rect 6788 37420 6837 37448
rect 6788 37408 6794 37420
rect 6825 37417 6837 37420
rect 6871 37417 6883 37451
rect 6825 37411 6883 37417
rect 7282 37408 7288 37460
rect 7340 37448 7346 37460
rect 7650 37448 7656 37460
rect 7340 37420 7656 37448
rect 7340 37408 7346 37420
rect 7650 37408 7656 37420
rect 7708 37448 7714 37460
rect 9490 37448 9496 37460
rect 7708 37420 9496 37448
rect 7708 37408 7714 37420
rect 9490 37408 9496 37420
rect 9548 37408 9554 37460
rect 10689 37451 10747 37457
rect 10689 37417 10701 37451
rect 10735 37448 10747 37451
rect 11054 37448 11060 37460
rect 10735 37420 11060 37448
rect 10735 37417 10747 37420
rect 10689 37411 10747 37417
rect 11054 37408 11060 37420
rect 11112 37408 11118 37460
rect 11149 37451 11207 37457
rect 11149 37417 11161 37451
rect 11195 37448 11207 37451
rect 11514 37448 11520 37460
rect 11195 37420 11520 37448
rect 11195 37417 11207 37420
rect 11149 37411 11207 37417
rect 11514 37408 11520 37420
rect 11572 37408 11578 37460
rect 14550 37408 14556 37460
rect 14608 37448 14614 37460
rect 14645 37451 14703 37457
rect 14645 37448 14657 37451
rect 14608 37420 14657 37448
rect 14608 37408 14614 37420
rect 14645 37417 14657 37420
rect 14691 37417 14703 37451
rect 15838 37448 15844 37460
rect 14645 37411 14703 37417
rect 15212 37420 15844 37448
rect 6564 37244 6592 37408
rect 8018 37340 8024 37392
rect 8076 37380 8082 37392
rect 14274 37380 14280 37392
rect 8076 37352 14280 37380
rect 8076 37340 8082 37352
rect 6914 37272 6920 37324
rect 6972 37312 6978 37324
rect 7009 37315 7067 37321
rect 7009 37312 7021 37315
rect 6972 37284 7021 37312
rect 6972 37272 6978 37284
rect 7009 37281 7021 37284
rect 7055 37281 7067 37315
rect 7009 37275 7067 37281
rect 10318 37272 10324 37324
rect 10376 37272 10382 37324
rect 13096 37321 13124 37352
rect 14274 37340 14280 37352
rect 14332 37340 14338 37392
rect 15212 37380 15240 37420
rect 15838 37408 15844 37420
rect 15896 37408 15902 37460
rect 17678 37408 17684 37460
rect 17736 37448 17742 37460
rect 18417 37451 18475 37457
rect 18417 37448 18429 37451
rect 17736 37420 18429 37448
rect 17736 37408 17742 37420
rect 18417 37417 18429 37420
rect 18463 37417 18475 37451
rect 18417 37411 18475 37417
rect 19242 37408 19248 37460
rect 19300 37448 19306 37460
rect 19613 37451 19671 37457
rect 19613 37448 19625 37451
rect 19300 37420 19625 37448
rect 19300 37408 19306 37420
rect 19613 37417 19625 37420
rect 19659 37417 19671 37451
rect 19613 37411 19671 37417
rect 23474 37408 23480 37460
rect 23532 37408 23538 37460
rect 26513 37451 26571 37457
rect 26513 37417 26525 37451
rect 26559 37448 26571 37451
rect 27246 37448 27252 37460
rect 26559 37420 27252 37448
rect 26559 37417 26571 37420
rect 26513 37411 26571 37417
rect 27246 37408 27252 37420
rect 27304 37408 27310 37460
rect 27890 37408 27896 37460
rect 27948 37408 27954 37460
rect 31941 37451 31999 37457
rect 31941 37448 31953 37451
rect 31726 37420 31953 37448
rect 14752 37352 15240 37380
rect 13081 37315 13139 37321
rect 13081 37281 13093 37315
rect 13127 37281 13139 37315
rect 14752 37312 14780 37352
rect 15286 37340 15292 37392
rect 15344 37340 15350 37392
rect 18156 37352 19380 37380
rect 13081 37275 13139 37281
rect 13832 37284 14780 37312
rect 6733 37247 6791 37253
rect 6733 37244 6745 37247
rect 6564 37216 6745 37244
rect 6733 37213 6745 37216
rect 6779 37244 6791 37247
rect 7098 37244 7104 37256
rect 6779 37216 7104 37244
rect 6779 37213 6791 37216
rect 6733 37207 6791 37213
rect 7098 37204 7104 37216
rect 7156 37204 7162 37256
rect 9950 37204 9956 37256
rect 10008 37244 10014 37256
rect 10413 37247 10471 37253
rect 10413 37244 10425 37247
rect 10008 37216 10425 37244
rect 10008 37204 10014 37216
rect 10413 37213 10425 37216
rect 10459 37213 10471 37247
rect 10413 37207 10471 37213
rect 10520 37216 10916 37244
rect 5534 37136 5540 37188
rect 5592 37176 5598 37188
rect 5592 37148 8340 37176
rect 5592 37136 5598 37148
rect 8312 37120 8340 37148
rect 7009 37111 7067 37117
rect 7009 37077 7021 37111
rect 7055 37108 7067 37111
rect 7190 37108 7196 37120
rect 7055 37080 7196 37108
rect 7055 37077 7067 37080
rect 7009 37071 7067 37077
rect 7190 37068 7196 37080
rect 7248 37068 7254 37120
rect 8294 37068 8300 37120
rect 8352 37068 8358 37120
rect 9030 37068 9036 37120
rect 9088 37108 9094 37120
rect 10520 37108 10548 37216
rect 10888 37176 10916 37216
rect 11054 37204 11060 37256
rect 11112 37244 11118 37256
rect 11149 37247 11207 37253
rect 11149 37244 11161 37247
rect 11112 37216 11161 37244
rect 11112 37204 11118 37216
rect 11149 37213 11161 37216
rect 11195 37213 11207 37247
rect 11149 37207 11207 37213
rect 11238 37204 11244 37256
rect 11296 37244 11302 37256
rect 11333 37247 11391 37253
rect 11333 37244 11345 37247
rect 11296 37216 11345 37244
rect 11296 37204 11302 37216
rect 11333 37213 11345 37216
rect 11379 37213 11391 37247
rect 12897 37247 12955 37253
rect 12897 37244 12909 37247
rect 11333 37207 11391 37213
rect 12406 37216 12909 37244
rect 12406 37176 12434 37216
rect 12897 37213 12909 37216
rect 12943 37213 12955 37247
rect 12897 37207 12955 37213
rect 13725 37247 13783 37253
rect 13725 37213 13737 37247
rect 13771 37244 13783 37247
rect 13832 37244 13860 37284
rect 13771 37216 13860 37244
rect 13909 37247 13967 37253
rect 13771 37213 13783 37216
rect 13725 37207 13783 37213
rect 13909 37213 13921 37247
rect 13955 37244 13967 37247
rect 14090 37244 14096 37256
rect 13955 37216 14096 37244
rect 13955 37213 13967 37216
rect 13909 37207 13967 37213
rect 10888 37148 12434 37176
rect 12912 37176 12940 37207
rect 13924 37176 13952 37207
rect 14090 37204 14096 37216
rect 14148 37244 14154 37256
rect 14752 37253 14780 37284
rect 14829 37315 14887 37321
rect 14829 37281 14841 37315
rect 14875 37312 14887 37315
rect 17037 37315 17095 37321
rect 17037 37312 17049 37315
rect 14875 37284 15516 37312
rect 14875 37281 14887 37284
rect 14829 37275 14887 37281
rect 15488 37253 15516 37284
rect 16408 37284 17049 37312
rect 14461 37247 14519 37253
rect 14461 37244 14473 37247
rect 14148 37216 14473 37244
rect 14148 37204 14154 37216
rect 14461 37213 14473 37216
rect 14507 37213 14519 37247
rect 14461 37207 14519 37213
rect 14737 37247 14795 37253
rect 14737 37213 14749 37247
rect 14783 37213 14795 37247
rect 14921 37247 14979 37253
rect 14921 37244 14933 37247
rect 14737 37207 14795 37213
rect 14844 37216 14933 37244
rect 12912 37148 13952 37176
rect 14274 37136 14280 37188
rect 14332 37136 14338 37188
rect 14476 37176 14504 37207
rect 14844 37176 14872 37216
rect 14921 37213 14933 37216
rect 14967 37213 14979 37247
rect 14921 37207 14979 37213
rect 15013 37247 15071 37253
rect 15013 37213 15025 37247
rect 15059 37213 15071 37247
rect 15013 37207 15071 37213
rect 15473 37247 15531 37253
rect 15473 37213 15485 37247
rect 15519 37213 15531 37247
rect 15473 37207 15531 37213
rect 15933 37247 15991 37253
rect 15933 37213 15945 37247
rect 15979 37213 15991 37247
rect 15933 37207 15991 37213
rect 15028 37176 15056 37207
rect 14476 37148 14872 37176
rect 14936 37148 15056 37176
rect 15948 37176 15976 37207
rect 16206 37204 16212 37256
rect 16264 37204 16270 37256
rect 16298 37204 16304 37256
rect 16356 37244 16362 37256
rect 16408 37253 16436 37284
rect 17037 37281 17049 37284
rect 17083 37281 17095 37315
rect 17037 37275 17095 37281
rect 16393 37247 16451 37253
rect 16393 37244 16405 37247
rect 16356 37216 16405 37244
rect 16356 37204 16362 37216
rect 16393 37213 16405 37216
rect 16439 37213 16451 37247
rect 16393 37207 16451 37213
rect 16482 37204 16488 37256
rect 16540 37244 16546 37256
rect 16945 37247 17003 37253
rect 16945 37244 16957 37247
rect 16540 37216 16957 37244
rect 16540 37204 16546 37216
rect 16945 37213 16957 37216
rect 16991 37244 17003 37247
rect 18156 37244 18184 37352
rect 18506 37272 18512 37324
rect 18564 37312 18570 37324
rect 18564 37284 19012 37312
rect 18564 37272 18570 37284
rect 16991 37216 18184 37244
rect 16991 37213 17003 37216
rect 16945 37207 17003 37213
rect 18230 37204 18236 37256
rect 18288 37244 18294 37256
rect 18984 37253 19012 37284
rect 19242 37272 19248 37324
rect 19300 37272 19306 37324
rect 18601 37247 18659 37253
rect 18601 37244 18613 37247
rect 18288 37216 18613 37244
rect 18288 37204 18294 37216
rect 18601 37213 18613 37216
rect 18647 37213 18659 37247
rect 18601 37207 18659 37213
rect 18969 37247 19027 37253
rect 18969 37213 18981 37247
rect 19015 37213 19027 37247
rect 18969 37207 19027 37213
rect 19058 37204 19064 37256
rect 19116 37204 19122 37256
rect 19260 37244 19288 37272
rect 19168 37216 19288 37244
rect 18693 37179 18751 37185
rect 18693 37176 18705 37179
rect 15948 37148 17356 37176
rect 9088 37080 10548 37108
rect 9088 37068 9094 37080
rect 12434 37068 12440 37120
rect 12492 37068 12498 37120
rect 12802 37068 12808 37120
rect 12860 37068 12866 37120
rect 13909 37111 13967 37117
rect 13909 37077 13921 37111
rect 13955 37108 13967 37111
rect 14734 37108 14740 37120
rect 13955 37080 14740 37108
rect 13955 37077 13967 37080
rect 13909 37071 13967 37077
rect 14734 37068 14740 37080
rect 14792 37108 14798 37120
rect 14936 37108 14964 37148
rect 17328 37120 17356 37148
rect 18064 37148 18705 37176
rect 18064 37120 18092 37148
rect 18693 37145 18705 37148
rect 18739 37145 18751 37179
rect 18693 37139 18751 37145
rect 18785 37179 18843 37185
rect 18785 37145 18797 37179
rect 18831 37176 18843 37179
rect 19168 37176 19196 37216
rect 18831 37148 19196 37176
rect 19245 37179 19303 37185
rect 18831 37145 18843 37148
rect 18785 37139 18843 37145
rect 19245 37145 19257 37179
rect 19291 37176 19303 37179
rect 19352 37176 19380 37352
rect 19426 37272 19432 37324
rect 19484 37272 19490 37324
rect 20162 37272 20168 37324
rect 20220 37272 20226 37324
rect 22281 37315 22339 37321
rect 22281 37281 22293 37315
rect 22327 37312 22339 37315
rect 22370 37312 22376 37324
rect 22327 37284 22376 37312
rect 22327 37281 22339 37284
rect 22281 37275 22339 37281
rect 22370 37272 22376 37284
rect 22428 37272 22434 37324
rect 23492 37312 23520 37408
rect 24946 37340 24952 37392
rect 25004 37340 25010 37392
rect 27614 37380 27620 37392
rect 25976 37352 27620 37380
rect 23492 37284 24808 37312
rect 19444 37185 19472 37272
rect 20180 37244 20208 37272
rect 22005 37247 22063 37253
rect 22005 37244 22017 37247
rect 20180 37216 22017 37244
rect 22005 37213 22017 37216
rect 22051 37213 22063 37247
rect 22005 37207 22063 37213
rect 23382 37204 23388 37256
rect 23440 37204 23446 37256
rect 23566 37204 23572 37256
rect 23624 37244 23630 37256
rect 24397 37247 24455 37253
rect 24397 37244 24409 37247
rect 23624 37216 24409 37244
rect 23624 37204 23630 37216
rect 24397 37213 24409 37216
rect 24443 37244 24455 37247
rect 24486 37244 24492 37256
rect 24443 37216 24492 37244
rect 24443 37213 24455 37216
rect 24397 37207 24455 37213
rect 24486 37204 24492 37216
rect 24544 37204 24550 37256
rect 24670 37204 24676 37256
rect 24728 37204 24734 37256
rect 24780 37253 24808 37284
rect 25222 37272 25228 37324
rect 25280 37312 25286 37324
rect 25409 37315 25467 37321
rect 25409 37312 25421 37315
rect 25280 37284 25421 37312
rect 25280 37272 25286 37284
rect 25409 37281 25421 37284
rect 25455 37281 25467 37315
rect 25409 37275 25467 37281
rect 25976 37256 26004 37352
rect 27614 37340 27620 37352
rect 27672 37340 27678 37392
rect 29549 37383 29607 37389
rect 29549 37349 29561 37383
rect 29595 37349 29607 37383
rect 29549 37343 29607 37349
rect 27522 37312 27528 37324
rect 27356 37284 27528 37312
rect 24765 37247 24823 37253
rect 24765 37213 24777 37247
rect 24811 37244 24823 37247
rect 24811 37216 25912 37244
rect 24811 37213 24823 37216
rect 24765 37207 24823 37213
rect 19291 37148 19380 37176
rect 19429 37179 19487 37185
rect 19291 37145 19303 37148
rect 19245 37139 19303 37145
rect 19429 37145 19441 37179
rect 19475 37145 19487 37179
rect 19429 37139 19487 37145
rect 14792 37080 14964 37108
rect 14792 37068 14798 37080
rect 17310 37068 17316 37120
rect 17368 37068 17374 37120
rect 18046 37068 18052 37120
rect 18104 37068 18110 37120
rect 18708 37108 18736 37139
rect 18966 37108 18972 37120
rect 18708 37080 18972 37108
rect 18966 37068 18972 37080
rect 19024 37068 19030 37120
rect 19260 37108 19288 37139
rect 19518 37136 19524 37188
rect 19576 37136 19582 37188
rect 24578 37136 24584 37188
rect 24636 37136 24642 37188
rect 25133 37179 25191 37185
rect 24918 37148 25084 37176
rect 19536 37108 19564 37136
rect 19260 37080 19564 37108
rect 23750 37068 23756 37120
rect 23808 37068 23814 37120
rect 24596 37108 24624 37136
rect 24918 37108 24946 37148
rect 24596 37080 24946 37108
rect 25056 37108 25084 37148
rect 25133 37145 25145 37179
rect 25179 37176 25191 37179
rect 25498 37176 25504 37188
rect 25179 37148 25504 37176
rect 25179 37145 25191 37148
rect 25133 37139 25191 37145
rect 25498 37136 25504 37148
rect 25556 37136 25562 37188
rect 25884 37176 25912 37216
rect 25958 37204 25964 37256
rect 26016 37204 26022 37256
rect 26050 37204 26056 37256
rect 26108 37244 26114 37256
rect 27356 37253 27384 37284
rect 27522 37272 27528 37284
rect 27580 37272 27586 37324
rect 29564 37312 29592 37343
rect 29564 37284 29960 37312
rect 26329 37247 26387 37253
rect 26329 37244 26341 37247
rect 26108 37216 26341 37244
rect 26108 37204 26114 37216
rect 26329 37213 26341 37216
rect 26375 37213 26387 37247
rect 26329 37207 26387 37213
rect 27341 37247 27399 37253
rect 27341 37213 27353 37247
rect 27387 37213 27399 37247
rect 27709 37247 27767 37253
rect 27709 37244 27721 37247
rect 27341 37207 27399 37213
rect 27448 37216 27721 37244
rect 26068 37176 26096 37204
rect 25884 37148 26096 37176
rect 26145 37179 26203 37185
rect 26145 37145 26157 37179
rect 26191 37145 26203 37179
rect 26145 37139 26203 37145
rect 25774 37108 25780 37120
rect 25056 37080 25780 37108
rect 25774 37068 25780 37080
rect 25832 37108 25838 37120
rect 26160 37108 26188 37139
rect 26234 37136 26240 37188
rect 26292 37136 26298 37188
rect 26344 37176 26372 37207
rect 27448 37188 27476 37216
rect 27709 37213 27721 37216
rect 27755 37213 27767 37247
rect 27709 37207 27767 37213
rect 28442 37204 28448 37256
rect 28500 37244 28506 37256
rect 29733 37247 29791 37253
rect 29733 37244 29745 37247
rect 28500 37216 29745 37244
rect 28500 37204 28506 37216
rect 29733 37213 29745 37216
rect 29779 37213 29791 37247
rect 29733 37207 29791 37213
rect 29825 37247 29883 37253
rect 29825 37213 29837 37247
rect 29871 37213 29883 37247
rect 29932 37244 29960 37284
rect 31202 37272 31208 37324
rect 31260 37312 31266 37324
rect 31726 37312 31754 37420
rect 31941 37417 31953 37420
rect 31987 37417 31999 37451
rect 31941 37411 31999 37417
rect 31260 37284 31754 37312
rect 31260 37272 31266 37284
rect 30193 37247 30251 37253
rect 30193 37244 30205 37247
rect 29932 37216 30205 37244
rect 29825 37207 29883 37213
rect 30193 37213 30205 37216
rect 30239 37213 30251 37247
rect 30193 37207 30251 37213
rect 27430 37176 27436 37188
rect 26344 37148 27436 37176
rect 27430 37136 27436 37148
rect 27488 37136 27494 37188
rect 27525 37179 27583 37185
rect 27525 37145 27537 37179
rect 27571 37145 27583 37179
rect 27525 37139 27583 37145
rect 27338 37108 27344 37120
rect 25832 37080 27344 37108
rect 25832 37068 25838 37080
rect 27338 37068 27344 37080
rect 27396 37108 27402 37120
rect 27540 37108 27568 37139
rect 27614 37136 27620 37188
rect 27672 37136 27678 37188
rect 27396 37080 27568 37108
rect 29840 37108 29868 37207
rect 31220 37162 31248 37272
rect 31312 37216 35664 37244
rect 31312 37108 31340 37216
rect 35636 37188 35664 37216
rect 40770 37204 40776 37256
rect 40828 37204 40834 37256
rect 31846 37136 31852 37188
rect 31904 37136 31910 37188
rect 35618 37136 35624 37188
rect 35676 37136 35682 37188
rect 29840 37080 31340 37108
rect 27396 37068 27402 37080
rect 31478 37068 31484 37120
rect 31536 37108 31542 37120
rect 31619 37111 31677 37117
rect 31619 37108 31631 37111
rect 31536 37080 31631 37108
rect 31536 37068 31542 37080
rect 31619 37077 31631 37080
rect 31665 37077 31677 37111
rect 31619 37071 31677 37077
rect 40954 37068 40960 37120
rect 41012 37068 41018 37120
rect 1104 37018 41400 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 41400 37018
rect 1104 36944 41400 36966
rect 5258 36904 5264 36916
rect 3712 36876 5264 36904
rect 3712 36836 3740 36876
rect 5258 36864 5264 36876
rect 5316 36904 5322 36916
rect 6914 36904 6920 36916
rect 5316 36876 6408 36904
rect 5316 36864 5322 36876
rect 3266 36808 3740 36836
rect 3786 36796 3792 36848
rect 3844 36796 3850 36848
rect 6380 36780 6408 36876
rect 6656 36876 6920 36904
rect 1762 36728 1768 36780
rect 1820 36728 1826 36780
rect 5718 36728 5724 36780
rect 5776 36728 5782 36780
rect 6362 36728 6368 36780
rect 6420 36728 6426 36780
rect 6656 36777 6684 36876
rect 6914 36864 6920 36876
rect 6972 36864 6978 36916
rect 7282 36864 7288 36916
rect 7340 36904 7346 36916
rect 8021 36907 8079 36913
rect 8021 36904 8033 36907
rect 7340 36876 8033 36904
rect 7340 36864 7346 36876
rect 8021 36873 8033 36876
rect 8067 36873 8079 36907
rect 8021 36867 8079 36873
rect 10321 36907 10379 36913
rect 10321 36873 10333 36907
rect 10367 36904 10379 36907
rect 10686 36904 10692 36916
rect 10367 36876 10692 36904
rect 10367 36873 10379 36876
rect 10321 36867 10379 36873
rect 10686 36864 10692 36876
rect 10744 36864 10750 36916
rect 22189 36907 22247 36913
rect 11900 36876 18092 36904
rect 6840 36808 7696 36836
rect 6641 36771 6699 36777
rect 6641 36737 6653 36771
rect 6687 36737 6699 36771
rect 6641 36731 6699 36737
rect 6730 36728 6736 36780
rect 6788 36768 6794 36780
rect 6840 36777 6868 36808
rect 6825 36771 6883 36777
rect 6825 36768 6837 36771
rect 6788 36740 6837 36768
rect 6788 36728 6794 36740
rect 6825 36737 6837 36740
rect 6871 36737 6883 36771
rect 6825 36731 6883 36737
rect 6917 36771 6975 36777
rect 6917 36737 6929 36771
rect 6963 36768 6975 36771
rect 7098 36768 7104 36780
rect 6963 36740 7104 36768
rect 6963 36737 6975 36740
rect 6917 36731 6975 36737
rect 7098 36728 7104 36740
rect 7156 36728 7162 36780
rect 7282 36768 7288 36780
rect 7244 36740 7288 36768
rect 7282 36728 7288 36740
rect 7340 36728 7346 36780
rect 7668 36777 7696 36808
rect 8294 36796 8300 36848
rect 8352 36836 8358 36848
rect 11900 36836 11928 36876
rect 12434 36836 12440 36848
rect 8352 36808 11928 36836
rect 11992 36808 12440 36836
rect 8352 36796 8358 36808
rect 7653 36771 7711 36777
rect 7653 36737 7665 36771
rect 7699 36737 7711 36771
rect 7653 36731 7711 36737
rect 7742 36728 7748 36780
rect 7800 36728 7806 36780
rect 9953 36771 10011 36777
rect 9953 36737 9965 36771
rect 9999 36768 10011 36771
rect 10226 36768 10232 36780
rect 9999 36740 10232 36768
rect 9999 36737 10011 36740
rect 9953 36731 10011 36737
rect 10226 36728 10232 36740
rect 10284 36728 10290 36780
rect 11992 36777 12020 36808
rect 12434 36796 12440 36808
rect 12492 36796 12498 36848
rect 14090 36796 14096 36848
rect 14148 36796 14154 36848
rect 17678 36836 17684 36848
rect 14476 36808 15792 36836
rect 11977 36771 12035 36777
rect 11977 36737 11989 36771
rect 12023 36737 12035 36771
rect 11977 36731 12035 36737
rect 2038 36660 2044 36712
rect 2096 36660 2102 36712
rect 4341 36703 4399 36709
rect 4341 36669 4353 36703
rect 4387 36669 4399 36703
rect 4341 36663 4399 36669
rect 4617 36703 4675 36709
rect 4617 36669 4629 36703
rect 4663 36700 4675 36703
rect 7009 36703 7067 36709
rect 7009 36700 7021 36703
rect 4663 36672 7021 36700
rect 4663 36669 4675 36672
rect 4617 36663 4675 36669
rect 7009 36669 7021 36672
rect 7055 36669 7067 36703
rect 7009 36663 7067 36669
rect 4062 36524 4068 36576
rect 4120 36564 4126 36576
rect 4356 36564 4384 36663
rect 7190 36660 7196 36712
rect 7248 36660 7254 36712
rect 7374 36660 7380 36712
rect 7432 36660 7438 36712
rect 7469 36703 7527 36709
rect 7469 36669 7481 36703
rect 7515 36700 7527 36703
rect 7558 36700 7564 36712
rect 7515 36672 7564 36700
rect 7515 36669 7527 36672
rect 7469 36663 7527 36669
rect 7558 36660 7564 36672
rect 7616 36660 7622 36712
rect 10045 36703 10103 36709
rect 10045 36669 10057 36703
rect 10091 36700 10103 36703
rect 10778 36700 10784 36712
rect 10091 36672 10784 36700
rect 10091 36669 10103 36672
rect 10045 36663 10103 36669
rect 10778 36660 10784 36672
rect 10836 36660 10842 36712
rect 12069 36703 12127 36709
rect 12069 36669 12081 36703
rect 12115 36669 12127 36703
rect 12345 36703 12403 36709
rect 12345 36700 12357 36703
rect 12069 36663 12127 36669
rect 12176 36672 12357 36700
rect 8662 36632 8668 36644
rect 5644 36604 8668 36632
rect 5644 36564 5672 36604
rect 8662 36592 8668 36604
rect 8720 36632 8726 36644
rect 12084 36632 12112 36663
rect 8720 36604 12112 36632
rect 8720 36592 8726 36604
rect 4120 36536 5672 36564
rect 4120 36524 4126 36536
rect 6086 36524 6092 36576
rect 6144 36524 6150 36576
rect 6454 36524 6460 36576
rect 6512 36524 6518 36576
rect 6914 36524 6920 36576
rect 6972 36564 6978 36576
rect 7653 36567 7711 36573
rect 7653 36564 7665 36567
rect 6972 36536 7665 36564
rect 6972 36524 6978 36536
rect 7653 36533 7665 36536
rect 7699 36533 7711 36567
rect 7653 36527 7711 36533
rect 11793 36567 11851 36573
rect 11793 36533 11805 36567
rect 11839 36564 11851 36567
rect 12176 36564 12204 36672
rect 12345 36669 12357 36672
rect 12391 36669 12403 36703
rect 13464 36700 13492 36754
rect 13906 36700 13912 36712
rect 13464 36672 13912 36700
rect 12345 36663 12403 36669
rect 13906 36660 13912 36672
rect 13964 36700 13970 36712
rect 14476 36700 14504 36808
rect 15764 36780 15792 36808
rect 17236 36808 17684 36836
rect 14553 36771 14611 36777
rect 14553 36737 14565 36771
rect 14599 36768 14611 36771
rect 15010 36768 15016 36780
rect 14599 36740 15016 36768
rect 14599 36737 14611 36740
rect 14553 36731 14611 36737
rect 15010 36728 15016 36740
rect 15068 36728 15074 36780
rect 15105 36771 15163 36777
rect 15105 36737 15117 36771
rect 15151 36737 15163 36771
rect 15105 36731 15163 36737
rect 13964 36672 14504 36700
rect 13964 36660 13970 36672
rect 14642 36660 14648 36712
rect 14700 36660 14706 36712
rect 15120 36700 15148 36731
rect 15746 36728 15752 36780
rect 15804 36728 15810 36780
rect 16025 36771 16083 36777
rect 16025 36737 16037 36771
rect 16071 36768 16083 36771
rect 16206 36768 16212 36780
rect 16071 36740 16212 36768
rect 16071 36737 16083 36740
rect 16025 36731 16083 36737
rect 16206 36728 16212 36740
rect 16264 36728 16270 36780
rect 16850 36728 16856 36780
rect 16908 36728 16914 36780
rect 17236 36777 17264 36808
rect 17678 36796 17684 36808
rect 17736 36796 17742 36848
rect 18064 36836 18092 36876
rect 19168 36876 21680 36904
rect 18064 36808 19104 36836
rect 17037 36771 17095 36777
rect 17037 36737 17049 36771
rect 17083 36768 17095 36771
rect 17221 36771 17279 36777
rect 17221 36768 17233 36771
rect 17083 36740 17233 36768
rect 17083 36737 17095 36740
rect 17037 36731 17095 36737
rect 17221 36737 17233 36740
rect 17267 36737 17279 36771
rect 17221 36731 17279 36737
rect 17405 36771 17463 36777
rect 17405 36737 17417 36771
rect 17451 36737 17463 36771
rect 17405 36731 17463 36737
rect 14936 36672 15148 36700
rect 16117 36703 16175 36709
rect 14274 36592 14280 36644
rect 14332 36632 14338 36644
rect 14936 36632 14964 36672
rect 16117 36669 16129 36703
rect 16163 36700 16175 36703
rect 16482 36700 16488 36712
rect 16163 36672 16488 36700
rect 16163 36669 16175 36672
rect 16117 36663 16175 36669
rect 16482 36660 16488 36672
rect 16540 36660 16546 36712
rect 17129 36703 17187 36709
rect 17129 36669 17141 36703
rect 17175 36700 17187 36703
rect 17420 36700 17448 36731
rect 18046 36728 18052 36780
rect 18104 36728 18110 36780
rect 18141 36771 18199 36777
rect 18141 36737 18153 36771
rect 18187 36768 18199 36771
rect 18187 36740 18276 36768
rect 18187 36737 18199 36740
rect 18141 36731 18199 36737
rect 17175 36672 17448 36700
rect 17175 36669 17187 36672
rect 17129 36663 17187 36669
rect 14332 36604 14964 36632
rect 14332 36592 14338 36604
rect 14936 36576 14964 36604
rect 16393 36635 16451 36641
rect 16393 36601 16405 36635
rect 16439 36632 16451 36635
rect 17144 36632 17172 36663
rect 18248 36644 18276 36740
rect 18322 36728 18328 36780
rect 18380 36728 18386 36780
rect 18414 36728 18420 36780
rect 18472 36728 18478 36780
rect 18693 36771 18751 36777
rect 18693 36737 18705 36771
rect 18739 36737 18751 36771
rect 18693 36731 18751 36737
rect 16439 36604 17172 36632
rect 17236 36604 17448 36632
rect 16439 36601 16451 36604
rect 16393 36595 16451 36601
rect 11839 36536 12204 36564
rect 11839 36533 11851 36536
rect 11793 36527 11851 36533
rect 14826 36524 14832 36576
rect 14884 36524 14890 36576
rect 14918 36524 14924 36576
rect 14976 36524 14982 36576
rect 15194 36524 15200 36576
rect 15252 36524 15258 36576
rect 15378 36524 15384 36576
rect 15436 36564 15442 36576
rect 16669 36567 16727 36573
rect 16669 36564 16681 36567
rect 15436 36536 16681 36564
rect 15436 36524 15442 36536
rect 16669 36533 16681 36536
rect 16715 36533 16727 36567
rect 16669 36527 16727 36533
rect 17034 36524 17040 36576
rect 17092 36564 17098 36576
rect 17236 36564 17264 36604
rect 17092 36536 17264 36564
rect 17092 36524 17098 36536
rect 17310 36524 17316 36576
rect 17368 36524 17374 36576
rect 17420 36564 17448 36604
rect 18230 36592 18236 36644
rect 18288 36592 18294 36644
rect 18340 36632 18368 36728
rect 18598 36660 18604 36712
rect 18656 36660 18662 36712
rect 18708 36632 18736 36731
rect 18340 36604 18736 36632
rect 18966 36592 18972 36644
rect 19024 36592 19030 36644
rect 19076 36632 19104 36808
rect 19168 36780 19196 36876
rect 20162 36836 20168 36848
rect 19628 36808 20168 36836
rect 19150 36728 19156 36780
rect 19208 36728 19214 36780
rect 19628 36777 19656 36808
rect 20162 36796 20168 36808
rect 20220 36796 20226 36848
rect 21652 36845 21680 36876
rect 22189 36873 22201 36907
rect 22235 36904 22247 36907
rect 22646 36904 22652 36916
rect 22235 36876 22652 36904
rect 22235 36873 22247 36876
rect 22189 36867 22247 36873
rect 22646 36864 22652 36876
rect 22704 36864 22710 36916
rect 24762 36864 24768 36916
rect 24820 36904 24826 36916
rect 25222 36904 25228 36916
rect 24820 36876 25228 36904
rect 24820 36864 24826 36876
rect 25222 36864 25228 36876
rect 25280 36864 25286 36916
rect 27430 36864 27436 36916
rect 27488 36864 27494 36916
rect 27801 36907 27859 36913
rect 27801 36873 27813 36907
rect 27847 36904 27859 36907
rect 28166 36904 28172 36916
rect 27847 36876 28172 36904
rect 27847 36873 27859 36876
rect 27801 36867 27859 36873
rect 28166 36864 28172 36876
rect 28224 36864 28230 36916
rect 31846 36904 31852 36916
rect 28552 36876 31852 36904
rect 21637 36839 21695 36845
rect 21637 36805 21649 36839
rect 21683 36805 21695 36839
rect 27448 36836 27476 36864
rect 27448 36808 27660 36836
rect 21637 36799 21695 36805
rect 19613 36771 19671 36777
rect 19613 36737 19625 36771
rect 19659 36737 19671 36771
rect 19613 36731 19671 36737
rect 20990 36728 20996 36780
rect 21048 36728 21054 36780
rect 22557 36771 22615 36777
rect 22557 36737 22569 36771
rect 22603 36768 22615 36771
rect 23750 36768 23756 36780
rect 22603 36740 23756 36768
rect 22603 36737 22615 36740
rect 22557 36731 22615 36737
rect 23750 36728 23756 36740
rect 23808 36728 23814 36780
rect 23934 36728 23940 36780
rect 23992 36768 23998 36780
rect 27246 36768 27252 36780
rect 23992 36740 27252 36768
rect 23992 36728 23998 36740
rect 27246 36728 27252 36740
rect 27304 36728 27310 36780
rect 27338 36728 27344 36780
rect 27396 36768 27402 36780
rect 27433 36771 27491 36777
rect 27433 36768 27445 36771
rect 27396 36740 27445 36768
rect 27396 36728 27402 36740
rect 27433 36737 27445 36740
rect 27479 36737 27491 36771
rect 27433 36731 27491 36737
rect 19245 36703 19303 36709
rect 19245 36669 19257 36703
rect 19291 36700 19303 36703
rect 19426 36700 19432 36712
rect 19291 36672 19432 36700
rect 19291 36669 19303 36672
rect 19245 36663 19303 36669
rect 19426 36660 19432 36672
rect 19484 36660 19490 36712
rect 19886 36660 19892 36712
rect 19944 36660 19950 36712
rect 22649 36703 22707 36709
rect 22649 36700 22661 36703
rect 22066 36672 22661 36700
rect 19610 36632 19616 36644
rect 19076 36604 19616 36632
rect 19610 36592 19616 36604
rect 19668 36592 19674 36644
rect 17586 36564 17592 36576
rect 17420 36536 17592 36564
rect 17586 36524 17592 36536
rect 17644 36564 17650 36576
rect 18417 36567 18475 36573
rect 18417 36564 18429 36567
rect 17644 36536 18429 36564
rect 17644 36524 17650 36536
rect 18417 36533 18429 36536
rect 18463 36533 18475 36567
rect 18417 36527 18475 36533
rect 18874 36524 18880 36576
rect 18932 36524 18938 36576
rect 18984 36564 19012 36592
rect 19521 36567 19579 36573
rect 19521 36564 19533 36567
rect 18984 36536 19533 36564
rect 19521 36533 19533 36536
rect 19567 36533 19579 36567
rect 19521 36527 19579 36533
rect 20530 36524 20536 36576
rect 20588 36564 20594 36576
rect 22066 36564 22094 36672
rect 22649 36669 22661 36672
rect 22695 36669 22707 36703
rect 22649 36663 22707 36669
rect 22830 36660 22836 36712
rect 22888 36660 22894 36712
rect 27448 36700 27476 36731
rect 27522 36728 27528 36780
rect 27580 36728 27586 36780
rect 27632 36777 27660 36808
rect 27706 36796 27712 36848
rect 27764 36836 27770 36848
rect 28552 36836 28580 36876
rect 31846 36864 31852 36876
rect 31904 36904 31910 36916
rect 40034 36904 40040 36916
rect 31904 36876 40040 36904
rect 31904 36864 31910 36876
rect 40034 36864 40040 36876
rect 40092 36864 40098 36916
rect 27764 36808 28658 36836
rect 27764 36796 27770 36808
rect 27617 36771 27675 36777
rect 27617 36737 27629 36771
rect 27663 36737 27675 36771
rect 27617 36731 27675 36737
rect 30006 36728 30012 36780
rect 30064 36728 30070 36780
rect 30193 36771 30251 36777
rect 30193 36768 30205 36771
rect 30116 36740 30205 36768
rect 27448 36672 27522 36700
rect 20588 36536 22094 36564
rect 27494 36564 27522 36672
rect 27798 36660 27804 36712
rect 27856 36700 27862 36712
rect 27893 36703 27951 36709
rect 27893 36700 27905 36703
rect 27856 36672 27905 36700
rect 27856 36660 27862 36672
rect 27893 36669 27905 36672
rect 27939 36669 27951 36703
rect 27893 36663 27951 36669
rect 28166 36660 28172 36712
rect 28224 36660 28230 36712
rect 29822 36660 29828 36712
rect 29880 36700 29886 36712
rect 29917 36703 29975 36709
rect 29917 36700 29929 36703
rect 29880 36672 29929 36700
rect 29880 36660 29886 36672
rect 29917 36669 29929 36672
rect 29963 36669 29975 36703
rect 29917 36663 29975 36669
rect 30116 36632 30144 36740
rect 30193 36737 30205 36740
rect 30239 36737 30251 36771
rect 30193 36731 30251 36737
rect 29380 36604 30144 36632
rect 29380 36576 29408 36604
rect 30190 36592 30196 36644
rect 30248 36632 30254 36644
rect 30285 36635 30343 36641
rect 30285 36632 30297 36635
rect 30248 36604 30297 36632
rect 30248 36592 30254 36604
rect 30285 36601 30297 36604
rect 30331 36601 30343 36635
rect 30285 36595 30343 36601
rect 28718 36564 28724 36576
rect 27494 36536 28724 36564
rect 20588 36524 20594 36536
rect 28718 36524 28724 36536
rect 28776 36524 28782 36576
rect 29362 36524 29368 36576
rect 29420 36524 29426 36576
rect 1104 36474 41400 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 41400 36474
rect 1104 36400 41400 36422
rect 2038 36320 2044 36372
rect 2096 36360 2102 36372
rect 2317 36363 2375 36369
rect 2317 36360 2329 36363
rect 2096 36332 2329 36360
rect 2096 36320 2102 36332
rect 2317 36329 2329 36332
rect 2363 36329 2375 36363
rect 4062 36360 4068 36372
rect 2317 36323 2375 36329
rect 3804 36332 4068 36360
rect 3418 36184 3424 36236
rect 3476 36184 3482 36236
rect 3804 36233 3832 36332
rect 4062 36320 4068 36332
rect 4120 36320 4126 36372
rect 6914 36320 6920 36372
rect 6972 36320 6978 36372
rect 7558 36320 7564 36372
rect 7616 36360 7622 36372
rect 8113 36363 8171 36369
rect 8113 36360 8125 36363
rect 7616 36332 8125 36360
rect 7616 36320 7622 36332
rect 8113 36329 8125 36332
rect 8159 36329 8171 36363
rect 8113 36323 8171 36329
rect 9861 36363 9919 36369
rect 9861 36329 9873 36363
rect 9907 36360 9919 36363
rect 10318 36360 10324 36372
rect 9907 36332 10324 36360
rect 9907 36329 9919 36332
rect 9861 36323 9919 36329
rect 10318 36320 10324 36332
rect 10376 36320 10382 36372
rect 10778 36320 10784 36372
rect 10836 36320 10842 36372
rect 12802 36320 12808 36372
rect 12860 36360 12866 36372
rect 13173 36363 13231 36369
rect 13173 36360 13185 36363
rect 12860 36332 13185 36360
rect 12860 36320 12866 36332
rect 13173 36329 13185 36332
rect 13219 36329 13231 36363
rect 13173 36323 13231 36329
rect 14826 36320 14832 36372
rect 14884 36320 14890 36372
rect 15010 36320 15016 36372
rect 15068 36360 15074 36372
rect 15381 36363 15439 36369
rect 15381 36360 15393 36363
rect 15068 36332 15393 36360
rect 15068 36320 15074 36332
rect 15381 36329 15393 36332
rect 15427 36329 15439 36363
rect 15381 36323 15439 36329
rect 16298 36320 16304 36372
rect 16356 36320 16362 36372
rect 16577 36363 16635 36369
rect 16577 36329 16589 36363
rect 16623 36360 16635 36363
rect 16850 36360 16856 36372
rect 16623 36332 16856 36360
rect 16623 36329 16635 36332
rect 16577 36323 16635 36329
rect 16850 36320 16856 36332
rect 16908 36320 16914 36372
rect 17310 36320 17316 36372
rect 17368 36320 17374 36372
rect 18414 36320 18420 36372
rect 18472 36360 18478 36372
rect 18785 36363 18843 36369
rect 18785 36360 18797 36363
rect 18472 36332 18797 36360
rect 18472 36320 18478 36332
rect 18785 36329 18797 36332
rect 18831 36329 18843 36363
rect 18785 36323 18843 36329
rect 19337 36363 19395 36369
rect 19337 36329 19349 36363
rect 19383 36360 19395 36363
rect 19886 36360 19892 36372
rect 19383 36332 19892 36360
rect 19383 36329 19395 36332
rect 19337 36323 19395 36329
rect 19886 36320 19892 36332
rect 19944 36320 19950 36372
rect 23750 36320 23756 36372
rect 23808 36360 23814 36372
rect 28261 36363 28319 36369
rect 23808 36332 28212 36360
rect 23808 36320 23814 36332
rect 5718 36292 5724 36304
rect 5184 36264 5724 36292
rect 3789 36227 3847 36233
rect 3789 36193 3801 36227
rect 3835 36193 3847 36227
rect 3789 36187 3847 36193
rect 2501 36159 2559 36165
rect 2501 36125 2513 36159
rect 2547 36156 2559 36159
rect 2547 36128 2820 36156
rect 5184 36142 5212 36264
rect 5718 36252 5724 36264
rect 5776 36292 5782 36304
rect 7926 36292 7932 36304
rect 5776 36264 7932 36292
rect 5776 36252 5782 36264
rect 7926 36252 7932 36264
rect 7984 36252 7990 36304
rect 10226 36292 10232 36304
rect 9600 36264 10232 36292
rect 6641 36227 6699 36233
rect 6641 36193 6653 36227
rect 6687 36224 6699 36227
rect 7006 36224 7012 36236
rect 6687 36196 7012 36224
rect 6687 36193 6699 36196
rect 6641 36187 6699 36193
rect 7006 36184 7012 36196
rect 7064 36184 7070 36236
rect 7576 36196 8340 36224
rect 2547 36125 2559 36128
rect 2501 36119 2559 36125
rect 2792 36029 2820 36128
rect 6086 36116 6092 36168
rect 6144 36156 6150 36168
rect 7576 36165 7604 36196
rect 8312 36168 8340 36196
rect 6549 36159 6607 36165
rect 6549 36156 6561 36159
rect 6144 36128 6561 36156
rect 6144 36116 6150 36128
rect 6549 36125 6561 36128
rect 6595 36125 6607 36159
rect 6549 36119 6607 36125
rect 7561 36159 7619 36165
rect 7561 36125 7573 36159
rect 7607 36125 7619 36159
rect 7561 36119 7619 36125
rect 7929 36159 7987 36165
rect 7929 36125 7941 36159
rect 7975 36156 7987 36159
rect 8202 36156 8208 36168
rect 7975 36128 8208 36156
rect 7975 36125 7987 36128
rect 7929 36119 7987 36125
rect 3145 36091 3203 36097
rect 3145 36057 3157 36091
rect 3191 36088 3203 36091
rect 3786 36088 3792 36100
rect 3191 36060 3792 36088
rect 3191 36057 3203 36060
rect 3145 36051 3203 36057
rect 3786 36048 3792 36060
rect 3844 36048 3850 36100
rect 4065 36091 4123 36097
rect 4065 36057 4077 36091
rect 4111 36088 4123 36091
rect 4154 36088 4160 36100
rect 4111 36060 4160 36088
rect 4111 36057 4123 36060
rect 4065 36051 4123 36057
rect 4154 36048 4160 36060
rect 4212 36048 4218 36100
rect 2777 36023 2835 36029
rect 2777 35989 2789 36023
rect 2823 35989 2835 36023
rect 2777 35983 2835 35989
rect 3237 36023 3295 36029
rect 3237 35989 3249 36023
rect 3283 36020 3295 36023
rect 3970 36020 3976 36032
rect 3283 35992 3976 36020
rect 3283 35989 3295 35992
rect 3237 35983 3295 35989
rect 3970 35980 3976 35992
rect 4028 35980 4034 36032
rect 5534 35980 5540 36032
rect 5592 35980 5598 36032
rect 6564 36020 6592 36119
rect 8202 36116 8208 36128
rect 8260 36116 8266 36168
rect 8294 36116 8300 36168
rect 8352 36116 8358 36168
rect 9600 36165 9628 36264
rect 10226 36252 10232 36264
rect 10284 36252 10290 36304
rect 14844 36292 14872 36320
rect 13648 36264 14872 36292
rect 15289 36295 15347 36301
rect 9677 36227 9735 36233
rect 9677 36193 9689 36227
rect 9723 36224 9735 36227
rect 10873 36227 10931 36233
rect 10873 36224 10885 36227
rect 9723 36196 10364 36224
rect 9723 36193 9735 36196
rect 9677 36187 9735 36193
rect 10336 36165 10364 36196
rect 10520 36196 10885 36224
rect 10520 36168 10548 36196
rect 10873 36193 10885 36196
rect 10919 36193 10931 36227
rect 10873 36187 10931 36193
rect 12710 36184 12716 36236
rect 12768 36184 12774 36236
rect 13648 36233 13676 36264
rect 15289 36261 15301 36295
rect 15335 36292 15347 36295
rect 15838 36292 15844 36304
rect 15335 36264 15844 36292
rect 15335 36261 15347 36264
rect 15289 36255 15347 36261
rect 15838 36252 15844 36264
rect 15896 36292 15902 36304
rect 16316 36292 16344 36320
rect 15896 36264 16344 36292
rect 15896 36252 15902 36264
rect 13633 36227 13691 36233
rect 13633 36193 13645 36227
rect 13679 36193 13691 36227
rect 13633 36187 13691 36193
rect 13722 36184 13728 36236
rect 13780 36224 13786 36236
rect 15473 36227 15531 36233
rect 13780 36196 15148 36224
rect 13780 36184 13786 36196
rect 9585 36159 9643 36165
rect 9585 36125 9597 36159
rect 9631 36125 9643 36159
rect 9585 36119 9643 36125
rect 9769 36159 9827 36165
rect 9769 36125 9781 36159
rect 9815 36156 9827 36159
rect 10137 36159 10195 36165
rect 10137 36156 10149 36159
rect 9815 36128 10149 36156
rect 9815 36125 9827 36128
rect 9769 36119 9827 36125
rect 10137 36125 10149 36128
rect 10183 36125 10195 36159
rect 10137 36119 10195 36125
rect 10229 36159 10287 36165
rect 10229 36125 10241 36159
rect 10275 36125 10287 36159
rect 10229 36119 10287 36125
rect 10321 36159 10379 36165
rect 10321 36125 10333 36159
rect 10367 36125 10379 36159
rect 10321 36119 10379 36125
rect 7742 36048 7748 36100
rect 7800 36048 7806 36100
rect 7837 36091 7895 36097
rect 7837 36057 7849 36091
rect 7883 36088 7895 36091
rect 8110 36088 8116 36100
rect 7883 36060 8116 36088
rect 7883 36057 7895 36060
rect 7837 36051 7895 36057
rect 7852 36020 7880 36051
rect 8110 36048 8116 36060
rect 8168 36048 8174 36100
rect 8220 36088 8248 36116
rect 8846 36088 8852 36100
rect 8220 36060 8852 36088
rect 8846 36048 8852 36060
rect 8904 36048 8910 36100
rect 6564 35992 7880 36020
rect 9784 36020 9812 36119
rect 10042 36048 10048 36100
rect 10100 36088 10106 36100
rect 10244 36088 10272 36119
rect 10502 36116 10508 36168
rect 10560 36116 10566 36168
rect 10597 36159 10655 36165
rect 10597 36125 10609 36159
rect 10643 36125 10655 36159
rect 10597 36119 10655 36125
rect 10689 36159 10747 36165
rect 10689 36125 10701 36159
rect 10735 36156 10747 36159
rect 10962 36156 10968 36168
rect 10735 36128 10968 36156
rect 10735 36125 10747 36128
rect 10689 36119 10747 36125
rect 10100 36060 10272 36088
rect 10612 36088 10640 36119
rect 10962 36116 10968 36128
rect 11020 36116 11026 36168
rect 12526 36116 12532 36168
rect 12584 36156 12590 36168
rect 12621 36159 12679 36165
rect 12621 36156 12633 36159
rect 12584 36128 12633 36156
rect 12584 36116 12590 36128
rect 12621 36125 12633 36128
rect 12667 36125 12679 36159
rect 12621 36119 12679 36125
rect 11054 36088 11060 36100
rect 10612 36060 11060 36088
rect 10100 36048 10106 36060
rect 10704 36032 10732 36060
rect 11054 36048 11060 36060
rect 11112 36048 11118 36100
rect 13541 36091 13599 36097
rect 13541 36088 13553 36091
rect 13004 36060 13553 36088
rect 10686 36020 10692 36032
rect 9784 35992 10692 36020
rect 10686 35980 10692 35992
rect 10744 35980 10750 36032
rect 13004 36029 13032 36060
rect 13541 36057 13553 36060
rect 13587 36057 13599 36091
rect 13541 36051 13599 36057
rect 12989 36023 13047 36029
rect 12989 35989 13001 36023
rect 13035 35989 13047 36023
rect 15120 36020 15148 36196
rect 15473 36193 15485 36227
rect 15519 36224 15531 36227
rect 16209 36227 16267 36233
rect 16209 36224 16221 36227
rect 15519 36196 16221 36224
rect 15519 36193 15531 36196
rect 15473 36187 15531 36193
rect 16209 36193 16221 36196
rect 16255 36224 16267 36227
rect 17328 36224 17356 36320
rect 18506 36252 18512 36304
rect 18564 36252 18570 36304
rect 19426 36292 19432 36304
rect 18616 36264 19432 36292
rect 18141 36227 18199 36233
rect 18141 36224 18153 36227
rect 16255 36196 17356 36224
rect 18064 36196 18153 36224
rect 16255 36193 16267 36196
rect 16209 36187 16267 36193
rect 18064 36168 18092 36196
rect 18141 36193 18153 36196
rect 18187 36193 18199 36227
rect 18141 36187 18199 36193
rect 15197 36159 15255 36165
rect 15197 36125 15209 36159
rect 15243 36125 15255 36159
rect 15197 36119 15255 36125
rect 15212 36088 15240 36119
rect 15930 36116 15936 36168
rect 15988 36156 15994 36168
rect 16393 36159 16451 36165
rect 16393 36156 16405 36159
rect 15988 36128 16405 36156
rect 15988 36116 15994 36128
rect 16393 36125 16405 36128
rect 16439 36156 16451 36159
rect 16482 36156 16488 36168
rect 16439 36128 16488 36156
rect 16439 36125 16451 36128
rect 16393 36119 16451 36125
rect 16482 36116 16488 36128
rect 16540 36116 16546 36168
rect 18046 36116 18052 36168
rect 18104 36116 18110 36168
rect 18325 36159 18383 36165
rect 18325 36125 18337 36159
rect 18371 36156 18383 36159
rect 18616 36156 18644 36264
rect 19426 36252 19432 36264
rect 19484 36252 19490 36304
rect 19610 36252 19616 36304
rect 19668 36292 19674 36304
rect 20162 36292 20168 36304
rect 19668 36264 20168 36292
rect 19668 36252 19674 36264
rect 20162 36252 20168 36264
rect 20220 36292 20226 36304
rect 22830 36292 22836 36304
rect 20220 36264 22836 36292
rect 20220 36252 20226 36264
rect 22830 36252 22836 36264
rect 22888 36252 22894 36304
rect 24210 36252 24216 36304
rect 24268 36292 24274 36304
rect 25958 36292 25964 36304
rect 24268 36264 25964 36292
rect 24268 36252 24274 36264
rect 25958 36252 25964 36264
rect 26016 36252 26022 36304
rect 27249 36295 27307 36301
rect 27249 36261 27261 36295
rect 27295 36292 27307 36295
rect 28184 36292 28212 36332
rect 28261 36329 28273 36363
rect 28307 36360 28319 36363
rect 28350 36360 28356 36372
rect 28307 36332 28356 36360
rect 28307 36329 28319 36332
rect 28261 36323 28319 36329
rect 28350 36320 28356 36332
rect 28408 36320 28414 36372
rect 28442 36320 28448 36372
rect 28500 36320 28506 36372
rect 28718 36320 28724 36372
rect 28776 36320 28782 36372
rect 29730 36320 29736 36372
rect 29788 36320 29794 36372
rect 40770 36360 40776 36372
rect 31726 36332 40776 36360
rect 31726 36292 31754 36332
rect 40770 36320 40776 36332
rect 40828 36320 40834 36372
rect 27295 36264 28120 36292
rect 28184 36264 31754 36292
rect 27295 36261 27307 36264
rect 27249 36255 27307 36261
rect 18874 36184 18880 36236
rect 18932 36224 18938 36236
rect 18932 36196 19472 36224
rect 18932 36184 18938 36196
rect 18371 36128 18644 36156
rect 18785 36159 18843 36165
rect 18371 36125 18383 36128
rect 18325 36119 18383 36125
rect 18785 36125 18797 36159
rect 18831 36125 18843 36159
rect 18785 36119 18843 36125
rect 16206 36088 16212 36100
rect 15212 36060 16212 36088
rect 16206 36048 16212 36060
rect 16264 36048 16270 36100
rect 17862 36048 17868 36100
rect 17920 36048 17926 36100
rect 18230 36048 18236 36100
rect 18288 36088 18294 36100
rect 18800 36088 18828 36119
rect 18966 36116 18972 36168
rect 19024 36116 19030 36168
rect 19242 36116 19248 36168
rect 19300 36116 19306 36168
rect 19444 36165 19472 36196
rect 22370 36184 22376 36236
rect 22428 36224 22434 36236
rect 27801 36227 27859 36233
rect 27801 36224 27813 36227
rect 22428 36196 27813 36224
rect 22428 36184 22434 36196
rect 27801 36193 27813 36196
rect 27847 36193 27859 36227
rect 27801 36187 27859 36193
rect 27982 36184 27988 36236
rect 28040 36184 28046 36236
rect 19429 36159 19487 36165
rect 19429 36125 19441 36159
rect 19475 36125 19487 36159
rect 19429 36119 19487 36125
rect 19978 36116 19984 36168
rect 20036 36116 20042 36168
rect 25590 36116 25596 36168
rect 25648 36156 25654 36168
rect 27522 36156 27528 36168
rect 25648 36128 27528 36156
rect 25648 36116 25654 36128
rect 27522 36116 27528 36128
rect 27580 36116 27586 36168
rect 27709 36159 27767 36165
rect 27709 36125 27721 36159
rect 27755 36156 27767 36159
rect 28000 36156 28028 36184
rect 28092 36165 28120 36264
rect 29362 36184 29368 36236
rect 29420 36224 29426 36236
rect 29420 36196 29960 36224
rect 29420 36184 29426 36196
rect 27755 36128 28028 36156
rect 28077 36159 28135 36165
rect 27755 36125 27767 36128
rect 27709 36119 27767 36125
rect 28077 36125 28089 36159
rect 28123 36125 28135 36159
rect 28077 36119 28135 36125
rect 19996 36088 20024 36116
rect 18288 36060 20024 36088
rect 25685 36091 25743 36097
rect 18288 36048 18294 36060
rect 25685 36057 25697 36091
rect 25731 36088 25743 36091
rect 25866 36088 25872 36100
rect 25731 36060 25872 36088
rect 25731 36057 25743 36060
rect 25685 36051 25743 36057
rect 25866 36048 25872 36060
rect 25924 36048 25930 36100
rect 25958 36048 25964 36100
rect 26016 36088 26022 36100
rect 26510 36088 26516 36100
rect 26016 36060 26516 36088
rect 26016 36048 26022 36060
rect 26510 36048 26516 36060
rect 26568 36088 26574 36100
rect 27724 36088 27752 36119
rect 28258 36116 28264 36168
rect 28316 36116 28322 36168
rect 28994 36116 29000 36168
rect 29052 36116 29058 36168
rect 29380 36156 29408 36184
rect 29549 36159 29607 36165
rect 29549 36156 29561 36159
rect 29380 36128 29561 36156
rect 29549 36125 29561 36128
rect 29595 36125 29607 36159
rect 29549 36119 29607 36125
rect 29641 36159 29699 36165
rect 29641 36125 29653 36159
rect 29687 36125 29699 36159
rect 29641 36119 29699 36125
rect 26568 36060 27752 36088
rect 26568 36048 26574 36060
rect 28626 36048 28632 36100
rect 28684 36048 28690 36100
rect 29012 36088 29040 36116
rect 29656 36088 29684 36119
rect 29822 36116 29828 36168
rect 29880 36116 29886 36168
rect 29932 36165 29960 36196
rect 30006 36184 30012 36236
rect 30064 36224 30070 36236
rect 33597 36227 33655 36233
rect 30064 36196 30420 36224
rect 30064 36184 30070 36196
rect 30392 36165 30420 36196
rect 33597 36193 33609 36227
rect 33643 36224 33655 36227
rect 33643 36196 34192 36224
rect 33643 36193 33655 36196
rect 33597 36187 33655 36193
rect 34164 36168 34192 36196
rect 29917 36159 29975 36165
rect 29917 36125 29929 36159
rect 29963 36125 29975 36159
rect 29917 36119 29975 36125
rect 30377 36159 30435 36165
rect 30377 36125 30389 36159
rect 30423 36125 30435 36159
rect 30377 36119 30435 36125
rect 31846 36116 31852 36168
rect 31904 36116 31910 36168
rect 31938 36116 31944 36168
rect 31996 36156 32002 36168
rect 33781 36159 33839 36165
rect 33781 36156 33793 36159
rect 31996 36128 33793 36156
rect 31996 36116 32002 36128
rect 33781 36125 33793 36128
rect 33827 36156 33839 36159
rect 33827 36128 33916 36156
rect 33827 36125 33839 36128
rect 33781 36119 33839 36125
rect 29012 36060 30512 36088
rect 17880 36020 17908 36048
rect 15120 35992 17908 36020
rect 12989 35983 13047 35989
rect 24118 35980 24124 36032
rect 24176 36020 24182 36032
rect 25777 36023 25835 36029
rect 25777 36020 25789 36023
rect 24176 35992 25789 36020
rect 24176 35980 24182 35992
rect 25777 35989 25789 35992
rect 25823 36020 25835 36023
rect 26234 36020 26240 36032
rect 25823 35992 26240 36020
rect 25823 35989 25835 35992
rect 25777 35983 25835 35989
rect 26234 35980 26240 35992
rect 26292 35980 26298 36032
rect 27246 35980 27252 36032
rect 27304 36020 27310 36032
rect 27617 36023 27675 36029
rect 27617 36020 27629 36023
rect 27304 35992 27629 36020
rect 27304 35980 27310 35992
rect 27617 35989 27629 35992
rect 27663 36020 27675 36023
rect 28074 36020 28080 36032
rect 27663 35992 28080 36020
rect 27663 35989 27675 35992
rect 27617 35983 27675 35989
rect 28074 35980 28080 35992
rect 28132 35980 28138 36032
rect 28902 35980 28908 36032
rect 28960 36020 28966 36032
rect 30484 36029 30512 36060
rect 31110 36048 31116 36100
rect 31168 36088 31174 36100
rect 31168 36060 33180 36088
rect 31168 36048 31174 36060
rect 33152 36032 33180 36060
rect 33888 36032 33916 36128
rect 34146 36116 34152 36168
rect 34204 36116 34210 36168
rect 30101 36023 30159 36029
rect 30101 36020 30113 36023
rect 28960 35992 30113 36020
rect 28960 35980 28966 35992
rect 30101 35989 30113 35992
rect 30147 35989 30159 36023
rect 30101 35983 30159 35989
rect 30469 36023 30527 36029
rect 30469 35989 30481 36023
rect 30515 35989 30527 36023
rect 30469 35983 30527 35989
rect 32122 35980 32128 36032
rect 32180 35980 32186 36032
rect 33134 35980 33140 36032
rect 33192 35980 33198 36032
rect 33870 35980 33876 36032
rect 33928 35980 33934 36032
rect 33962 35980 33968 36032
rect 34020 35980 34026 36032
rect 1104 35930 41400 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 41400 35930
rect 1104 35856 41400 35878
rect 4154 35776 4160 35828
rect 4212 35816 4218 35828
rect 4249 35819 4307 35825
rect 4249 35816 4261 35819
rect 4212 35788 4261 35816
rect 4212 35776 4218 35788
rect 4249 35785 4261 35788
rect 4295 35785 4307 35819
rect 4249 35779 4307 35785
rect 7009 35819 7067 35825
rect 7009 35785 7021 35819
rect 7055 35816 7067 35819
rect 8110 35816 8116 35828
rect 7055 35788 8116 35816
rect 7055 35785 7067 35788
rect 7009 35779 7067 35785
rect 8110 35776 8116 35788
rect 8168 35776 8174 35828
rect 10962 35816 10968 35828
rect 10152 35788 10968 35816
rect 4433 35683 4491 35689
rect 4433 35649 4445 35683
rect 4479 35680 4491 35683
rect 4479 35652 4752 35680
rect 4479 35649 4491 35652
rect 4433 35643 4491 35649
rect 4724 35553 4752 35652
rect 5074 35640 5080 35692
rect 5132 35640 5138 35692
rect 5169 35683 5227 35689
rect 5169 35649 5181 35683
rect 5215 35680 5227 35683
rect 5534 35680 5540 35692
rect 5215 35652 5540 35680
rect 5215 35649 5227 35652
rect 5169 35643 5227 35649
rect 5534 35640 5540 35652
rect 5592 35680 5598 35692
rect 5592 35652 6408 35680
rect 5592 35640 5598 35652
rect 5350 35572 5356 35624
rect 5408 35572 5414 35624
rect 6380 35612 6408 35652
rect 6454 35640 6460 35692
rect 6512 35680 6518 35692
rect 6825 35683 6883 35689
rect 6825 35680 6837 35683
rect 6512 35652 6837 35680
rect 6512 35640 6518 35652
rect 6825 35649 6837 35652
rect 6871 35649 6883 35683
rect 6825 35643 6883 35649
rect 7006 35640 7012 35692
rect 7064 35680 7070 35692
rect 10152 35689 10180 35788
rect 10962 35776 10968 35788
rect 11020 35776 11026 35828
rect 14458 35776 14464 35828
rect 14516 35776 14522 35828
rect 15657 35819 15715 35825
rect 15657 35785 15669 35819
rect 15703 35816 15715 35819
rect 16206 35816 16212 35828
rect 15703 35788 16212 35816
rect 15703 35785 15715 35788
rect 15657 35779 15715 35785
rect 16206 35776 16212 35788
rect 16264 35776 16270 35828
rect 17221 35819 17279 35825
rect 17221 35785 17233 35819
rect 17267 35785 17279 35819
rect 17221 35779 17279 35785
rect 10410 35708 10416 35760
rect 10468 35748 10474 35760
rect 14476 35748 14504 35776
rect 17236 35748 17264 35779
rect 19426 35776 19432 35828
rect 19484 35816 19490 35828
rect 19981 35819 20039 35825
rect 19981 35816 19993 35819
rect 19484 35788 19993 35816
rect 19484 35776 19490 35788
rect 19981 35785 19993 35788
rect 20027 35785 20039 35819
rect 23474 35816 23480 35828
rect 19981 35779 20039 35785
rect 23308 35788 23480 35816
rect 17310 35748 17316 35760
rect 10468 35720 11100 35748
rect 14476 35720 17316 35748
rect 10468 35708 10474 35720
rect 7101 35683 7159 35689
rect 7101 35680 7113 35683
rect 7064 35652 7113 35680
rect 7064 35640 7070 35652
rect 7101 35649 7113 35652
rect 7147 35649 7159 35683
rect 7101 35643 7159 35649
rect 10137 35683 10195 35689
rect 10137 35649 10149 35683
rect 10183 35649 10195 35683
rect 10137 35643 10195 35649
rect 6546 35612 6552 35624
rect 6380 35584 6552 35612
rect 6546 35572 6552 35584
rect 6604 35572 6610 35624
rect 9950 35572 9956 35624
rect 10008 35612 10014 35624
rect 10045 35615 10103 35621
rect 10045 35612 10057 35615
rect 10008 35584 10057 35612
rect 10008 35572 10014 35584
rect 10045 35581 10057 35584
rect 10091 35581 10103 35615
rect 10045 35575 10103 35581
rect 10226 35572 10232 35624
rect 10284 35572 10290 35624
rect 10321 35615 10379 35621
rect 10321 35581 10333 35615
rect 10367 35612 10379 35615
rect 10428 35612 10456 35708
rect 10689 35683 10747 35689
rect 10689 35649 10701 35683
rect 10735 35680 10747 35683
rect 10962 35680 10968 35692
rect 10735 35652 10968 35680
rect 10735 35649 10747 35652
rect 10689 35643 10747 35649
rect 10962 35640 10968 35652
rect 11020 35640 11026 35692
rect 11072 35680 11100 35720
rect 17310 35708 17316 35720
rect 17368 35708 17374 35760
rect 14918 35680 14924 35692
rect 11072 35652 14924 35680
rect 14918 35640 14924 35652
rect 14976 35640 14982 35692
rect 15557 35683 15615 35689
rect 15557 35680 15569 35683
rect 15488 35652 15569 35680
rect 10367 35584 10456 35612
rect 10505 35615 10563 35621
rect 10367 35581 10379 35584
rect 10321 35575 10379 35581
rect 10505 35581 10517 35615
rect 10551 35581 10563 35615
rect 10505 35575 10563 35581
rect 4709 35547 4767 35553
rect 4709 35513 4721 35547
rect 4755 35513 4767 35547
rect 10244 35544 10272 35572
rect 10520 35544 10548 35575
rect 13630 35572 13636 35624
rect 13688 35612 13694 35624
rect 14461 35615 14519 35621
rect 14461 35612 14473 35615
rect 13688 35584 14473 35612
rect 13688 35572 13694 35584
rect 14461 35581 14473 35584
rect 14507 35612 14519 35615
rect 15488 35612 15516 35652
rect 15557 35649 15569 35652
rect 15603 35649 15615 35683
rect 15557 35643 15615 35649
rect 15930 35640 15936 35692
rect 15988 35680 15994 35692
rect 17162 35683 17220 35689
rect 17162 35680 17174 35683
rect 15988 35652 17174 35680
rect 15988 35640 15994 35652
rect 17162 35649 17174 35652
rect 17208 35680 17220 35683
rect 18046 35680 18052 35692
rect 17208 35652 18052 35680
rect 17208 35649 17220 35652
rect 17162 35643 17220 35649
rect 18046 35640 18052 35652
rect 18104 35680 18110 35692
rect 19150 35680 19156 35692
rect 18104 35652 19156 35680
rect 18104 35640 18110 35652
rect 19150 35640 19156 35652
rect 19208 35640 19214 35692
rect 19797 35683 19855 35689
rect 19797 35649 19809 35683
rect 19843 35680 19855 35683
rect 20622 35680 20628 35692
rect 19843 35652 20628 35680
rect 19843 35649 19855 35652
rect 19797 35643 19855 35649
rect 20622 35640 20628 35652
rect 20680 35640 20686 35692
rect 21910 35640 21916 35692
rect 21968 35680 21974 35692
rect 22005 35683 22063 35689
rect 22005 35680 22017 35683
rect 21968 35652 22017 35680
rect 21968 35640 21974 35652
rect 22005 35649 22017 35652
rect 22051 35649 22063 35683
rect 22005 35643 22063 35649
rect 22281 35683 22339 35689
rect 22281 35649 22293 35683
rect 22327 35680 22339 35683
rect 22370 35680 22376 35692
rect 22327 35652 22376 35680
rect 22327 35649 22339 35652
rect 22281 35643 22339 35649
rect 22370 35640 22376 35652
rect 22428 35640 22434 35692
rect 23308 35689 23336 35788
rect 23474 35776 23480 35788
rect 23532 35816 23538 35828
rect 24670 35816 24676 35828
rect 23532 35788 24676 35816
rect 23532 35776 23538 35788
rect 24670 35776 24676 35788
rect 24728 35776 24734 35828
rect 24946 35776 24952 35828
rect 25004 35776 25010 35828
rect 25314 35776 25320 35828
rect 25372 35816 25378 35828
rect 25593 35819 25651 35825
rect 25593 35816 25605 35819
rect 25372 35788 25605 35816
rect 25372 35776 25378 35788
rect 25593 35785 25605 35788
rect 25639 35785 25651 35819
rect 26053 35819 26111 35825
rect 26053 35816 26065 35819
rect 25593 35779 25651 35785
rect 25700 35788 26065 35816
rect 23569 35751 23627 35757
rect 23569 35717 23581 35751
rect 23615 35748 23627 35751
rect 23934 35748 23940 35760
rect 23615 35720 23940 35748
rect 23615 35717 23627 35720
rect 23569 35711 23627 35717
rect 23934 35708 23940 35720
rect 23992 35708 23998 35760
rect 24964 35748 24992 35776
rect 24044 35720 24992 35748
rect 24044 35689 24072 35720
rect 22465 35683 22523 35689
rect 22465 35649 22477 35683
rect 22511 35680 22523 35683
rect 23201 35683 23259 35689
rect 23201 35680 23213 35683
rect 22511 35652 23213 35680
rect 22511 35649 22523 35652
rect 22465 35643 22523 35649
rect 23201 35649 23213 35652
rect 23247 35649 23259 35683
rect 23201 35643 23259 35649
rect 23293 35683 23351 35689
rect 23293 35649 23305 35683
rect 23339 35649 23351 35683
rect 23293 35643 23351 35649
rect 24029 35683 24087 35689
rect 24029 35649 24041 35683
rect 24075 35649 24087 35683
rect 24029 35643 24087 35649
rect 24118 35640 24124 35692
rect 24176 35640 24182 35692
rect 24305 35683 24363 35689
rect 24305 35649 24317 35683
rect 24351 35649 24363 35683
rect 24305 35643 24363 35649
rect 24397 35683 24455 35689
rect 24397 35649 24409 35683
rect 24443 35680 24455 35683
rect 24578 35680 24584 35692
rect 24443 35652 24584 35680
rect 24443 35649 24455 35652
rect 24397 35643 24455 35649
rect 14507 35584 15516 35612
rect 14507 35581 14519 35584
rect 14461 35575 14519 35581
rect 10244 35516 10548 35544
rect 4709 35507 4767 35513
rect 14274 35504 14280 35556
rect 14332 35544 14338 35556
rect 15378 35544 15384 35556
rect 14332 35516 15384 35544
rect 14332 35504 14338 35516
rect 15378 35504 15384 35516
rect 15436 35504 15442 35556
rect 15488 35544 15516 35584
rect 17402 35572 17408 35624
rect 17460 35612 17466 35624
rect 17681 35615 17739 35621
rect 17681 35612 17693 35615
rect 17460 35584 17693 35612
rect 17460 35572 17466 35584
rect 17681 35581 17693 35584
rect 17727 35581 17739 35615
rect 17681 35575 17739 35581
rect 19242 35572 19248 35624
rect 19300 35572 19306 35624
rect 22554 35572 22560 35624
rect 22612 35572 22618 35624
rect 23106 35612 23112 35624
rect 22664 35584 23112 35612
rect 15562 35544 15568 35556
rect 15488 35516 15568 35544
rect 15562 35504 15568 35516
rect 15620 35504 15626 35556
rect 17037 35547 17095 35553
rect 17037 35513 17049 35547
rect 17083 35544 17095 35547
rect 19260 35544 19288 35572
rect 17083 35516 19288 35544
rect 17083 35513 17095 35516
rect 17037 35507 17095 35513
rect 22664 35488 22692 35584
rect 23106 35572 23112 35584
rect 23164 35612 23170 35624
rect 24136 35612 24164 35640
rect 23164 35584 24164 35612
rect 24320 35612 24348 35643
rect 24578 35640 24584 35652
rect 24636 35640 24642 35692
rect 24670 35640 24676 35692
rect 24728 35640 24734 35692
rect 24489 35615 24547 35621
rect 24489 35612 24501 35615
rect 24320 35584 24501 35612
rect 23164 35572 23170 35584
rect 24489 35581 24501 35584
rect 24535 35581 24547 35615
rect 24489 35575 24547 35581
rect 24762 35572 24768 35624
rect 24820 35572 24826 35624
rect 24854 35572 24860 35624
rect 24912 35572 24918 35624
rect 24964 35621 24992 35720
rect 25222 35708 25228 35760
rect 25280 35748 25286 35760
rect 25700 35748 25728 35788
rect 26053 35785 26065 35788
rect 26099 35785 26111 35819
rect 26053 35779 26111 35785
rect 26234 35776 26240 35828
rect 26292 35816 26298 35828
rect 31941 35819 31999 35825
rect 31941 35816 31953 35819
rect 26292 35788 31953 35816
rect 26292 35776 26298 35788
rect 31941 35785 31953 35788
rect 31987 35785 31999 35819
rect 31941 35779 31999 35785
rect 25280 35720 25728 35748
rect 25280 35708 25286 35720
rect 27522 35708 27528 35760
rect 27580 35748 27586 35760
rect 28166 35748 28172 35760
rect 27580 35720 28172 35748
rect 27580 35708 27586 35720
rect 28166 35708 28172 35720
rect 28224 35708 28230 35760
rect 29730 35708 29736 35760
rect 29788 35748 29794 35760
rect 31297 35751 31355 35757
rect 29788 35720 30052 35748
rect 29788 35708 29794 35720
rect 25133 35683 25191 35689
rect 25133 35649 25145 35683
rect 25179 35649 25191 35683
rect 25133 35643 25191 35649
rect 25409 35683 25467 35689
rect 25409 35649 25421 35683
rect 25455 35680 25467 35683
rect 25590 35680 25596 35692
rect 25455 35652 25596 35680
rect 25455 35649 25467 35652
rect 25409 35643 25467 35649
rect 24949 35615 25007 35621
rect 24949 35581 24961 35615
rect 24995 35581 25007 35615
rect 24949 35575 25007 35581
rect 23290 35504 23296 35556
rect 23348 35544 23354 35556
rect 25148 35544 25176 35643
rect 25590 35640 25596 35652
rect 25648 35640 25654 35692
rect 25682 35640 25688 35692
rect 25740 35680 25746 35692
rect 26418 35680 26424 35692
rect 25740 35652 26424 35680
rect 25740 35640 25746 35652
rect 26418 35640 26424 35652
rect 26476 35640 26482 35692
rect 29914 35640 29920 35692
rect 29972 35640 29978 35692
rect 30024 35689 30052 35720
rect 30300 35720 31064 35748
rect 30300 35692 30328 35720
rect 30009 35683 30067 35689
rect 30009 35649 30021 35683
rect 30055 35649 30067 35683
rect 30009 35643 30067 35649
rect 30098 35640 30104 35692
rect 30156 35689 30162 35692
rect 30156 35683 30180 35689
rect 30168 35680 30180 35683
rect 30168 35652 30236 35680
rect 30168 35649 30180 35652
rect 30156 35643 30180 35649
rect 30156 35640 30162 35643
rect 25777 35615 25835 35621
rect 25777 35581 25789 35615
rect 25823 35612 25835 35615
rect 25866 35612 25872 35624
rect 25823 35584 25872 35612
rect 25823 35581 25835 35584
rect 25777 35575 25835 35581
rect 25866 35572 25872 35584
rect 25924 35612 25930 35624
rect 26050 35612 26056 35624
rect 25924 35584 26056 35612
rect 25924 35572 25930 35584
rect 26050 35572 26056 35584
rect 26108 35612 26114 35624
rect 27522 35612 27528 35624
rect 26108 35584 27528 35612
rect 26108 35572 26114 35584
rect 27522 35572 27528 35584
rect 27580 35572 27586 35624
rect 29270 35572 29276 35624
rect 29328 35612 29334 35624
rect 29822 35612 29828 35624
rect 29328 35584 29828 35612
rect 29328 35572 29334 35584
rect 29822 35572 29828 35584
rect 29880 35572 29886 35624
rect 30208 35612 30236 35652
rect 30282 35640 30288 35692
rect 30340 35640 30346 35692
rect 30929 35683 30987 35689
rect 30929 35649 30941 35683
rect 30975 35649 30987 35683
rect 31036 35680 31064 35720
rect 31297 35717 31309 35751
rect 31343 35748 31355 35751
rect 31846 35748 31852 35760
rect 31343 35720 31852 35748
rect 31343 35717 31355 35720
rect 31297 35711 31355 35717
rect 31846 35708 31852 35720
rect 31904 35748 31910 35760
rect 31904 35720 31984 35748
rect 31904 35708 31910 35720
rect 31110 35689 31116 35692
rect 31104 35680 31116 35689
rect 31036 35652 31116 35680
rect 30929 35643 30987 35649
rect 31104 35643 31116 35652
rect 30944 35612 30972 35643
rect 31110 35640 31116 35643
rect 31168 35640 31174 35692
rect 31205 35683 31263 35689
rect 31205 35649 31217 35683
rect 31251 35680 31263 35683
rect 31389 35683 31447 35689
rect 31251 35652 31340 35680
rect 31251 35649 31263 35652
rect 31205 35643 31263 35649
rect 31312 35612 31340 35652
rect 31389 35649 31401 35683
rect 31435 35680 31447 35683
rect 31754 35680 31760 35692
rect 31435 35652 31760 35680
rect 31435 35649 31447 35652
rect 31389 35643 31447 35649
rect 31754 35640 31760 35652
rect 31812 35640 31818 35692
rect 31956 35680 31984 35720
rect 32122 35708 32128 35760
rect 32180 35748 32186 35760
rect 32217 35751 32275 35757
rect 32217 35748 32229 35751
rect 32180 35720 32229 35748
rect 32180 35708 32186 35720
rect 32217 35717 32229 35720
rect 32263 35717 32275 35751
rect 32217 35711 32275 35717
rect 33134 35708 33140 35760
rect 33192 35748 33198 35760
rect 33192 35720 34560 35748
rect 33192 35708 33198 35720
rect 34532 35692 34560 35720
rect 32769 35683 32827 35689
rect 32769 35680 32781 35683
rect 31956 35652 32781 35680
rect 32769 35649 32781 35652
rect 32815 35649 32827 35683
rect 32769 35643 32827 35649
rect 33505 35683 33563 35689
rect 33505 35649 33517 35683
rect 33551 35680 33563 35683
rect 34149 35683 34207 35689
rect 34149 35680 34161 35683
rect 33551 35652 34161 35680
rect 33551 35649 33563 35652
rect 33505 35643 33563 35649
rect 34149 35649 34161 35652
rect 34195 35680 34207 35683
rect 34195 35652 34284 35680
rect 34195 35649 34207 35652
rect 34149 35643 34207 35649
rect 31481 35615 31539 35621
rect 31481 35612 31493 35615
rect 30208 35584 31248 35612
rect 31312 35584 31493 35612
rect 29641 35547 29699 35553
rect 23348 35516 25820 35544
rect 23348 35504 23354 35516
rect 6641 35479 6699 35485
rect 6641 35445 6653 35479
rect 6687 35476 6699 35479
rect 6822 35476 6828 35488
rect 6687 35448 6828 35476
rect 6687 35445 6699 35448
rect 6641 35439 6699 35445
rect 6822 35436 6828 35448
rect 6880 35436 6886 35488
rect 9858 35436 9864 35488
rect 9916 35436 9922 35488
rect 10134 35436 10140 35488
rect 10192 35476 10198 35488
rect 10873 35479 10931 35485
rect 10873 35476 10885 35479
rect 10192 35448 10885 35476
rect 10192 35436 10198 35448
rect 10873 35445 10885 35448
rect 10919 35445 10931 35479
rect 10873 35439 10931 35445
rect 15102 35436 15108 35488
rect 15160 35436 15166 35488
rect 16482 35436 16488 35488
rect 16540 35476 16546 35488
rect 17218 35476 17224 35488
rect 16540 35448 17224 35476
rect 16540 35436 16546 35448
rect 17218 35436 17224 35448
rect 17276 35436 17282 35488
rect 17589 35479 17647 35485
rect 17589 35445 17601 35479
rect 17635 35476 17647 35479
rect 17954 35476 17960 35488
rect 17635 35448 17960 35476
rect 17635 35445 17647 35448
rect 17589 35439 17647 35445
rect 17954 35436 17960 35448
rect 18012 35436 18018 35488
rect 21818 35436 21824 35488
rect 21876 35436 21882 35488
rect 22646 35436 22652 35488
rect 22704 35436 22710 35488
rect 23845 35479 23903 35485
rect 23845 35445 23857 35479
rect 23891 35476 23903 35479
rect 24394 35476 24400 35488
rect 23891 35448 24400 35476
rect 23891 35445 23903 35448
rect 23845 35439 23903 35445
rect 24394 35436 24400 35448
rect 24452 35436 24458 35488
rect 24578 35436 24584 35488
rect 24636 35476 24642 35488
rect 25130 35476 25136 35488
rect 24636 35448 25136 35476
rect 24636 35436 24642 35448
rect 25130 35436 25136 35448
rect 25188 35436 25194 35488
rect 25682 35436 25688 35488
rect 25740 35436 25746 35488
rect 25792 35476 25820 35516
rect 29641 35513 29653 35547
rect 29687 35544 29699 35547
rect 31110 35544 31116 35556
rect 29687 35516 31116 35544
rect 29687 35513 29699 35516
rect 29641 35507 29699 35513
rect 31110 35504 31116 35516
rect 31168 35504 31174 35556
rect 31220 35544 31248 35584
rect 31481 35581 31493 35584
rect 31527 35612 31539 35615
rect 32122 35612 32128 35624
rect 31527 35584 32128 35612
rect 31527 35581 31539 35584
rect 31481 35575 31539 35581
rect 32122 35572 32128 35584
rect 32180 35612 32186 35624
rect 33520 35612 33548 35643
rect 34256 35624 34284 35652
rect 34514 35640 34520 35692
rect 34572 35640 34578 35692
rect 34701 35683 34759 35689
rect 34701 35680 34713 35683
rect 34624 35652 34713 35680
rect 32180 35584 33548 35612
rect 32180 35572 32186 35584
rect 34238 35572 34244 35624
rect 34296 35572 34302 35624
rect 34624 35621 34652 35652
rect 34701 35649 34713 35652
rect 34747 35649 34759 35683
rect 34701 35643 34759 35649
rect 34609 35615 34667 35621
rect 34609 35581 34621 35615
rect 34655 35581 34667 35615
rect 34885 35615 34943 35621
rect 34885 35612 34897 35615
rect 34609 35575 34667 35581
rect 34716 35584 34897 35612
rect 31849 35547 31907 35553
rect 31849 35544 31861 35547
rect 31220 35516 31861 35544
rect 31849 35513 31861 35516
rect 31895 35544 31907 35547
rect 31938 35544 31944 35556
rect 31895 35516 31944 35544
rect 31895 35513 31907 35516
rect 31849 35507 31907 35513
rect 31938 35504 31944 35516
rect 31996 35504 32002 35556
rect 33778 35504 33784 35556
rect 33836 35504 33842 35556
rect 34716 35488 34744 35584
rect 34885 35581 34897 35584
rect 34931 35581 34943 35615
rect 34885 35575 34943 35581
rect 30466 35476 30472 35488
rect 25792 35448 30472 35476
rect 30466 35436 30472 35448
rect 30524 35436 30530 35488
rect 31018 35436 31024 35488
rect 31076 35436 31082 35488
rect 31386 35436 31392 35488
rect 31444 35476 31450 35488
rect 32309 35479 32367 35485
rect 32309 35476 32321 35479
rect 31444 35448 32321 35476
rect 31444 35436 31450 35448
rect 32309 35445 32321 35448
rect 32355 35445 32367 35479
rect 32309 35439 32367 35445
rect 33965 35479 34023 35485
rect 33965 35445 33977 35479
rect 34011 35476 34023 35479
rect 34146 35476 34152 35488
rect 34011 35448 34152 35476
rect 34011 35445 34023 35448
rect 33965 35439 34023 35445
rect 34146 35436 34152 35448
rect 34204 35436 34210 35488
rect 34330 35436 34336 35488
rect 34388 35436 34394 35488
rect 34698 35436 34704 35488
rect 34756 35436 34762 35488
rect 1104 35386 41400 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 41400 35386
rect 1104 35312 41400 35334
rect 7193 35275 7251 35281
rect 7193 35241 7205 35275
rect 7239 35272 7251 35275
rect 7742 35272 7748 35284
rect 7239 35244 7748 35272
rect 7239 35241 7251 35244
rect 7193 35235 7251 35241
rect 7742 35232 7748 35244
rect 7800 35232 7806 35284
rect 8665 35275 8723 35281
rect 8665 35241 8677 35275
rect 8711 35272 8723 35275
rect 8754 35272 8760 35284
rect 8711 35244 8760 35272
rect 8711 35241 8723 35244
rect 8665 35235 8723 35241
rect 8754 35232 8760 35244
rect 8812 35232 8818 35284
rect 9769 35275 9827 35281
rect 9769 35241 9781 35275
rect 9815 35272 9827 35275
rect 9858 35272 9864 35284
rect 9815 35244 9864 35272
rect 9815 35241 9827 35244
rect 9769 35235 9827 35241
rect 9858 35232 9864 35244
rect 9916 35232 9922 35284
rect 13538 35272 13544 35284
rect 12406 35244 13544 35272
rect 9953 35207 10011 35213
rect 9953 35173 9965 35207
rect 9999 35173 10011 35207
rect 9953 35167 10011 35173
rect 4706 35096 4712 35148
rect 4764 35136 4770 35148
rect 7009 35139 7067 35145
rect 7009 35136 7021 35139
rect 4764 35108 7021 35136
rect 4764 35096 4770 35108
rect 7009 35105 7021 35108
rect 7055 35136 7067 35139
rect 7558 35136 7564 35148
rect 7055 35108 7564 35136
rect 7055 35105 7067 35108
rect 7009 35099 7067 35105
rect 7558 35096 7564 35108
rect 7616 35096 7622 35148
rect 8389 35139 8447 35145
rect 8389 35105 8401 35139
rect 8435 35136 8447 35139
rect 9968 35136 9996 35167
rect 8435 35108 9996 35136
rect 8435 35105 8447 35108
rect 8389 35099 8447 35105
rect 11514 35096 11520 35148
rect 11572 35136 11578 35148
rect 12250 35136 12256 35148
rect 11572 35108 12256 35136
rect 11572 35096 11578 35108
rect 12250 35096 12256 35108
rect 12308 35096 12314 35148
rect 4062 35028 4068 35080
rect 4120 35068 4126 35080
rect 6917 35071 6975 35077
rect 6917 35068 6929 35071
rect 4120 35040 6929 35068
rect 4120 35028 4126 35040
rect 6917 35037 6929 35040
rect 6963 35068 6975 35071
rect 7282 35068 7288 35080
rect 6963 35040 7288 35068
rect 6963 35037 6975 35040
rect 6917 35031 6975 35037
rect 7282 35028 7288 35040
rect 7340 35028 7346 35080
rect 8297 35071 8355 35077
rect 8297 35037 8309 35071
rect 8343 35068 8355 35071
rect 10042 35068 10048 35080
rect 8343 35040 10048 35068
rect 8343 35037 8355 35040
rect 8297 35031 8355 35037
rect 10042 35028 10048 35040
rect 10100 35028 10106 35080
rect 10134 35028 10140 35080
rect 10192 35028 10198 35080
rect 10413 35071 10471 35077
rect 10413 35037 10425 35071
rect 10459 35068 10471 35071
rect 10594 35068 10600 35080
rect 10459 35040 10600 35068
rect 10459 35037 10471 35040
rect 10413 35031 10471 35037
rect 10594 35028 10600 35040
rect 10652 35068 10658 35080
rect 11057 35071 11115 35077
rect 11057 35068 11069 35071
rect 10652 35040 11069 35068
rect 10652 35028 10658 35040
rect 11057 35037 11069 35040
rect 11103 35037 11115 35071
rect 11057 35031 11115 35037
rect 9585 35003 9643 35009
rect 9585 34969 9597 35003
rect 9631 35000 9643 35003
rect 10502 35000 10508 35012
rect 9631 34972 10508 35000
rect 9631 34969 9643 34972
rect 9585 34963 9643 34969
rect 10502 34960 10508 34972
rect 10560 35000 10566 35012
rect 10873 35003 10931 35009
rect 10873 35000 10885 35003
rect 10560 34972 10885 35000
rect 10560 34960 10566 34972
rect 10873 34969 10885 34972
rect 10919 34969 10931 35003
rect 11072 35000 11100 35031
rect 11238 35028 11244 35080
rect 11296 35068 11302 35080
rect 11333 35071 11391 35077
rect 11333 35068 11345 35071
rect 11296 35040 11345 35068
rect 11296 35028 11302 35040
rect 11333 35037 11345 35040
rect 11379 35037 11391 35071
rect 11333 35031 11391 35037
rect 11698 35028 11704 35080
rect 11756 35028 11762 35080
rect 11885 35071 11943 35077
rect 11885 35037 11897 35071
rect 11931 35068 11943 35071
rect 12406 35068 12434 35244
rect 13538 35232 13544 35244
rect 13596 35272 13602 35284
rect 13596 35244 15516 35272
rect 13596 35232 13602 35244
rect 15488 35204 15516 35244
rect 15562 35232 15568 35284
rect 15620 35272 15626 35284
rect 15933 35275 15991 35281
rect 15933 35272 15945 35275
rect 15620 35244 15945 35272
rect 15620 35232 15626 35244
rect 15933 35241 15945 35244
rect 15979 35241 15991 35275
rect 15933 35235 15991 35241
rect 16761 35275 16819 35281
rect 16761 35241 16773 35275
rect 16807 35272 16819 35275
rect 17494 35272 17500 35284
rect 16807 35244 17500 35272
rect 16807 35241 16819 35244
rect 16761 35235 16819 35241
rect 17494 35232 17500 35244
rect 17552 35232 17558 35284
rect 21082 35232 21088 35284
rect 21140 35272 21146 35284
rect 23014 35272 23020 35284
rect 21140 35244 23020 35272
rect 21140 35232 21146 35244
rect 23014 35232 23020 35244
rect 23072 35232 23078 35284
rect 23201 35275 23259 35281
rect 23201 35241 23213 35275
rect 23247 35272 23259 35275
rect 23477 35275 23535 35281
rect 23477 35272 23489 35275
rect 23247 35244 23489 35272
rect 23247 35241 23259 35244
rect 23201 35235 23259 35241
rect 23477 35241 23489 35244
rect 23523 35241 23535 35275
rect 23477 35235 23535 35241
rect 23845 35275 23903 35281
rect 23845 35241 23857 35275
rect 23891 35272 23903 35275
rect 23891 35244 24946 35272
rect 23891 35241 23903 35244
rect 23845 35235 23903 35241
rect 15838 35204 15844 35216
rect 15488 35176 15844 35204
rect 15838 35164 15844 35176
rect 15896 35164 15902 35216
rect 23382 35204 23388 35216
rect 22204 35176 23388 35204
rect 14185 35139 14243 35145
rect 14185 35105 14197 35139
rect 14231 35136 14243 35139
rect 16298 35136 16304 35148
rect 14231 35108 16304 35136
rect 14231 35105 14243 35108
rect 14185 35099 14243 35105
rect 16298 35096 16304 35108
rect 16356 35096 16362 35148
rect 16393 35139 16451 35145
rect 16393 35105 16405 35139
rect 16439 35105 16451 35139
rect 20809 35139 20867 35145
rect 20809 35136 20821 35139
rect 16393 35099 16451 35105
rect 19904 35108 20821 35136
rect 15746 35068 15752 35080
rect 11931 35040 12434 35068
rect 15594 35040 15752 35068
rect 11931 35037 11943 35040
rect 11885 35031 11943 35037
rect 11900 35000 11928 35031
rect 15746 35028 15752 35040
rect 15804 35068 15810 35080
rect 16206 35068 16212 35080
rect 15804 35040 16212 35068
rect 15804 35028 15810 35040
rect 16206 35028 16212 35040
rect 16264 35028 16270 35080
rect 11072 34972 11928 35000
rect 14461 35003 14519 35009
rect 10873 34963 10931 34969
rect 14461 34969 14473 35003
rect 14507 35000 14519 35003
rect 14550 35000 14556 35012
rect 14507 34972 14556 35000
rect 14507 34969 14519 34972
rect 14461 34963 14519 34969
rect 14550 34960 14556 34972
rect 14608 34960 14614 35012
rect 16408 35000 16436 35099
rect 16482 35028 16488 35080
rect 16540 35028 16546 35080
rect 19426 35028 19432 35080
rect 19484 35068 19490 35080
rect 19904 35077 19932 35108
rect 20809 35105 20821 35108
rect 20855 35105 20867 35139
rect 20809 35099 20867 35105
rect 21085 35139 21143 35145
rect 21085 35105 21097 35139
rect 21131 35136 21143 35139
rect 21818 35136 21824 35148
rect 21131 35108 21824 35136
rect 21131 35105 21143 35108
rect 21085 35099 21143 35105
rect 21818 35096 21824 35108
rect 21876 35096 21882 35148
rect 19889 35071 19947 35077
rect 19889 35068 19901 35071
rect 19484 35040 19901 35068
rect 19484 35028 19490 35040
rect 19889 35037 19901 35040
rect 19935 35037 19947 35071
rect 19889 35031 19947 35037
rect 20073 35071 20131 35077
rect 20073 35037 20085 35071
rect 20119 35068 20131 35071
rect 20119 35040 20392 35068
rect 22204 35054 22232 35176
rect 23382 35164 23388 35176
rect 23440 35164 23446 35216
rect 23566 35164 23572 35216
rect 23624 35204 23630 35216
rect 24578 35204 24584 35216
rect 23624 35176 24584 35204
rect 23624 35164 23630 35176
rect 24578 35164 24584 35176
rect 24636 35164 24642 35216
rect 24918 35204 24946 35244
rect 25130 35232 25136 35284
rect 25188 35272 25194 35284
rect 25777 35275 25835 35281
rect 25777 35272 25789 35275
rect 25188 35244 25789 35272
rect 25188 35232 25194 35244
rect 25777 35241 25789 35244
rect 25823 35241 25835 35275
rect 25777 35235 25835 35241
rect 26418 35232 26424 35284
rect 26476 35232 26482 35284
rect 26786 35232 26792 35284
rect 26844 35232 26850 35284
rect 27062 35232 27068 35284
rect 27120 35232 27126 35284
rect 27154 35232 27160 35284
rect 27212 35232 27218 35284
rect 29178 35232 29184 35284
rect 29236 35232 29242 35284
rect 31018 35232 31024 35284
rect 31076 35232 31082 35284
rect 31110 35232 31116 35284
rect 31168 35232 31174 35284
rect 32125 35275 32183 35281
rect 32125 35241 32137 35275
rect 32171 35241 32183 35275
rect 32125 35235 32183 35241
rect 26436 35204 26464 35232
rect 27338 35204 27344 35216
rect 24918 35176 25324 35204
rect 26436 35176 27344 35204
rect 23937 35139 23995 35145
rect 23937 35136 23949 35139
rect 22388 35108 23949 35136
rect 20119 35037 20131 35040
rect 20073 35031 20131 35037
rect 20364 35012 20392 35040
rect 15764 34972 16436 35000
rect 9766 34892 9772 34944
rect 9824 34941 9830 34944
rect 9824 34935 9843 34941
rect 9831 34901 9843 34935
rect 9824 34895 9843 34901
rect 9824 34892 9830 34895
rect 9950 34892 9956 34944
rect 10008 34932 10014 34944
rect 10229 34935 10287 34941
rect 10229 34932 10241 34935
rect 10008 34904 10241 34932
rect 10008 34892 10014 34904
rect 10229 34901 10241 34904
rect 10275 34901 10287 34935
rect 10229 34895 10287 34901
rect 10318 34892 10324 34944
rect 10376 34892 10382 34944
rect 11241 34935 11299 34941
rect 11241 34901 11253 34935
rect 11287 34932 11299 34935
rect 11606 34932 11612 34944
rect 11287 34904 11612 34932
rect 11287 34901 11299 34904
rect 11241 34895 11299 34901
rect 11606 34892 11612 34904
rect 11664 34892 11670 34944
rect 11882 34892 11888 34944
rect 11940 34892 11946 34944
rect 14090 34892 14096 34944
rect 14148 34932 14154 34944
rect 15764 34932 15792 34972
rect 20346 34960 20352 35012
rect 20404 34960 20410 35012
rect 14148 34904 15792 34932
rect 14148 34892 14154 34904
rect 20254 34892 20260 34944
rect 20312 34892 20318 34944
rect 21726 34892 21732 34944
rect 21784 34932 21790 34944
rect 22388 34932 22416 35108
rect 23937 35105 23949 35108
rect 23983 35136 23995 35139
rect 24210 35136 24216 35148
rect 23983 35108 24216 35136
rect 23983 35105 23995 35108
rect 23937 35099 23995 35105
rect 24210 35096 24216 35108
rect 24268 35096 24274 35148
rect 24320 35108 24716 35136
rect 23106 35028 23112 35080
rect 23164 35028 23170 35080
rect 23198 35028 23204 35080
rect 23256 35028 23262 35080
rect 23661 35071 23719 35077
rect 23661 35037 23673 35071
rect 23707 35037 23719 35071
rect 23661 35031 23719 35037
rect 22922 34960 22928 35012
rect 22980 34960 22986 35012
rect 23676 35000 23704 35031
rect 24118 35028 24124 35080
rect 24176 35028 24182 35080
rect 24136 35000 24164 35028
rect 23676 34972 24164 35000
rect 24320 34944 24348 35108
rect 24394 35028 24400 35080
rect 24452 35028 24458 35080
rect 24578 35077 24584 35080
rect 24545 35071 24584 35077
rect 24545 35037 24557 35071
rect 24545 35031 24584 35037
rect 24578 35028 24584 35031
rect 24636 35028 24642 35080
rect 24688 35077 24716 35108
rect 25296 35080 25324 35176
rect 27338 35164 27344 35176
rect 27396 35204 27402 35216
rect 27525 35207 27583 35213
rect 27525 35204 27537 35207
rect 27396 35176 27537 35204
rect 27396 35164 27402 35176
rect 27525 35173 27537 35176
rect 27571 35173 27583 35207
rect 31036 35204 31064 35232
rect 27525 35167 27583 35173
rect 30944 35176 31064 35204
rect 25958 35136 25964 35148
rect 25516 35108 25964 35136
rect 25516 35080 25544 35108
rect 25958 35096 25964 35108
rect 26016 35096 26022 35148
rect 26053 35139 26111 35145
rect 26053 35105 26065 35139
rect 26099 35136 26111 35139
rect 26697 35139 26755 35145
rect 26697 35136 26709 35139
rect 26099 35108 26709 35136
rect 26099 35105 26111 35108
rect 26053 35099 26111 35105
rect 26697 35105 26709 35108
rect 26743 35105 26755 35139
rect 29546 35136 29552 35148
rect 26697 35099 26755 35105
rect 26804 35108 29552 35136
rect 24673 35071 24731 35077
rect 24673 35037 24685 35071
rect 24719 35037 24731 35071
rect 24673 35031 24731 35037
rect 24903 35071 24961 35077
rect 24903 35037 24915 35071
rect 24949 35068 24961 35071
rect 25038 35068 25044 35080
rect 24949 35040 25044 35068
rect 24949 35037 24961 35040
rect 24903 35031 24961 35037
rect 25038 35028 25044 35040
rect 25096 35028 25102 35080
rect 25130 35028 25136 35080
rect 25188 35028 25194 35080
rect 25296 35077 25320 35080
rect 25281 35071 25320 35077
rect 25281 35037 25293 35071
rect 25281 35031 25320 35037
rect 25314 35028 25320 35031
rect 25372 35028 25378 35080
rect 25406 35028 25412 35080
rect 25464 35028 25470 35080
rect 25498 35028 25504 35080
rect 25556 35028 25562 35080
rect 25639 35071 25697 35077
rect 25639 35037 25651 35071
rect 25685 35068 25697 35071
rect 26142 35068 26148 35080
rect 25685 35040 26148 35068
rect 25685 35037 25697 35040
rect 25639 35031 25697 35037
rect 26142 35028 26148 35040
rect 26200 35028 26206 35080
rect 26234 35028 26240 35080
rect 26292 35028 26298 35080
rect 26513 35071 26571 35077
rect 26513 35037 26525 35071
rect 26559 35068 26571 35071
rect 26804 35068 26832 35108
rect 29546 35096 29552 35108
rect 29604 35096 29610 35148
rect 26559 35040 26832 35068
rect 26881 35071 26939 35077
rect 26559 35037 26571 35040
rect 26513 35031 26571 35037
rect 26881 35037 26893 35071
rect 26927 35037 26939 35071
rect 26881 35031 26939 35037
rect 24765 35003 24823 35009
rect 24765 34969 24777 35003
rect 24811 35000 24823 35003
rect 24811 34972 25452 35000
rect 24811 34969 24823 34972
rect 24765 34963 24823 34969
rect 25424 34944 25452 34972
rect 25774 34960 25780 35012
rect 25832 35000 25838 35012
rect 26528 35000 26556 35031
rect 25832 34972 26556 35000
rect 25832 34960 25838 34972
rect 26602 34960 26608 35012
rect 26660 34960 26666 35012
rect 21784 34904 22416 34932
rect 21784 34892 21790 34904
rect 22554 34892 22560 34944
rect 22612 34892 22618 34944
rect 23385 34935 23443 34941
rect 23385 34901 23397 34935
rect 23431 34932 23443 34935
rect 23658 34932 23664 34944
rect 23431 34904 23664 34932
rect 23431 34901 23443 34904
rect 23385 34895 23443 34901
rect 23658 34892 23664 34904
rect 23716 34892 23722 34944
rect 24302 34892 24308 34944
rect 24360 34892 24366 34944
rect 25038 34892 25044 34944
rect 25096 34892 25102 34944
rect 25406 34892 25412 34944
rect 25464 34932 25470 34944
rect 26234 34932 26240 34944
rect 25464 34904 26240 34932
rect 25464 34892 25470 34904
rect 26234 34892 26240 34904
rect 26292 34892 26298 34944
rect 26326 34892 26332 34944
rect 26384 34932 26390 34944
rect 26896 34932 26924 35031
rect 26970 35028 26976 35080
rect 27028 35068 27034 35080
rect 27341 35071 27399 35077
rect 27341 35068 27353 35071
rect 27028 35040 27353 35068
rect 27028 35028 27034 35040
rect 27341 35037 27353 35040
rect 27387 35037 27399 35071
rect 27341 35031 27399 35037
rect 27522 35028 27528 35080
rect 27580 35068 27586 35080
rect 27617 35071 27675 35077
rect 27617 35068 27629 35071
rect 27580 35040 27629 35068
rect 27580 35028 27586 35040
rect 27617 35037 27629 35040
rect 27663 35068 27675 35071
rect 28902 35068 28908 35080
rect 27663 35040 28908 35068
rect 27663 35037 27675 35040
rect 27617 35031 27675 35037
rect 28902 35028 28908 35040
rect 28960 35028 28966 35080
rect 28994 35028 29000 35080
rect 29052 35068 29058 35080
rect 30944 35077 30972 35176
rect 31018 35096 31024 35148
rect 31076 35096 31082 35148
rect 29089 35071 29147 35077
rect 29089 35068 29101 35071
rect 29052 35040 29101 35068
rect 29052 35028 29058 35040
rect 29089 35037 29101 35040
rect 29135 35037 29147 35071
rect 29089 35031 29147 35037
rect 30837 35071 30895 35077
rect 30837 35037 30849 35071
rect 30883 35037 30895 35071
rect 30837 35031 30895 35037
rect 30929 35071 30987 35077
rect 30929 35037 30941 35071
rect 30975 35037 30987 35071
rect 31128 35068 31156 35232
rect 32140 35204 32168 35235
rect 33502 35232 33508 35284
rect 33560 35232 33566 35284
rect 34698 35272 34704 35284
rect 33612 35244 34704 35272
rect 33612 35204 33640 35244
rect 34698 35232 34704 35244
rect 34756 35232 34762 35284
rect 36078 35232 36084 35284
rect 36136 35232 36142 35284
rect 32140 35176 33640 35204
rect 34238 35164 34244 35216
rect 34296 35204 34302 35216
rect 36096 35204 36124 35232
rect 34296 35176 36124 35204
rect 34296 35164 34302 35176
rect 32033 35139 32091 35145
rect 32033 35136 32045 35139
rect 31588 35108 32045 35136
rect 31205 35071 31263 35077
rect 31205 35068 31217 35071
rect 31128 35040 31217 35068
rect 30929 35031 30987 35037
rect 31205 35037 31217 35040
rect 31251 35037 31263 35071
rect 31205 35031 31263 35037
rect 28810 34960 28816 35012
rect 28868 35000 28874 35012
rect 29730 35000 29736 35012
rect 28868 34972 29736 35000
rect 28868 34960 28874 34972
rect 29730 34960 29736 34972
rect 29788 34960 29794 35012
rect 30852 35000 30880 35031
rect 31386 35028 31392 35080
rect 31444 35028 31450 35080
rect 31588 35012 31616 35108
rect 32033 35105 32045 35108
rect 32079 35105 32091 35139
rect 32033 35099 32091 35105
rect 32582 35096 32588 35148
rect 32640 35136 32646 35148
rect 33778 35136 33784 35148
rect 32640 35108 33784 35136
rect 32640 35096 32646 35108
rect 33778 35096 33784 35108
rect 33836 35136 33842 35148
rect 33873 35139 33931 35145
rect 33873 35136 33885 35139
rect 33836 35108 33885 35136
rect 33836 35096 33842 35108
rect 33873 35105 33885 35108
rect 33919 35136 33931 35139
rect 33919 35108 34100 35136
rect 33919 35105 33931 35108
rect 33873 35099 33931 35105
rect 31941 35071 31999 35077
rect 31941 35037 31953 35071
rect 31987 35068 31999 35071
rect 32858 35068 32864 35080
rect 31987 35040 32864 35068
rect 31987 35037 31999 35040
rect 31941 35031 31999 35037
rect 32858 35028 32864 35040
rect 32916 35028 32922 35080
rect 33413 35071 33471 35077
rect 33413 35037 33425 35071
rect 33459 35068 33471 35071
rect 33962 35068 33968 35080
rect 33459 35040 33968 35068
rect 33459 35037 33471 35040
rect 33413 35031 33471 35037
rect 33962 35028 33968 35040
rect 34020 35028 34026 35080
rect 34072 35068 34100 35108
rect 34330 35068 34336 35080
rect 34072 35040 34336 35068
rect 34330 35028 34336 35040
rect 34388 35068 34394 35080
rect 35989 35071 36047 35077
rect 35989 35068 36001 35071
rect 34388 35040 36001 35068
rect 34388 35028 34394 35040
rect 35989 35037 36001 35040
rect 36035 35068 36047 35071
rect 36035 35040 36860 35068
rect 36035 35037 36047 35040
rect 35989 35031 36047 35037
rect 30852 34972 31340 35000
rect 26384 34904 26924 34932
rect 26384 34892 26390 34904
rect 27246 34892 27252 34944
rect 27304 34932 27310 34944
rect 29454 34932 29460 34944
rect 27304 34904 29460 34932
rect 27304 34892 27310 34904
rect 29454 34892 29460 34904
rect 29512 34932 29518 34944
rect 30006 34932 30012 34944
rect 29512 34904 30012 34932
rect 29512 34892 29518 34904
rect 30006 34892 30012 34904
rect 30064 34892 30070 34944
rect 31110 34892 31116 34944
rect 31168 34892 31174 34944
rect 31312 34932 31340 34972
rect 31570 34960 31576 35012
rect 31628 34960 31634 35012
rect 31662 34960 31668 35012
rect 31720 34960 31726 35012
rect 31754 34960 31760 35012
rect 31812 35000 31818 35012
rect 32582 35000 32588 35012
rect 31812 34972 32588 35000
rect 31812 34960 31818 34972
rect 32582 34960 32588 34972
rect 32640 34960 32646 35012
rect 36832 34944 36860 35040
rect 32309 34935 32367 34941
rect 32309 34932 32321 34935
rect 31312 34904 32321 34932
rect 32309 34901 32321 34904
rect 32355 34901 32367 34935
rect 32309 34895 32367 34901
rect 34054 34892 34060 34944
rect 34112 34932 34118 34944
rect 34333 34935 34391 34941
rect 34333 34932 34345 34935
rect 34112 34904 34345 34932
rect 34112 34892 34118 34904
rect 34333 34901 34345 34904
rect 34379 34901 34391 34935
rect 34333 34895 34391 34901
rect 36354 34892 36360 34944
rect 36412 34932 36418 34944
rect 36449 34935 36507 34941
rect 36449 34932 36461 34935
rect 36412 34904 36461 34932
rect 36412 34892 36418 34904
rect 36449 34901 36461 34904
rect 36495 34901 36507 34935
rect 36449 34895 36507 34901
rect 36814 34892 36820 34944
rect 36872 34892 36878 34944
rect 1104 34842 41400 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 41400 34842
rect 1104 34768 41400 34790
rect 1026 34688 1032 34740
rect 1084 34728 1090 34740
rect 2041 34731 2099 34737
rect 2041 34728 2053 34731
rect 1084 34700 2053 34728
rect 1084 34688 1090 34700
rect 2041 34697 2053 34700
rect 2087 34697 2099 34731
rect 2041 34691 2099 34697
rect 7558 34688 7564 34740
rect 7616 34728 7622 34740
rect 8757 34731 8815 34737
rect 8757 34728 8769 34731
rect 7616 34700 8769 34728
rect 7616 34688 7622 34700
rect 8757 34697 8769 34700
rect 8803 34697 8815 34731
rect 8757 34691 8815 34697
rect 9674 34688 9680 34740
rect 9732 34688 9738 34740
rect 10318 34688 10324 34740
rect 10376 34688 10382 34740
rect 10962 34688 10968 34740
rect 11020 34688 11026 34740
rect 11238 34688 11244 34740
rect 11296 34728 11302 34740
rect 11885 34731 11943 34737
rect 11885 34728 11897 34731
rect 11296 34700 11897 34728
rect 11296 34688 11302 34700
rect 11885 34697 11897 34700
rect 11931 34697 11943 34731
rect 11885 34691 11943 34697
rect 11977 34731 12035 34737
rect 11977 34697 11989 34731
rect 12023 34728 12035 34731
rect 12023 34700 12848 34728
rect 12023 34697 12035 34700
rect 11977 34691 12035 34697
rect 6546 34620 6552 34672
rect 6604 34660 6610 34672
rect 7009 34663 7067 34669
rect 7009 34660 7021 34663
rect 6604 34632 7021 34660
rect 6604 34620 6610 34632
rect 7009 34629 7021 34632
rect 7055 34660 7067 34663
rect 9217 34663 9275 34669
rect 7055 34632 7512 34660
rect 7055 34629 7067 34632
rect 7009 34623 7067 34629
rect 1854 34552 1860 34604
rect 1912 34552 1918 34604
rect 6825 34595 6883 34601
rect 6825 34561 6837 34595
rect 6871 34592 6883 34595
rect 6914 34592 6920 34604
rect 6871 34564 6920 34592
rect 6871 34561 6883 34564
rect 6825 34555 6883 34561
rect 6914 34552 6920 34564
rect 6972 34592 6978 34604
rect 7484 34601 7512 34632
rect 9217 34629 9229 34663
rect 9263 34660 9275 34663
rect 10336 34660 10364 34688
rect 9263 34632 10364 34660
rect 9263 34629 9275 34632
rect 9217 34623 9275 34629
rect 9600 34601 9628 34632
rect 11514 34620 11520 34672
rect 11572 34620 11578 34672
rect 11733 34663 11791 34669
rect 11733 34629 11745 34663
rect 11779 34660 11791 34663
rect 12066 34660 12072 34672
rect 11779 34632 12072 34660
rect 11779 34629 11791 34632
rect 11733 34623 11791 34629
rect 12066 34620 12072 34632
rect 12124 34620 12130 34672
rect 12820 34660 12848 34700
rect 13078 34688 13084 34740
rect 13136 34728 13142 34740
rect 13173 34731 13231 34737
rect 13173 34728 13185 34731
rect 13136 34700 13185 34728
rect 13136 34688 13142 34700
rect 13173 34697 13185 34700
rect 13219 34697 13231 34731
rect 14274 34728 14280 34740
rect 13173 34691 13231 34697
rect 14200 34700 14280 34728
rect 12176 34632 12756 34660
rect 12820 34632 13308 34660
rect 7285 34595 7343 34601
rect 7285 34592 7297 34595
rect 6972 34564 7297 34592
rect 6972 34552 6978 34564
rect 7285 34561 7297 34564
rect 7331 34561 7343 34595
rect 7285 34555 7343 34561
rect 7469 34595 7527 34601
rect 7469 34561 7481 34595
rect 7515 34592 7527 34595
rect 9125 34595 9183 34601
rect 7515 34564 7604 34592
rect 7515 34561 7527 34564
rect 7469 34555 7527 34561
rect 7576 34536 7604 34564
rect 9125 34561 9137 34595
rect 9171 34592 9183 34595
rect 9585 34595 9643 34601
rect 9171 34564 9536 34592
rect 9171 34561 9183 34564
rect 9125 34555 9183 34561
rect 7558 34484 7564 34536
rect 7616 34484 7622 34536
rect 9309 34527 9367 34533
rect 9309 34493 9321 34527
rect 9355 34493 9367 34527
rect 9508 34524 9536 34564
rect 9585 34561 9597 34595
rect 9631 34561 9643 34595
rect 9585 34555 9643 34561
rect 9769 34595 9827 34601
rect 9769 34561 9781 34595
rect 9815 34592 9827 34595
rect 10410 34592 10416 34604
rect 9815 34564 10416 34592
rect 9815 34561 9827 34564
rect 9769 34555 9827 34561
rect 9784 34524 9812 34555
rect 10410 34552 10416 34564
rect 10468 34552 10474 34604
rect 10873 34595 10931 34601
rect 10873 34561 10885 34595
rect 10919 34561 10931 34595
rect 10873 34555 10931 34561
rect 11057 34595 11115 34601
rect 11057 34561 11069 34595
rect 11103 34592 11115 34595
rect 11606 34592 11612 34604
rect 11103 34564 11612 34592
rect 11103 34561 11115 34564
rect 11057 34555 11115 34561
rect 9508 34496 9812 34524
rect 10888 34524 10916 34555
rect 11606 34552 11612 34564
rect 11664 34552 11670 34604
rect 11882 34552 11888 34604
rect 11940 34592 11946 34604
rect 12176 34601 12204 34632
rect 12161 34595 12219 34601
rect 12161 34592 12173 34595
rect 11940 34564 12173 34592
rect 11940 34552 11946 34564
rect 12161 34561 12173 34564
rect 12207 34561 12219 34595
rect 12161 34555 12219 34561
rect 12342 34552 12348 34604
rect 12400 34552 12406 34604
rect 12437 34595 12495 34601
rect 12437 34561 12449 34595
rect 12483 34592 12495 34595
rect 12618 34592 12624 34604
rect 12483 34564 12624 34592
rect 12483 34561 12495 34564
rect 12437 34555 12495 34561
rect 12618 34552 12624 34564
rect 12676 34552 12682 34604
rect 12728 34601 12756 34632
rect 12713 34595 12771 34601
rect 12713 34561 12725 34595
rect 12759 34561 12771 34595
rect 12713 34555 12771 34561
rect 12802 34552 12808 34604
rect 12860 34592 12866 34604
rect 13280 34601 13308 34632
rect 13081 34595 13139 34601
rect 13081 34592 13093 34595
rect 12860 34564 13093 34592
rect 12860 34552 12866 34564
rect 13081 34561 13093 34564
rect 13127 34561 13139 34595
rect 13081 34555 13139 34561
rect 13265 34595 13323 34601
rect 13265 34561 13277 34595
rect 13311 34561 13323 34595
rect 13265 34555 13323 34561
rect 13538 34552 13544 34604
rect 13596 34552 13602 34604
rect 14200 34601 14228 34700
rect 14274 34688 14280 34700
rect 14332 34688 14338 34740
rect 17678 34728 17684 34740
rect 17328 34700 17684 34728
rect 14458 34620 14464 34672
rect 14516 34620 14522 34672
rect 14553 34663 14611 34669
rect 14553 34629 14565 34663
rect 14599 34660 14611 34663
rect 15102 34660 15108 34672
rect 14599 34632 15108 34660
rect 14599 34629 14611 34632
rect 14553 34623 14611 34629
rect 15102 34620 15108 34632
rect 15160 34620 15166 34672
rect 17328 34669 17356 34700
rect 17678 34688 17684 34700
rect 17736 34688 17742 34740
rect 19705 34731 19763 34737
rect 19705 34697 19717 34731
rect 19751 34728 19763 34731
rect 19978 34728 19984 34740
rect 19751 34700 19984 34728
rect 19751 34697 19763 34700
rect 19705 34691 19763 34697
rect 19978 34688 19984 34700
rect 20036 34688 20042 34740
rect 20070 34688 20076 34740
rect 20128 34688 20134 34740
rect 20622 34688 20628 34740
rect 20680 34688 20686 34740
rect 22557 34731 22615 34737
rect 22557 34697 22569 34731
rect 22603 34728 22615 34731
rect 22922 34728 22928 34740
rect 22603 34700 22928 34728
rect 22603 34697 22615 34700
rect 22557 34691 22615 34697
rect 22922 34688 22928 34700
rect 22980 34688 22986 34740
rect 23106 34688 23112 34740
rect 23164 34728 23170 34740
rect 23385 34731 23443 34737
rect 23385 34728 23397 34731
rect 23164 34700 23397 34728
rect 23164 34688 23170 34700
rect 23385 34697 23397 34700
rect 23431 34697 23443 34731
rect 23385 34691 23443 34697
rect 23474 34688 23480 34740
rect 23532 34688 23538 34740
rect 24762 34728 24768 34740
rect 23584 34700 24768 34728
rect 17313 34663 17371 34669
rect 17313 34629 17325 34663
rect 17359 34629 17371 34663
rect 20088 34660 20116 34688
rect 17313 34623 17371 34629
rect 18892 34632 20116 34660
rect 14185 34595 14243 34601
rect 14185 34561 14197 34595
rect 14231 34561 14243 34595
rect 14185 34555 14243 34561
rect 14278 34595 14336 34601
rect 14278 34561 14290 34595
rect 14324 34592 14336 34595
rect 14324 34564 14504 34592
rect 14324 34561 14336 34564
rect 14278 34555 14336 34561
rect 11698 34524 11704 34536
rect 10888 34496 11704 34524
rect 9309 34487 9367 34493
rect 4982 34416 4988 34468
rect 5040 34456 5046 34468
rect 6178 34456 6184 34468
rect 5040 34428 6184 34456
rect 5040 34416 5046 34428
rect 6178 34416 6184 34428
rect 6236 34456 6242 34468
rect 7650 34456 7656 34468
rect 6236 34428 7656 34456
rect 6236 34416 6242 34428
rect 7650 34416 7656 34428
rect 7708 34416 7714 34468
rect 8938 34416 8944 34468
rect 8996 34456 9002 34468
rect 9324 34456 9352 34487
rect 11698 34484 11704 34496
rect 11756 34484 11762 34536
rect 12897 34527 12955 34533
rect 12897 34524 12909 34527
rect 11808 34496 12909 34524
rect 11330 34456 11336 34468
rect 8996 34428 11336 34456
rect 8996 34416 9002 34428
rect 11330 34416 11336 34428
rect 11388 34416 11394 34468
rect 11808 34456 11836 34496
rect 12897 34493 12909 34496
rect 12943 34493 12955 34527
rect 12897 34487 12955 34493
rect 12989 34527 13047 34533
rect 12989 34493 13001 34527
rect 13035 34524 13047 34527
rect 13556 34524 13584 34552
rect 13035 34496 13584 34524
rect 13035 34493 13047 34496
rect 12989 34487 13047 34493
rect 14090 34484 14096 34536
rect 14148 34484 14154 34536
rect 11630 34428 11836 34456
rect 12529 34459 12587 34465
rect 6914 34348 6920 34400
rect 6972 34388 6978 34400
rect 7193 34391 7251 34397
rect 7193 34388 7205 34391
rect 6972 34360 7205 34388
rect 6972 34348 6978 34360
rect 7193 34357 7205 34360
rect 7239 34357 7251 34391
rect 7193 34351 7251 34357
rect 7374 34348 7380 34400
rect 7432 34348 7438 34400
rect 11146 34348 11152 34400
rect 11204 34388 11210 34400
rect 11630 34388 11658 34428
rect 12529 34425 12541 34459
rect 12575 34456 12587 34459
rect 14108 34456 14136 34484
rect 12575 34428 14136 34456
rect 12575 34425 12587 34428
rect 12529 34419 12587 34425
rect 11204 34360 11658 34388
rect 11723 34391 11781 34397
rect 11204 34348 11210 34360
rect 11723 34357 11735 34391
rect 11769 34388 11781 34391
rect 12342 34388 12348 34400
rect 11769 34360 12348 34388
rect 11769 34357 11781 34360
rect 11723 34351 11781 34357
rect 12342 34348 12348 34360
rect 12400 34348 12406 34400
rect 14476 34388 14504 34564
rect 14642 34552 14648 34604
rect 14700 34601 14706 34604
rect 14700 34592 14708 34601
rect 17129 34595 17187 34601
rect 14700 34564 14745 34592
rect 14700 34555 14708 34564
rect 17129 34561 17141 34595
rect 17175 34561 17187 34595
rect 17129 34555 17187 34561
rect 14700 34552 14706 34555
rect 14550 34484 14556 34536
rect 14608 34524 14614 34536
rect 14608 34496 14780 34524
rect 14608 34484 14614 34496
rect 14752 34456 14780 34496
rect 14829 34459 14887 34465
rect 14829 34456 14841 34459
rect 14752 34428 14841 34456
rect 14829 34425 14841 34428
rect 14875 34425 14887 34459
rect 17144 34456 17172 34555
rect 17218 34552 17224 34604
rect 17276 34552 17282 34604
rect 17431 34595 17489 34601
rect 17431 34561 17443 34595
rect 17477 34561 17489 34595
rect 17431 34555 17489 34561
rect 17681 34595 17739 34601
rect 17681 34561 17693 34595
rect 17727 34561 17739 34595
rect 17681 34555 17739 34561
rect 17144 34428 17205 34456
rect 14829 34419 14887 34425
rect 16114 34388 16120 34400
rect 14476 34360 16120 34388
rect 16114 34348 16120 34360
rect 16172 34348 16178 34400
rect 16758 34348 16764 34400
rect 16816 34388 16822 34400
rect 16945 34391 17003 34397
rect 16945 34388 16957 34391
rect 16816 34360 16957 34388
rect 16816 34348 16822 34360
rect 16945 34357 16957 34360
rect 16991 34357 17003 34391
rect 17177 34388 17205 34428
rect 17310 34416 17316 34468
rect 17368 34456 17374 34468
rect 17446 34456 17474 34555
rect 17586 34484 17592 34536
rect 17644 34484 17650 34536
rect 17696 34524 17724 34555
rect 17862 34552 17868 34604
rect 17920 34592 17926 34604
rect 18892 34592 18920 34632
rect 20438 34620 20444 34672
rect 20496 34620 20502 34672
rect 23492 34660 23520 34688
rect 21560 34632 23152 34660
rect 21560 34604 21588 34632
rect 17920 34564 18920 34592
rect 19153 34595 19211 34601
rect 17920 34552 17926 34564
rect 19153 34561 19165 34595
rect 19199 34592 19211 34595
rect 19886 34592 19892 34604
rect 19199 34564 19892 34592
rect 19199 34561 19211 34564
rect 19153 34555 19211 34561
rect 19886 34552 19892 34564
rect 19944 34552 19950 34604
rect 20165 34595 20223 34601
rect 20165 34561 20177 34595
rect 20211 34561 20223 34595
rect 20165 34555 20223 34561
rect 20257 34595 20315 34601
rect 20257 34561 20269 34595
rect 20303 34561 20315 34595
rect 20257 34555 20315 34561
rect 17770 34524 17776 34536
rect 17696 34496 17776 34524
rect 17770 34484 17776 34496
rect 17828 34524 17834 34536
rect 19613 34527 19671 34533
rect 19613 34524 19625 34527
rect 17828 34496 19625 34524
rect 17828 34484 17834 34496
rect 19613 34493 19625 34496
rect 19659 34493 19671 34527
rect 19613 34487 19671 34493
rect 17368 34428 17474 34456
rect 17604 34456 17632 34484
rect 17604 34428 19012 34456
rect 17368 34416 17374 34428
rect 18984 34400 19012 34428
rect 19058 34416 19064 34468
rect 19116 34456 19122 34468
rect 19426 34456 19432 34468
rect 19116 34428 19432 34456
rect 19116 34416 19122 34428
rect 19426 34416 19432 34428
rect 19484 34416 19490 34468
rect 19521 34459 19579 34465
rect 19521 34425 19533 34459
rect 19567 34456 19579 34459
rect 20180 34456 20208 34555
rect 20272 34468 20300 34555
rect 21542 34552 21548 34604
rect 21600 34552 21606 34604
rect 22830 34552 22836 34604
rect 22888 34552 22894 34604
rect 23124 34601 23152 34632
rect 23308 34632 23520 34660
rect 23308 34601 23336 34632
rect 23584 34601 23612 34700
rect 24762 34688 24768 34700
rect 24820 34688 24826 34740
rect 26142 34728 26148 34740
rect 24872 34700 26148 34728
rect 23934 34660 23940 34672
rect 23860 34632 23940 34660
rect 23860 34601 23888 34632
rect 23934 34620 23940 34632
rect 23992 34660 23998 34672
rect 24872 34660 24900 34700
rect 26142 34688 26148 34700
rect 26200 34688 26206 34740
rect 26418 34688 26424 34740
rect 26476 34688 26482 34740
rect 26786 34688 26792 34740
rect 26844 34688 26850 34740
rect 27614 34688 27620 34740
rect 27672 34688 27678 34740
rect 29086 34728 29092 34740
rect 29012 34700 29092 34728
rect 23992 34632 24900 34660
rect 24949 34663 25007 34669
rect 23992 34620 23998 34632
rect 24949 34629 24961 34663
rect 24995 34660 25007 34663
rect 26436 34660 26464 34688
rect 28258 34660 28264 34672
rect 24995 34632 26464 34660
rect 27264 34632 28264 34660
rect 24995 34629 25007 34632
rect 24949 34623 25007 34629
rect 23109 34595 23167 34601
rect 23109 34561 23121 34595
rect 23155 34561 23167 34595
rect 23109 34555 23167 34561
rect 23293 34595 23351 34601
rect 23293 34561 23305 34595
rect 23339 34561 23351 34595
rect 23293 34555 23351 34561
rect 23569 34595 23627 34601
rect 23569 34561 23581 34595
rect 23615 34561 23627 34595
rect 23569 34555 23627 34561
rect 23845 34595 23903 34601
rect 23845 34561 23857 34595
rect 23891 34561 23903 34595
rect 23845 34555 23903 34561
rect 24765 34595 24823 34601
rect 24765 34561 24777 34595
rect 24811 34592 24823 34595
rect 25498 34592 25504 34604
rect 24811 34564 25504 34592
rect 24811 34561 24823 34564
rect 24765 34555 24823 34561
rect 23017 34527 23075 34533
rect 23017 34524 23029 34527
rect 22664 34496 23029 34524
rect 19567 34428 20208 34456
rect 19567 34425 19579 34428
rect 19521 34419 19579 34425
rect 18049 34391 18107 34397
rect 18049 34388 18061 34391
rect 17177 34360 18061 34388
rect 16945 34351 17003 34357
rect 18049 34357 18061 34360
rect 18095 34357 18107 34391
rect 18049 34351 18107 34357
rect 18966 34348 18972 34400
rect 19024 34388 19030 34400
rect 19978 34388 19984 34400
rect 19024 34360 19984 34388
rect 19024 34348 19030 34360
rect 19978 34348 19984 34360
rect 20036 34348 20042 34400
rect 20180 34388 20208 34428
rect 20254 34416 20260 34468
rect 20312 34416 20318 34468
rect 22664 34400 22692 34496
rect 23017 34493 23029 34496
rect 23063 34493 23075 34527
rect 23124 34524 23152 34555
rect 23584 34524 23612 34555
rect 25498 34552 25504 34564
rect 25556 34552 25562 34604
rect 26237 34595 26295 34601
rect 26237 34561 26249 34595
rect 26283 34561 26295 34595
rect 26237 34555 26295 34561
rect 23124 34496 23612 34524
rect 23753 34527 23811 34533
rect 23017 34487 23075 34493
rect 23753 34493 23765 34527
rect 23799 34524 23811 34527
rect 24302 34524 24308 34536
rect 23799 34496 24308 34524
rect 23799 34493 23811 34496
rect 23753 34487 23811 34493
rect 24302 34484 24308 34496
rect 24360 34524 24366 34536
rect 25133 34527 25191 34533
rect 25133 34524 25145 34527
rect 24360 34496 25145 34524
rect 24360 34484 24366 34496
rect 25133 34493 25145 34496
rect 25179 34493 25191 34527
rect 26252 34524 26280 34555
rect 26418 34552 26424 34604
rect 26476 34552 26482 34604
rect 26510 34552 26516 34604
rect 26568 34552 26574 34604
rect 26605 34595 26663 34601
rect 26605 34561 26617 34595
rect 26651 34592 26663 34595
rect 26694 34592 26700 34604
rect 26651 34564 26700 34592
rect 26651 34561 26663 34564
rect 26605 34555 26663 34561
rect 26694 34552 26700 34564
rect 26752 34552 26758 34604
rect 26878 34552 26884 34604
rect 26936 34592 26942 34604
rect 27264 34601 27292 34632
rect 28258 34620 28264 34632
rect 28316 34620 28322 34672
rect 28902 34620 28908 34672
rect 28960 34660 28966 34672
rect 29012 34660 29040 34700
rect 29086 34688 29092 34700
rect 29144 34688 29150 34740
rect 29546 34688 29552 34740
rect 29604 34688 29610 34740
rect 29851 34731 29909 34737
rect 29851 34697 29863 34731
rect 29897 34728 29909 34731
rect 30098 34728 30104 34740
rect 29897 34700 30104 34728
rect 29897 34697 29909 34700
rect 29851 34691 29909 34697
rect 30098 34688 30104 34700
rect 30156 34688 30162 34740
rect 30466 34688 30472 34740
rect 30524 34728 30530 34740
rect 31113 34731 31171 34737
rect 31113 34728 31125 34731
rect 30524 34700 31125 34728
rect 30524 34688 30530 34700
rect 31113 34697 31125 34700
rect 31159 34697 31171 34731
rect 31113 34691 31171 34697
rect 32766 34688 32772 34740
rect 32824 34688 32830 34740
rect 33962 34688 33968 34740
rect 34020 34728 34026 34740
rect 35342 34728 35348 34740
rect 34020 34700 35348 34728
rect 34020 34688 34026 34700
rect 35342 34688 35348 34700
rect 35400 34688 35406 34740
rect 28960 34632 29040 34660
rect 28960 34620 28966 34632
rect 29270 34620 29276 34672
rect 29328 34620 29334 34672
rect 29564 34660 29592 34688
rect 29641 34663 29699 34669
rect 29641 34660 29653 34663
rect 29564 34632 29653 34660
rect 29641 34629 29653 34632
rect 29687 34629 29699 34663
rect 29641 34623 29699 34629
rect 26973 34595 27031 34601
rect 26973 34592 26985 34595
rect 26936 34564 26985 34592
rect 26936 34552 26942 34564
rect 26973 34561 26985 34564
rect 27019 34561 27031 34595
rect 26973 34555 27031 34561
rect 27121 34595 27179 34601
rect 27121 34561 27133 34595
rect 27167 34561 27179 34595
rect 27121 34555 27179 34561
rect 27249 34595 27307 34601
rect 27249 34561 27261 34595
rect 27295 34561 27307 34595
rect 27249 34555 27307 34561
rect 27136 34524 27164 34555
rect 27338 34552 27344 34604
rect 27396 34592 27402 34604
rect 27479 34595 27537 34601
rect 27396 34564 27438 34592
rect 27396 34552 27402 34564
rect 27479 34561 27491 34595
rect 27525 34592 27537 34595
rect 28810 34592 28816 34604
rect 27525 34564 28816 34592
rect 27525 34561 27537 34564
rect 27479 34555 27537 34561
rect 28810 34552 28816 34564
rect 28868 34552 28874 34604
rect 29089 34595 29147 34601
rect 29089 34561 29101 34595
rect 29135 34592 29147 34595
rect 29288 34592 29316 34620
rect 29135 34564 29316 34592
rect 29365 34595 29423 34601
rect 29135 34561 29147 34564
rect 29089 34555 29147 34561
rect 29365 34561 29377 34595
rect 29411 34582 29423 34595
rect 29454 34582 29460 34604
rect 29411 34561 29460 34582
rect 29365 34555 29460 34561
rect 29380 34554 29460 34555
rect 29454 34552 29460 34554
rect 29512 34552 29518 34604
rect 29546 34552 29552 34604
rect 29604 34552 29610 34604
rect 28902 34524 28908 34536
rect 26252 34496 26740 34524
rect 27136 34496 27200 34524
rect 25133 34487 25191 34493
rect 23661 34459 23719 34465
rect 23661 34425 23673 34459
rect 23707 34456 23719 34459
rect 24578 34456 24584 34468
rect 23707 34428 24584 34456
rect 23707 34425 23719 34428
rect 23661 34419 23719 34425
rect 24578 34416 24584 34428
rect 24636 34416 24642 34468
rect 20530 34388 20536 34400
rect 20180 34360 20536 34388
rect 20530 34348 20536 34360
rect 20588 34348 20594 34400
rect 22646 34348 22652 34400
rect 22704 34348 22710 34400
rect 22925 34391 22983 34397
rect 22925 34357 22937 34391
rect 22971 34388 22983 34391
rect 23842 34388 23848 34400
rect 22971 34360 23848 34388
rect 22971 34357 22983 34360
rect 22925 34351 22983 34357
rect 23842 34348 23848 34360
rect 23900 34348 23906 34400
rect 24394 34348 24400 34400
rect 24452 34388 24458 34400
rect 26602 34388 26608 34400
rect 24452 34360 26608 34388
rect 24452 34348 24458 34360
rect 26602 34348 26608 34360
rect 26660 34348 26666 34400
rect 26712 34388 26740 34496
rect 27172 34456 27200 34496
rect 28460 34496 28908 34524
rect 28460 34456 28488 34496
rect 28902 34484 28908 34496
rect 28960 34484 28966 34536
rect 29656 34524 29684 34623
rect 29730 34620 29736 34672
rect 29788 34620 29794 34672
rect 30006 34620 30012 34672
rect 30064 34660 30070 34672
rect 30190 34660 30196 34672
rect 30064 34632 30196 34660
rect 30064 34620 30070 34632
rect 30190 34620 30196 34632
rect 30248 34660 30254 34672
rect 31570 34660 31576 34672
rect 30248 34632 31576 34660
rect 30248 34620 30254 34632
rect 31570 34620 31576 34632
rect 31628 34620 31634 34672
rect 32306 34620 32312 34672
rect 32364 34620 32370 34672
rect 32784 34660 32812 34688
rect 32861 34663 32919 34669
rect 32861 34660 32873 34663
rect 32784 34632 32873 34660
rect 32861 34629 32873 34632
rect 32907 34629 32919 34663
rect 32861 34623 32919 34629
rect 32968 34632 34192 34660
rect 29748 34592 29776 34620
rect 31021 34595 31079 34601
rect 31021 34592 31033 34595
rect 29748 34564 31033 34592
rect 31021 34561 31033 34564
rect 31067 34592 31079 34595
rect 31294 34592 31300 34604
rect 31067 34564 31300 34592
rect 31067 34561 31079 34564
rect 31021 34555 31079 34561
rect 31294 34552 31300 34564
rect 31352 34552 31358 34604
rect 32674 34552 32680 34604
rect 32732 34552 32738 34604
rect 32769 34595 32827 34601
rect 32769 34561 32781 34595
rect 32815 34592 32827 34595
rect 32968 34592 32996 34632
rect 34164 34604 34192 34632
rect 34256 34632 37780 34660
rect 32815 34564 32996 34592
rect 33137 34595 33195 34601
rect 32815 34561 32827 34564
rect 32769 34555 32827 34561
rect 33137 34561 33149 34595
rect 33183 34592 33195 34595
rect 33686 34592 33692 34604
rect 33183 34564 33692 34592
rect 33183 34561 33195 34564
rect 33137 34555 33195 34561
rect 29288 34496 29684 34524
rect 27172 34428 28488 34456
rect 28534 34416 28540 34468
rect 28592 34456 28598 34468
rect 29288 34465 29316 34496
rect 32214 34484 32220 34536
rect 32272 34484 32278 34536
rect 29181 34459 29239 34465
rect 29181 34456 29193 34459
rect 28592 34428 29193 34456
rect 28592 34416 28598 34428
rect 29181 34425 29193 34428
rect 29227 34425 29239 34459
rect 29181 34419 29239 34425
rect 29273 34459 29331 34465
rect 29273 34425 29285 34459
rect 29319 34425 29331 34459
rect 29273 34419 29331 34425
rect 27154 34388 27160 34400
rect 26712 34360 27160 34388
rect 27154 34348 27160 34360
rect 27212 34348 27218 34400
rect 28718 34348 28724 34400
rect 28776 34388 28782 34400
rect 28905 34391 28963 34397
rect 28905 34388 28917 34391
rect 28776 34360 28917 34388
rect 28776 34348 28782 34360
rect 28905 34357 28917 34360
rect 28951 34357 28963 34391
rect 29196 34388 29224 34419
rect 29362 34416 29368 34468
rect 29420 34416 29426 34468
rect 29730 34416 29736 34468
rect 29788 34456 29794 34468
rect 30009 34459 30067 34465
rect 30009 34456 30021 34459
rect 29788 34428 30021 34456
rect 29788 34416 29794 34428
rect 30009 34425 30021 34428
rect 30055 34425 30067 34459
rect 30009 34419 30067 34425
rect 30558 34416 30564 34468
rect 30616 34456 30622 34468
rect 32784 34456 32812 34555
rect 33686 34552 33692 34564
rect 33744 34552 33750 34604
rect 34146 34552 34152 34604
rect 34204 34552 34210 34604
rect 33410 34484 33416 34536
rect 33468 34524 33474 34536
rect 34256 34524 34284 34632
rect 35253 34595 35311 34601
rect 35253 34561 35265 34595
rect 35299 34561 35311 34595
rect 35253 34555 35311 34561
rect 35437 34595 35495 34601
rect 35437 34561 35449 34595
rect 35483 34592 35495 34595
rect 35710 34592 35716 34604
rect 35483 34564 35716 34592
rect 35483 34561 35495 34564
rect 35437 34555 35495 34561
rect 33468 34496 34284 34524
rect 35268 34524 35296 34555
rect 35710 34552 35716 34564
rect 35768 34552 35774 34604
rect 36265 34595 36323 34601
rect 36265 34561 36277 34595
rect 36311 34592 36323 34595
rect 36354 34592 36360 34604
rect 36311 34564 36360 34592
rect 36311 34561 36323 34564
rect 36265 34555 36323 34561
rect 36354 34552 36360 34564
rect 36412 34552 36418 34604
rect 37752 34536 37780 34632
rect 35268 34496 35388 34524
rect 33468 34484 33474 34496
rect 30616 34428 32812 34456
rect 30616 34416 30622 34428
rect 34790 34416 34796 34468
rect 34848 34456 34854 34468
rect 35069 34459 35127 34465
rect 35069 34456 35081 34459
rect 34848 34428 35081 34456
rect 34848 34416 34854 34428
rect 35069 34425 35081 34428
rect 35115 34425 35127 34459
rect 35360 34456 35388 34496
rect 35526 34484 35532 34536
rect 35584 34524 35590 34536
rect 35621 34527 35679 34533
rect 35621 34524 35633 34527
rect 35584 34496 35633 34524
rect 35584 34484 35590 34496
rect 35621 34493 35633 34496
rect 35667 34493 35679 34527
rect 35621 34487 35679 34493
rect 36446 34484 36452 34536
rect 36504 34484 36510 34536
rect 37734 34484 37740 34536
rect 37792 34484 37798 34536
rect 35434 34456 35440 34468
rect 35360 34428 35440 34456
rect 35069 34419 35127 34425
rect 35434 34416 35440 34428
rect 35492 34456 35498 34468
rect 36354 34456 36360 34468
rect 35492 34428 36360 34456
rect 35492 34416 35498 34428
rect 36354 34416 36360 34428
rect 36412 34416 36418 34468
rect 29380 34388 29408 34416
rect 29196 34360 29408 34388
rect 29825 34391 29883 34397
rect 28905 34351 28963 34357
rect 29825 34357 29837 34391
rect 29871 34388 29883 34391
rect 30282 34388 30288 34400
rect 29871 34360 30288 34388
rect 29871 34357 29883 34360
rect 29825 34351 29883 34357
rect 30282 34348 30288 34360
rect 30340 34348 30346 34400
rect 33870 34348 33876 34400
rect 33928 34388 33934 34400
rect 37458 34388 37464 34400
rect 33928 34360 37464 34388
rect 33928 34348 33934 34360
rect 37458 34348 37464 34360
rect 37516 34348 37522 34400
rect 1104 34298 41400 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 41400 34298
rect 1104 34224 41400 34246
rect 5074 34144 5080 34196
rect 5132 34184 5138 34196
rect 5169 34187 5227 34193
rect 5169 34184 5181 34187
rect 5132 34156 5181 34184
rect 5132 34144 5138 34156
rect 5169 34153 5181 34156
rect 5215 34153 5227 34187
rect 5169 34147 5227 34153
rect 8294 34144 8300 34196
rect 8352 34144 8358 34196
rect 9766 34144 9772 34196
rect 9824 34144 9830 34196
rect 11609 34187 11667 34193
rect 11609 34153 11621 34187
rect 11655 34184 11667 34187
rect 11698 34184 11704 34196
rect 11655 34156 11704 34184
rect 11655 34153 11667 34156
rect 11609 34147 11667 34153
rect 11698 34144 11704 34156
rect 11756 34144 11762 34196
rect 11808 34156 12112 34184
rect 4801 34119 4859 34125
rect 4801 34085 4813 34119
rect 4847 34116 4859 34119
rect 5258 34116 5264 34128
rect 4847 34088 5264 34116
rect 4847 34085 4859 34088
rect 4801 34079 4859 34085
rect 5258 34076 5264 34088
rect 5316 34076 5322 34128
rect 5810 34116 5816 34128
rect 5460 34088 5816 34116
rect 4062 34008 4068 34060
rect 4120 34008 4126 34060
rect 5353 34051 5411 34057
rect 5353 34017 5365 34051
rect 5399 34048 5411 34051
rect 5460 34048 5488 34088
rect 5810 34076 5816 34088
rect 5868 34076 5874 34128
rect 6914 34076 6920 34128
rect 6972 34116 6978 34128
rect 6972 34088 7696 34116
rect 6972 34076 6978 34088
rect 7285 34051 7343 34057
rect 7285 34048 7297 34051
rect 5399 34020 5488 34048
rect 5644 34020 7297 34048
rect 5399 34017 5411 34020
rect 5353 34011 5411 34017
rect 3973 33983 4031 33989
rect 3973 33949 3985 33983
rect 4019 33980 4031 33983
rect 4430 33980 4436 33992
rect 4019 33952 4436 33980
rect 4019 33949 4031 33952
rect 3973 33943 4031 33949
rect 4430 33940 4436 33952
rect 4488 33940 4494 33992
rect 4525 33983 4583 33989
rect 4525 33949 4537 33983
rect 4571 33949 4583 33983
rect 4525 33943 4583 33949
rect 4540 33856 4568 33943
rect 4706 33940 4712 33992
rect 4764 33940 4770 33992
rect 4801 33983 4859 33989
rect 4801 33949 4813 33983
rect 4847 33980 4859 33983
rect 4982 33980 4988 33992
rect 4847 33952 4988 33980
rect 4847 33949 4859 33952
rect 4801 33943 4859 33949
rect 4982 33940 4988 33952
rect 5040 33940 5046 33992
rect 5077 33983 5135 33989
rect 5077 33949 5089 33983
rect 5123 33980 5135 33983
rect 5445 33983 5503 33989
rect 5123 33952 5304 33980
rect 5123 33949 5135 33952
rect 5077 33943 5135 33949
rect 4724 33912 4752 33940
rect 5276 33924 5304 33952
rect 5445 33949 5457 33983
rect 5491 33980 5503 33983
rect 5644 33980 5672 34020
rect 7285 34017 7297 34020
rect 7331 34017 7343 34051
rect 7285 34011 7343 34017
rect 7374 34008 7380 34060
rect 7432 34048 7438 34060
rect 7668 34057 7696 34088
rect 9674 34076 9680 34128
rect 9732 34116 9738 34128
rect 11808 34116 11836 34156
rect 9732 34088 9996 34116
rect 9732 34076 9738 34088
rect 7561 34051 7619 34057
rect 7561 34048 7573 34051
rect 7432 34020 7573 34048
rect 7432 34008 7438 34020
rect 7561 34017 7573 34020
rect 7607 34017 7619 34051
rect 7561 34011 7619 34017
rect 7653 34051 7711 34057
rect 7653 34017 7665 34051
rect 7699 34017 7711 34051
rect 7653 34011 7711 34017
rect 8036 34020 9812 34048
rect 5491 33952 5672 33980
rect 5491 33949 5503 33952
rect 5445 33943 5503 33949
rect 5718 33940 5724 33992
rect 5776 33940 5782 33992
rect 5813 33983 5871 33989
rect 5813 33949 5825 33983
rect 5859 33980 5871 33983
rect 6273 33983 6331 33989
rect 6273 33980 6285 33983
rect 5859 33952 6285 33980
rect 5859 33949 5871 33952
rect 5813 33943 5871 33949
rect 6273 33949 6285 33952
rect 6319 33949 6331 33983
rect 6273 33943 6331 33949
rect 6822 33940 6828 33992
rect 6880 33980 6886 33992
rect 6917 33983 6975 33989
rect 6917 33980 6929 33983
rect 6880 33952 6929 33980
rect 6880 33940 6886 33952
rect 6917 33949 6929 33952
rect 6963 33949 6975 33983
rect 6917 33943 6975 33949
rect 7006 33940 7012 33992
rect 7064 33980 7070 33992
rect 7469 33983 7527 33989
rect 7469 33980 7481 33983
rect 7064 33952 7481 33980
rect 7064 33940 7070 33952
rect 7469 33949 7481 33952
rect 7515 33949 7527 33983
rect 7469 33943 7527 33949
rect 4890 33912 4896 33924
rect 4724 33884 4896 33912
rect 4890 33872 4896 33884
rect 4948 33872 4954 33924
rect 5258 33872 5264 33924
rect 5316 33872 5322 33924
rect 5902 33872 5908 33924
rect 5960 33872 5966 33924
rect 6089 33915 6147 33921
rect 6089 33881 6101 33915
rect 6135 33881 6147 33915
rect 6089 33875 6147 33881
rect 6549 33915 6607 33921
rect 6549 33881 6561 33915
rect 6595 33912 6607 33915
rect 7576 33912 7604 34011
rect 8036 33989 8064 34020
rect 7745 33983 7803 33989
rect 7745 33949 7757 33983
rect 7791 33980 7803 33983
rect 8021 33983 8079 33989
rect 8021 33980 8033 33983
rect 7791 33952 8033 33980
rect 7791 33949 7803 33952
rect 7745 33943 7803 33949
rect 8021 33949 8033 33952
rect 8067 33949 8079 33983
rect 8021 33943 8079 33949
rect 9674 33940 9680 33992
rect 9732 33940 9738 33992
rect 6595 33884 7604 33912
rect 6595 33881 6607 33884
rect 6549 33875 6607 33881
rect 4341 33847 4399 33853
rect 4341 33813 4353 33847
rect 4387 33844 4399 33847
rect 4522 33844 4528 33856
rect 4387 33816 4528 33844
rect 4387 33813 4399 33816
rect 4341 33807 4399 33813
rect 4522 33804 4528 33816
rect 4580 33804 4586 33856
rect 4617 33847 4675 33853
rect 4617 33813 4629 33847
rect 4663 33844 4675 33847
rect 4985 33847 5043 33853
rect 4985 33844 4997 33847
rect 4663 33816 4997 33844
rect 4663 33813 4675 33816
rect 4617 33807 4675 33813
rect 4985 33813 4997 33816
rect 5031 33844 5043 33847
rect 6104 33844 6132 33875
rect 6932 33856 6960 33884
rect 5031 33816 6132 33844
rect 5031 33813 5043 33816
rect 4985 33807 5043 33813
rect 6914 33804 6920 33856
rect 6972 33804 6978 33856
rect 7190 33804 7196 33856
rect 7248 33804 7254 33856
rect 9784 33844 9812 34020
rect 9861 33985 9919 33991
rect 9861 33951 9873 33985
rect 9907 33980 9919 33985
rect 9968 33980 9996 34088
rect 10981 34088 11836 34116
rect 11977 34119 12035 34125
rect 10686 33980 10692 33992
rect 9907 33952 10692 33980
rect 9907 33951 9919 33952
rect 9861 33945 9919 33951
rect 10686 33940 10692 33952
rect 10744 33980 10750 33992
rect 10981 33980 11009 34088
rect 11977 34085 11989 34119
rect 12023 34085 12035 34119
rect 11977 34079 12035 34085
rect 12084 34116 12112 34156
rect 12710 34144 12716 34196
rect 12768 34184 12774 34196
rect 12897 34187 12955 34193
rect 12897 34184 12909 34187
rect 12768 34156 12909 34184
rect 12768 34144 12774 34156
rect 12897 34153 12909 34156
rect 12943 34153 12955 34187
rect 12897 34147 12955 34153
rect 13725 34187 13783 34193
rect 13725 34153 13737 34187
rect 13771 34184 13783 34187
rect 14458 34184 14464 34196
rect 13771 34156 14464 34184
rect 13771 34153 13783 34156
rect 13725 34147 13783 34153
rect 14458 34144 14464 34156
rect 14516 34144 14522 34196
rect 16206 34144 16212 34196
rect 16264 34184 16270 34196
rect 16264 34156 18276 34184
rect 16264 34144 16270 34156
rect 18248 34128 18276 34156
rect 19886 34144 19892 34196
rect 19944 34144 19950 34196
rect 20438 34144 20444 34196
rect 20496 34144 20502 34196
rect 20530 34144 20536 34196
rect 20588 34184 20594 34196
rect 20809 34187 20867 34193
rect 20809 34184 20821 34187
rect 20588 34156 20821 34184
rect 20588 34144 20594 34156
rect 20809 34153 20821 34156
rect 20855 34153 20867 34187
rect 22554 34184 22560 34196
rect 20809 34147 20867 34153
rect 22444 34156 22560 34184
rect 12084 34088 14320 34116
rect 11146 34008 11152 34060
rect 11204 34048 11210 34060
rect 11204 34020 11836 34048
rect 11204 34008 11210 34020
rect 10744 33952 11009 33980
rect 10744 33940 10750 33952
rect 11054 33940 11060 33992
rect 11112 33980 11118 33992
rect 11808 33989 11836 34020
rect 11425 33983 11483 33989
rect 11425 33980 11437 33983
rect 11112 33952 11437 33980
rect 11112 33940 11118 33952
rect 11425 33949 11437 33952
rect 11471 33949 11483 33983
rect 11425 33943 11483 33949
rect 11793 33983 11851 33989
rect 11793 33949 11805 33983
rect 11839 33949 11851 33983
rect 11793 33943 11851 33949
rect 11882 33940 11888 33992
rect 11940 33940 11946 33992
rect 11992 33980 12020 34079
rect 12084 34057 12112 34088
rect 12069 34051 12127 34057
rect 12069 34017 12081 34051
rect 12115 34017 12127 34051
rect 12069 34011 12127 34017
rect 13449 34051 13507 34057
rect 13449 34017 13461 34051
rect 13495 34048 13507 34051
rect 14093 34051 14151 34057
rect 14093 34048 14105 34051
rect 13495 34020 14105 34048
rect 13495 34017 13507 34020
rect 13449 34011 13507 34017
rect 14093 34017 14105 34020
rect 14139 34017 14151 34051
rect 14093 34011 14151 34017
rect 12802 33980 12808 33992
rect 11992 33952 12808 33980
rect 12802 33940 12808 33952
rect 12860 33940 12866 33992
rect 13081 33983 13139 33989
rect 13081 33949 13093 33983
rect 13127 33949 13139 33983
rect 13081 33943 13139 33949
rect 11241 33915 11299 33921
rect 11241 33881 11253 33915
rect 11287 33912 11299 33915
rect 12618 33912 12624 33924
rect 11287 33884 12624 33912
rect 11287 33881 11299 33884
rect 11241 33875 11299 33881
rect 12618 33872 12624 33884
rect 12676 33872 12682 33924
rect 13096 33912 13124 33943
rect 13170 33940 13176 33992
rect 13228 33980 13234 33992
rect 13265 33983 13323 33989
rect 13265 33980 13277 33983
rect 13228 33952 13277 33980
rect 13228 33940 13234 33952
rect 13265 33949 13277 33952
rect 13311 33949 13323 33983
rect 13265 33943 13323 33949
rect 13357 33983 13415 33989
rect 13357 33949 13369 33983
rect 13403 33980 13415 33983
rect 13538 33980 13544 33992
rect 13403 33952 13544 33980
rect 13403 33949 13415 33952
rect 13357 33943 13415 33949
rect 13538 33940 13544 33952
rect 13596 33940 13602 33992
rect 13725 33983 13783 33989
rect 13725 33949 13737 33983
rect 13771 33949 13783 33983
rect 13725 33943 13783 33949
rect 13446 33912 13452 33924
rect 13096 33884 13452 33912
rect 13446 33872 13452 33884
rect 13504 33912 13510 33924
rect 13740 33912 13768 33943
rect 13906 33940 13912 33992
rect 13964 33940 13970 33992
rect 14292 33989 14320 34088
rect 18230 34076 18236 34128
rect 18288 34076 18294 34128
rect 20456 34116 20484 34144
rect 20180 34088 20484 34116
rect 16298 34008 16304 34060
rect 16356 34048 16362 34060
rect 16945 34051 17003 34057
rect 16945 34048 16957 34051
rect 16356 34020 16957 34048
rect 16356 34008 16362 34020
rect 16945 34017 16957 34020
rect 16991 34048 17003 34051
rect 18690 34048 18696 34060
rect 16991 34020 18696 34048
rect 16991 34017 17003 34020
rect 16945 34011 17003 34017
rect 18690 34008 18696 34020
rect 18748 34048 18754 34060
rect 19058 34048 19064 34060
rect 18748 34020 19064 34048
rect 18748 34008 18754 34020
rect 19058 34008 19064 34020
rect 19116 34008 19122 34060
rect 19797 34051 19855 34057
rect 19797 34017 19809 34051
rect 19843 34048 19855 34051
rect 20180 34048 20208 34088
rect 20349 34051 20407 34057
rect 20349 34048 20361 34051
rect 19843 34020 20361 34048
rect 19843 34017 19855 34020
rect 19797 34011 19855 34017
rect 20349 34017 20361 34020
rect 20395 34017 20407 34051
rect 20349 34011 20407 34017
rect 20530 34008 20536 34060
rect 20588 34048 20594 34060
rect 21177 34051 21235 34057
rect 21177 34048 21189 34051
rect 20588 34020 21189 34048
rect 20588 34008 20594 34020
rect 21177 34017 21189 34020
rect 21223 34017 21235 34051
rect 21177 34011 21235 34017
rect 21450 34008 21456 34060
rect 21508 34008 21514 34060
rect 21545 34051 21603 34057
rect 21545 34017 21557 34051
rect 21591 34048 21603 34051
rect 22094 34048 22100 34060
rect 21591 34020 22100 34048
rect 21591 34017 21603 34020
rect 21545 34011 21603 34017
rect 22094 34008 22100 34020
rect 22152 34008 22158 34060
rect 14277 33983 14335 33989
rect 14277 33949 14289 33983
rect 14323 33949 14335 33983
rect 14277 33943 14335 33949
rect 13504 33884 13768 33912
rect 14292 33912 14320 33943
rect 14458 33940 14464 33992
rect 14516 33940 14522 33992
rect 14550 33940 14556 33992
rect 14608 33940 14614 33992
rect 15746 33940 15752 33992
rect 15804 33940 15810 33992
rect 16577 33983 16635 33989
rect 16577 33949 16589 33983
rect 16623 33980 16635 33983
rect 16758 33980 16764 33992
rect 16623 33952 16764 33980
rect 16623 33949 16635 33952
rect 16577 33943 16635 33949
rect 16758 33940 16764 33952
rect 16816 33940 16822 33992
rect 16850 33940 16856 33992
rect 16908 33940 16914 33992
rect 19337 33983 19395 33989
rect 19337 33980 19349 33983
rect 18524 33952 19349 33980
rect 15194 33912 15200 33924
rect 14292 33884 15200 33912
rect 13504 33872 13510 33884
rect 15194 33872 15200 33884
rect 15252 33912 15258 33924
rect 15764 33912 15792 33940
rect 15252 33884 15792 33912
rect 15252 33872 15258 33884
rect 16114 33872 16120 33924
rect 16172 33912 16178 33924
rect 16393 33915 16451 33921
rect 16172 33884 16344 33912
rect 16172 33872 16178 33884
rect 16206 33844 16212 33856
rect 9784 33816 16212 33844
rect 16206 33804 16212 33816
rect 16264 33804 16270 33856
rect 16316 33844 16344 33884
rect 16393 33881 16405 33915
rect 16439 33912 16451 33915
rect 17221 33915 17279 33921
rect 17221 33912 17233 33915
rect 16439 33884 17233 33912
rect 16439 33881 16451 33884
rect 16393 33875 16451 33881
rect 17221 33881 17233 33884
rect 17267 33881 17279 33915
rect 17221 33875 17279 33881
rect 18230 33872 18236 33924
rect 18288 33872 18294 33924
rect 16761 33847 16819 33853
rect 16761 33844 16773 33847
rect 16316 33816 16773 33844
rect 16761 33813 16773 33816
rect 16807 33844 16819 33847
rect 17034 33844 17040 33856
rect 16807 33816 17040 33844
rect 16807 33813 16819 33816
rect 16761 33807 16819 33813
rect 17034 33804 17040 33816
rect 17092 33804 17098 33856
rect 17126 33804 17132 33856
rect 17184 33844 17190 33856
rect 18524 33844 18552 33952
rect 19337 33949 19349 33952
rect 19383 33980 19395 33983
rect 19610 33980 19616 33992
rect 19383 33952 19616 33980
rect 19383 33949 19395 33952
rect 19337 33943 19395 33949
rect 19610 33940 19616 33952
rect 19668 33940 19674 33992
rect 19978 33940 19984 33992
rect 20036 33980 20042 33992
rect 20073 33983 20131 33989
rect 20073 33980 20085 33983
rect 20036 33952 20085 33980
rect 20036 33940 20042 33952
rect 20073 33949 20085 33952
rect 20119 33949 20131 33983
rect 20073 33943 20131 33949
rect 20254 33940 20260 33992
rect 20312 33980 20318 33992
rect 20441 33983 20499 33989
rect 20441 33980 20453 33983
rect 20312 33952 20453 33980
rect 20312 33940 20318 33952
rect 18966 33872 18972 33924
rect 19024 33872 19030 33924
rect 19058 33872 19064 33924
rect 19116 33912 19122 33924
rect 19116 33884 20116 33912
rect 19116 33872 19122 33884
rect 20088 33856 20116 33884
rect 17184 33816 18552 33844
rect 17184 33804 17190 33816
rect 18598 33804 18604 33856
rect 18656 33844 18662 33856
rect 19337 33847 19395 33853
rect 19337 33844 19349 33847
rect 18656 33816 19349 33844
rect 18656 33804 18662 33816
rect 19337 33813 19349 33816
rect 19383 33813 19395 33847
rect 19337 33807 19395 33813
rect 20070 33804 20076 33856
rect 20128 33804 20134 33856
rect 20364 33844 20392 33952
rect 20441 33949 20453 33952
rect 20487 33949 20499 33983
rect 20441 33943 20499 33949
rect 20625 33983 20683 33989
rect 20625 33949 20637 33983
rect 20671 33949 20683 33983
rect 20625 33943 20683 33949
rect 20530 33872 20536 33924
rect 20588 33912 20594 33924
rect 20640 33912 20668 33943
rect 21358 33940 21364 33992
rect 21416 33940 21422 33992
rect 21637 33983 21695 33989
rect 21637 33980 21649 33983
rect 21468 33952 21649 33980
rect 20588 33884 20668 33912
rect 20588 33872 20594 33884
rect 21468 33844 21496 33952
rect 21637 33949 21649 33952
rect 21683 33949 21695 33983
rect 21637 33943 21695 33949
rect 22278 33940 22284 33992
rect 22336 33940 22342 33992
rect 22444 33989 22472 34156
rect 22554 34144 22560 34156
rect 22612 34144 22618 34196
rect 24029 34187 24087 34193
rect 24029 34153 24041 34187
rect 24075 34184 24087 34187
rect 25038 34184 25044 34196
rect 24075 34156 25044 34184
rect 24075 34153 24087 34156
rect 24029 34147 24087 34153
rect 25038 34144 25044 34156
rect 25096 34144 25102 34196
rect 27614 34184 27620 34196
rect 25700 34156 27620 34184
rect 22830 34116 22836 34128
rect 22572 34088 22836 34116
rect 22572 33989 22600 34088
rect 22830 34076 22836 34088
rect 22888 34076 22894 34128
rect 24854 34116 24860 34128
rect 23860 34088 24860 34116
rect 23860 34048 23888 34088
rect 24854 34076 24860 34088
rect 24912 34116 24918 34128
rect 25590 34116 25596 34128
rect 24912 34088 25596 34116
rect 24912 34076 24918 34088
rect 25590 34076 25596 34088
rect 25648 34076 25654 34128
rect 22664 34020 23888 34048
rect 23937 34051 23995 34057
rect 22664 33992 22692 34020
rect 23937 34017 23949 34051
rect 23983 34048 23995 34051
rect 24397 34051 24455 34057
rect 24397 34048 24409 34051
rect 23983 34020 24409 34048
rect 23983 34017 23995 34020
rect 23937 34011 23995 34017
rect 24397 34017 24409 34020
rect 24443 34017 24455 34051
rect 24397 34011 24455 34017
rect 25222 34008 25228 34060
rect 25280 34048 25286 34060
rect 25700 34048 25728 34156
rect 27614 34144 27620 34156
rect 27672 34144 27678 34196
rect 28534 34144 28540 34196
rect 28592 34144 28598 34196
rect 30837 34187 30895 34193
rect 30837 34184 30849 34187
rect 28644 34156 30849 34184
rect 27430 34116 27436 34128
rect 25280 34020 25728 34048
rect 26804 34088 27436 34116
rect 25280 34008 25286 34020
rect 22429 33983 22487 33989
rect 22429 33949 22441 33983
rect 22475 33949 22487 33983
rect 22429 33943 22487 33949
rect 22557 33983 22615 33989
rect 22557 33949 22569 33983
rect 22603 33949 22615 33983
rect 22557 33943 22615 33949
rect 22646 33940 22652 33992
rect 22704 33940 22710 33992
rect 22787 33983 22845 33989
rect 22787 33949 22799 33983
rect 22833 33980 22845 33983
rect 23566 33980 23572 33992
rect 22833 33952 23572 33980
rect 22833 33949 22845 33952
rect 22787 33943 22845 33949
rect 20364 33816 21496 33844
rect 21634 33804 21640 33856
rect 21692 33844 21698 33856
rect 22802 33844 22830 33943
rect 23566 33940 23572 33952
rect 23624 33940 23630 33992
rect 24029 33983 24087 33989
rect 24029 33949 24041 33983
rect 24075 33949 24087 33983
rect 24029 33943 24087 33949
rect 23198 33872 23204 33924
rect 23256 33912 23262 33924
rect 23753 33915 23811 33921
rect 23753 33912 23765 33915
rect 23256 33884 23765 33912
rect 23256 33872 23262 33884
rect 23753 33881 23765 33884
rect 23799 33881 23811 33915
rect 24044 33912 24072 33943
rect 24118 33940 24124 33992
rect 24176 33980 24182 33992
rect 24581 33983 24639 33989
rect 24581 33980 24593 33983
rect 24176 33952 24593 33980
rect 24176 33940 24182 33952
rect 24581 33949 24593 33952
rect 24627 33949 24639 33983
rect 24581 33943 24639 33949
rect 24673 33983 24731 33989
rect 24673 33949 24685 33983
rect 24719 33980 24731 33983
rect 24719 33952 24808 33980
rect 24719 33949 24731 33952
rect 24673 33943 24731 33949
rect 24780 33912 24808 33952
rect 24854 33940 24860 33992
rect 24912 33980 24918 33992
rect 24949 33983 25007 33989
rect 24949 33980 24961 33983
rect 24912 33952 24961 33980
rect 24912 33940 24918 33952
rect 24949 33949 24961 33952
rect 24995 33980 25007 33983
rect 25682 33980 25688 33992
rect 24995 33952 25688 33980
rect 24995 33949 25007 33952
rect 24949 33943 25007 33949
rect 25682 33940 25688 33952
rect 25740 33940 25746 33992
rect 26804 33989 26832 34088
rect 27430 34076 27436 34088
rect 27488 34076 27494 34128
rect 27709 34119 27767 34125
rect 27709 34085 27721 34119
rect 27755 34085 27767 34119
rect 28552 34116 28580 34144
rect 27709 34079 27767 34085
rect 28460 34088 28580 34116
rect 27724 34048 27752 34079
rect 26988 34020 27752 34048
rect 26988 33989 27016 34020
rect 26697 33983 26755 33989
rect 26697 33949 26709 33983
rect 26743 33949 26755 33983
rect 26697 33943 26755 33949
rect 26789 33983 26847 33989
rect 26789 33949 26801 33983
rect 26835 33949 26847 33983
rect 26789 33943 26847 33949
rect 26973 33983 27031 33989
rect 26973 33949 26985 33983
rect 27019 33949 27031 33983
rect 26973 33943 27031 33949
rect 27065 33983 27123 33989
rect 27065 33949 27077 33983
rect 27111 33949 27123 33983
rect 27065 33943 27123 33949
rect 24044 33884 24716 33912
rect 24780 33884 25728 33912
rect 23753 33875 23811 33881
rect 24688 33856 24716 33884
rect 25700 33856 25728 33884
rect 26712 33856 26740 33943
rect 27080 33912 27108 33943
rect 27154 33940 27160 33992
rect 27212 33940 27218 33992
rect 27341 33983 27399 33989
rect 27341 33949 27353 33983
rect 27387 33949 27399 33983
rect 27341 33943 27399 33949
rect 26804 33884 27108 33912
rect 26804 33856 26832 33884
rect 27356 33856 27384 33943
rect 27522 33940 27528 33992
rect 27580 33940 27586 33992
rect 27430 33872 27436 33924
rect 27488 33912 27494 33924
rect 27893 33915 27951 33921
rect 27893 33912 27905 33915
rect 27488 33884 27905 33912
rect 27488 33872 27494 33884
rect 27893 33881 27905 33884
rect 27939 33881 27951 33915
rect 28460 33912 28488 34088
rect 28644 34048 28672 34156
rect 30837 34153 30849 34156
rect 30883 34153 30895 34187
rect 30837 34147 30895 34153
rect 33778 34144 33784 34196
rect 33836 34184 33842 34196
rect 36909 34187 36967 34193
rect 36909 34184 36921 34187
rect 33836 34156 36921 34184
rect 33836 34144 33842 34156
rect 36909 34153 36921 34156
rect 36955 34153 36967 34187
rect 36909 34147 36967 34153
rect 37458 34144 37464 34196
rect 37516 34144 37522 34196
rect 28718 34076 28724 34128
rect 28776 34076 28782 34128
rect 29270 34076 29276 34128
rect 29328 34116 29334 34128
rect 31481 34119 31539 34125
rect 29328 34088 30236 34116
rect 29328 34076 29334 34088
rect 28552 34020 28672 34048
rect 28736 34048 28764 34076
rect 28736 34020 29592 34048
rect 28552 33992 28580 34020
rect 28534 33940 28540 33992
rect 28592 33940 28598 33992
rect 28630 33983 28688 33989
rect 28630 33949 28642 33983
rect 28676 33949 28688 33983
rect 28630 33943 28688 33949
rect 28644 33912 28672 33943
rect 28810 33940 28816 33992
rect 28868 33940 28874 33992
rect 28994 33940 29000 33992
rect 29052 33989 29058 33992
rect 29564 33989 29592 34020
rect 29657 33992 29685 34088
rect 29052 33980 29060 33989
rect 29549 33983 29607 33989
rect 29052 33952 29097 33980
rect 29052 33943 29060 33952
rect 29549 33949 29561 33983
rect 29595 33949 29607 33983
rect 29549 33943 29607 33949
rect 29052 33940 29058 33943
rect 29638 33940 29644 33992
rect 29696 33940 29702 33992
rect 29917 33983 29975 33989
rect 29917 33980 29929 33983
rect 29748 33952 29929 33980
rect 28460 33884 28672 33912
rect 27893 33875 27951 33881
rect 28902 33872 28908 33924
rect 28960 33872 28966 33924
rect 29454 33872 29460 33924
rect 29512 33912 29518 33924
rect 29748 33912 29776 33952
rect 29917 33949 29929 33952
rect 29963 33949 29975 33983
rect 29917 33943 29975 33949
rect 30006 33940 30012 33992
rect 30064 33989 30070 33992
rect 30064 33980 30072 33989
rect 30208 33980 30236 34088
rect 31481 34085 31493 34119
rect 31527 34116 31539 34119
rect 32214 34116 32220 34128
rect 31527 34088 32220 34116
rect 31527 34085 31539 34088
rect 31481 34079 31539 34085
rect 30282 34008 30288 34060
rect 30340 34008 30346 34060
rect 31680 34057 31708 34088
rect 32214 34076 32220 34088
rect 32272 34116 32278 34128
rect 32950 34116 32956 34128
rect 32272 34088 32956 34116
rect 32272 34076 32278 34088
rect 32950 34076 32956 34088
rect 33008 34116 33014 34128
rect 35434 34116 35440 34128
rect 33008 34088 33364 34116
rect 33008 34076 33014 34088
rect 31665 34051 31723 34057
rect 31665 34017 31677 34051
rect 31711 34017 31723 34051
rect 31665 34011 31723 34017
rect 32033 34051 32091 34057
rect 32033 34017 32045 34051
rect 32079 34048 32091 34051
rect 32582 34048 32588 34060
rect 32079 34020 32588 34048
rect 32079 34017 32091 34020
rect 32033 34011 32091 34017
rect 32582 34008 32588 34020
rect 32640 34008 32646 34060
rect 33042 34008 33048 34060
rect 33100 34048 33106 34060
rect 33137 34051 33195 34057
rect 33137 34048 33149 34051
rect 33100 34020 33149 34048
rect 33100 34008 33106 34020
rect 33137 34017 33149 34020
rect 33183 34017 33195 34051
rect 33336 34048 33364 34088
rect 34072 34088 35440 34116
rect 33336 34020 33456 34048
rect 33137 34011 33195 34017
rect 30469 33983 30527 33989
rect 30469 33980 30481 33983
rect 30064 33952 30109 33980
rect 30208 33952 30481 33980
rect 30064 33943 30072 33952
rect 30469 33949 30481 33952
rect 30515 33949 30527 33983
rect 30469 33943 30527 33949
rect 30064 33940 30070 33943
rect 30558 33940 30564 33992
rect 30616 33940 30622 33992
rect 30650 33940 30656 33992
rect 30708 33940 30714 33992
rect 32766 33980 32772 33992
rect 31956 33952 32772 33980
rect 29512 33884 29776 33912
rect 29825 33915 29883 33921
rect 29512 33872 29518 33884
rect 29825 33881 29837 33915
rect 29871 33912 29883 33915
rect 30668 33912 30696 33940
rect 31956 33921 31984 33952
rect 32766 33940 32772 33952
rect 32824 33980 32830 33992
rect 33428 33989 33456 34020
rect 32861 33983 32919 33989
rect 32861 33980 32873 33983
rect 32824 33952 32873 33980
rect 32824 33940 32830 33952
rect 32861 33949 32873 33952
rect 32907 33949 32919 33983
rect 32861 33943 32919 33949
rect 33413 33983 33471 33989
rect 33413 33949 33425 33983
rect 33459 33949 33471 33983
rect 33413 33943 33471 33949
rect 33594 33940 33600 33992
rect 33652 33980 33658 33992
rect 34072 33989 34100 34088
rect 35434 34076 35440 34088
rect 35492 34076 35498 34128
rect 34790 34048 34796 34060
rect 34348 34020 34796 34048
rect 34348 33989 34376 34020
rect 34790 34008 34796 34020
rect 34848 34048 34854 34060
rect 35345 34051 35403 34057
rect 35345 34048 35357 34051
rect 34848 34020 35357 34048
rect 34848 34008 34854 34020
rect 35345 34017 35357 34020
rect 35391 34048 35403 34051
rect 36170 34048 36176 34060
rect 35391 34020 36176 34048
rect 35391 34017 35403 34020
rect 35345 34011 35403 34017
rect 36170 34008 36176 34020
rect 36228 34048 36234 34060
rect 36265 34051 36323 34057
rect 36265 34048 36277 34051
rect 36228 34020 36277 34048
rect 36228 34008 36234 34020
rect 36265 34017 36277 34020
rect 36311 34017 36323 34051
rect 36265 34011 36323 34017
rect 34057 33983 34115 33989
rect 34057 33980 34069 33983
rect 33652 33952 34069 33980
rect 33652 33940 33658 33952
rect 34057 33949 34069 33952
rect 34103 33949 34115 33983
rect 34057 33943 34115 33949
rect 34333 33983 34391 33989
rect 34333 33949 34345 33983
rect 34379 33949 34391 33983
rect 34333 33943 34391 33949
rect 31113 33915 31171 33921
rect 29871 33884 30512 33912
rect 30668 33884 30972 33912
rect 29871 33881 29883 33884
rect 29825 33875 29883 33881
rect 30484 33856 30512 33884
rect 21692 33816 22830 33844
rect 21692 33804 21698 33816
rect 22922 33804 22928 33856
rect 22980 33804 22986 33856
rect 24210 33804 24216 33856
rect 24268 33804 24274 33856
rect 24670 33804 24676 33856
rect 24728 33804 24734 33856
rect 25682 33804 25688 33856
rect 25740 33804 25746 33856
rect 26510 33804 26516 33856
rect 26568 33804 26574 33856
rect 26694 33804 26700 33856
rect 26752 33804 26758 33856
rect 26786 33804 26792 33856
rect 26844 33804 26850 33856
rect 27338 33804 27344 33856
rect 27396 33804 27402 33856
rect 27706 33804 27712 33856
rect 27764 33844 27770 33856
rect 27985 33847 28043 33853
rect 27985 33844 27997 33847
rect 27764 33816 27997 33844
rect 27764 33804 27770 33816
rect 27985 33813 27997 33816
rect 28031 33813 28043 33847
rect 27985 33807 28043 33813
rect 29178 33804 29184 33856
rect 29236 33804 29242 33856
rect 29362 33804 29368 33856
rect 29420 33844 29426 33856
rect 30193 33847 30251 33853
rect 30193 33844 30205 33847
rect 29420 33816 30205 33844
rect 29420 33804 29426 33816
rect 30193 33813 30205 33816
rect 30239 33813 30251 33847
rect 30193 33807 30251 33813
rect 30466 33804 30472 33856
rect 30524 33804 30530 33856
rect 30944 33844 30972 33884
rect 31113 33881 31125 33915
rect 31159 33912 31171 33915
rect 31941 33915 31999 33921
rect 31941 33912 31953 33915
rect 31159 33884 31953 33912
rect 31159 33881 31171 33884
rect 31113 33875 31171 33881
rect 31941 33881 31953 33884
rect 31987 33881 31999 33915
rect 31941 33875 31999 33881
rect 32122 33872 32128 33924
rect 32180 33921 32186 33924
rect 32180 33915 32208 33921
rect 32196 33881 32208 33915
rect 32180 33875 32208 33881
rect 32180 33872 32186 33875
rect 31573 33847 31631 33853
rect 31573 33844 31585 33847
rect 30944 33816 31585 33844
rect 31573 33813 31585 33816
rect 31619 33813 31631 33847
rect 31573 33807 31631 33813
rect 32306 33804 32312 33856
rect 32364 33804 32370 33856
rect 32674 33804 32680 33856
rect 32732 33844 32738 33856
rect 33778 33844 33784 33856
rect 32732 33816 33784 33844
rect 32732 33804 32738 33816
rect 33778 33804 33784 33816
rect 33836 33844 33842 33856
rect 34348 33844 34376 33943
rect 34514 33940 34520 33992
rect 34572 33980 34578 33992
rect 34701 33983 34759 33989
rect 34701 33980 34713 33983
rect 34572 33952 34713 33980
rect 34572 33940 34578 33952
rect 34701 33949 34713 33952
rect 34747 33949 34759 33983
rect 34701 33943 34759 33949
rect 34882 33940 34888 33992
rect 34940 33940 34946 33992
rect 36633 33983 36691 33989
rect 36633 33980 36645 33983
rect 35912 33952 36645 33980
rect 35912 33921 35940 33952
rect 36633 33949 36645 33952
rect 36679 33949 36691 33983
rect 38105 33983 38163 33989
rect 38105 33980 38117 33983
rect 36633 33943 36691 33949
rect 37246 33952 38117 33980
rect 35897 33915 35955 33921
rect 35897 33912 35909 33915
rect 35360 33884 35909 33912
rect 35360 33856 35388 33884
rect 35897 33881 35909 33884
rect 35943 33881 35955 33915
rect 35897 33875 35955 33881
rect 36081 33915 36139 33921
rect 36081 33881 36093 33915
rect 36127 33912 36139 33915
rect 36354 33912 36360 33924
rect 36127 33884 36360 33912
rect 36127 33881 36139 33884
rect 36081 33875 36139 33881
rect 36354 33872 36360 33884
rect 36412 33912 36418 33924
rect 36541 33915 36599 33921
rect 36541 33912 36553 33915
rect 36412 33884 36553 33912
rect 36412 33872 36418 33884
rect 36541 33881 36553 33884
rect 36587 33881 36599 33915
rect 36541 33875 36599 33881
rect 36725 33915 36783 33921
rect 36725 33881 36737 33915
rect 36771 33912 36783 33915
rect 37246 33912 37274 33952
rect 38105 33949 38117 33952
rect 38151 33949 38163 33983
rect 38105 33943 38163 33949
rect 36771 33884 37274 33912
rect 36771 33881 36783 33884
rect 36725 33875 36783 33881
rect 33836 33816 34376 33844
rect 33836 33804 33842 33816
rect 34606 33804 34612 33856
rect 34664 33844 34670 33856
rect 35069 33847 35127 33853
rect 35069 33844 35081 33847
rect 34664 33816 35081 33844
rect 34664 33804 34670 33816
rect 35069 33813 35081 33816
rect 35115 33813 35127 33847
rect 35069 33807 35127 33813
rect 35342 33804 35348 33856
rect 35400 33804 35406 33856
rect 35434 33804 35440 33856
rect 35492 33844 35498 33856
rect 35529 33847 35587 33853
rect 35529 33844 35541 33847
rect 35492 33816 35541 33844
rect 35492 33804 35498 33816
rect 35529 33813 35541 33816
rect 35575 33813 35587 33847
rect 35529 33807 35587 33813
rect 35710 33804 35716 33856
rect 35768 33844 35774 33856
rect 35989 33847 36047 33853
rect 35989 33844 36001 33847
rect 35768 33816 36001 33844
rect 35768 33804 35774 33816
rect 35989 33813 36001 33816
rect 36035 33844 36047 33847
rect 36740 33844 36768 33875
rect 37366 33872 37372 33924
rect 37424 33872 37430 33924
rect 37826 33872 37832 33924
rect 37884 33912 37890 33924
rect 37921 33915 37979 33921
rect 37921 33912 37933 33915
rect 37884 33884 37933 33912
rect 37884 33872 37890 33884
rect 37921 33881 37933 33884
rect 37967 33881 37979 33915
rect 37921 33875 37979 33881
rect 36035 33816 36768 33844
rect 36035 33813 36047 33816
rect 35989 33807 36047 33813
rect 1104 33754 41400 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 41400 33754
rect 1104 33680 41400 33702
rect 6549 33643 6607 33649
rect 4264 33612 5304 33640
rect 4264 33513 4292 33612
rect 4341 33575 4399 33581
rect 4341 33541 4353 33575
rect 4387 33572 4399 33575
rect 4525 33575 4583 33581
rect 4525 33572 4537 33575
rect 4387 33544 4537 33572
rect 4387 33541 4399 33544
rect 4341 33535 4399 33541
rect 4525 33541 4537 33544
rect 4571 33541 4583 33575
rect 5276 33572 5304 33612
rect 6549 33609 6561 33643
rect 6595 33640 6607 33643
rect 6822 33640 6828 33652
rect 6595 33612 6828 33640
rect 6595 33609 6607 33612
rect 6549 33603 6607 33609
rect 6822 33600 6828 33612
rect 6880 33600 6886 33652
rect 6914 33600 6920 33652
rect 6972 33600 6978 33652
rect 9674 33600 9680 33652
rect 9732 33640 9738 33652
rect 9861 33643 9919 33649
rect 9861 33640 9873 33643
rect 9732 33612 9873 33640
rect 9732 33600 9738 33612
rect 9861 33609 9873 33612
rect 9907 33640 9919 33643
rect 11615 33643 11673 33649
rect 9907 33612 10180 33640
rect 9907 33609 9919 33612
rect 9861 33603 9919 33609
rect 5902 33572 5908 33584
rect 4525 33535 4583 33541
rect 4724 33544 5120 33572
rect 4249 33507 4307 33513
rect 4249 33473 4261 33507
rect 4295 33473 4307 33507
rect 4249 33467 4307 33473
rect 4430 33464 4436 33516
rect 4488 33504 4494 33516
rect 4724 33504 4752 33544
rect 4488 33476 4752 33504
rect 4801 33507 4859 33513
rect 4488 33464 4494 33476
rect 4801 33473 4813 33507
rect 4847 33504 4859 33507
rect 4890 33504 4896 33516
rect 4847 33476 4896 33504
rect 4847 33473 4859 33476
rect 4801 33467 4859 33473
rect 4890 33464 4896 33476
rect 4948 33464 4954 33516
rect 5092 33445 5120 33544
rect 5276 33544 5908 33572
rect 5276 33516 5304 33544
rect 5902 33532 5908 33544
rect 5960 33532 5966 33584
rect 6365 33575 6423 33581
rect 6365 33541 6377 33575
rect 6411 33572 6423 33575
rect 6730 33572 6736 33584
rect 6411 33544 6736 33572
rect 6411 33541 6423 33544
rect 6365 33535 6423 33541
rect 6730 33532 6736 33544
rect 6788 33532 6794 33584
rect 5258 33464 5264 33516
rect 5316 33464 5322 33516
rect 6270 33464 6276 33516
rect 6328 33464 6334 33516
rect 6641 33507 6699 33513
rect 6641 33473 6653 33507
rect 6687 33504 6699 33507
rect 6932 33504 6960 33600
rect 7466 33532 7472 33584
rect 7524 33572 7530 33584
rect 7837 33575 7895 33581
rect 7837 33572 7849 33575
rect 7524 33544 7849 33572
rect 7524 33532 7530 33544
rect 7837 33541 7849 33544
rect 7883 33572 7895 33575
rect 7883 33544 9628 33572
rect 7883 33541 7895 33544
rect 7837 33535 7895 33541
rect 6687 33476 6960 33504
rect 6687 33473 6699 33476
rect 6641 33467 6699 33473
rect 8662 33464 8668 33516
rect 8720 33504 8726 33516
rect 9122 33504 9128 33516
rect 8720 33476 9128 33504
rect 8720 33464 8726 33476
rect 9122 33464 9128 33476
rect 9180 33464 9186 33516
rect 9493 33507 9551 33513
rect 9493 33473 9505 33507
rect 9539 33473 9551 33507
rect 9493 33467 9551 33473
rect 4709 33439 4767 33445
rect 4709 33405 4721 33439
rect 4755 33405 4767 33439
rect 4709 33399 4767 33405
rect 5077 33439 5135 33445
rect 5077 33405 5089 33439
rect 5123 33436 5135 33439
rect 6288 33436 6316 33464
rect 5123 33408 6316 33436
rect 5123 33405 5135 33408
rect 5077 33399 5135 33405
rect 4724 33368 4752 33399
rect 5445 33371 5503 33377
rect 5445 33368 5457 33371
rect 4724 33340 5457 33368
rect 5445 33337 5457 33340
rect 5491 33337 5503 33371
rect 5445 33331 5503 33337
rect 5810 33328 5816 33380
rect 5868 33368 5874 33380
rect 6365 33371 6423 33377
rect 6365 33368 6377 33371
rect 5868 33340 6377 33368
rect 5868 33328 5874 33340
rect 6365 33337 6377 33340
rect 6411 33337 6423 33371
rect 6365 33331 6423 33337
rect 4522 33260 4528 33312
rect 4580 33260 4586 33312
rect 4982 33260 4988 33312
rect 5040 33260 5046 33312
rect 9508 33300 9536 33467
rect 9600 33436 9628 33544
rect 9692 33544 10089 33572
rect 9692 33516 9720 33544
rect 9674 33464 9680 33516
rect 9732 33464 9738 33516
rect 9953 33507 10011 33513
rect 9953 33473 9965 33507
rect 9999 33473 10011 33507
rect 9953 33467 10011 33473
rect 9858 33436 9864 33448
rect 9600 33408 9864 33436
rect 9858 33396 9864 33408
rect 9916 33396 9922 33448
rect 9968 33368 9996 33467
rect 10061 33436 10089 33544
rect 10152 33513 10180 33612
rect 11615 33609 11627 33643
rect 11661 33640 11673 33643
rect 11882 33640 11888 33652
rect 11661 33612 11888 33640
rect 11661 33609 11673 33612
rect 11615 33603 11673 33609
rect 11882 33600 11888 33612
rect 11940 33600 11946 33652
rect 12066 33600 12072 33652
rect 12124 33600 12130 33652
rect 12618 33600 12624 33652
rect 12676 33600 12682 33652
rect 13265 33643 13323 33649
rect 13265 33609 13277 33643
rect 13311 33640 13323 33643
rect 13446 33640 13452 33652
rect 13311 33612 13452 33640
rect 13311 33609 13323 33612
rect 13265 33603 13323 33609
rect 13446 33600 13452 33612
rect 13504 33600 13510 33652
rect 14458 33600 14464 33652
rect 14516 33640 14522 33652
rect 14651 33643 14709 33649
rect 14651 33640 14663 33643
rect 14516 33612 14663 33640
rect 14516 33600 14522 33612
rect 14651 33609 14663 33612
rect 14697 33609 14709 33643
rect 14651 33603 14709 33609
rect 14737 33643 14795 33649
rect 14737 33609 14749 33643
rect 14783 33640 14795 33643
rect 16485 33643 16543 33649
rect 14783 33612 16436 33640
rect 14783 33609 14795 33612
rect 14737 33603 14795 33609
rect 11514 33532 11520 33584
rect 11572 33532 11578 33584
rect 12084 33572 12112 33600
rect 13170 33572 13176 33584
rect 12084 33544 13176 33572
rect 10137 33507 10195 33513
rect 10137 33473 10149 33507
rect 10183 33473 10195 33507
rect 10137 33467 10195 33473
rect 10229 33507 10287 33513
rect 10229 33473 10241 33507
rect 10275 33504 10287 33507
rect 11330 33504 11336 33516
rect 10275 33476 11336 33504
rect 10275 33473 10287 33476
rect 10229 33467 10287 33473
rect 11330 33464 11336 33476
rect 11388 33464 11394 33516
rect 11701 33507 11759 33513
rect 11701 33473 11713 33507
rect 11747 33473 11759 33507
rect 11701 33467 11759 33473
rect 11793 33507 11851 33513
rect 11793 33473 11805 33507
rect 11839 33504 11851 33507
rect 12084 33504 12112 33544
rect 13170 33532 13176 33544
rect 13228 33532 13234 33584
rect 13998 33532 14004 33584
rect 14056 33572 14062 33584
rect 14119 33575 14177 33581
rect 14119 33572 14131 33575
rect 14056 33544 14131 33572
rect 14056 33532 14062 33544
rect 14108 33541 14131 33544
rect 14165 33541 14177 33575
rect 14108 33535 14177 33541
rect 14309 33575 14367 33581
rect 14309 33541 14321 33575
rect 14355 33572 14367 33575
rect 14355 33544 14872 33572
rect 14355 33541 14367 33544
rect 14309 33535 14367 33541
rect 11839 33476 12112 33504
rect 12161 33507 12219 33513
rect 11839 33473 11851 33476
rect 11793 33467 11851 33473
rect 12161 33473 12173 33507
rect 12207 33504 12219 33507
rect 12618 33504 12624 33516
rect 12207 33476 12624 33504
rect 12207 33473 12219 33476
rect 12161 33467 12219 33473
rect 10318 33436 10324 33448
rect 10061 33408 10324 33436
rect 10318 33396 10324 33408
rect 10376 33396 10382 33448
rect 10870 33396 10876 33448
rect 10928 33436 10934 33448
rect 11716 33436 11744 33467
rect 12618 33464 12624 33476
rect 12676 33504 12682 33516
rect 12897 33507 12955 33513
rect 12897 33504 12909 33507
rect 12676 33476 12909 33504
rect 12676 33464 12682 33476
rect 12897 33473 12909 33476
rect 12943 33473 12955 33507
rect 12897 33467 12955 33473
rect 13078 33464 13084 33516
rect 13136 33464 13142 33516
rect 10928 33408 11744 33436
rect 10928 33396 10934 33408
rect 11146 33368 11152 33380
rect 9968 33340 11152 33368
rect 11146 33328 11152 33340
rect 11204 33328 11210 33380
rect 13188 33368 13216 33532
rect 14108 33504 14136 33535
rect 14844 33516 14872 33544
rect 14553 33507 14611 33513
rect 14553 33504 14565 33507
rect 14108 33476 14565 33504
rect 14553 33473 14565 33476
rect 14599 33504 14611 33507
rect 14642 33504 14648 33516
rect 14599 33476 14648 33504
rect 14599 33473 14611 33476
rect 14553 33467 14611 33473
rect 14642 33464 14648 33476
rect 14700 33464 14706 33516
rect 14826 33464 14832 33516
rect 14884 33464 14890 33516
rect 14461 33371 14519 33377
rect 14461 33368 14473 33371
rect 13188 33340 14473 33368
rect 14461 33337 14473 33340
rect 14507 33368 14519 33371
rect 14550 33368 14556 33380
rect 14507 33340 14556 33368
rect 14507 33337 14519 33340
rect 14461 33331 14519 33337
rect 14550 33328 14556 33340
rect 14608 33328 14614 33380
rect 10042 33300 10048 33312
rect 9508 33272 10048 33300
rect 10042 33260 10048 33272
rect 10100 33260 10106 33312
rect 10226 33260 10232 33312
rect 10284 33260 10290 33312
rect 10410 33260 10416 33312
rect 10468 33260 10474 33312
rect 12342 33260 12348 33312
rect 12400 33260 12406 33312
rect 14277 33303 14335 33309
rect 14277 33269 14289 33303
rect 14323 33300 14335 33303
rect 14936 33300 14964 33612
rect 16408 33572 16436 33612
rect 16485 33609 16497 33643
rect 16531 33640 16543 33643
rect 16850 33640 16856 33652
rect 16531 33612 16856 33640
rect 16531 33609 16543 33612
rect 16485 33603 16543 33609
rect 16850 33600 16856 33612
rect 16908 33600 16914 33652
rect 17126 33600 17132 33652
rect 17184 33600 17190 33652
rect 17678 33600 17684 33652
rect 17736 33600 17742 33652
rect 17770 33600 17776 33652
rect 17828 33600 17834 33652
rect 17862 33600 17868 33652
rect 17920 33600 17926 33652
rect 19996 33612 21036 33640
rect 17144 33572 17172 33600
rect 17788 33572 17816 33600
rect 16408 33544 17172 33572
rect 17604 33544 17816 33572
rect 16114 33464 16120 33516
rect 16172 33464 16178 33516
rect 16206 33464 16212 33516
rect 16264 33504 16270 33516
rect 16758 33504 16764 33516
rect 16264 33476 16764 33504
rect 16264 33464 16270 33476
rect 16758 33464 16764 33476
rect 16816 33464 16822 33516
rect 17310 33464 17316 33516
rect 17368 33504 17374 33516
rect 17604 33513 17632 33544
rect 17589 33507 17647 33513
rect 17368 33476 17540 33504
rect 17368 33464 17374 33476
rect 16022 33396 16028 33448
rect 16080 33396 16086 33448
rect 17218 33396 17224 33448
rect 17276 33396 17282 33448
rect 17512 33436 17540 33476
rect 17589 33473 17601 33507
rect 17635 33473 17647 33507
rect 17589 33467 17647 33473
rect 17773 33507 17831 33513
rect 17773 33473 17785 33507
rect 17819 33504 17831 33507
rect 17880 33504 17908 33600
rect 18230 33532 18236 33584
rect 18288 33572 18294 33584
rect 19996 33572 20024 33612
rect 18288 33544 20024 33572
rect 18288 33532 18294 33544
rect 17819 33476 17908 33504
rect 17819 33473 17831 33476
rect 17773 33467 17831 33473
rect 19426 33464 19432 33516
rect 19484 33464 19490 33516
rect 19518 33464 19524 33516
rect 19576 33464 19582 33516
rect 21008 33504 21036 33612
rect 22278 33600 22284 33652
rect 22336 33640 22342 33652
rect 23937 33643 23995 33649
rect 23937 33640 23949 33643
rect 22336 33612 23949 33640
rect 22336 33600 22342 33612
rect 23937 33609 23949 33612
rect 23983 33609 23995 33643
rect 23937 33603 23995 33609
rect 25130 33600 25136 33652
rect 25188 33600 25194 33652
rect 26694 33600 26700 33652
rect 26752 33600 26758 33652
rect 27522 33600 27528 33652
rect 27580 33640 27586 33652
rect 27982 33640 27988 33652
rect 27580 33612 27988 33640
rect 27580 33600 27586 33612
rect 27982 33600 27988 33612
rect 28040 33640 28046 33652
rect 30006 33640 30012 33652
rect 28040 33612 30012 33640
rect 28040 33600 28046 33612
rect 30006 33600 30012 33612
rect 30064 33600 30070 33652
rect 33226 33600 33232 33652
rect 33284 33600 33290 33652
rect 34333 33643 34391 33649
rect 34333 33609 34345 33643
rect 34379 33640 34391 33643
rect 34882 33640 34888 33652
rect 34379 33612 34888 33640
rect 34379 33609 34391 33612
rect 34333 33603 34391 33609
rect 34882 33600 34888 33612
rect 34940 33600 34946 33652
rect 35342 33600 35348 33652
rect 35400 33640 35406 33652
rect 35529 33643 35587 33649
rect 35529 33640 35541 33643
rect 35400 33612 35541 33640
rect 35400 33600 35406 33612
rect 35529 33609 35541 33612
rect 35575 33609 35587 33643
rect 36725 33643 36783 33649
rect 36725 33640 36737 33643
rect 35529 33603 35587 33609
rect 36188 33612 36737 33640
rect 23014 33572 23020 33584
rect 22296 33544 23020 33572
rect 21174 33504 21180 33516
rect 21008 33490 21180 33504
rect 21022 33476 21180 33490
rect 21174 33464 21180 33476
rect 21232 33464 21238 33516
rect 21913 33507 21971 33513
rect 21913 33473 21925 33507
rect 21959 33504 21971 33507
rect 22002 33504 22008 33516
rect 21959 33476 22008 33504
rect 21959 33473 21971 33476
rect 21913 33467 21971 33473
rect 22002 33464 22008 33476
rect 22060 33464 22066 33516
rect 22296 33513 22324 33544
rect 23014 33532 23020 33544
rect 23072 33572 23078 33584
rect 25148 33572 25176 33600
rect 23072 33544 25176 33572
rect 26712 33572 26740 33600
rect 28994 33572 29000 33584
rect 26712 33544 29000 33572
rect 23072 33532 23078 33544
rect 28994 33532 29000 33544
rect 29052 33532 29058 33584
rect 33594 33572 33600 33584
rect 32508 33544 33600 33572
rect 22281 33507 22339 33513
rect 22281 33473 22293 33507
rect 22327 33473 22339 33507
rect 22281 33467 22339 33473
rect 24121 33507 24179 33513
rect 24121 33473 24133 33507
rect 24167 33504 24179 33507
rect 24854 33504 24860 33516
rect 24167 33476 24860 33504
rect 24167 33473 24179 33476
rect 24121 33467 24179 33473
rect 24854 33464 24860 33476
rect 24912 33464 24918 33516
rect 25501 33507 25559 33513
rect 25501 33473 25513 33507
rect 25547 33473 25559 33507
rect 25501 33467 25559 33473
rect 18598 33436 18604 33448
rect 17512 33408 18604 33436
rect 18598 33396 18604 33408
rect 18656 33396 18662 33448
rect 19444 33436 19472 33464
rect 19613 33439 19671 33445
rect 19613 33436 19625 33439
rect 19444 33408 19625 33436
rect 19613 33405 19625 33408
rect 19659 33405 19671 33439
rect 20254 33436 20260 33448
rect 19613 33399 19671 33405
rect 19720 33408 20260 33436
rect 17862 33328 17868 33380
rect 17920 33368 17926 33380
rect 19720 33368 19748 33408
rect 20254 33396 20260 33408
rect 20312 33396 20318 33448
rect 24026 33436 24032 33448
rect 22388 33408 24032 33436
rect 22388 33380 22416 33408
rect 24026 33396 24032 33408
rect 24084 33436 24090 33448
rect 24397 33439 24455 33445
rect 24397 33436 24409 33439
rect 24084 33408 24409 33436
rect 24084 33396 24090 33408
rect 24397 33405 24409 33408
rect 24443 33436 24455 33439
rect 25516 33436 25544 33467
rect 25590 33464 25596 33516
rect 25648 33504 25654 33516
rect 25777 33507 25835 33513
rect 25777 33504 25789 33507
rect 25648 33476 25789 33504
rect 25648 33464 25654 33476
rect 25777 33473 25789 33476
rect 25823 33473 25835 33507
rect 25777 33467 25835 33473
rect 27249 33507 27307 33513
rect 27249 33473 27261 33507
rect 27295 33473 27307 33507
rect 27249 33467 27307 33473
rect 26970 33436 26976 33448
rect 24443 33408 26976 33436
rect 24443 33405 24455 33408
rect 24397 33399 24455 33405
rect 26970 33396 26976 33408
rect 27028 33396 27034 33448
rect 27264 33436 27292 33467
rect 27338 33464 27344 33516
rect 27396 33504 27402 33516
rect 30466 33504 30472 33516
rect 27396 33476 30472 33504
rect 27396 33464 27402 33476
rect 30466 33464 30472 33476
rect 30524 33464 30530 33516
rect 32214 33464 32220 33516
rect 32272 33504 32278 33516
rect 32508 33513 32536 33544
rect 33594 33532 33600 33544
rect 33652 33532 33658 33584
rect 33778 33532 33784 33584
rect 33836 33572 33842 33584
rect 35544 33572 35572 33603
rect 36188 33584 36216 33612
rect 36725 33609 36737 33612
rect 36771 33609 36783 33643
rect 36725 33603 36783 33609
rect 33836 33544 34100 33572
rect 35544 33544 35903 33572
rect 33836 33532 33842 33544
rect 32309 33507 32367 33513
rect 32309 33504 32321 33507
rect 32272 33476 32321 33504
rect 32272 33464 32278 33476
rect 32309 33473 32321 33476
rect 32355 33473 32367 33507
rect 32309 33467 32367 33473
rect 32493 33507 32551 33513
rect 32493 33473 32505 33507
rect 32539 33473 32551 33507
rect 32493 33467 32551 33473
rect 32950 33464 32956 33516
rect 33008 33504 33014 33516
rect 33045 33507 33103 33513
rect 33045 33504 33057 33507
rect 33008 33476 33057 33504
rect 33008 33464 33014 33476
rect 33045 33473 33057 33476
rect 33091 33504 33103 33507
rect 33962 33504 33968 33516
rect 33091 33476 33968 33504
rect 33091 33473 33103 33476
rect 33045 33467 33103 33473
rect 33962 33464 33968 33476
rect 34020 33464 34026 33516
rect 34072 33504 34100 33544
rect 34174 33507 34232 33513
rect 34174 33504 34186 33507
rect 34072 33476 34186 33504
rect 34174 33473 34186 33476
rect 34220 33473 34232 33507
rect 34174 33467 34232 33473
rect 35345 33507 35403 33513
rect 35345 33473 35357 33507
rect 35391 33473 35403 33507
rect 35345 33467 35403 33473
rect 28902 33436 28908 33448
rect 27264 33408 28908 33436
rect 28902 33396 28908 33408
rect 28960 33436 28966 33448
rect 29454 33436 29460 33448
rect 28960 33408 29460 33436
rect 28960 33396 28966 33408
rect 29454 33396 29460 33408
rect 29512 33396 29518 33448
rect 30282 33396 30288 33448
rect 30340 33436 30346 33448
rect 32585 33439 32643 33445
rect 32585 33436 32597 33439
rect 30340 33408 32597 33436
rect 30340 33396 30346 33408
rect 32585 33405 32597 33408
rect 32631 33436 32643 33439
rect 32674 33436 32680 33448
rect 32631 33408 32680 33436
rect 32631 33405 32643 33408
rect 32585 33399 32643 33405
rect 32674 33396 32680 33408
rect 32732 33436 32738 33448
rect 33413 33439 33471 33445
rect 33413 33436 33425 33439
rect 32732 33408 33425 33436
rect 32732 33396 32738 33408
rect 33413 33405 33425 33408
rect 33459 33405 33471 33439
rect 33413 33399 33471 33405
rect 33594 33396 33600 33448
rect 33652 33436 33658 33448
rect 33689 33439 33747 33445
rect 33689 33436 33701 33439
rect 33652 33408 33701 33436
rect 33652 33396 33658 33408
rect 33689 33405 33701 33408
rect 33735 33405 33747 33439
rect 33689 33399 33747 33405
rect 34057 33439 34115 33445
rect 34057 33405 34069 33439
rect 34103 33405 34115 33439
rect 35366 33436 35394 33467
rect 35710 33464 35716 33516
rect 35768 33464 35774 33516
rect 35875 33513 35903 33544
rect 36170 33532 36176 33584
rect 36228 33532 36234 33584
rect 37844 33544 38608 33572
rect 35860 33507 35918 33513
rect 35860 33473 35872 33507
rect 35906 33473 35918 33507
rect 35860 33467 35918 33473
rect 35986 33436 35992 33448
rect 35366 33408 35992 33436
rect 34057 33399 34115 33405
rect 17920 33340 19748 33368
rect 17920 33328 17926 33340
rect 22094 33328 22100 33380
rect 22152 33328 22158 33380
rect 22370 33328 22376 33380
rect 22428 33328 22434 33380
rect 24305 33371 24363 33377
rect 24305 33337 24317 33371
rect 24351 33368 24363 33371
rect 24351 33340 25452 33368
rect 24351 33337 24363 33340
rect 24305 33331 24363 33337
rect 14323 33272 14964 33300
rect 14323 33269 14335 33272
rect 14277 33263 14335 33269
rect 15654 33260 15660 33312
rect 15712 33300 15718 33312
rect 16942 33300 16948 33312
rect 15712 33272 16948 33300
rect 15712 33260 15718 33272
rect 16942 33260 16948 33272
rect 17000 33260 17006 33312
rect 19337 33303 19395 33309
rect 19337 33269 19349 33303
rect 19383 33300 19395 33303
rect 19870 33303 19928 33309
rect 19870 33300 19882 33303
rect 19383 33272 19882 33300
rect 19383 33269 19395 33272
rect 19337 33263 19395 33269
rect 19870 33269 19882 33272
rect 19916 33269 19928 33303
rect 19870 33263 19928 33269
rect 20254 33260 20260 33312
rect 20312 33300 20318 33312
rect 20898 33300 20904 33312
rect 20312 33272 20904 33300
rect 20312 33260 20318 33272
rect 20898 33260 20904 33272
rect 20956 33260 20962 33312
rect 21358 33260 21364 33312
rect 21416 33260 21422 33312
rect 22112 33300 22140 33328
rect 25222 33300 25228 33312
rect 22112 33272 25228 33300
rect 25222 33260 25228 33272
rect 25280 33260 25286 33312
rect 25314 33260 25320 33312
rect 25372 33260 25378 33312
rect 25424 33300 25452 33340
rect 25498 33328 25504 33380
rect 25556 33368 25562 33380
rect 25593 33371 25651 33377
rect 25593 33368 25605 33371
rect 25556 33340 25605 33368
rect 25556 33328 25562 33340
rect 25593 33337 25605 33340
rect 25639 33337 25651 33371
rect 25593 33331 25651 33337
rect 25682 33328 25688 33380
rect 25740 33368 25746 33380
rect 28810 33368 28816 33380
rect 25740 33340 28816 33368
rect 25740 33328 25746 33340
rect 28810 33328 28816 33340
rect 28868 33328 28874 33380
rect 34072 33368 34100 33399
rect 35986 33396 35992 33408
rect 36044 33396 36050 33448
rect 36081 33439 36139 33445
rect 36081 33405 36093 33439
rect 36127 33436 36139 33439
rect 36188 33436 36216 33532
rect 37844 33516 37872 33544
rect 36541 33507 36599 33513
rect 36541 33473 36553 33507
rect 36587 33504 36599 33507
rect 37274 33504 37280 33516
rect 36587 33476 37280 33504
rect 36587 33473 36599 33476
rect 36541 33467 36599 33473
rect 37274 33464 37280 33476
rect 37332 33464 37338 33516
rect 37826 33464 37832 33516
rect 37884 33464 37890 33516
rect 37921 33507 37979 33513
rect 37921 33473 37933 33507
rect 37967 33473 37979 33507
rect 37921 33467 37979 33473
rect 36127 33408 36216 33436
rect 36127 33405 36139 33408
rect 36081 33399 36139 33405
rect 36630 33396 36636 33448
rect 36688 33436 36694 33448
rect 37553 33439 37611 33445
rect 37553 33436 37565 33439
rect 36688 33408 37565 33436
rect 36688 33396 36694 33408
rect 37553 33405 37565 33408
rect 37599 33405 37611 33439
rect 37553 33399 37611 33405
rect 37936 33436 37964 33467
rect 38010 33464 38016 33516
rect 38068 33504 38074 33516
rect 38289 33507 38347 33513
rect 38289 33504 38301 33507
rect 38068 33476 38301 33504
rect 38068 33464 38074 33476
rect 38289 33473 38301 33476
rect 38335 33473 38347 33507
rect 38580 33504 38608 33544
rect 38657 33507 38715 33513
rect 38657 33504 38669 33507
rect 38580 33476 38669 33504
rect 38289 33467 38347 33473
rect 38657 33473 38669 33476
rect 38703 33473 38715 33507
rect 38657 33467 38715 33473
rect 40586 33464 40592 33516
rect 40644 33464 40650 33516
rect 37936 33408 38424 33436
rect 33428 33340 34100 33368
rect 25700 33300 25728 33328
rect 25424 33272 25728 33300
rect 25774 33260 25780 33312
rect 25832 33300 25838 33312
rect 26326 33300 26332 33312
rect 25832 33272 26332 33300
rect 25832 33260 25838 33272
rect 26326 33260 26332 33272
rect 26384 33260 26390 33312
rect 26786 33260 26792 33312
rect 26844 33300 26850 33312
rect 27430 33300 27436 33312
rect 26844 33272 27436 33300
rect 26844 33260 26850 33272
rect 27430 33260 27436 33272
rect 27488 33260 27494 33312
rect 27614 33260 27620 33312
rect 27672 33300 27678 33312
rect 30558 33300 30564 33312
rect 27672 33272 30564 33300
rect 27672 33260 27678 33272
rect 30558 33260 30564 33272
rect 30616 33260 30622 33312
rect 32122 33260 32128 33312
rect 32180 33260 32186 33312
rect 32766 33260 32772 33312
rect 32824 33300 32830 33312
rect 33428 33309 33456 33340
rect 33413 33303 33471 33309
rect 33413 33300 33425 33303
rect 32824 33272 33425 33300
rect 32824 33260 32830 33272
rect 33413 33269 33425 33272
rect 33459 33269 33471 33303
rect 34072 33300 34100 33340
rect 34330 33328 34336 33380
rect 34388 33368 34394 33380
rect 36173 33371 36231 33377
rect 36173 33368 36185 33371
rect 34388 33340 36185 33368
rect 34388 33328 34394 33340
rect 36173 33337 36185 33340
rect 36219 33337 36231 33371
rect 36173 33331 36231 33337
rect 36354 33328 36360 33380
rect 36412 33368 36418 33380
rect 37936 33368 37964 33408
rect 38396 33380 38424 33408
rect 39206 33396 39212 33448
rect 39264 33396 39270 33448
rect 39485 33439 39543 33445
rect 39485 33405 39497 33439
rect 39531 33436 39543 33439
rect 41046 33436 41052 33448
rect 39531 33408 41052 33436
rect 39531 33405 39543 33408
rect 39485 33399 39543 33405
rect 41046 33396 41052 33408
rect 41104 33396 41110 33448
rect 36412 33340 37964 33368
rect 36412 33328 36418 33340
rect 38378 33328 38384 33380
rect 38436 33328 38442 33380
rect 35710 33300 35716 33312
rect 34072 33272 35716 33300
rect 33413 33263 33471 33269
rect 35710 33260 35716 33272
rect 35768 33260 35774 33312
rect 35989 33303 36047 33309
rect 35989 33269 36001 33303
rect 36035 33300 36047 33303
rect 36372 33300 36400 33328
rect 36035 33272 36400 33300
rect 36035 33269 36047 33272
rect 35989 33263 36047 33269
rect 40954 33260 40960 33312
rect 41012 33260 41018 33312
rect 1104 33210 41400 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 41400 33210
rect 1104 33136 41400 33158
rect 7282 33056 7288 33108
rect 7340 33056 7346 33108
rect 11146 33056 11152 33108
rect 11204 33056 11210 33108
rect 12069 33099 12127 33105
rect 12069 33065 12081 33099
rect 12115 33096 12127 33099
rect 14550 33096 14556 33108
rect 12115 33068 14556 33096
rect 12115 33065 12127 33068
rect 12069 33059 12127 33065
rect 14550 33056 14556 33068
rect 14608 33056 14614 33108
rect 15838 33056 15844 33108
rect 15896 33056 15902 33108
rect 15933 33099 15991 33105
rect 15933 33065 15945 33099
rect 15979 33096 15991 33099
rect 16114 33096 16120 33108
rect 15979 33068 16120 33096
rect 15979 33065 15991 33068
rect 15933 33059 15991 33065
rect 16114 33056 16120 33068
rect 16172 33056 16178 33108
rect 16758 33056 16764 33108
rect 16816 33096 16822 33108
rect 17589 33099 17647 33105
rect 17589 33096 17601 33099
rect 16816 33068 17601 33096
rect 16816 33056 16822 33068
rect 17589 33065 17601 33068
rect 17635 33065 17647 33099
rect 17589 33059 17647 33065
rect 19518 33056 19524 33108
rect 19576 33056 19582 33108
rect 20438 33056 20444 33108
rect 20496 33096 20502 33108
rect 22649 33099 22707 33105
rect 22649 33096 22661 33099
rect 20496 33068 22661 33096
rect 20496 33056 20502 33068
rect 22649 33065 22661 33068
rect 22695 33065 22707 33099
rect 22649 33059 22707 33065
rect 24762 33056 24768 33108
rect 24820 33056 24826 33108
rect 26053 33099 26111 33105
rect 26053 33065 26065 33099
rect 26099 33096 26111 33099
rect 26510 33096 26516 33108
rect 26099 33068 26516 33096
rect 26099 33065 26111 33068
rect 26053 33059 26111 33065
rect 26510 33056 26516 33068
rect 26568 33056 26574 33108
rect 30653 33099 30711 33105
rect 30653 33096 30665 33099
rect 27540 33068 30665 33096
rect 7098 32988 7104 33040
rect 7156 33028 7162 33040
rect 8018 33028 8024 33040
rect 7156 33000 8024 33028
rect 7156 32988 7162 33000
rect 8018 32988 8024 33000
rect 8076 32988 8082 33040
rect 11164 33028 11192 33056
rect 12253 33031 12311 33037
rect 12253 33028 12265 33031
rect 11164 33000 12265 33028
rect 12253 32997 12265 33000
rect 12299 32997 12311 33031
rect 14568 33028 14596 33056
rect 14568 33000 16068 33028
rect 12253 32991 12311 32997
rect 10778 32920 10784 32972
rect 10836 32960 10842 32972
rect 15930 32960 15936 32972
rect 10836 32932 15936 32960
rect 10836 32920 10842 32932
rect 15930 32920 15936 32932
rect 15988 32920 15994 32972
rect 16040 32969 16068 33000
rect 23382 32988 23388 33040
rect 23440 33028 23446 33040
rect 24489 33031 24547 33037
rect 24489 33028 24501 33031
rect 23440 33000 24501 33028
rect 23440 32988 23446 33000
rect 24489 32997 24501 33000
rect 24535 32997 24547 33031
rect 24780 33028 24808 33056
rect 24489 32991 24547 32997
rect 24596 33000 24808 33028
rect 16025 32963 16083 32969
rect 16025 32929 16037 32963
rect 16071 32960 16083 32963
rect 16485 32963 16543 32969
rect 16485 32960 16497 32963
rect 16071 32932 16497 32960
rect 16071 32929 16083 32932
rect 16025 32923 16083 32929
rect 16485 32929 16497 32932
rect 16531 32929 16543 32963
rect 16485 32923 16543 32929
rect 20162 32920 20168 32972
rect 20220 32920 20226 32972
rect 21358 32960 21364 32972
rect 20732 32932 21364 32960
rect 7190 32852 7196 32904
rect 7248 32852 7254 32904
rect 11606 32852 11612 32904
rect 11664 32852 11670 32904
rect 11701 32895 11759 32901
rect 11701 32861 11713 32895
rect 11747 32892 11759 32895
rect 11747 32864 12020 32892
rect 11747 32861 11759 32864
rect 11701 32855 11759 32861
rect 11992 32836 12020 32864
rect 12066 32852 12072 32904
rect 12124 32852 12130 32904
rect 15654 32852 15660 32904
rect 15712 32892 15718 32904
rect 15749 32895 15807 32901
rect 15749 32892 15761 32895
rect 15712 32864 15761 32892
rect 15712 32852 15718 32864
rect 15749 32861 15761 32864
rect 15795 32861 15807 32895
rect 15749 32855 15807 32861
rect 16135 32895 16193 32901
rect 16135 32861 16147 32895
rect 16181 32892 16193 32895
rect 17310 32892 17316 32904
rect 16181 32864 17316 32892
rect 16181 32861 16193 32864
rect 16135 32855 16193 32861
rect 11974 32784 11980 32836
rect 12032 32824 12038 32836
rect 13998 32824 14004 32836
rect 12032 32796 14004 32824
rect 12032 32784 12038 32796
rect 13998 32784 14004 32796
rect 14056 32784 14062 32836
rect 15764 32824 15792 32855
rect 17310 32852 17316 32864
rect 17368 32852 17374 32904
rect 17497 32895 17555 32901
rect 17497 32861 17509 32895
rect 17543 32892 17555 32895
rect 19889 32895 19947 32901
rect 17543 32864 18092 32892
rect 17543 32861 17555 32864
rect 17497 32855 17555 32861
rect 15930 32824 15936 32836
rect 15764 32796 15936 32824
rect 15930 32784 15936 32796
rect 15988 32784 15994 32836
rect 16301 32827 16359 32833
rect 16301 32824 16313 32827
rect 16040 32796 16313 32824
rect 7650 32716 7656 32768
rect 7708 32716 7714 32768
rect 9858 32716 9864 32768
rect 9916 32756 9922 32768
rect 15654 32756 15660 32768
rect 9916 32728 15660 32756
rect 9916 32716 9922 32728
rect 15654 32716 15660 32728
rect 15712 32716 15718 32768
rect 15838 32716 15844 32768
rect 15896 32756 15902 32768
rect 16040 32756 16068 32796
rect 16301 32793 16313 32796
rect 16347 32793 16359 32827
rect 16301 32787 16359 32793
rect 18064 32768 18092 32864
rect 19889 32861 19901 32895
rect 19935 32892 19947 32895
rect 20732 32892 20760 32932
rect 21358 32920 21364 32932
rect 21416 32920 21422 32972
rect 19935 32864 20760 32892
rect 20809 32895 20867 32901
rect 19935 32861 19947 32864
rect 19889 32855 19947 32861
rect 20809 32861 20821 32895
rect 20855 32892 20867 32895
rect 20990 32892 20996 32904
rect 20855 32864 20996 32892
rect 20855 32861 20867 32864
rect 20809 32855 20867 32861
rect 20990 32852 20996 32864
rect 21048 32852 21054 32904
rect 21085 32895 21143 32901
rect 21085 32861 21097 32895
rect 21131 32892 21143 32895
rect 21174 32892 21180 32904
rect 21131 32864 21180 32892
rect 21131 32861 21143 32864
rect 21085 32855 21143 32861
rect 21174 32852 21180 32864
rect 21232 32852 21238 32904
rect 22833 32895 22891 32901
rect 22833 32892 22845 32895
rect 22296 32864 22845 32892
rect 22296 32768 22324 32864
rect 22833 32861 22845 32864
rect 22879 32861 22891 32895
rect 22833 32855 22891 32861
rect 24489 32895 24547 32901
rect 24489 32861 24501 32895
rect 24535 32892 24547 32895
rect 24596 32892 24624 33000
rect 24670 32920 24676 32972
rect 24728 32920 24734 32972
rect 25866 32920 25872 32972
rect 25924 32960 25930 32972
rect 27246 32960 27252 32972
rect 25924 32932 27252 32960
rect 25924 32920 25930 32932
rect 27246 32920 27252 32932
rect 27304 32920 27310 32972
rect 27540 32904 27568 33068
rect 30653 33065 30665 33068
rect 30699 33065 30711 33099
rect 30653 33059 30711 33065
rect 35986 33056 35992 33108
rect 36044 33096 36050 33108
rect 36449 33099 36507 33105
rect 36449 33096 36461 33099
rect 36044 33068 36461 33096
rect 36044 33056 36050 33068
rect 36449 33065 36461 33068
rect 36495 33065 36507 33099
rect 36449 33059 36507 33065
rect 30282 32988 30288 33040
rect 30340 33028 30346 33040
rect 34149 33031 34207 33037
rect 34149 33028 34161 33031
rect 30340 33000 34161 33028
rect 30340 32988 30346 33000
rect 34149 32997 34161 33000
rect 34195 32997 34207 33031
rect 34149 32991 34207 32997
rect 36354 32988 36360 33040
rect 36412 32988 36418 33040
rect 24765 32895 24823 32901
rect 24765 32892 24777 32895
rect 24535 32864 24624 32892
rect 24688 32864 24777 32892
rect 24535 32861 24547 32864
rect 24489 32855 24547 32861
rect 22557 32827 22615 32833
rect 22557 32793 22569 32827
rect 22603 32793 22615 32827
rect 22557 32787 22615 32793
rect 15896 32728 16068 32756
rect 15896 32716 15902 32728
rect 18046 32716 18052 32768
rect 18104 32716 18110 32768
rect 19978 32716 19984 32768
rect 20036 32716 20042 32768
rect 20070 32716 20076 32768
rect 20128 32756 20134 32768
rect 21818 32756 21824 32768
rect 20128 32728 21824 32756
rect 20128 32716 20134 32728
rect 21818 32716 21824 32728
rect 21876 32716 21882 32768
rect 22278 32716 22284 32768
rect 22336 32716 22342 32768
rect 22572 32756 22600 32787
rect 22738 32784 22744 32836
rect 22796 32784 22802 32836
rect 24688 32768 24716 32864
rect 24765 32861 24777 32864
rect 24811 32861 24823 32895
rect 24765 32855 24823 32861
rect 25314 32852 25320 32904
rect 25372 32892 25378 32904
rect 25777 32895 25835 32901
rect 25777 32892 25789 32895
rect 25372 32864 25789 32892
rect 25372 32852 25378 32864
rect 25777 32861 25789 32864
rect 25823 32861 25835 32895
rect 25777 32855 25835 32861
rect 25961 32895 26019 32901
rect 25961 32861 25973 32895
rect 26007 32861 26019 32895
rect 25961 32855 26019 32861
rect 24854 32784 24860 32836
rect 24912 32784 24918 32836
rect 25976 32824 26004 32855
rect 26050 32852 26056 32904
rect 26108 32852 26114 32904
rect 26694 32852 26700 32904
rect 26752 32892 26758 32904
rect 27154 32892 27160 32904
rect 26752 32864 27160 32892
rect 26752 32852 26758 32864
rect 27154 32852 27160 32864
rect 27212 32892 27218 32904
rect 27522 32892 27528 32904
rect 27212 32864 27528 32892
rect 27212 32852 27218 32864
rect 27522 32852 27528 32864
rect 27580 32852 27586 32904
rect 28074 32852 28080 32904
rect 28132 32892 28138 32904
rect 30374 32892 30380 32904
rect 28132 32864 30380 32892
rect 28132 32852 28138 32864
rect 30374 32852 30380 32864
rect 30432 32852 30438 32904
rect 30561 32895 30619 32901
rect 30561 32861 30573 32895
rect 30607 32892 30619 32895
rect 30650 32892 30656 32904
rect 30607 32864 30656 32892
rect 30607 32861 30619 32864
rect 30561 32855 30619 32861
rect 30650 32852 30656 32864
rect 30708 32852 30714 32904
rect 33873 32895 33931 32901
rect 33873 32861 33885 32895
rect 33919 32861 33931 32895
rect 33873 32855 33931 32861
rect 33965 32895 34023 32901
rect 33965 32861 33977 32895
rect 34011 32861 34023 32895
rect 33965 32855 34023 32861
rect 25976 32796 26372 32824
rect 26344 32768 26372 32796
rect 26602 32784 26608 32836
rect 26660 32824 26666 32836
rect 27430 32824 27436 32836
rect 26660 32796 27436 32824
rect 26660 32784 26666 32796
rect 27430 32784 27436 32796
rect 27488 32784 27494 32836
rect 28258 32784 28264 32836
rect 28316 32824 28322 32836
rect 28316 32796 30880 32824
rect 28316 32784 28322 32796
rect 30852 32768 30880 32796
rect 23474 32756 23480 32768
rect 22572 32728 23480 32756
rect 23474 32716 23480 32728
rect 23532 32716 23538 32768
rect 24670 32716 24676 32768
rect 24728 32716 24734 32768
rect 26234 32716 26240 32768
rect 26292 32716 26298 32768
rect 26326 32716 26332 32768
rect 26384 32716 26390 32768
rect 26878 32716 26884 32768
rect 26936 32756 26942 32768
rect 29270 32756 29276 32768
rect 26936 32728 29276 32756
rect 26936 32716 26942 32728
rect 29270 32716 29276 32728
rect 29328 32716 29334 32768
rect 30834 32716 30840 32768
rect 30892 32716 30898 32768
rect 33888 32756 33916 32855
rect 33980 32824 34008 32855
rect 34146 32852 34152 32904
rect 34204 32892 34210 32904
rect 34701 32895 34759 32901
rect 34701 32892 34713 32895
rect 34204 32864 34713 32892
rect 34204 32852 34210 32864
rect 34701 32861 34713 32864
rect 34747 32861 34759 32895
rect 34701 32855 34759 32861
rect 34790 32852 34796 32904
rect 34848 32892 34854 32904
rect 36372 32901 36400 32988
rect 36464 32960 36492 33059
rect 37366 33056 37372 33108
rect 37424 33096 37430 33108
rect 37737 33099 37795 33105
rect 37737 33096 37749 33099
rect 37424 33068 37749 33096
rect 37424 33056 37430 33068
rect 37737 33065 37749 33068
rect 37783 33065 37795 33099
rect 37737 33059 37795 33065
rect 38010 33056 38016 33108
rect 38068 33096 38074 33108
rect 38289 33099 38347 33105
rect 38289 33096 38301 33099
rect 38068 33068 38301 33096
rect 38068 33056 38074 33068
rect 38289 33065 38301 33068
rect 38335 33065 38347 33099
rect 38289 33059 38347 33065
rect 38378 33056 38384 33108
rect 38436 33096 38442 33108
rect 38841 33099 38899 33105
rect 38841 33096 38853 33099
rect 38436 33068 38853 33096
rect 38436 33056 38442 33068
rect 38841 33065 38853 33068
rect 38887 33065 38899 33099
rect 38841 33059 38899 33065
rect 41046 33056 41052 33108
rect 41104 33056 41110 33108
rect 37090 32960 37096 32972
rect 36464 32932 37096 32960
rect 37090 32920 37096 32932
rect 37148 32920 37154 32972
rect 37274 32960 37280 32972
rect 37200 32932 37280 32960
rect 34885 32895 34943 32901
rect 34885 32892 34897 32895
rect 34848 32864 34897 32892
rect 34848 32852 34854 32864
rect 34885 32861 34897 32864
rect 34931 32861 34943 32895
rect 34885 32855 34943 32861
rect 36357 32895 36415 32901
rect 36357 32861 36369 32895
rect 36403 32861 36415 32895
rect 36357 32855 36415 32861
rect 36725 32895 36783 32901
rect 36725 32861 36737 32895
rect 36771 32861 36783 32895
rect 36725 32855 36783 32861
rect 36817 32895 36875 32901
rect 36817 32861 36829 32895
rect 36863 32892 36875 32895
rect 37200 32892 37228 32932
rect 37274 32920 37280 32932
rect 37332 32920 37338 32972
rect 37844 32932 38056 32960
rect 36863 32864 37228 32892
rect 37578 32895 37636 32901
rect 36863 32861 36875 32864
rect 36817 32855 36875 32861
rect 37578 32861 37590 32895
rect 37624 32892 37636 32895
rect 37844 32892 37872 32932
rect 38028 32901 38056 32932
rect 38470 32920 38476 32972
rect 38528 32960 38534 32972
rect 39393 32963 39451 32969
rect 39393 32960 39405 32963
rect 38528 32932 39405 32960
rect 38528 32920 38534 32932
rect 39393 32929 39405 32932
rect 39439 32929 39451 32963
rect 39393 32923 39451 32929
rect 37624 32864 37872 32892
rect 37921 32895 37979 32901
rect 37624 32861 37636 32864
rect 37578 32855 37636 32861
rect 37921 32861 37933 32895
rect 37967 32861 37979 32895
rect 37921 32855 37979 32861
rect 38013 32895 38071 32901
rect 38013 32861 38025 32895
rect 38059 32861 38071 32895
rect 38013 32855 38071 32861
rect 34808 32824 34836 32852
rect 33980 32796 34836 32824
rect 36740 32824 36768 32855
rect 37369 32827 37427 32833
rect 37369 32824 37381 32827
rect 36740 32796 37381 32824
rect 37369 32793 37381 32796
rect 37415 32824 37427 32827
rect 37826 32824 37832 32836
rect 37415 32796 37832 32824
rect 37415 32793 37427 32796
rect 37369 32787 37427 32793
rect 37568 32768 37596 32796
rect 37826 32784 37832 32796
rect 37884 32824 37890 32836
rect 37936 32824 37964 32855
rect 37884 32796 37964 32824
rect 38028 32824 38056 32855
rect 38102 32852 38108 32904
rect 38160 32892 38166 32904
rect 38381 32895 38439 32901
rect 38381 32892 38393 32895
rect 38160 32864 38393 32892
rect 38160 32852 38166 32864
rect 38381 32861 38393 32864
rect 38427 32861 38439 32895
rect 38381 32855 38439 32861
rect 38654 32852 38660 32904
rect 38712 32892 38718 32904
rect 39209 32895 39267 32901
rect 39209 32892 39221 32895
rect 38712 32864 39221 32892
rect 38712 32852 38718 32864
rect 39209 32861 39221 32864
rect 39255 32861 39267 32895
rect 39209 32855 39267 32861
rect 39850 32852 39856 32904
rect 39908 32852 39914 32904
rect 40494 32852 40500 32904
rect 40552 32852 40558 32904
rect 38749 32827 38807 32833
rect 38749 32824 38761 32827
rect 38028 32796 38761 32824
rect 37884 32784 37890 32796
rect 34054 32756 34060 32768
rect 33888 32728 34060 32756
rect 34054 32716 34060 32728
rect 34112 32716 34118 32768
rect 35069 32759 35127 32765
rect 35069 32725 35081 32759
rect 35115 32756 35127 32759
rect 35342 32756 35348 32768
rect 35115 32728 35348 32756
rect 35115 32725 35127 32728
rect 35069 32719 35127 32725
rect 35342 32716 35348 32728
rect 35400 32716 35406 32768
rect 36998 32716 37004 32768
rect 37056 32716 37062 32768
rect 37274 32716 37280 32768
rect 37332 32756 37338 32768
rect 37461 32759 37519 32765
rect 37461 32756 37473 32759
rect 37332 32728 37473 32756
rect 37332 32716 37338 32728
rect 37461 32725 37473 32728
rect 37507 32725 37519 32759
rect 37461 32719 37519 32725
rect 37550 32716 37556 32768
rect 37608 32716 37614 32768
rect 37642 32716 37648 32768
rect 37700 32756 37706 32768
rect 38028 32756 38056 32796
rect 38749 32793 38761 32796
rect 38795 32793 38807 32827
rect 38749 32787 38807 32793
rect 37700 32728 38056 32756
rect 37700 32716 37706 32728
rect 38562 32716 38568 32768
rect 38620 32716 38626 32768
rect 39574 32716 39580 32768
rect 39632 32756 39638 32768
rect 39945 32759 40003 32765
rect 39945 32756 39957 32759
rect 39632 32728 39957 32756
rect 39632 32716 39638 32728
rect 39945 32725 39957 32728
rect 39991 32725 40003 32759
rect 39945 32719 40003 32725
rect 1104 32666 41400 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 41400 32666
rect 1104 32592 41400 32614
rect 5718 32512 5724 32564
rect 5776 32552 5782 32564
rect 6822 32552 6828 32564
rect 5776 32524 6828 32552
rect 5776 32512 5782 32524
rect 6822 32512 6828 32524
rect 6880 32512 6886 32564
rect 6914 32512 6920 32564
rect 6972 32552 6978 32564
rect 7282 32552 7288 32564
rect 6972 32524 7288 32552
rect 6972 32512 6978 32524
rect 7282 32512 7288 32524
rect 7340 32512 7346 32564
rect 7650 32512 7656 32564
rect 7708 32552 7714 32564
rect 7929 32555 7987 32561
rect 7929 32552 7941 32555
rect 7708 32524 7941 32552
rect 7708 32512 7714 32524
rect 7929 32521 7941 32524
rect 7975 32521 7987 32555
rect 7929 32515 7987 32521
rect 8018 32512 8024 32564
rect 8076 32552 8082 32564
rect 9766 32552 9772 32564
rect 8076 32524 9168 32552
rect 8076 32512 8082 32524
rect 4982 32444 4988 32496
rect 5040 32444 5046 32496
rect 5077 32487 5135 32493
rect 5077 32453 5089 32487
rect 5123 32484 5135 32487
rect 6086 32484 6092 32496
rect 5123 32456 6092 32484
rect 5123 32453 5135 32456
rect 5077 32447 5135 32453
rect 6086 32444 6092 32456
rect 6144 32444 6150 32496
rect 8294 32484 8300 32496
rect 7208 32456 8300 32484
rect 4801 32419 4859 32425
rect 4801 32385 4813 32419
rect 4847 32416 4859 32419
rect 5000 32416 5028 32444
rect 4847 32388 5028 32416
rect 4847 32385 4859 32388
rect 4801 32379 4859 32385
rect 5994 32376 6000 32428
rect 6052 32376 6058 32428
rect 6178 32376 6184 32428
rect 6236 32376 6242 32428
rect 7208 32425 7236 32456
rect 8294 32444 8300 32456
rect 8352 32444 8358 32496
rect 9140 32425 9168 32524
rect 9232 32524 9772 32552
rect 6549 32419 6607 32425
rect 6549 32385 6561 32419
rect 6595 32416 6607 32419
rect 7193 32419 7251 32425
rect 7193 32416 7205 32419
rect 6595 32388 7205 32416
rect 6595 32385 6607 32388
rect 6549 32379 6607 32385
rect 7193 32385 7205 32388
rect 7239 32385 7251 32419
rect 9033 32419 9091 32425
rect 9033 32416 9045 32419
rect 7193 32379 7251 32385
rect 7484 32388 9045 32416
rect 5074 32308 5080 32360
rect 5132 32308 5138 32360
rect 6270 32308 6276 32360
rect 6328 32348 6334 32360
rect 6457 32351 6515 32357
rect 6457 32348 6469 32351
rect 6328 32320 6469 32348
rect 6328 32308 6334 32320
rect 6457 32317 6469 32320
rect 6503 32317 6515 32351
rect 6457 32311 6515 32317
rect 7484 32280 7512 32388
rect 9033 32385 9045 32388
rect 9079 32385 9091 32419
rect 9033 32379 9091 32385
rect 9126 32419 9184 32425
rect 9126 32385 9138 32419
rect 9172 32385 9184 32419
rect 9126 32379 9184 32385
rect 8294 32308 8300 32360
rect 8352 32308 8358 32360
rect 8389 32351 8447 32357
rect 8389 32317 8401 32351
rect 8435 32348 8447 32351
rect 9232 32348 9260 32524
rect 9766 32512 9772 32524
rect 9824 32512 9830 32564
rect 10321 32555 10379 32561
rect 10321 32521 10333 32555
rect 10367 32521 10379 32555
rect 10321 32515 10379 32521
rect 9309 32487 9367 32493
rect 9309 32453 9321 32487
rect 9355 32484 9367 32487
rect 10336 32484 10364 32515
rect 11330 32512 11336 32564
rect 11388 32512 11394 32564
rect 11977 32555 12035 32561
rect 11977 32521 11989 32555
rect 12023 32552 12035 32555
rect 12066 32552 12072 32564
rect 12023 32524 12072 32552
rect 12023 32521 12035 32524
rect 11977 32515 12035 32521
rect 12066 32512 12072 32524
rect 12124 32512 12130 32564
rect 13541 32555 13599 32561
rect 13541 32552 13553 32555
rect 12406 32524 13553 32552
rect 9355 32456 10364 32484
rect 11348 32484 11376 32512
rect 12406 32484 12434 32524
rect 13541 32521 13553 32524
rect 13587 32521 13599 32555
rect 13541 32515 13599 32521
rect 13817 32555 13875 32561
rect 13817 32521 13829 32555
rect 13863 32552 13875 32555
rect 13906 32552 13912 32564
rect 13863 32524 13912 32552
rect 13863 32521 13875 32524
rect 13817 32515 13875 32521
rect 13906 32512 13912 32524
rect 13964 32512 13970 32564
rect 14550 32512 14556 32564
rect 14608 32552 14614 32564
rect 14737 32555 14795 32561
rect 14608 32524 14694 32552
rect 14608 32512 14614 32524
rect 14666 32484 14694 32524
rect 14737 32521 14749 32555
rect 14783 32552 14795 32555
rect 14826 32552 14832 32564
rect 14783 32524 14832 32552
rect 14783 32521 14795 32524
rect 14737 32515 14795 32521
rect 14826 32512 14832 32524
rect 14884 32512 14890 32564
rect 16022 32512 16028 32564
rect 16080 32512 16086 32564
rect 17954 32512 17960 32564
rect 18012 32552 18018 32564
rect 18141 32555 18199 32561
rect 18141 32552 18153 32555
rect 18012 32524 18153 32552
rect 18012 32512 18018 32524
rect 18141 32521 18153 32524
rect 18187 32521 18199 32555
rect 18141 32515 18199 32521
rect 22738 32512 22744 32564
rect 22796 32552 22802 32564
rect 24673 32555 24731 32561
rect 24673 32552 24685 32555
rect 22796 32524 24685 32552
rect 22796 32512 22802 32524
rect 24673 32521 24685 32524
rect 24719 32521 24731 32555
rect 24673 32515 24731 32521
rect 24762 32512 24768 32564
rect 24820 32552 24826 32564
rect 26973 32555 27031 32561
rect 26973 32552 26985 32555
rect 24820 32524 26985 32552
rect 24820 32512 24826 32524
rect 26973 32521 26985 32524
rect 27019 32521 27031 32555
rect 26973 32515 27031 32521
rect 27062 32512 27068 32564
rect 27120 32552 27126 32564
rect 30745 32555 30803 32561
rect 30745 32552 30757 32555
rect 27120 32524 30757 32552
rect 27120 32512 27126 32524
rect 30745 32521 30757 32524
rect 30791 32521 30803 32555
rect 30745 32515 30803 32521
rect 31202 32512 31208 32564
rect 31260 32552 31266 32564
rect 31260 32524 32536 32552
rect 31260 32512 31266 32524
rect 15562 32484 15568 32496
rect 11348 32456 12434 32484
rect 13464 32456 14596 32484
rect 14666 32456 15568 32484
rect 9355 32453 9367 32456
rect 9309 32447 9367 32453
rect 9398 32376 9404 32428
rect 9456 32376 9462 32428
rect 9498 32419 9556 32425
rect 9498 32385 9510 32419
rect 9544 32385 9556 32419
rect 9498 32379 9556 32385
rect 9953 32419 10011 32425
rect 9953 32385 9965 32419
rect 9999 32416 10011 32419
rect 10594 32416 10600 32428
rect 9999 32388 10600 32416
rect 9999 32385 10011 32388
rect 9953 32379 10011 32385
rect 9508 32348 9536 32379
rect 10594 32376 10600 32388
rect 10652 32376 10658 32428
rect 11793 32419 11851 32425
rect 11793 32385 11805 32419
rect 11839 32385 11851 32419
rect 11793 32379 11851 32385
rect 8435 32320 9260 32348
rect 9324 32320 9536 32348
rect 8435 32317 8447 32320
rect 8389 32311 8447 32317
rect 8404 32280 8432 32311
rect 9324 32280 9352 32320
rect 9858 32308 9864 32360
rect 9916 32308 9922 32360
rect 11808 32348 11836 32379
rect 11882 32376 11888 32428
rect 11940 32416 11946 32428
rect 13464 32425 13492 32456
rect 11977 32419 12035 32425
rect 11977 32416 11989 32419
rect 11940 32388 11989 32416
rect 11940 32376 11946 32388
rect 11977 32385 11989 32388
rect 12023 32385 12035 32419
rect 11977 32379 12035 32385
rect 13449 32419 13507 32425
rect 13449 32385 13461 32419
rect 13495 32385 13507 32419
rect 13449 32379 13507 32385
rect 13633 32419 13691 32425
rect 13633 32385 13645 32419
rect 13679 32385 13691 32419
rect 13633 32379 13691 32385
rect 12342 32348 12348 32360
rect 11808 32320 12348 32348
rect 12342 32308 12348 32320
rect 12400 32308 12406 32360
rect 13648 32348 13676 32379
rect 13998 32376 14004 32428
rect 14056 32376 14062 32428
rect 14568 32425 14596 32456
rect 15562 32444 15568 32456
rect 15620 32444 15626 32496
rect 18046 32444 18052 32496
rect 18104 32484 18110 32496
rect 21818 32484 21824 32496
rect 18104 32456 21824 32484
rect 18104 32444 18110 32456
rect 21818 32444 21824 32456
rect 21876 32444 21882 32496
rect 22278 32444 22284 32496
rect 22336 32444 22342 32496
rect 22462 32444 22468 32496
rect 22520 32484 22526 32496
rect 22649 32487 22707 32493
rect 22649 32484 22661 32487
rect 22520 32456 22661 32484
rect 22520 32444 22526 32456
rect 22649 32453 22661 32456
rect 22695 32484 22707 32487
rect 22830 32484 22836 32496
rect 22695 32456 22836 32484
rect 22695 32453 22707 32456
rect 22649 32447 22707 32453
rect 22830 32444 22836 32456
rect 22888 32444 22894 32496
rect 24210 32444 24216 32496
rect 24268 32444 24274 32496
rect 24854 32484 24860 32496
rect 24504 32456 24860 32484
rect 14553 32419 14611 32425
rect 14553 32385 14565 32419
rect 14599 32416 14611 32419
rect 15841 32419 15899 32425
rect 14599 32388 15240 32416
rect 14599 32385 14611 32388
rect 14553 32379 14611 32385
rect 14274 32348 14280 32360
rect 12544 32320 14280 32348
rect 12544 32292 12572 32320
rect 14274 32308 14280 32320
rect 14332 32348 14338 32360
rect 14369 32351 14427 32357
rect 14369 32348 14381 32351
rect 14332 32320 14381 32348
rect 14332 32308 14338 32320
rect 14369 32317 14381 32320
rect 14415 32317 14427 32351
rect 14369 32311 14427 32317
rect 5920 32252 7512 32280
rect 7668 32252 8432 32280
rect 8496 32252 9352 32280
rect 5920 32224 5948 32252
rect 4890 32172 4896 32224
rect 4948 32172 4954 32224
rect 5902 32172 5908 32224
rect 5960 32172 5966 32224
rect 5997 32215 6055 32221
rect 5997 32181 6009 32215
rect 6043 32212 6055 32215
rect 6638 32212 6644 32224
rect 6043 32184 6644 32212
rect 6043 32181 6055 32184
rect 5997 32175 6055 32181
rect 6638 32172 6644 32184
rect 6696 32172 6702 32224
rect 6822 32172 6828 32224
rect 6880 32212 6886 32224
rect 7668 32212 7696 32252
rect 6880 32184 7696 32212
rect 6880 32172 6886 32184
rect 7742 32172 7748 32224
rect 7800 32172 7806 32224
rect 8202 32172 8208 32224
rect 8260 32212 8266 32224
rect 8496 32212 8524 32252
rect 12526 32240 12532 32292
rect 12584 32240 12590 32292
rect 15212 32224 15240 32388
rect 15841 32385 15853 32419
rect 15887 32385 15899 32419
rect 15841 32379 15899 32385
rect 16025 32419 16083 32425
rect 16025 32385 16037 32419
rect 16071 32416 16083 32419
rect 16071 32388 16344 32416
rect 16071 32385 16083 32388
rect 16025 32379 16083 32385
rect 15856 32348 15884 32379
rect 16206 32348 16212 32360
rect 15856 32320 16212 32348
rect 16206 32308 16212 32320
rect 16264 32308 16270 32360
rect 16316 32292 16344 32388
rect 21174 32376 21180 32428
rect 21232 32416 21238 32428
rect 21634 32416 21640 32428
rect 21232 32388 21640 32416
rect 21232 32376 21238 32388
rect 21634 32376 21640 32388
rect 21692 32416 21698 32428
rect 22005 32419 22063 32425
rect 22005 32416 22017 32419
rect 21692 32388 22017 32416
rect 21692 32376 21698 32388
rect 22005 32385 22017 32388
rect 22051 32385 22063 32419
rect 22296 32416 22324 32444
rect 24504 32425 24532 32456
rect 24854 32444 24860 32456
rect 24912 32484 24918 32496
rect 24912 32456 27660 32484
rect 24912 32444 24918 32456
rect 27632 32428 27660 32456
rect 28258 32444 28264 32496
rect 28316 32484 28322 32496
rect 28353 32487 28411 32493
rect 28353 32484 28365 32487
rect 28316 32456 28365 32484
rect 28316 32444 28322 32456
rect 28353 32453 28365 32456
rect 28399 32453 28411 32487
rect 28353 32447 28411 32453
rect 28445 32487 28503 32493
rect 28445 32453 28457 32487
rect 28491 32484 28503 32487
rect 28626 32484 28632 32496
rect 28491 32456 28632 32484
rect 28491 32453 28503 32456
rect 28445 32447 28503 32453
rect 28626 32444 28632 32456
rect 28684 32484 28690 32496
rect 30101 32487 30159 32493
rect 30101 32484 30113 32487
rect 28684 32456 30113 32484
rect 28684 32444 28690 32456
rect 30101 32453 30113 32456
rect 30147 32484 30159 32487
rect 30650 32484 30656 32496
rect 30147 32456 30656 32484
rect 30147 32453 30159 32456
rect 30101 32447 30159 32453
rect 30650 32444 30656 32456
rect 30708 32484 30714 32496
rect 30708 32456 31064 32484
rect 30708 32444 30714 32456
rect 22373 32419 22431 32425
rect 22373 32416 22385 32419
rect 22005 32379 22063 32385
rect 22112 32388 22385 32416
rect 19150 32308 19156 32360
rect 19208 32348 19214 32360
rect 22112 32348 22140 32388
rect 22373 32385 22385 32388
rect 22419 32385 22431 32419
rect 22373 32379 22431 32385
rect 24489 32419 24547 32425
rect 24489 32385 24501 32419
rect 24535 32385 24547 32419
rect 24489 32379 24547 32385
rect 25406 32376 25412 32428
rect 25464 32416 25470 32428
rect 26513 32419 26571 32425
rect 26513 32416 26525 32419
rect 25464 32388 26525 32416
rect 25464 32376 25470 32388
rect 26513 32385 26525 32388
rect 26559 32385 26571 32419
rect 26513 32379 26571 32385
rect 19208 32320 22140 32348
rect 22281 32351 22339 32357
rect 19208 32308 19214 32320
rect 22281 32317 22293 32351
rect 22327 32348 22339 32351
rect 22646 32348 22652 32360
rect 22327 32320 22652 32348
rect 22327 32317 22339 32320
rect 22281 32311 22339 32317
rect 16298 32240 16304 32292
rect 16356 32240 16362 32292
rect 21358 32240 21364 32292
rect 21416 32280 21422 32292
rect 22296 32280 22324 32311
rect 22646 32308 22652 32320
rect 22704 32308 22710 32360
rect 24394 32308 24400 32360
rect 24452 32308 24458 32360
rect 26528 32348 26556 32379
rect 26694 32376 26700 32428
rect 26752 32376 26758 32428
rect 26789 32419 26847 32425
rect 26789 32385 26801 32419
rect 26835 32416 26847 32419
rect 26835 32388 27476 32416
rect 26835 32385 26847 32388
rect 26789 32379 26847 32385
rect 26602 32348 26608 32360
rect 26528 32320 26608 32348
rect 26602 32308 26608 32320
rect 26660 32348 26666 32360
rect 27249 32351 27307 32357
rect 27249 32348 27261 32351
rect 26660 32320 27261 32348
rect 26660 32308 26666 32320
rect 27249 32317 27261 32320
rect 27295 32317 27307 32351
rect 27448 32348 27476 32388
rect 27522 32376 27528 32428
rect 27580 32376 27586 32428
rect 27614 32376 27620 32428
rect 27672 32376 27678 32428
rect 27709 32419 27767 32425
rect 27709 32385 27721 32419
rect 27755 32385 27767 32419
rect 27709 32379 27767 32385
rect 28169 32419 28227 32425
rect 28169 32385 28181 32419
rect 28215 32385 28227 32419
rect 28169 32379 28227 32385
rect 28537 32419 28595 32425
rect 28537 32385 28549 32419
rect 28583 32416 28595 32419
rect 28810 32416 28816 32428
rect 28583 32388 28816 32416
rect 28583 32385 28595 32388
rect 28537 32379 28595 32385
rect 27724 32348 27752 32379
rect 27982 32348 27988 32360
rect 27448 32320 27988 32348
rect 27249 32311 27307 32317
rect 27982 32308 27988 32320
rect 28040 32308 28046 32360
rect 28184 32348 28212 32379
rect 28810 32376 28816 32388
rect 28868 32376 28874 32428
rect 28994 32416 29000 32428
rect 29052 32425 29058 32428
rect 29052 32419 29075 32425
rect 28966 32376 29000 32416
rect 29063 32416 29075 32419
rect 29181 32419 29239 32425
rect 29063 32388 29145 32416
rect 29063 32385 29075 32388
rect 29052 32379 29075 32385
rect 29181 32385 29193 32419
rect 29227 32385 29239 32419
rect 29181 32379 29239 32385
rect 29052 32376 29058 32379
rect 28966 32348 28994 32376
rect 28184 32320 28994 32348
rect 29196 32348 29224 32379
rect 29270 32376 29276 32428
rect 29328 32376 29334 32428
rect 29365 32419 29423 32425
rect 29365 32385 29377 32419
rect 29411 32416 29423 32419
rect 29454 32416 29460 32428
rect 29411 32388 29460 32416
rect 29411 32385 29423 32388
rect 29365 32379 29423 32385
rect 29454 32376 29460 32388
rect 29512 32376 29518 32428
rect 29638 32376 29644 32428
rect 29696 32416 29702 32428
rect 29733 32419 29791 32425
rect 29733 32416 29745 32419
rect 29696 32388 29745 32416
rect 29696 32376 29702 32388
rect 29733 32385 29745 32388
rect 29779 32385 29791 32419
rect 29733 32379 29791 32385
rect 30282 32376 30288 32428
rect 30340 32376 30346 32428
rect 30374 32376 30380 32428
rect 30432 32376 30438 32428
rect 31036 32425 31064 32456
rect 31726 32456 32444 32484
rect 31021 32419 31079 32425
rect 31021 32385 31033 32419
rect 31067 32385 31079 32419
rect 31481 32419 31539 32425
rect 31481 32416 31493 32419
rect 31021 32379 31079 32385
rect 31128 32388 31493 32416
rect 29914 32348 29920 32360
rect 29196 32320 29920 32348
rect 29914 32308 29920 32320
rect 29972 32348 29978 32360
rect 30300 32348 30328 32376
rect 30561 32351 30619 32357
rect 30561 32348 30573 32351
rect 29972 32320 30573 32348
rect 29972 32308 29978 32320
rect 30561 32317 30573 32320
rect 30607 32317 30619 32351
rect 30561 32311 30619 32317
rect 30653 32351 30711 32357
rect 30653 32317 30665 32351
rect 30699 32348 30711 32351
rect 31128 32348 31156 32388
rect 31481 32385 31493 32388
rect 31527 32416 31539 32419
rect 31726 32416 31754 32456
rect 32416 32425 32444 32456
rect 32508 32450 32536 32524
rect 32582 32512 32588 32564
rect 32640 32512 32646 32564
rect 32858 32512 32864 32564
rect 32916 32512 32922 32564
rect 33870 32512 33876 32564
rect 33928 32552 33934 32564
rect 34790 32552 34796 32564
rect 33928 32524 34796 32552
rect 33928 32512 33934 32524
rect 34790 32512 34796 32524
rect 34848 32512 34854 32564
rect 35986 32512 35992 32564
rect 36044 32552 36050 32564
rect 36173 32555 36231 32561
rect 36173 32552 36185 32555
rect 36044 32524 36185 32552
rect 36044 32512 36050 32524
rect 36173 32521 36185 32524
rect 36219 32521 36231 32555
rect 36173 32515 36231 32521
rect 37090 32512 37096 32564
rect 37148 32552 37154 32564
rect 38010 32552 38016 32564
rect 37148 32524 38016 32552
rect 37148 32512 37154 32524
rect 38010 32512 38016 32524
rect 38068 32512 38074 32564
rect 38289 32555 38347 32561
rect 38289 32521 38301 32555
rect 38335 32552 38347 32555
rect 38654 32552 38660 32564
rect 38335 32524 38660 32552
rect 38335 32521 38347 32524
rect 38289 32515 38347 32521
rect 38654 32512 38660 32524
rect 38712 32512 38718 32564
rect 40494 32512 40500 32564
rect 40552 32552 40558 32564
rect 40589 32555 40647 32561
rect 40589 32552 40601 32555
rect 40552 32524 40601 32552
rect 40552 32512 40558 32524
rect 40589 32521 40601 32524
rect 40635 32521 40647 32555
rect 40589 32515 40647 32521
rect 40954 32512 40960 32564
rect 41012 32512 41018 32564
rect 32600 32456 34376 32484
rect 32600 32450 32628 32456
rect 31527 32388 31754 32416
rect 32125 32419 32183 32425
rect 31527 32385 31539 32388
rect 31481 32379 31539 32385
rect 32125 32385 32137 32419
rect 32171 32416 32183 32419
rect 32401 32419 32459 32425
rect 32508 32422 32628 32450
rect 32171 32388 32352 32416
rect 32171 32385 32183 32388
rect 32125 32379 32183 32385
rect 30699 32320 31156 32348
rect 31205 32351 31263 32357
rect 30699 32317 30711 32320
rect 30653 32311 30711 32317
rect 31205 32317 31217 32351
rect 31251 32348 31263 32351
rect 32214 32348 32220 32360
rect 31251 32320 32220 32348
rect 31251 32317 31263 32320
rect 31205 32311 31263 32317
rect 32214 32308 32220 32320
rect 32272 32308 32278 32360
rect 21416 32252 22324 32280
rect 21416 32240 21422 32252
rect 23750 32240 23756 32292
rect 23808 32280 23814 32292
rect 24210 32280 24216 32292
rect 23808 32252 24216 32280
rect 23808 32240 23814 32252
rect 24210 32240 24216 32252
rect 24268 32240 24274 32292
rect 24762 32240 24768 32292
rect 24820 32280 24826 32292
rect 24820 32252 25452 32280
rect 24820 32240 24826 32252
rect 8260 32184 8524 32212
rect 8260 32172 8266 32184
rect 8570 32172 8576 32224
rect 8628 32172 8634 32224
rect 9674 32172 9680 32224
rect 9732 32172 9738 32224
rect 12434 32172 12440 32224
rect 12492 32212 12498 32224
rect 14182 32212 14188 32224
rect 12492 32184 14188 32212
rect 12492 32172 12498 32184
rect 14182 32172 14188 32184
rect 14240 32172 14246 32224
rect 15194 32172 15200 32224
rect 15252 32172 15258 32224
rect 15930 32172 15936 32224
rect 15988 32212 15994 32224
rect 16482 32212 16488 32224
rect 15988 32184 16488 32212
rect 15988 32172 15994 32184
rect 16482 32172 16488 32184
rect 16540 32172 16546 32224
rect 21450 32172 21456 32224
rect 21508 32212 21514 32224
rect 21821 32215 21879 32221
rect 21821 32212 21833 32215
rect 21508 32184 21833 32212
rect 21508 32172 21514 32184
rect 21821 32181 21833 32184
rect 21867 32181 21879 32215
rect 21821 32175 21879 32181
rect 22189 32215 22247 32221
rect 22189 32181 22201 32215
rect 22235 32212 22247 32215
rect 24302 32212 24308 32224
rect 22235 32184 24308 32212
rect 22235 32181 22247 32184
rect 22189 32175 22247 32181
rect 24302 32172 24308 32184
rect 24360 32172 24366 32224
rect 24489 32215 24547 32221
rect 24489 32181 24501 32215
rect 24535 32212 24547 32215
rect 24670 32212 24676 32224
rect 24535 32184 24676 32212
rect 24535 32181 24547 32184
rect 24489 32175 24547 32181
rect 24670 32172 24676 32184
rect 24728 32212 24734 32224
rect 25314 32212 25320 32224
rect 24728 32184 25320 32212
rect 24728 32172 24734 32184
rect 25314 32172 25320 32184
rect 25372 32172 25378 32224
rect 25424 32212 25452 32252
rect 26326 32240 26332 32292
rect 26384 32280 26390 32292
rect 27433 32283 27491 32289
rect 26384 32252 27200 32280
rect 26384 32240 26390 32252
rect 27172 32224 27200 32252
rect 27433 32249 27445 32283
rect 27479 32280 27491 32283
rect 27890 32280 27896 32292
rect 27479 32252 27896 32280
rect 27479 32249 27491 32252
rect 27433 32243 27491 32249
rect 27890 32240 27896 32252
rect 27948 32280 27954 32292
rect 29549 32283 29607 32289
rect 29549 32280 29561 32283
rect 27948 32252 29561 32280
rect 27948 32240 27954 32252
rect 29549 32249 29561 32252
rect 29595 32249 29607 32283
rect 32324 32280 32352 32388
rect 32401 32385 32413 32419
rect 32447 32385 32459 32419
rect 32401 32379 32459 32385
rect 29549 32243 29607 32249
rect 31128 32252 32352 32280
rect 32416 32280 32444 32379
rect 32674 32376 32680 32428
rect 32732 32376 32738 32428
rect 32953 32419 33011 32425
rect 32953 32385 32965 32419
rect 32999 32416 33011 32419
rect 33042 32416 33048 32428
rect 32999 32388 33048 32416
rect 32999 32385 33011 32388
rect 32953 32379 33011 32385
rect 33042 32376 33048 32388
rect 33100 32376 33106 32428
rect 32692 32348 32720 32376
rect 34238 32348 34244 32360
rect 32692 32320 34244 32348
rect 34238 32308 34244 32320
rect 34296 32308 34302 32360
rect 34348 32348 34376 32456
rect 34422 32444 34428 32496
rect 34480 32484 34486 32496
rect 37826 32484 37832 32496
rect 34480 32456 37832 32484
rect 34480 32444 34486 32456
rect 36262 32376 36268 32428
rect 36320 32416 36326 32428
rect 36357 32419 36415 32425
rect 36357 32416 36369 32419
rect 36320 32388 36369 32416
rect 36320 32376 36326 32388
rect 36357 32385 36369 32388
rect 36403 32416 36415 32419
rect 36446 32416 36452 32428
rect 36403 32388 36452 32416
rect 36403 32385 36415 32388
rect 36357 32379 36415 32385
rect 36446 32376 36452 32388
rect 36504 32376 36510 32428
rect 36648 32425 36676 32456
rect 37826 32444 37832 32456
rect 37884 32484 37890 32496
rect 39206 32484 39212 32496
rect 37884 32456 38516 32484
rect 37884 32444 37890 32456
rect 38488 32428 38516 32456
rect 38856 32456 39212 32484
rect 36633 32419 36691 32425
rect 36633 32385 36645 32419
rect 36679 32385 36691 32419
rect 37458 32416 37464 32428
rect 36633 32379 36691 32385
rect 37200 32388 37464 32416
rect 37200 32348 37228 32388
rect 37458 32376 37464 32388
rect 37516 32376 37522 32428
rect 37737 32419 37795 32425
rect 37737 32385 37749 32419
rect 37783 32385 37795 32419
rect 37737 32379 37795 32385
rect 34348 32320 37228 32348
rect 37274 32308 37280 32360
rect 37332 32348 37338 32360
rect 37645 32351 37703 32357
rect 37645 32348 37657 32351
rect 37332 32320 37657 32348
rect 37332 32308 37338 32320
rect 37645 32317 37657 32320
rect 37691 32317 37703 32351
rect 37752 32348 37780 32379
rect 38010 32376 38016 32428
rect 38068 32416 38074 32428
rect 38105 32419 38163 32425
rect 38105 32416 38117 32419
rect 38068 32388 38117 32416
rect 38068 32376 38074 32388
rect 38105 32385 38117 32388
rect 38151 32385 38163 32419
rect 38105 32379 38163 32385
rect 38378 32376 38384 32428
rect 38436 32376 38442 32428
rect 38470 32376 38476 32428
rect 38528 32376 38534 32428
rect 38856 32425 38884 32456
rect 39206 32444 39212 32456
rect 39264 32444 39270 32496
rect 38841 32419 38899 32425
rect 38841 32385 38853 32419
rect 38887 32385 38899 32419
rect 40328 32416 40356 32470
rect 40586 32416 40592 32428
rect 40328 32388 40592 32416
rect 38841 32379 38899 32385
rect 40586 32376 40592 32388
rect 40644 32376 40650 32428
rect 40770 32376 40776 32428
rect 40828 32376 40834 32428
rect 38396 32348 38424 32376
rect 37752 32320 38424 32348
rect 39117 32351 39175 32357
rect 37645 32311 37703 32317
rect 39117 32317 39129 32351
rect 39163 32348 39175 32351
rect 39574 32348 39580 32360
rect 39163 32320 39580 32348
rect 39163 32317 39175 32320
rect 39117 32311 39175 32317
rect 32677 32283 32735 32289
rect 32677 32280 32689 32283
rect 32416 32252 32689 32280
rect 27062 32212 27068 32224
rect 25424 32184 27068 32212
rect 27062 32172 27068 32184
rect 27120 32172 27126 32224
rect 27154 32172 27160 32224
rect 27212 32172 27218 32224
rect 27338 32172 27344 32224
rect 27396 32172 27402 32224
rect 27522 32172 27528 32224
rect 27580 32212 27586 32224
rect 28721 32215 28779 32221
rect 28721 32212 28733 32215
rect 27580 32184 28733 32212
rect 27580 32172 27586 32184
rect 28721 32181 28733 32184
rect 28767 32181 28779 32215
rect 28721 32175 28779 32181
rect 28994 32172 29000 32224
rect 29052 32212 29058 32224
rect 29638 32212 29644 32224
rect 29052 32184 29644 32212
rect 29052 32172 29058 32184
rect 29638 32172 29644 32184
rect 29696 32172 29702 32224
rect 30190 32172 30196 32224
rect 30248 32172 30254 32224
rect 30742 32172 30748 32224
rect 30800 32212 30806 32224
rect 31128 32221 31156 32252
rect 31113 32215 31171 32221
rect 31113 32212 31125 32215
rect 30800 32184 31125 32212
rect 30800 32172 30806 32184
rect 31113 32181 31125 32184
rect 31159 32181 31171 32215
rect 31113 32175 31171 32181
rect 31297 32215 31355 32221
rect 31297 32181 31309 32215
rect 31343 32212 31355 32215
rect 32030 32212 32036 32224
rect 31343 32184 32036 32212
rect 31343 32181 31355 32184
rect 31297 32175 31355 32181
rect 32030 32172 32036 32184
rect 32088 32212 32094 32224
rect 32125 32215 32183 32221
rect 32125 32212 32137 32215
rect 32088 32184 32137 32212
rect 32088 32172 32094 32184
rect 32125 32181 32137 32184
rect 32171 32181 32183 32215
rect 32324 32212 32352 32252
rect 32677 32249 32689 32252
rect 32723 32249 32735 32283
rect 37660 32280 37688 32311
rect 39574 32308 39580 32320
rect 39632 32308 39638 32360
rect 38102 32280 38108 32292
rect 37660 32252 38108 32280
rect 32677 32243 32735 32249
rect 38102 32240 38108 32252
rect 38160 32240 38166 32292
rect 33134 32212 33140 32224
rect 32324 32184 33140 32212
rect 32125 32175 32183 32181
rect 33134 32172 33140 32184
rect 33192 32172 33198 32224
rect 33318 32172 33324 32224
rect 33376 32212 33382 32224
rect 34606 32212 34612 32224
rect 33376 32184 34612 32212
rect 33376 32172 33382 32184
rect 34606 32172 34612 32184
rect 34664 32172 34670 32224
rect 37550 32172 37556 32224
rect 37608 32212 37614 32224
rect 38013 32215 38071 32221
rect 38013 32212 38025 32215
rect 37608 32184 38025 32212
rect 37608 32172 37614 32184
rect 38013 32181 38025 32184
rect 38059 32181 38071 32215
rect 38013 32175 38071 32181
rect 1104 32122 41400 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 41400 32122
rect 1104 32048 41400 32070
rect 4798 31968 4804 32020
rect 4856 31968 4862 32020
rect 4890 31968 4896 32020
rect 4948 31968 4954 32020
rect 5169 32011 5227 32017
rect 5169 31977 5181 32011
rect 5215 32008 5227 32011
rect 5994 32008 6000 32020
rect 5215 31980 6000 32008
rect 5215 31977 5227 31980
rect 5169 31971 5227 31977
rect 5994 31968 6000 31980
rect 6052 31968 6058 32020
rect 6086 31968 6092 32020
rect 6144 31968 6150 32020
rect 7190 32008 7196 32020
rect 6472 31980 7196 32008
rect 4816 31872 4844 31968
rect 4908 31940 4936 31968
rect 5813 31943 5871 31949
rect 5813 31940 5825 31943
rect 4908 31912 5825 31940
rect 5813 31909 5825 31912
rect 5859 31909 5871 31943
rect 5813 31903 5871 31909
rect 5902 31900 5908 31952
rect 5960 31900 5966 31952
rect 4893 31875 4951 31881
rect 4893 31872 4905 31875
rect 4816 31844 4905 31872
rect 4893 31841 4905 31844
rect 4939 31872 4951 31875
rect 5350 31872 5356 31884
rect 4939 31844 5356 31872
rect 4939 31841 4951 31844
rect 4893 31835 4951 31841
rect 5350 31832 5356 31844
rect 5408 31832 5414 31884
rect 2958 31764 2964 31816
rect 3016 31764 3022 31816
rect 4801 31807 4859 31813
rect 4801 31773 4813 31807
rect 4847 31804 4859 31807
rect 4982 31804 4988 31816
rect 4847 31776 4988 31804
rect 4847 31773 4859 31776
rect 4801 31767 4859 31773
rect 4982 31764 4988 31776
rect 5040 31764 5046 31816
rect 5445 31807 5503 31813
rect 5445 31773 5457 31807
rect 5491 31804 5503 31807
rect 5718 31804 5724 31816
rect 5491 31776 5724 31804
rect 5491 31773 5503 31776
rect 5445 31767 5503 31773
rect 5718 31764 5724 31776
rect 5776 31764 5782 31816
rect 5905 31807 5963 31813
rect 5905 31773 5917 31807
rect 5951 31804 5963 31807
rect 5994 31804 6000 31816
rect 5951 31776 6000 31804
rect 5951 31773 5963 31776
rect 5905 31767 5963 31773
rect 5994 31764 6000 31776
rect 6052 31764 6058 31816
rect 6104 31813 6132 31968
rect 6472 31881 6500 31980
rect 7190 31968 7196 31980
rect 7248 31968 7254 32020
rect 7926 31968 7932 32020
rect 7984 32008 7990 32020
rect 7984 31980 10272 32008
rect 7984 31968 7990 31980
rect 6457 31875 6515 31881
rect 6457 31841 6469 31875
rect 6503 31841 6515 31875
rect 6457 31835 6515 31841
rect 6638 31832 6644 31884
rect 6696 31872 6702 31884
rect 7742 31872 7748 31884
rect 6696 31844 7052 31872
rect 6696 31832 6702 31844
rect 6089 31807 6147 31813
rect 6089 31773 6101 31807
rect 6135 31773 6147 31807
rect 6089 31767 6147 31773
rect 6178 31764 6184 31816
rect 6236 31764 6242 31816
rect 6549 31807 6607 31813
rect 6549 31773 6561 31807
rect 6595 31804 6607 31807
rect 6914 31804 6920 31816
rect 6595 31776 6920 31804
rect 6595 31773 6607 31776
rect 6549 31767 6607 31773
rect 6914 31764 6920 31776
rect 6972 31764 6978 31816
rect 7024 31813 7052 31844
rect 7392 31844 7748 31872
rect 7009 31807 7067 31813
rect 7009 31773 7021 31807
rect 7055 31773 7067 31807
rect 7009 31767 7067 31773
rect 7098 31764 7104 31816
rect 7156 31804 7162 31816
rect 7392 31813 7420 31844
rect 7742 31832 7748 31844
rect 7800 31832 7806 31884
rect 9217 31875 9275 31881
rect 9217 31841 9229 31875
rect 9263 31872 9275 31875
rect 9674 31872 9680 31884
rect 9263 31844 9680 31872
rect 9263 31841 9275 31844
rect 9217 31835 9275 31841
rect 9674 31832 9680 31844
rect 9732 31832 9738 31884
rect 10244 31872 10272 31980
rect 12618 31968 12624 32020
rect 12676 31968 12682 32020
rect 13078 31968 13084 32020
rect 13136 32008 13142 32020
rect 14918 32008 14924 32020
rect 13136 31980 14924 32008
rect 13136 31968 13142 31980
rect 14918 31968 14924 31980
rect 14976 31968 14982 32020
rect 15194 31968 15200 32020
rect 15252 31968 15258 32020
rect 15654 31968 15660 32020
rect 15712 32008 15718 32020
rect 15712 31980 17908 32008
rect 15712 31968 15718 31980
rect 16025 31943 16083 31949
rect 16025 31909 16037 31943
rect 16071 31940 16083 31943
rect 16853 31943 16911 31949
rect 16071 31912 16436 31940
rect 16071 31909 16083 31912
rect 16025 31903 16083 31909
rect 10244 31844 10364 31872
rect 7285 31807 7343 31813
rect 7156 31776 7201 31804
rect 7156 31764 7162 31776
rect 7285 31773 7297 31807
rect 7331 31773 7343 31807
rect 7285 31767 7343 31773
rect 7390 31807 7448 31813
rect 7390 31773 7402 31807
rect 7436 31773 7448 31807
rect 7390 31767 7448 31773
rect 7515 31807 7573 31813
rect 7515 31773 7527 31807
rect 7561 31804 7573 31807
rect 8202 31804 8208 31816
rect 7561 31776 8208 31804
rect 7561 31773 7573 31776
rect 7515 31767 7573 31773
rect 2774 31628 2780 31680
rect 2832 31628 2838 31680
rect 6917 31671 6975 31677
rect 6917 31637 6929 31671
rect 6963 31668 6975 31671
rect 7300 31668 7328 31767
rect 8202 31764 8208 31776
rect 8260 31764 8266 31816
rect 8941 31807 8999 31813
rect 8941 31773 8953 31807
rect 8987 31773 8999 31807
rect 10336 31790 10364 31844
rect 11606 31832 11612 31884
rect 11664 31872 11670 31884
rect 12713 31875 12771 31881
rect 12713 31872 12725 31875
rect 11664 31844 12725 31872
rect 11664 31832 11670 31844
rect 12713 31841 12725 31844
rect 12759 31841 12771 31875
rect 12713 31835 12771 31841
rect 14550 31832 14556 31884
rect 14608 31872 14614 31884
rect 14829 31875 14887 31881
rect 14829 31872 14841 31875
rect 14608 31844 14841 31872
rect 14608 31832 14614 31844
rect 14829 31841 14841 31844
rect 14875 31841 14887 31875
rect 14829 31835 14887 31841
rect 14918 31832 14924 31884
rect 14976 31832 14982 31884
rect 16408 31881 16436 31912
rect 16853 31909 16865 31943
rect 16899 31940 16911 31943
rect 17402 31940 17408 31952
rect 16899 31912 17408 31940
rect 16899 31909 16911 31912
rect 16853 31903 16911 31909
rect 17402 31900 17408 31912
rect 17460 31900 17466 31952
rect 16393 31875 16451 31881
rect 15028 31844 15884 31872
rect 8941 31767 8999 31773
rect 8956 31680 8984 31767
rect 12434 31764 12440 31816
rect 12492 31764 12498 31816
rect 12526 31764 12532 31816
rect 12584 31764 12590 31816
rect 14182 31764 14188 31816
rect 14240 31764 14246 31816
rect 14642 31764 14648 31816
rect 14700 31764 14706 31816
rect 14737 31807 14795 31813
rect 14737 31773 14749 31807
rect 14783 31804 14795 31807
rect 14783 31798 14872 31804
rect 15028 31798 15056 31844
rect 15212 31813 15240 31844
rect 14783 31776 15056 31798
rect 14783 31773 14795 31776
rect 14737 31767 14795 31773
rect 14844 31770 15056 31776
rect 15105 31807 15163 31813
rect 15105 31773 15117 31807
rect 15151 31773 15163 31807
rect 15105 31767 15163 31773
rect 15197 31807 15255 31813
rect 15197 31773 15209 31807
rect 15243 31773 15255 31807
rect 15197 31767 15255 31773
rect 15381 31807 15439 31813
rect 15381 31773 15393 31807
rect 15427 31773 15439 31807
rect 15381 31767 15439 31773
rect 15473 31807 15531 31813
rect 15473 31773 15485 31807
rect 15519 31804 15531 31807
rect 15562 31804 15568 31816
rect 15519 31776 15568 31804
rect 15519 31773 15531 31776
rect 15473 31767 15531 31773
rect 12544 31736 12572 31764
rect 12452 31708 12572 31736
rect 14200 31736 14228 31764
rect 15120 31736 15148 31767
rect 14200 31708 15148 31736
rect 12452 31680 12480 31708
rect 6963 31640 7328 31668
rect 6963 31637 6975 31640
rect 6917 31631 6975 31637
rect 7650 31628 7656 31680
rect 7708 31628 7714 31680
rect 8938 31628 8944 31680
rect 8996 31628 9002 31680
rect 9398 31628 9404 31680
rect 9456 31668 9462 31680
rect 10689 31671 10747 31677
rect 10689 31668 10701 31671
rect 9456 31640 10701 31668
rect 9456 31628 9462 31640
rect 10689 31637 10701 31640
rect 10735 31637 10747 31671
rect 10689 31631 10747 31637
rect 12434 31628 12440 31680
rect 12492 31628 12498 31680
rect 14458 31628 14464 31680
rect 14516 31628 14522 31680
rect 14642 31628 14648 31680
rect 14700 31668 14706 31680
rect 15397 31668 15425 31767
rect 15562 31764 15568 31776
rect 15620 31764 15626 31816
rect 15746 31764 15752 31816
rect 15804 31764 15810 31816
rect 15856 31813 15884 31844
rect 16393 31841 16405 31875
rect 16439 31841 16451 31875
rect 16393 31835 16451 31841
rect 15841 31807 15899 31813
rect 15841 31773 15853 31807
rect 15887 31804 15899 31807
rect 16298 31804 16304 31816
rect 15887 31776 16304 31804
rect 15887 31773 15899 31776
rect 15841 31767 15899 31773
rect 16298 31764 16304 31776
rect 16356 31764 16362 31816
rect 17880 31813 17908 31980
rect 22186 31968 22192 32020
rect 22244 32008 22250 32020
rect 22557 32011 22615 32017
rect 22557 32008 22569 32011
rect 22244 31980 22569 32008
rect 22244 31968 22250 31980
rect 22557 31977 22569 31980
rect 22603 31977 22615 32011
rect 22557 31971 22615 31977
rect 23658 31968 23664 32020
rect 23716 31968 23722 32020
rect 23845 32011 23903 32017
rect 23845 31977 23857 32011
rect 23891 32008 23903 32011
rect 24118 32008 24124 32020
rect 23891 31980 24124 32008
rect 23891 31977 23903 31980
rect 23845 31971 23903 31977
rect 24118 31968 24124 31980
rect 24176 31968 24182 32020
rect 24210 31968 24216 32020
rect 24268 32008 24274 32020
rect 24397 32011 24455 32017
rect 24397 32008 24409 32011
rect 24268 31980 24409 32008
rect 24268 31968 24274 31980
rect 24397 31977 24409 31980
rect 24443 31977 24455 32011
rect 24397 31971 24455 31977
rect 25314 31968 25320 32020
rect 25372 31968 25378 32020
rect 25866 31968 25872 32020
rect 25924 32008 25930 32020
rect 26513 32011 26571 32017
rect 26513 32008 26525 32011
rect 25924 31980 26525 32008
rect 25924 31968 25930 31980
rect 26513 31977 26525 31980
rect 26559 31977 26571 32011
rect 26513 31971 26571 31977
rect 26602 31968 26608 32020
rect 26660 32008 26666 32020
rect 26697 32011 26755 32017
rect 26697 32008 26709 32011
rect 26660 31980 26709 32008
rect 26660 31968 26666 31980
rect 26697 31977 26709 31980
rect 26743 31977 26755 32011
rect 26697 31971 26755 31977
rect 27246 31968 27252 32020
rect 27304 31968 27310 32020
rect 27338 31968 27344 32020
rect 27396 31968 27402 32020
rect 27890 31968 27896 32020
rect 27948 31968 27954 32020
rect 27982 31968 27988 32020
rect 28040 32008 28046 32020
rect 33318 32008 33324 32020
rect 28040 31980 33324 32008
rect 28040 31968 28046 31980
rect 33318 31968 33324 31980
rect 33376 31968 33382 32020
rect 34606 31968 34612 32020
rect 34664 31968 34670 32020
rect 34885 32011 34943 32017
rect 34885 31977 34897 32011
rect 34931 32008 34943 32011
rect 35342 32008 35348 32020
rect 34931 31980 35348 32008
rect 34931 31977 34943 31980
rect 34885 31971 34943 31977
rect 35342 31968 35348 31980
rect 35400 32008 35406 32020
rect 35400 31980 35756 32008
rect 35400 31968 35406 31980
rect 19334 31900 19340 31952
rect 19392 31940 19398 31952
rect 25958 31940 25964 31952
rect 19392 31912 25964 31940
rect 19392 31900 19398 31912
rect 25958 31900 25964 31912
rect 26016 31900 26022 31952
rect 26326 31900 26332 31952
rect 26384 31940 26390 31952
rect 26878 31940 26884 31952
rect 26384 31912 26884 31940
rect 26384 31900 26390 31912
rect 18690 31832 18696 31884
rect 18748 31832 18754 31884
rect 23293 31875 23351 31881
rect 23293 31872 23305 31875
rect 20916 31844 21588 31872
rect 20916 31816 20944 31844
rect 21560 31816 21588 31844
rect 21744 31844 22692 31872
rect 16563 31807 16621 31813
rect 16563 31773 16575 31807
rect 16609 31773 16621 31807
rect 16563 31767 16621 31773
rect 17865 31807 17923 31813
rect 17865 31773 17877 31807
rect 17911 31804 17923 31807
rect 19334 31804 19340 31816
rect 17911 31776 19340 31804
rect 17911 31773 17923 31776
rect 17865 31767 17923 31773
rect 15654 31696 15660 31748
rect 15712 31736 15718 31748
rect 16206 31736 16212 31748
rect 15712 31708 16212 31736
rect 15712 31696 15718 31708
rect 16206 31696 16212 31708
rect 16264 31696 16270 31748
rect 14700 31640 15425 31668
rect 14700 31628 14706 31640
rect 16114 31628 16120 31680
rect 16172 31668 16178 31680
rect 16592 31668 16620 31767
rect 19334 31764 19340 31776
rect 19392 31764 19398 31816
rect 20898 31764 20904 31816
rect 20956 31764 20962 31816
rect 21450 31764 21456 31816
rect 21508 31764 21514 31816
rect 21542 31764 21548 31816
rect 21600 31764 21606 31816
rect 21744 31813 21772 31844
rect 21729 31807 21787 31813
rect 21729 31773 21741 31807
rect 21775 31773 21787 31807
rect 21729 31767 21787 31773
rect 21918 31807 21976 31813
rect 21918 31773 21930 31807
rect 21964 31773 21976 31807
rect 21918 31767 21976 31773
rect 20162 31696 20168 31748
rect 20220 31736 20226 31748
rect 20346 31736 20352 31748
rect 20220 31708 20352 31736
rect 20220 31696 20226 31708
rect 20346 31696 20352 31708
rect 20404 31696 20410 31748
rect 21821 31739 21879 31745
rect 21821 31736 21833 31739
rect 21744 31708 21833 31736
rect 21744 31680 21772 31708
rect 21821 31705 21833 31708
rect 21867 31705 21879 31739
rect 21933 31736 21961 31767
rect 22370 31736 22376 31748
rect 21933 31708 22376 31736
rect 21821 31699 21879 31705
rect 22370 31696 22376 31708
rect 22428 31696 22434 31748
rect 22664 31736 22692 31844
rect 22756 31844 23305 31872
rect 22756 31813 22784 31844
rect 23293 31841 23305 31844
rect 23339 31841 23351 31875
rect 23293 31835 23351 31841
rect 23753 31875 23811 31881
rect 23753 31841 23765 31875
rect 23799 31872 23811 31875
rect 23799 31844 24440 31872
rect 23799 31841 23811 31844
rect 23753 31835 23811 31841
rect 22741 31807 22799 31813
rect 22741 31773 22753 31807
rect 22787 31773 22799 31807
rect 22741 31767 22799 31773
rect 22830 31764 22836 31816
rect 22888 31804 22894 31816
rect 23017 31807 23075 31813
rect 23017 31804 23029 31807
rect 22888 31776 23029 31804
rect 22888 31764 22894 31776
rect 23017 31773 23029 31776
rect 23063 31773 23075 31807
rect 23017 31767 23075 31773
rect 23474 31764 23480 31816
rect 23532 31804 23538 31816
rect 24412 31813 24440 31844
rect 24486 31832 24492 31884
rect 24544 31832 24550 31884
rect 24854 31872 24860 31884
rect 24596 31844 24860 31872
rect 23569 31807 23627 31813
rect 23569 31804 23581 31807
rect 23532 31776 23581 31804
rect 23532 31764 23538 31776
rect 23569 31773 23581 31776
rect 23615 31773 23627 31807
rect 24029 31807 24087 31813
rect 24029 31804 24041 31807
rect 23569 31767 23627 31773
rect 23952 31776 24041 31804
rect 23290 31736 23296 31748
rect 22664 31708 23296 31736
rect 23290 31696 23296 31708
rect 23348 31696 23354 31748
rect 23952 31736 23980 31776
rect 24029 31773 24041 31776
rect 24075 31773 24087 31807
rect 24029 31767 24087 31773
rect 24397 31807 24455 31813
rect 24397 31773 24409 31807
rect 24443 31804 24455 31807
rect 24596 31804 24624 31844
rect 24854 31832 24860 31844
rect 24912 31832 24918 31884
rect 25314 31832 25320 31884
rect 25372 31872 25378 31884
rect 25866 31872 25872 31884
rect 25372 31844 25872 31872
rect 25372 31832 25378 31844
rect 25866 31832 25872 31844
rect 25924 31832 25930 31884
rect 26804 31881 26832 31912
rect 26878 31900 26884 31912
rect 26936 31900 26942 31952
rect 26970 31900 26976 31952
rect 27028 31900 27034 31952
rect 27157 31943 27215 31949
rect 27157 31909 27169 31943
rect 27203 31940 27215 31943
rect 27356 31940 27384 31968
rect 27203 31912 27384 31940
rect 27617 31943 27675 31949
rect 27203 31909 27215 31912
rect 27157 31903 27215 31909
rect 27617 31909 27629 31943
rect 27663 31909 27675 31943
rect 28902 31940 28908 31952
rect 27617 31903 27675 31909
rect 28460 31912 28908 31940
rect 26789 31875 26847 31881
rect 26789 31841 26801 31875
rect 26835 31841 26847 31875
rect 26988 31872 27016 31900
rect 26789 31835 26847 31841
rect 26896 31844 27016 31872
rect 24443 31776 24624 31804
rect 24673 31807 24731 31813
rect 24443 31773 24455 31776
rect 24397 31767 24455 31773
rect 24673 31773 24685 31807
rect 24719 31804 24731 31807
rect 24762 31804 24768 31816
rect 24719 31776 24768 31804
rect 24719 31773 24731 31776
rect 24673 31767 24731 31773
rect 24688 31736 24716 31767
rect 24762 31764 24768 31776
rect 24820 31764 24826 31816
rect 26418 31764 26424 31816
rect 26476 31804 26482 31816
rect 26694 31804 26700 31816
rect 26476 31776 26700 31804
rect 26476 31764 26482 31776
rect 26694 31764 26700 31776
rect 26752 31764 26758 31816
rect 23584 31708 24716 31736
rect 23584 31680 23612 31708
rect 24946 31696 24952 31748
rect 25004 31696 25010 31748
rect 25133 31739 25191 31745
rect 25133 31705 25145 31739
rect 25179 31705 25191 31739
rect 25133 31699 25191 31705
rect 16172 31640 16620 31668
rect 16172 31628 16178 31640
rect 16850 31628 16856 31680
rect 16908 31668 16914 31680
rect 21082 31668 21088 31680
rect 16908 31640 21088 31668
rect 16908 31628 16914 31640
rect 21082 31628 21088 31640
rect 21140 31628 21146 31680
rect 21726 31628 21732 31680
rect 21784 31628 21790 31680
rect 22094 31628 22100 31680
rect 22152 31628 22158 31680
rect 23566 31628 23572 31680
rect 23624 31628 23630 31680
rect 24854 31628 24860 31680
rect 24912 31628 24918 31680
rect 25148 31668 25176 31699
rect 26326 31696 26332 31748
rect 26384 31696 26390 31748
rect 26418 31668 26424 31680
rect 25148 31640 26424 31668
rect 26418 31628 26424 31640
rect 26476 31628 26482 31680
rect 26539 31671 26597 31677
rect 26539 31637 26551 31671
rect 26585 31668 26597 31671
rect 26896 31668 26924 31844
rect 26973 31807 27031 31813
rect 26973 31773 26985 31807
rect 27019 31773 27031 31807
rect 26973 31767 27031 31773
rect 26988 31680 27016 31767
rect 27246 31764 27252 31816
rect 27304 31764 27310 31816
rect 27433 31807 27491 31813
rect 27433 31773 27445 31807
rect 27479 31804 27491 31807
rect 27522 31804 27528 31816
rect 27479 31776 27528 31804
rect 27479 31773 27491 31776
rect 27433 31767 27491 31773
rect 27522 31764 27528 31776
rect 27580 31764 27586 31816
rect 27632 31804 27660 31903
rect 27709 31807 27767 31813
rect 27709 31804 27721 31807
rect 27632 31776 27721 31804
rect 27709 31773 27721 31776
rect 27755 31773 27767 31807
rect 27709 31767 27767 31773
rect 27801 31807 27859 31813
rect 27801 31773 27813 31807
rect 27847 31804 27859 31807
rect 27847 31776 27881 31804
rect 27847 31773 27859 31776
rect 27801 31767 27859 31773
rect 27154 31696 27160 31748
rect 27212 31736 27218 31748
rect 27816 31736 27844 31767
rect 28074 31764 28080 31816
rect 28132 31804 28138 31816
rect 28460 31813 28488 31912
rect 28902 31900 28908 31912
rect 28960 31900 28966 31952
rect 29086 31900 29092 31952
rect 29144 31940 29150 31952
rect 29181 31943 29239 31949
rect 29181 31940 29193 31943
rect 29144 31912 29193 31940
rect 29144 31900 29150 31912
rect 29181 31909 29193 31912
rect 29227 31940 29239 31943
rect 30006 31940 30012 31952
rect 29227 31912 30012 31940
rect 29227 31909 29239 31912
rect 29181 31903 29239 31909
rect 30006 31900 30012 31912
rect 30064 31900 30070 31952
rect 31849 31943 31907 31949
rect 31849 31940 31861 31943
rect 30300 31912 31861 31940
rect 30300 31884 30328 31912
rect 31849 31909 31861 31912
rect 31895 31909 31907 31943
rect 31849 31903 31907 31909
rect 28552 31844 29224 31872
rect 28445 31807 28503 31813
rect 28445 31804 28457 31807
rect 28132 31776 28457 31804
rect 28132 31764 28138 31776
rect 28445 31773 28457 31776
rect 28491 31773 28503 31807
rect 28445 31767 28503 31773
rect 27212 31708 27844 31736
rect 27212 31696 27218 31708
rect 28166 31696 28172 31748
rect 28224 31736 28230 31748
rect 28552 31736 28580 31844
rect 28629 31807 28687 31813
rect 28629 31773 28641 31807
rect 28675 31804 28687 31807
rect 28675 31776 28948 31804
rect 28675 31773 28687 31776
rect 28629 31767 28687 31773
rect 28813 31739 28871 31745
rect 28813 31736 28825 31739
rect 28224 31708 28825 31736
rect 28224 31696 28230 31708
rect 28813 31705 28825 31708
rect 28859 31705 28871 31739
rect 28920 31736 28948 31776
rect 28994 31764 29000 31816
rect 29052 31764 29058 31816
rect 29196 31804 29224 31844
rect 29638 31832 29644 31884
rect 29696 31872 29702 31884
rect 29917 31875 29975 31881
rect 29917 31872 29929 31875
rect 29696 31844 29929 31872
rect 29696 31832 29702 31844
rect 29917 31841 29929 31844
rect 29963 31841 29975 31875
rect 29917 31835 29975 31841
rect 30282 31832 30288 31884
rect 30340 31832 30346 31884
rect 31573 31875 31631 31881
rect 31573 31872 31585 31875
rect 30668 31844 31585 31872
rect 30374 31804 30380 31816
rect 29196 31798 29408 31804
rect 29472 31798 30380 31804
rect 29196 31776 30380 31798
rect 29380 31770 29500 31776
rect 30374 31764 30380 31776
rect 30432 31764 30438 31816
rect 29086 31736 29092 31748
rect 28920 31708 29092 31736
rect 28813 31699 28871 31705
rect 29086 31696 29092 31708
rect 29144 31736 29150 31748
rect 29546 31736 29552 31748
rect 29144 31708 29552 31736
rect 29144 31696 29150 31708
rect 29546 31696 29552 31708
rect 29604 31696 29610 31748
rect 29733 31739 29791 31745
rect 29733 31705 29745 31739
rect 29779 31736 29791 31739
rect 30558 31736 30564 31748
rect 29779 31708 30564 31736
rect 29779 31705 29791 31708
rect 29733 31699 29791 31705
rect 30558 31696 30564 31708
rect 30616 31736 30622 31748
rect 30668 31736 30696 31844
rect 31573 31841 31585 31844
rect 31619 31872 31631 31875
rect 31754 31872 31760 31884
rect 31619 31844 31760 31872
rect 31619 31841 31631 31844
rect 31573 31835 31631 31841
rect 31754 31832 31760 31844
rect 31812 31832 31818 31884
rect 31864 31872 31892 31903
rect 34422 31900 34428 31952
rect 34480 31940 34486 31952
rect 34624 31940 34652 31968
rect 35069 31943 35127 31949
rect 35069 31940 35081 31943
rect 34480 31912 34560 31940
rect 34624 31912 35081 31940
rect 34480 31900 34486 31912
rect 33594 31872 33600 31884
rect 31864 31844 33600 31872
rect 33594 31832 33600 31844
rect 33652 31832 33658 31884
rect 34532 31872 34560 31912
rect 35069 31909 35081 31912
rect 35115 31909 35127 31943
rect 35728 31940 35756 31980
rect 36630 31968 36636 32020
rect 36688 31968 36694 32020
rect 36722 31968 36728 32020
rect 36780 32008 36786 32020
rect 37090 32008 37096 32020
rect 36780 31980 37096 32008
rect 36780 31968 36786 31980
rect 37090 31968 37096 31980
rect 37148 32008 37154 32020
rect 37277 32011 37335 32017
rect 37277 32008 37289 32011
rect 37148 31980 37289 32008
rect 37148 31968 37154 31980
rect 37277 31977 37289 31980
rect 37323 31977 37335 32011
rect 37277 31971 37335 31977
rect 37458 31968 37464 32020
rect 37516 32008 37522 32020
rect 38657 32011 38715 32017
rect 38657 32008 38669 32011
rect 37516 31980 38669 32008
rect 37516 31968 37522 31980
rect 38657 31977 38669 31980
rect 38703 31977 38715 32011
rect 38657 31971 38715 31977
rect 37829 31943 37887 31949
rect 35728 31912 37412 31940
rect 35069 31903 35127 31909
rect 35710 31872 35716 31884
rect 34164 31844 34560 31872
rect 34716 31844 35716 31872
rect 30837 31807 30895 31813
rect 30837 31773 30849 31807
rect 30883 31773 30895 31807
rect 30837 31767 30895 31773
rect 31021 31807 31079 31813
rect 31021 31773 31033 31807
rect 31067 31804 31079 31807
rect 31202 31804 31208 31816
rect 31067 31776 31208 31804
rect 31067 31773 31079 31776
rect 31021 31767 31079 31773
rect 30616 31708 30696 31736
rect 30852 31736 30880 31767
rect 31202 31764 31208 31776
rect 31260 31764 31266 31816
rect 31297 31807 31355 31813
rect 31297 31773 31309 31807
rect 31343 31804 31355 31807
rect 31478 31804 31484 31816
rect 31343 31776 31484 31804
rect 31343 31773 31355 31776
rect 31297 31767 31355 31773
rect 31478 31764 31484 31776
rect 31536 31804 31542 31816
rect 31849 31807 31907 31813
rect 31849 31804 31861 31807
rect 31536 31776 31861 31804
rect 31536 31764 31542 31776
rect 31849 31773 31861 31776
rect 31895 31773 31907 31807
rect 31849 31767 31907 31773
rect 32122 31764 32128 31816
rect 32180 31764 32186 31816
rect 32398 31764 32404 31816
rect 32456 31804 32462 31816
rect 33226 31804 33232 31816
rect 32456 31776 33232 31804
rect 32456 31764 32462 31776
rect 33226 31764 33232 31776
rect 33284 31804 33290 31816
rect 33505 31807 33563 31813
rect 33505 31804 33517 31807
rect 33284 31776 33517 31804
rect 33284 31764 33290 31776
rect 33505 31773 33517 31776
rect 33551 31773 33563 31807
rect 33505 31767 33563 31773
rect 33962 31764 33968 31816
rect 34020 31764 34026 31816
rect 34164 31813 34192 31844
rect 34149 31807 34207 31813
rect 34149 31773 34161 31807
rect 34195 31773 34207 31807
rect 34149 31767 34207 31773
rect 34238 31764 34244 31816
rect 34296 31804 34302 31816
rect 34333 31807 34391 31813
rect 34333 31804 34345 31807
rect 34296 31776 34345 31804
rect 34296 31764 34302 31776
rect 34333 31773 34345 31776
rect 34379 31773 34391 31807
rect 34333 31767 34391 31773
rect 34425 31807 34483 31813
rect 34425 31773 34437 31807
rect 34471 31804 34483 31807
rect 34606 31804 34612 31816
rect 34471 31776 34612 31804
rect 34471 31773 34483 31776
rect 34425 31767 34483 31773
rect 32140 31736 32168 31764
rect 30852 31708 32168 31736
rect 30616 31696 30622 31708
rect 32674 31696 32680 31748
rect 32732 31736 32738 31748
rect 33321 31739 33379 31745
rect 33321 31736 33333 31739
rect 32732 31708 33333 31736
rect 32732 31696 32738 31708
rect 33321 31705 33333 31708
rect 33367 31705 33379 31739
rect 33321 31699 33379 31705
rect 34057 31739 34115 31745
rect 34057 31705 34069 31739
rect 34103 31705 34115 31739
rect 34348 31736 34376 31767
rect 34606 31764 34612 31776
rect 34664 31764 34670 31816
rect 34716 31813 34744 31844
rect 35710 31832 35716 31844
rect 35768 31832 35774 31884
rect 36814 31872 36820 31884
rect 36372 31844 36820 31872
rect 34701 31807 34759 31813
rect 34701 31773 34713 31807
rect 34747 31773 34759 31807
rect 34701 31767 34759 31773
rect 34882 31764 34888 31816
rect 34940 31764 34946 31816
rect 35342 31764 35348 31816
rect 35400 31804 35406 31816
rect 36372 31813 36400 31844
rect 36814 31832 36820 31844
rect 36872 31832 36878 31884
rect 36998 31832 37004 31884
rect 37056 31832 37062 31884
rect 35621 31807 35679 31813
rect 35621 31804 35633 31807
rect 35400 31776 35633 31804
rect 35400 31764 35406 31776
rect 35621 31773 35633 31776
rect 35667 31773 35679 31807
rect 35621 31767 35679 31773
rect 35989 31807 36047 31813
rect 35989 31773 36001 31807
rect 36035 31773 36047 31807
rect 35989 31767 36047 31773
rect 36357 31807 36415 31813
rect 36357 31773 36369 31807
rect 36403 31773 36415 31807
rect 36357 31767 36415 31773
rect 36541 31807 36599 31813
rect 36541 31773 36553 31807
rect 36587 31804 36599 31807
rect 37016 31804 37044 31832
rect 36587 31776 37044 31804
rect 36587 31773 36599 31776
rect 36541 31767 36599 31773
rect 34974 31736 34980 31748
rect 34348 31708 34980 31736
rect 34057 31699 34115 31705
rect 26585 31640 26924 31668
rect 26585 31637 26597 31640
rect 26539 31631 26597 31637
rect 26970 31628 26976 31680
rect 27028 31628 27034 31680
rect 27890 31628 27896 31680
rect 27948 31668 27954 31680
rect 28077 31671 28135 31677
rect 28077 31668 28089 31671
rect 27948 31640 28089 31668
rect 27948 31628 27954 31640
rect 28077 31637 28089 31640
rect 28123 31637 28135 31671
rect 28077 31631 28135 31637
rect 29454 31628 29460 31680
rect 29512 31668 29518 31680
rect 30837 31671 30895 31677
rect 30837 31668 30849 31671
rect 29512 31640 30849 31668
rect 29512 31628 29518 31640
rect 30837 31637 30849 31640
rect 30883 31637 30895 31671
rect 30837 31631 30895 31637
rect 31478 31628 31484 31680
rect 31536 31668 31542 31680
rect 32490 31668 32496 31680
rect 31536 31640 32496 31668
rect 31536 31628 31542 31640
rect 32490 31628 32496 31640
rect 32548 31628 32554 31680
rect 33502 31628 33508 31680
rect 33560 31668 33566 31680
rect 33689 31671 33747 31677
rect 33689 31668 33701 31671
rect 33560 31640 33701 31668
rect 33560 31628 33566 31640
rect 33689 31637 33701 31640
rect 33735 31637 33747 31671
rect 33689 31631 33747 31637
rect 33778 31628 33784 31680
rect 33836 31628 33842 31680
rect 33870 31628 33876 31680
rect 33928 31668 33934 31680
rect 34072 31668 34100 31699
rect 34974 31696 34980 31708
rect 35032 31736 35038 31748
rect 36004 31736 36032 31767
rect 35032 31708 36032 31736
rect 37185 31739 37243 31745
rect 35032 31696 35038 31708
rect 35728 31680 35756 31708
rect 37185 31705 37197 31739
rect 37231 31736 37243 31739
rect 37274 31736 37280 31748
rect 37231 31708 37280 31736
rect 37231 31705 37243 31708
rect 37185 31699 37243 31705
rect 37274 31696 37280 31708
rect 37332 31696 37338 31748
rect 37384 31736 37412 31912
rect 37829 31909 37841 31943
rect 37875 31909 37887 31943
rect 37829 31903 37887 31909
rect 37550 31764 37556 31816
rect 37608 31764 37614 31816
rect 37642 31764 37648 31816
rect 37700 31764 37706 31816
rect 37844 31804 37872 31903
rect 38562 31900 38568 31952
rect 38620 31900 38626 31952
rect 38028 31844 38516 31872
rect 37921 31807 37979 31813
rect 37921 31804 37933 31807
rect 37844 31776 37933 31804
rect 37921 31773 37933 31776
rect 37967 31773 37979 31807
rect 37921 31767 37979 31773
rect 38028 31736 38056 31844
rect 37384 31708 38056 31736
rect 38194 31696 38200 31748
rect 38252 31696 38258 31748
rect 38488 31736 38516 31844
rect 38580 31813 38608 31900
rect 38672 31844 41644 31872
rect 38565 31807 38623 31813
rect 38565 31773 38577 31807
rect 38611 31773 38623 31807
rect 38565 31767 38623 31773
rect 38672 31736 38700 31844
rect 41616 31816 41644 31844
rect 41598 31764 41604 31816
rect 41656 31764 41662 31816
rect 38488 31708 38700 31736
rect 33928 31640 34100 31668
rect 33928 31628 33934 31640
rect 34514 31628 34520 31680
rect 34572 31668 34578 31680
rect 35342 31668 35348 31680
rect 34572 31640 35348 31668
rect 34572 31628 34578 31640
rect 35342 31628 35348 31640
rect 35400 31628 35406 31680
rect 35710 31628 35716 31680
rect 35768 31628 35774 31680
rect 1104 31578 41400 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 41400 31578
rect 1104 31504 41400 31526
rect 8938 31464 8944 31476
rect 2240 31436 8944 31464
rect 2038 31288 2044 31340
rect 2096 31288 2102 31340
rect 2240 31337 2268 31436
rect 2501 31399 2559 31405
rect 2501 31365 2513 31399
rect 2547 31396 2559 31399
rect 2774 31396 2780 31408
rect 2547 31368 2780 31396
rect 2547 31365 2559 31368
rect 2501 31359 2559 31365
rect 2774 31356 2780 31368
rect 2832 31356 2838 31408
rect 3050 31356 3056 31408
rect 3108 31356 3114 31408
rect 2225 31331 2283 31337
rect 2225 31297 2237 31331
rect 2271 31297 2283 31331
rect 2225 31291 2283 31297
rect 4890 31288 4896 31340
rect 4948 31288 4954 31340
rect 4982 31288 4988 31340
rect 5040 31288 5046 31340
rect 6656 31337 6684 31436
rect 8938 31424 8944 31436
rect 8996 31424 9002 31476
rect 10042 31424 10048 31476
rect 10100 31464 10106 31476
rect 14366 31464 14372 31476
rect 10100 31436 14372 31464
rect 10100 31424 10106 31436
rect 14366 31424 14372 31436
rect 14424 31424 14430 31476
rect 15470 31464 15476 31476
rect 15304 31436 15476 31464
rect 7190 31356 7196 31408
rect 7248 31396 7254 31408
rect 8956 31396 8984 31424
rect 15102 31396 15108 31408
rect 7248 31368 7406 31396
rect 8956 31368 11560 31396
rect 13018 31368 15108 31396
rect 7248 31356 7254 31368
rect 6641 31331 6699 31337
rect 6641 31297 6653 31331
rect 6687 31297 6699 31331
rect 6641 31291 6699 31297
rect 8941 31331 8999 31337
rect 8941 31297 8953 31331
rect 8987 31328 8999 31331
rect 9490 31328 9496 31340
rect 8987 31300 9496 31328
rect 8987 31297 8999 31300
rect 8941 31291 8999 31297
rect 9490 31288 9496 31300
rect 9548 31288 9554 31340
rect 11532 31337 11560 31368
rect 15102 31356 15108 31368
rect 15160 31356 15166 31408
rect 15304 31405 15332 31436
rect 15470 31424 15476 31436
rect 15528 31424 15534 31476
rect 16206 31424 16212 31476
rect 16264 31424 16270 31476
rect 16298 31424 16304 31476
rect 16356 31464 16362 31476
rect 16761 31467 16819 31473
rect 16761 31464 16773 31467
rect 16356 31436 16773 31464
rect 16356 31424 16362 31436
rect 16761 31433 16773 31436
rect 16807 31433 16819 31467
rect 20990 31464 20996 31476
rect 16761 31427 16819 31433
rect 17604 31436 18552 31464
rect 15289 31399 15347 31405
rect 15289 31365 15301 31399
rect 15335 31365 15347 31399
rect 15841 31399 15899 31405
rect 15841 31396 15853 31399
rect 15289 31359 15347 31365
rect 15396 31368 15853 31396
rect 11517 31331 11575 31337
rect 11517 31297 11529 31331
rect 11563 31297 11575 31331
rect 11517 31291 11575 31297
rect 14274 31288 14280 31340
rect 14332 31328 14338 31340
rect 14369 31331 14427 31337
rect 14369 31328 14381 31331
rect 14332 31300 14381 31328
rect 14332 31288 14338 31300
rect 14369 31297 14381 31300
rect 14415 31297 14427 31331
rect 14369 31291 14427 31297
rect 15194 31288 15200 31340
rect 15252 31328 15258 31340
rect 15396 31328 15424 31368
rect 15841 31365 15853 31368
rect 15887 31396 15899 31399
rect 15930 31396 15936 31408
rect 15887 31368 15936 31396
rect 15887 31365 15899 31368
rect 15841 31359 15899 31365
rect 15930 31356 15936 31368
rect 15988 31356 15994 31408
rect 16025 31399 16083 31405
rect 16025 31365 16037 31399
rect 16071 31396 16083 31399
rect 16942 31396 16948 31408
rect 16071 31368 16948 31396
rect 16071 31365 16083 31368
rect 16025 31359 16083 31365
rect 16942 31356 16948 31368
rect 17000 31356 17006 31408
rect 17494 31356 17500 31408
rect 17552 31396 17558 31408
rect 17604 31396 17632 31436
rect 18524 31396 18552 31436
rect 19444 31436 20996 31464
rect 19444 31396 19472 31436
rect 20990 31424 20996 31436
rect 21048 31424 21054 31476
rect 21082 31424 21088 31476
rect 21140 31464 21146 31476
rect 22186 31464 22192 31476
rect 21140 31436 22192 31464
rect 21140 31424 21146 31436
rect 22186 31424 22192 31436
rect 22244 31424 22250 31476
rect 22554 31464 22560 31476
rect 22296 31436 22560 31464
rect 17552 31368 17710 31396
rect 18524 31368 19550 31396
rect 17552 31356 17558 31368
rect 15252 31300 15424 31328
rect 15473 31331 15531 31337
rect 15252 31288 15258 31300
rect 15473 31297 15485 31331
rect 15519 31328 15531 31331
rect 16114 31328 16120 31340
rect 15519 31300 16120 31328
rect 15519 31297 15531 31300
rect 15473 31291 15531 31297
rect 16114 31288 16120 31300
rect 16172 31328 16178 31340
rect 16301 31331 16359 31337
rect 16301 31328 16313 31331
rect 16172 31300 16313 31328
rect 16172 31288 16178 31300
rect 16301 31297 16313 31300
rect 16347 31297 16359 31331
rect 16301 31291 16359 31297
rect 16482 31288 16488 31340
rect 16540 31328 16546 31340
rect 16669 31331 16727 31337
rect 16669 31328 16681 31331
rect 16540 31300 16681 31328
rect 16540 31288 16546 31300
rect 16669 31297 16681 31300
rect 16715 31297 16727 31331
rect 16669 31291 16727 31297
rect 16853 31331 16911 31337
rect 16853 31297 16865 31331
rect 16899 31328 16911 31331
rect 16960 31328 16988 31356
rect 22296 31337 22324 31436
rect 22554 31424 22560 31436
rect 22612 31464 22618 31476
rect 22922 31464 22928 31476
rect 22612 31436 22928 31464
rect 22612 31424 22618 31436
rect 22922 31424 22928 31436
rect 22980 31424 22986 31476
rect 23109 31467 23167 31473
rect 23109 31433 23121 31467
rect 23155 31464 23167 31467
rect 23750 31464 23756 31476
rect 23155 31436 23756 31464
rect 23155 31433 23167 31436
rect 23109 31427 23167 31433
rect 23750 31424 23756 31436
rect 23808 31424 23814 31476
rect 24026 31464 24032 31476
rect 23952 31436 24032 31464
rect 23952 31405 23980 31436
rect 24026 31424 24032 31436
rect 24084 31424 24090 31476
rect 24118 31424 24124 31476
rect 24176 31424 24182 31476
rect 24305 31467 24363 31473
rect 24305 31433 24317 31467
rect 24351 31464 24363 31467
rect 24946 31464 24952 31476
rect 24351 31436 24952 31464
rect 24351 31433 24363 31436
rect 24305 31427 24363 31433
rect 24946 31424 24952 31436
rect 25004 31424 25010 31476
rect 26973 31467 27031 31473
rect 26973 31433 26985 31467
rect 27019 31464 27031 31467
rect 27246 31464 27252 31476
rect 27019 31436 27252 31464
rect 27019 31433 27031 31436
rect 26973 31427 27031 31433
rect 27246 31424 27252 31436
rect 27304 31424 27310 31476
rect 27338 31424 27344 31476
rect 27396 31464 27402 31476
rect 27617 31467 27675 31473
rect 27617 31464 27629 31467
rect 27396 31436 27629 31464
rect 27396 31424 27402 31436
rect 27617 31433 27629 31436
rect 27663 31464 27675 31467
rect 27663 31436 27936 31464
rect 27663 31433 27675 31436
rect 27617 31427 27675 31433
rect 23937 31399 23995 31405
rect 23937 31365 23949 31399
rect 23983 31365 23995 31399
rect 24136 31396 24164 31424
rect 24670 31396 24676 31408
rect 24136 31368 24676 31396
rect 23937 31359 23995 31365
rect 24670 31356 24676 31368
rect 24728 31396 24734 31408
rect 24765 31399 24823 31405
rect 24765 31396 24777 31399
rect 24728 31368 24777 31396
rect 24728 31356 24734 31368
rect 24765 31365 24777 31368
rect 24811 31365 24823 31399
rect 24765 31359 24823 31365
rect 26697 31399 26755 31405
rect 26697 31365 26709 31399
rect 26743 31396 26755 31399
rect 27798 31396 27804 31408
rect 26743 31368 27804 31396
rect 26743 31365 26755 31368
rect 26697 31359 26755 31365
rect 27798 31356 27804 31368
rect 27856 31356 27862 31408
rect 27908 31396 27936 31436
rect 28994 31424 29000 31476
rect 29052 31464 29058 31476
rect 29362 31464 29368 31476
rect 29052 31436 29368 31464
rect 29052 31424 29058 31436
rect 29362 31424 29368 31436
rect 29420 31424 29426 31476
rect 29730 31424 29736 31476
rect 29788 31464 29794 31476
rect 30926 31464 30932 31476
rect 29788 31436 30932 31464
rect 29788 31424 29794 31436
rect 30926 31424 30932 31436
rect 30984 31424 30990 31476
rect 31018 31424 31024 31476
rect 31076 31464 31082 31476
rect 32493 31467 32551 31473
rect 32493 31464 32505 31467
rect 31076 31436 32505 31464
rect 31076 31424 31082 31436
rect 32493 31433 32505 31436
rect 32539 31433 32551 31467
rect 33502 31464 33508 31476
rect 32493 31427 32551 31433
rect 33336 31436 33508 31464
rect 33137 31399 33195 31405
rect 33137 31396 33149 31399
rect 27908 31368 29776 31396
rect 16899 31300 16988 31328
rect 21361 31331 21419 31337
rect 16899 31297 16911 31300
rect 16853 31291 16911 31297
rect 21361 31297 21373 31331
rect 21407 31297 21419 31331
rect 21361 31291 21419 31297
rect 21545 31331 21603 31337
rect 21545 31297 21557 31331
rect 21591 31297 21603 31331
rect 21545 31291 21603 31297
rect 21821 31331 21879 31337
rect 21821 31297 21833 31331
rect 21867 31297 21879 31331
rect 21821 31291 21879 31297
rect 22281 31331 22339 31337
rect 22281 31297 22293 31331
rect 22327 31297 22339 31331
rect 22281 31291 22339 31297
rect 22480 31300 22876 31328
rect 3694 31220 3700 31272
rect 3752 31260 3758 31272
rect 4249 31263 4307 31269
rect 4249 31260 4261 31263
rect 3752 31232 4261 31260
rect 3752 31220 3758 31232
rect 4249 31229 4261 31232
rect 4295 31229 4307 31263
rect 4249 31223 4307 31229
rect 6917 31263 6975 31269
rect 6917 31229 6929 31263
rect 6963 31260 6975 31263
rect 7650 31260 7656 31272
rect 6963 31232 7656 31260
rect 6963 31229 6975 31232
rect 6917 31223 6975 31229
rect 7650 31220 7656 31232
rect 7708 31220 7714 31272
rect 8570 31220 8576 31272
rect 8628 31260 8634 31272
rect 8849 31263 8907 31269
rect 8849 31260 8861 31263
rect 8628 31232 8861 31260
rect 8628 31220 8634 31232
rect 8849 31229 8861 31232
rect 8895 31229 8907 31263
rect 8849 31223 8907 31229
rect 9309 31263 9367 31269
rect 9309 31229 9321 31263
rect 9355 31260 9367 31263
rect 9858 31260 9864 31272
rect 9355 31232 9864 31260
rect 9355 31229 9367 31232
rect 9309 31223 9367 31229
rect 9858 31220 9864 31232
rect 9916 31220 9922 31272
rect 11790 31220 11796 31272
rect 11848 31220 11854 31272
rect 13538 31220 13544 31272
rect 13596 31220 13602 31272
rect 14182 31220 14188 31272
rect 14240 31220 14246 31272
rect 14458 31220 14464 31272
rect 14516 31220 14522 31272
rect 14734 31220 14740 31272
rect 14792 31260 14798 31272
rect 16945 31263 17003 31269
rect 16945 31260 16957 31263
rect 14792 31232 16957 31260
rect 14792 31220 14798 31232
rect 16945 31229 16957 31232
rect 16991 31229 17003 31263
rect 16945 31223 17003 31229
rect 5261 31195 5319 31201
rect 5261 31161 5273 31195
rect 5307 31192 5319 31195
rect 6178 31192 6184 31204
rect 5307 31164 6184 31192
rect 5307 31161 5319 31164
rect 5261 31155 5319 31161
rect 6178 31152 6184 31164
rect 6236 31152 6242 31204
rect 14200 31192 14228 31220
rect 15657 31195 15715 31201
rect 15657 31192 15669 31195
rect 14200 31164 15669 31192
rect 15657 31161 15669 31164
rect 15703 31161 15715 31195
rect 16574 31192 16580 31204
rect 15657 31155 15715 31161
rect 16224 31164 16580 31192
rect 1762 31084 1768 31136
rect 1820 31124 1826 31136
rect 1857 31127 1915 31133
rect 1857 31124 1869 31127
rect 1820 31096 1869 31124
rect 1820 31084 1826 31096
rect 1857 31093 1869 31096
rect 1903 31093 1915 31127
rect 1857 31087 1915 31093
rect 5074 31084 5080 31136
rect 5132 31124 5138 31136
rect 6730 31124 6736 31136
rect 5132 31096 6736 31124
rect 5132 31084 5138 31096
rect 6730 31084 6736 31096
rect 6788 31084 6794 31136
rect 7282 31084 7288 31136
rect 7340 31124 7346 31136
rect 7926 31124 7932 31136
rect 7340 31096 7932 31124
rect 7340 31084 7346 31096
rect 7926 31084 7932 31096
rect 7984 31084 7990 31136
rect 8386 31084 8392 31136
rect 8444 31084 8450 31136
rect 14737 31127 14795 31133
rect 14737 31093 14749 31127
rect 14783 31124 14795 31127
rect 16224 31124 16252 31164
rect 16574 31152 16580 31164
rect 16632 31152 16638 31204
rect 14783 31096 16252 31124
rect 14783 31093 14795 31096
rect 14737 31087 14795 31093
rect 16390 31084 16396 31136
rect 16448 31084 16454 31136
rect 16960 31124 16988 31223
rect 17218 31220 17224 31272
rect 17276 31220 17282 31272
rect 18690 31260 18696 31272
rect 18248 31232 18696 31260
rect 18248 31124 18276 31232
rect 18690 31220 18696 31232
rect 18748 31260 18754 31272
rect 18785 31263 18843 31269
rect 18785 31260 18797 31263
rect 18748 31232 18797 31260
rect 18748 31220 18754 31232
rect 18785 31229 18797 31232
rect 18831 31229 18843 31263
rect 18785 31223 18843 31229
rect 19058 31220 19064 31272
rect 19116 31220 19122 31272
rect 20625 31263 20683 31269
rect 20625 31260 20637 31263
rect 20548 31232 20637 31260
rect 16960 31096 18276 31124
rect 18693 31127 18751 31133
rect 18693 31093 18705 31127
rect 18739 31124 18751 31127
rect 19242 31124 19248 31136
rect 18739 31096 19248 31124
rect 18739 31093 18751 31096
rect 18693 31087 18751 31093
rect 19242 31084 19248 31096
rect 19300 31084 19306 31136
rect 20438 31084 20444 31136
rect 20496 31124 20502 31136
rect 20548 31133 20576 31232
rect 20625 31229 20637 31232
rect 20671 31260 20683 31263
rect 21376 31260 21404 31291
rect 20671 31232 21404 31260
rect 20671 31229 20683 31232
rect 20625 31223 20683 31229
rect 21560 31192 21588 31291
rect 20640 31164 21588 31192
rect 21836 31192 21864 31291
rect 21913 31263 21971 31269
rect 21913 31229 21925 31263
rect 21959 31260 21971 31263
rect 22002 31260 22008 31272
rect 21959 31232 22008 31260
rect 21959 31229 21971 31232
rect 21913 31223 21971 31229
rect 22002 31220 22008 31232
rect 22060 31260 22066 31272
rect 22186 31260 22192 31272
rect 22060 31232 22192 31260
rect 22060 31220 22066 31232
rect 22186 31220 22192 31232
rect 22244 31260 22250 31272
rect 22373 31263 22431 31269
rect 22373 31260 22385 31263
rect 22244 31232 22385 31260
rect 22244 31220 22250 31232
rect 22373 31229 22385 31232
rect 22419 31229 22431 31263
rect 22373 31223 22431 31229
rect 22480 31192 22508 31300
rect 22557 31263 22615 31269
rect 22557 31229 22569 31263
rect 22603 31260 22615 31263
rect 22603 31232 22784 31260
rect 22603 31229 22615 31232
rect 22557 31223 22615 31229
rect 21836 31164 22508 31192
rect 20640 31136 20668 31164
rect 20533 31127 20591 31133
rect 20533 31124 20545 31127
rect 20496 31096 20545 31124
rect 20496 31084 20502 31096
rect 20533 31093 20545 31096
rect 20579 31093 20591 31127
rect 20533 31087 20591 31093
rect 20622 31084 20628 31136
rect 20680 31084 20686 31136
rect 21266 31084 21272 31136
rect 21324 31084 21330 31136
rect 21361 31127 21419 31133
rect 21361 31093 21373 31127
rect 21407 31124 21419 31127
rect 21726 31124 21732 31136
rect 21407 31096 21732 31124
rect 21407 31093 21419 31096
rect 21361 31087 21419 31093
rect 21726 31084 21732 31096
rect 21784 31084 21790 31136
rect 22005 31127 22063 31133
rect 22005 31093 22017 31127
rect 22051 31124 22063 31127
rect 22094 31124 22100 31136
rect 22051 31096 22100 31124
rect 22051 31093 22063 31096
rect 22005 31087 22063 31093
rect 22094 31084 22100 31096
rect 22152 31084 22158 31136
rect 22186 31084 22192 31136
rect 22244 31084 22250 31136
rect 22278 31084 22284 31136
rect 22336 31084 22342 31136
rect 22756 31124 22784 31232
rect 22848 31192 22876 31300
rect 22922 31288 22928 31340
rect 22980 31328 22986 31340
rect 23017 31331 23075 31337
rect 23017 31328 23029 31331
rect 22980 31300 23029 31328
rect 22980 31288 22986 31300
rect 23017 31297 23029 31300
rect 23063 31297 23075 31331
rect 23017 31291 23075 31297
rect 23566 31288 23572 31340
rect 23624 31328 23630 31340
rect 23842 31337 23848 31340
rect 23661 31331 23719 31337
rect 23661 31328 23673 31331
rect 23624 31300 23673 31328
rect 23624 31288 23630 31300
rect 23661 31297 23673 31300
rect 23707 31297 23719 31331
rect 23661 31291 23719 31297
rect 23809 31331 23848 31337
rect 23809 31297 23821 31331
rect 23809 31291 23848 31297
rect 23842 31288 23848 31291
rect 23900 31288 23906 31340
rect 24029 31331 24087 31337
rect 24029 31328 24041 31331
rect 23952 31300 24041 31328
rect 23952 31272 23980 31300
rect 24029 31297 24041 31300
rect 24075 31297 24087 31331
rect 24029 31291 24087 31297
rect 24123 31288 24129 31340
rect 24181 31288 24187 31340
rect 24228 31300 24532 31328
rect 23934 31220 23940 31272
rect 23992 31260 23998 31272
rect 24228 31260 24256 31300
rect 23992 31232 24256 31260
rect 23992 31220 23998 31232
rect 24302 31220 24308 31272
rect 24360 31260 24366 31272
rect 24397 31263 24455 31269
rect 24397 31260 24409 31263
rect 24360 31232 24409 31260
rect 24360 31220 24366 31232
rect 24397 31229 24409 31232
rect 24443 31229 24455 31263
rect 24504 31260 24532 31300
rect 24578 31288 24584 31340
rect 24636 31288 24642 31340
rect 25222 31288 25228 31340
rect 25280 31328 25286 31340
rect 25409 31331 25467 31337
rect 25409 31328 25421 31331
rect 25280 31300 25421 31328
rect 25280 31288 25286 31300
rect 25409 31297 25421 31300
rect 25455 31297 25467 31331
rect 25409 31291 25467 31297
rect 25501 31331 25559 31337
rect 25501 31297 25513 31331
rect 25547 31297 25559 31331
rect 25501 31291 25559 31297
rect 25685 31331 25743 31337
rect 25685 31297 25697 31331
rect 25731 31297 25743 31331
rect 25685 31291 25743 31297
rect 24762 31260 24768 31272
rect 24504 31232 24768 31260
rect 24397 31223 24455 31229
rect 24762 31220 24768 31232
rect 24820 31220 24826 31272
rect 25225 31195 25283 31201
rect 25225 31192 25237 31195
rect 22848 31164 25237 31192
rect 25225 31161 25237 31164
rect 25271 31161 25283 31195
rect 25225 31155 25283 31161
rect 25406 31152 25412 31204
rect 25464 31152 25470 31204
rect 25516 31192 25544 31291
rect 25700 31260 25728 31291
rect 25774 31288 25780 31340
rect 25832 31288 25838 31340
rect 25866 31288 25872 31340
rect 25924 31288 25930 31340
rect 26510 31288 26516 31340
rect 26568 31328 26574 31340
rect 27341 31331 27399 31337
rect 27341 31328 27353 31331
rect 26568 31300 27353 31328
rect 26568 31288 26574 31300
rect 27341 31297 27353 31300
rect 27387 31297 27399 31331
rect 27341 31291 27399 31297
rect 27709 31331 27767 31337
rect 27709 31297 27721 31331
rect 27755 31328 27767 31331
rect 27890 31328 27896 31340
rect 27755 31300 27896 31328
rect 27755 31297 27767 31300
rect 27709 31291 27767 31297
rect 27890 31288 27896 31300
rect 27948 31288 27954 31340
rect 29086 31288 29092 31340
rect 29144 31328 29150 31340
rect 29273 31331 29331 31337
rect 29273 31328 29285 31331
rect 29144 31300 29285 31328
rect 29144 31288 29150 31300
rect 29273 31297 29285 31300
rect 29319 31328 29331 31331
rect 29641 31331 29699 31337
rect 29641 31328 29653 31331
rect 29319 31300 29653 31328
rect 29319 31297 29331 31300
rect 29273 31291 29331 31297
rect 29641 31297 29653 31300
rect 29687 31297 29699 31331
rect 29641 31291 29699 31297
rect 27433 31263 27491 31269
rect 27433 31260 27445 31263
rect 25700 31232 27445 31260
rect 27433 31229 27445 31232
rect 27479 31260 27491 31263
rect 28534 31260 28540 31272
rect 27479 31232 28540 31260
rect 27479 31229 27491 31232
rect 27433 31223 27491 31229
rect 28534 31220 28540 31232
rect 28592 31220 28598 31272
rect 29546 31220 29552 31272
rect 29604 31220 29610 31272
rect 29748 31260 29776 31368
rect 29932 31368 33149 31396
rect 29932 31337 29960 31368
rect 33137 31365 33149 31368
rect 33183 31365 33195 31399
rect 33137 31359 33195 31365
rect 29917 31331 29975 31337
rect 29917 31297 29929 31331
rect 29963 31297 29975 31331
rect 31386 31328 31392 31340
rect 29917 31291 29975 31297
rect 30024 31300 31392 31328
rect 30024 31260 30052 31300
rect 31386 31288 31392 31300
rect 31444 31288 31450 31340
rect 31478 31288 31484 31340
rect 31536 31288 31542 31340
rect 31665 31331 31723 31337
rect 31665 31297 31677 31331
rect 31711 31328 31723 31331
rect 31754 31328 31760 31340
rect 31711 31300 31760 31328
rect 31711 31297 31723 31300
rect 31665 31291 31723 31297
rect 31754 31288 31760 31300
rect 31812 31288 31818 31340
rect 32125 31331 32183 31337
rect 32125 31297 32137 31331
rect 32171 31328 32183 31331
rect 32398 31328 32404 31340
rect 32171 31300 32404 31328
rect 32171 31297 32183 31300
rect 32125 31291 32183 31297
rect 32398 31288 32404 31300
rect 32456 31288 32462 31340
rect 32490 31288 32496 31340
rect 32548 31328 32554 31340
rect 33336 31337 33364 31436
rect 33502 31424 33508 31436
rect 33560 31424 33566 31476
rect 33870 31424 33876 31476
rect 33928 31464 33934 31476
rect 34882 31464 34888 31476
rect 33928 31436 34888 31464
rect 33928 31424 33934 31436
rect 34882 31424 34888 31436
rect 34940 31464 34946 31476
rect 35069 31467 35127 31473
rect 35069 31464 35081 31467
rect 34940 31436 35081 31464
rect 34940 31424 34946 31436
rect 35069 31433 35081 31436
rect 35115 31433 35127 31467
rect 35069 31427 35127 31433
rect 35802 31424 35808 31476
rect 35860 31464 35866 31476
rect 36906 31464 36912 31476
rect 35860 31436 36912 31464
rect 35860 31424 35866 31436
rect 36906 31424 36912 31436
rect 36964 31464 36970 31476
rect 41046 31464 41052 31476
rect 36964 31436 41052 31464
rect 36964 31424 36970 31436
rect 41046 31424 41052 31436
rect 41104 31424 41110 31476
rect 33643 31399 33701 31405
rect 33643 31365 33655 31399
rect 33689 31396 33701 31399
rect 33778 31396 33784 31408
rect 33689 31368 33784 31396
rect 33689 31365 33701 31368
rect 33643 31359 33701 31365
rect 33778 31356 33784 31368
rect 33836 31356 33842 31408
rect 34698 31356 34704 31408
rect 34756 31396 34762 31408
rect 35526 31396 35532 31408
rect 34756 31368 35532 31396
rect 34756 31356 34762 31368
rect 35526 31356 35532 31368
rect 35584 31356 35590 31408
rect 37737 31399 37795 31405
rect 37737 31365 37749 31399
rect 37783 31396 37795 31399
rect 37783 31368 38516 31396
rect 37783 31365 37795 31368
rect 37737 31359 37795 31365
rect 32585 31331 32643 31337
rect 32585 31328 32597 31331
rect 32548 31300 32597 31328
rect 32548 31288 32554 31300
rect 32585 31297 32597 31300
rect 32631 31297 32643 31331
rect 32585 31291 32643 31297
rect 33321 31331 33379 31337
rect 33321 31297 33333 31331
rect 33367 31297 33379 31331
rect 33321 31291 33379 31297
rect 29748 31232 30052 31260
rect 30377 31263 30435 31269
rect 30377 31229 30389 31263
rect 30423 31229 30435 31263
rect 30377 31223 30435 31229
rect 25516 31164 25728 31192
rect 25424 31124 25452 31152
rect 25700 31136 25728 31164
rect 25958 31152 25964 31204
rect 26016 31192 26022 31204
rect 26326 31192 26332 31204
rect 26016 31164 26332 31192
rect 26016 31152 26022 31164
rect 26326 31152 26332 31164
rect 26384 31152 26390 31204
rect 26418 31152 26424 31204
rect 26476 31192 26482 31204
rect 27522 31192 27528 31204
rect 26476 31164 27528 31192
rect 26476 31152 26482 31164
rect 27522 31152 27528 31164
rect 27580 31192 27586 31204
rect 30392 31192 30420 31223
rect 30926 31220 30932 31272
rect 30984 31260 30990 31272
rect 32217 31263 32275 31269
rect 32217 31260 32229 31263
rect 30984 31232 32229 31260
rect 30984 31220 30990 31232
rect 32217 31229 32229 31232
rect 32263 31229 32275 31263
rect 32600 31260 32628 31291
rect 33410 31288 33416 31340
rect 33468 31288 33474 31340
rect 33505 31331 33563 31337
rect 33505 31297 33517 31331
rect 33551 31297 33563 31331
rect 33505 31291 33563 31297
rect 33520 31260 33548 31291
rect 34054 31288 34060 31340
rect 34112 31328 34118 31340
rect 34885 31331 34943 31337
rect 34885 31328 34897 31331
rect 34112 31300 34897 31328
rect 34112 31288 34118 31300
rect 34885 31297 34897 31300
rect 34931 31297 34943 31331
rect 34885 31291 34943 31297
rect 34974 31288 34980 31340
rect 35032 31288 35038 31340
rect 38010 31288 38016 31340
rect 38068 31288 38074 31340
rect 38488 31337 38516 31368
rect 40034 31356 40040 31408
rect 40092 31356 40098 31408
rect 38473 31331 38531 31337
rect 38473 31297 38485 31331
rect 38519 31328 38531 31331
rect 38562 31328 38568 31340
rect 38519 31300 38568 31328
rect 38519 31297 38531 31300
rect 38473 31291 38531 31297
rect 38562 31288 38568 31300
rect 38620 31288 38626 31340
rect 38749 31331 38807 31337
rect 38749 31297 38761 31331
rect 38795 31328 38807 31331
rect 38930 31328 38936 31340
rect 38795 31300 38936 31328
rect 38795 31297 38807 31300
rect 38749 31291 38807 31297
rect 38930 31288 38936 31300
rect 38988 31288 38994 31340
rect 32600 31232 33548 31260
rect 32217 31223 32275 31229
rect 27580 31164 30420 31192
rect 32232 31192 32260 31223
rect 33520 31192 33548 31232
rect 33594 31220 33600 31272
rect 33652 31260 33658 31272
rect 33781 31263 33839 31269
rect 33781 31260 33793 31263
rect 33652 31232 33793 31260
rect 33652 31220 33658 31232
rect 33781 31229 33793 31232
rect 33827 31229 33839 31263
rect 33781 31223 33839 31229
rect 33962 31220 33968 31272
rect 34020 31260 34026 31272
rect 34238 31260 34244 31272
rect 34020 31232 34244 31260
rect 34020 31220 34026 31232
rect 34238 31220 34244 31232
rect 34296 31220 34302 31272
rect 34330 31220 34336 31272
rect 34388 31220 34394 31272
rect 34422 31220 34428 31272
rect 34480 31220 34486 31272
rect 34517 31263 34575 31269
rect 34517 31229 34529 31263
rect 34563 31229 34575 31263
rect 34517 31223 34575 31229
rect 34701 31263 34759 31269
rect 34701 31229 34713 31263
rect 34747 31260 34759 31263
rect 34790 31260 34796 31272
rect 34747 31232 34796 31260
rect 34747 31229 34759 31232
rect 34701 31223 34759 31229
rect 34057 31195 34115 31201
rect 34057 31192 34069 31195
rect 32232 31164 32812 31192
rect 33520 31164 34069 31192
rect 27580 31152 27586 31164
rect 22756 31096 25452 31124
rect 25682 31084 25688 31136
rect 25740 31084 25746 31136
rect 25774 31084 25780 31136
rect 25832 31124 25838 31136
rect 26786 31124 26792 31136
rect 25832 31096 26792 31124
rect 25832 31084 25838 31096
rect 26786 31084 26792 31096
rect 26844 31084 26850 31136
rect 27246 31084 27252 31136
rect 27304 31084 27310 31136
rect 28258 31084 28264 31136
rect 28316 31124 28322 31136
rect 28534 31124 28540 31136
rect 28316 31096 28540 31124
rect 28316 31084 28322 31096
rect 28534 31084 28540 31096
rect 28592 31084 28598 31136
rect 29089 31127 29147 31133
rect 29089 31093 29101 31127
rect 29135 31124 29147 31127
rect 29270 31124 29276 31136
rect 29135 31096 29276 31124
rect 29135 31093 29147 31096
rect 29089 31087 29147 31093
rect 29270 31084 29276 31096
rect 29328 31084 29334 31136
rect 29454 31084 29460 31136
rect 29512 31084 29518 31136
rect 30098 31084 30104 31136
rect 30156 31084 30162 31136
rect 31478 31084 31484 31136
rect 31536 31124 31542 31136
rect 31849 31127 31907 31133
rect 31849 31124 31861 31127
rect 31536 31096 31861 31124
rect 31536 31084 31542 31096
rect 31849 31093 31861 31096
rect 31895 31093 31907 31127
rect 31849 31087 31907 31093
rect 32122 31084 32128 31136
rect 32180 31084 32186 31136
rect 32674 31084 32680 31136
rect 32732 31084 32738 31136
rect 32784 31124 32812 31164
rect 34057 31161 34069 31164
rect 34103 31161 34115 31195
rect 34532 31192 34560 31223
rect 34790 31220 34796 31232
rect 34848 31220 34854 31272
rect 34992 31192 35020 31288
rect 38194 31220 38200 31272
rect 38252 31260 38258 31272
rect 38289 31263 38347 31269
rect 38289 31260 38301 31263
rect 38252 31232 38301 31260
rect 38252 31220 38258 31232
rect 38289 31229 38301 31232
rect 38335 31260 38347 31263
rect 38335 31232 38976 31260
rect 38335 31229 38347 31232
rect 38289 31223 38347 31229
rect 38948 31201 38976 31232
rect 39022 31220 39028 31272
rect 39080 31260 39086 31272
rect 39301 31263 39359 31269
rect 39301 31260 39313 31263
rect 39080 31232 39313 31260
rect 39080 31220 39086 31232
rect 39301 31229 39313 31232
rect 39347 31229 39359 31263
rect 39301 31223 39359 31229
rect 39574 31220 39580 31272
rect 39632 31220 39638 31272
rect 38933 31195 38991 31201
rect 34532 31164 35020 31192
rect 38488 31164 38792 31192
rect 34057 31155 34115 31161
rect 33594 31124 33600 31136
rect 32784 31096 33600 31124
rect 33594 31084 33600 31096
rect 33652 31084 33658 31136
rect 37274 31084 37280 31136
rect 37332 31124 37338 31136
rect 37829 31127 37887 31133
rect 37829 31124 37841 31127
rect 37332 31096 37841 31124
rect 37332 31084 37338 31096
rect 37829 31093 37841 31096
rect 37875 31124 37887 31127
rect 38378 31124 38384 31136
rect 37875 31096 38384 31124
rect 37875 31093 37887 31096
rect 37829 31087 37887 31093
rect 38378 31084 38384 31096
rect 38436 31084 38442 31136
rect 38488 31133 38516 31164
rect 38764 31136 38792 31164
rect 38933 31161 38945 31195
rect 38979 31161 38991 31195
rect 38933 31155 38991 31161
rect 38473 31127 38531 31133
rect 38473 31093 38485 31127
rect 38519 31093 38531 31127
rect 38473 31087 38531 31093
rect 38654 31084 38660 31136
rect 38712 31084 38718 31136
rect 38746 31084 38752 31136
rect 38804 31084 38810 31136
rect 41049 31127 41107 31133
rect 41049 31093 41061 31127
rect 41095 31124 41107 31127
rect 41095 31096 41460 31124
rect 41095 31093 41107 31096
rect 41049 31087 41107 31093
rect 1104 31034 41400 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 41400 31034
rect 1104 30960 41400 30982
rect 2958 30880 2964 30932
rect 3016 30920 3022 30932
rect 3789 30923 3847 30929
rect 3789 30920 3801 30923
rect 3016 30892 3801 30920
rect 3016 30880 3022 30892
rect 3789 30889 3801 30892
rect 3835 30889 3847 30923
rect 3789 30883 3847 30889
rect 11790 30880 11796 30932
rect 11848 30920 11854 30932
rect 12897 30923 12955 30929
rect 12897 30920 12909 30923
rect 11848 30892 12909 30920
rect 11848 30880 11854 30892
rect 12897 30889 12909 30892
rect 12943 30889 12955 30923
rect 12897 30883 12955 30889
rect 13538 30880 13544 30932
rect 13596 30880 13602 30932
rect 15102 30880 15108 30932
rect 15160 30880 15166 30932
rect 17218 30880 17224 30932
rect 17276 30920 17282 30932
rect 17589 30923 17647 30929
rect 17589 30920 17601 30923
rect 17276 30892 17601 30920
rect 17276 30880 17282 30892
rect 17589 30889 17601 30892
rect 17635 30889 17647 30923
rect 17589 30883 17647 30889
rect 19058 30880 19064 30932
rect 19116 30920 19122 30932
rect 20533 30923 20591 30929
rect 20533 30920 20545 30923
rect 19116 30892 20545 30920
rect 19116 30880 19122 30892
rect 20533 30889 20545 30892
rect 20579 30889 20591 30923
rect 20533 30883 20591 30889
rect 21266 30880 21272 30932
rect 21324 30880 21330 30932
rect 21818 30880 21824 30932
rect 21876 30920 21882 30932
rect 22189 30923 22247 30929
rect 22189 30920 22201 30923
rect 21876 30892 22201 30920
rect 21876 30880 21882 30892
rect 22189 30889 22201 30892
rect 22235 30889 22247 30923
rect 22189 30883 22247 30889
rect 22278 30880 22284 30932
rect 22336 30880 22342 30932
rect 22830 30880 22836 30932
rect 22888 30880 22894 30932
rect 23106 30880 23112 30932
rect 23164 30920 23170 30932
rect 24210 30920 24216 30932
rect 23164 30892 24216 30920
rect 23164 30880 23170 30892
rect 24210 30880 24216 30892
rect 24268 30880 24274 30932
rect 24394 30880 24400 30932
rect 24452 30880 24458 30932
rect 26053 30923 26111 30929
rect 26053 30920 26065 30923
rect 24780 30892 26065 30920
rect 11606 30812 11612 30864
rect 11664 30852 11670 30864
rect 12342 30852 12348 30864
rect 11664 30824 12348 30852
rect 11664 30812 11670 30824
rect 12342 30812 12348 30824
rect 12400 30812 12406 30864
rect 12452 30824 13032 30852
rect 1673 30787 1731 30793
rect 1673 30753 1685 30787
rect 1719 30784 1731 30787
rect 1762 30784 1768 30796
rect 1719 30756 1768 30784
rect 1719 30753 1731 30756
rect 1673 30747 1731 30753
rect 1762 30744 1768 30756
rect 1820 30744 1826 30796
rect 3418 30744 3424 30796
rect 3476 30784 3482 30796
rect 4341 30787 4399 30793
rect 4341 30784 4353 30787
rect 3476 30756 4353 30784
rect 3476 30744 3482 30756
rect 4341 30753 4353 30756
rect 4387 30753 4399 30787
rect 4341 30747 4399 30753
rect 5074 30744 5080 30796
rect 5132 30744 5138 30796
rect 10965 30787 11023 30793
rect 10965 30753 10977 30787
rect 11011 30784 11023 30787
rect 11011 30756 12204 30784
rect 11011 30753 11023 30756
rect 10965 30747 11023 30753
rect 1394 30676 1400 30728
rect 1452 30676 1458 30728
rect 3050 30716 3056 30728
rect 2806 30688 3056 30716
rect 3050 30676 3056 30688
rect 3108 30676 3114 30728
rect 4249 30719 4307 30725
rect 4249 30685 4261 30719
rect 4295 30716 4307 30719
rect 5092 30716 5120 30744
rect 10870 30716 10876 30728
rect 4295 30688 5120 30716
rect 10612 30688 10876 30716
rect 4295 30685 4307 30688
rect 4249 30679 4307 30685
rect 2958 30608 2964 30660
rect 3016 30648 3022 30660
rect 3421 30651 3479 30657
rect 3421 30648 3433 30651
rect 3016 30620 3433 30648
rect 3016 30608 3022 30620
rect 3421 30617 3433 30620
rect 3467 30617 3479 30651
rect 3421 30611 3479 30617
rect 4062 30608 4068 30660
rect 4120 30648 4126 30660
rect 4120 30620 4292 30648
rect 4120 30608 4126 30620
rect 3694 30540 3700 30592
rect 3752 30580 3758 30592
rect 4157 30583 4215 30589
rect 4157 30580 4169 30583
rect 3752 30552 4169 30580
rect 3752 30540 3758 30552
rect 4157 30549 4169 30552
rect 4203 30549 4215 30583
rect 4264 30580 4292 30620
rect 10226 30608 10232 30660
rect 10284 30648 10290 30660
rect 10612 30657 10640 30688
rect 10870 30676 10876 30688
rect 10928 30676 10934 30728
rect 11241 30719 11299 30725
rect 11241 30716 11253 30719
rect 10981 30688 11253 30716
rect 10597 30651 10655 30657
rect 10597 30648 10609 30651
rect 10284 30620 10609 30648
rect 10284 30608 10290 30620
rect 10597 30617 10609 30620
rect 10643 30617 10655 30651
rect 10597 30611 10655 30617
rect 10781 30651 10839 30657
rect 10781 30617 10793 30651
rect 10827 30648 10839 30651
rect 10981 30648 11009 30688
rect 11241 30685 11253 30688
rect 11287 30716 11299 30719
rect 11701 30719 11759 30725
rect 11701 30716 11713 30719
rect 11287 30688 11713 30716
rect 11287 30685 11299 30688
rect 11241 30679 11299 30685
rect 11701 30685 11713 30688
rect 11747 30716 11759 30719
rect 12066 30716 12072 30728
rect 11747 30688 12072 30716
rect 11747 30685 11759 30688
rect 11701 30679 11759 30685
rect 12066 30676 12072 30688
rect 12124 30676 12130 30728
rect 12176 30725 12204 30756
rect 12452 30728 12480 30824
rect 12621 30787 12679 30793
rect 12621 30753 12633 30787
rect 12667 30784 12679 30787
rect 12667 30756 12848 30784
rect 12667 30753 12679 30756
rect 12621 30747 12679 30753
rect 12161 30719 12219 30725
rect 12161 30685 12173 30719
rect 12207 30685 12219 30719
rect 12161 30679 12219 30685
rect 12434 30676 12440 30728
rect 12492 30676 12498 30728
rect 12526 30676 12532 30728
rect 12584 30676 12590 30728
rect 12820 30725 12848 30756
rect 13004 30725 13032 30824
rect 12713 30719 12771 30725
rect 12713 30685 12725 30719
rect 12759 30685 12771 30719
rect 12713 30679 12771 30685
rect 12805 30719 12863 30725
rect 12805 30685 12817 30719
rect 12851 30685 12863 30719
rect 12805 30679 12863 30685
rect 12989 30719 13047 30725
rect 12989 30685 13001 30719
rect 13035 30685 13047 30719
rect 12989 30679 13047 30685
rect 10827 30620 11009 30648
rect 11057 30651 11115 30657
rect 10827 30617 10839 30620
rect 10781 30611 10839 30617
rect 11057 30617 11069 30651
rect 11103 30648 11115 30651
rect 11146 30648 11152 30660
rect 11103 30620 11152 30648
rect 11103 30617 11115 30620
rect 11057 30611 11115 30617
rect 11146 30608 11152 30620
rect 11204 30608 11210 30660
rect 11422 30608 11428 30660
rect 11480 30608 11486 30660
rect 11514 30608 11520 30660
rect 11572 30608 11578 30660
rect 12728 30648 12756 30679
rect 13556 30648 13584 30880
rect 15120 30852 15148 30880
rect 17126 30852 17132 30864
rect 15120 30824 17132 30852
rect 17126 30812 17132 30824
rect 17184 30852 17190 30864
rect 17494 30852 17500 30864
rect 17184 30824 17500 30852
rect 17184 30812 17190 30824
rect 17494 30812 17500 30824
rect 17552 30812 17558 30864
rect 19150 30852 19156 30864
rect 17788 30824 19156 30852
rect 14642 30744 14648 30796
rect 14700 30784 14706 30796
rect 16390 30784 16396 30796
rect 14700 30756 16396 30784
rect 14700 30744 14706 30756
rect 16390 30744 16396 30756
rect 16448 30744 16454 30796
rect 16574 30744 16580 30796
rect 16632 30784 16638 30796
rect 17586 30784 17592 30796
rect 16632 30756 17592 30784
rect 16632 30744 16638 30756
rect 17586 30744 17592 30756
rect 17644 30744 17650 30796
rect 17788 30793 17816 30824
rect 19150 30812 19156 30824
rect 19208 30852 19214 30864
rect 19208 30824 20024 30852
rect 19208 30812 19214 30824
rect 17773 30787 17831 30793
rect 17773 30753 17785 30787
rect 17819 30753 17831 30787
rect 17773 30747 17831 30753
rect 18141 30787 18199 30793
rect 18141 30753 18153 30787
rect 18187 30784 18199 30787
rect 19889 30787 19947 30793
rect 19889 30784 19901 30787
rect 18187 30756 19901 30784
rect 18187 30753 18199 30756
rect 18141 30747 18199 30753
rect 19889 30753 19901 30756
rect 19935 30753 19947 30787
rect 19889 30747 19947 30753
rect 17865 30719 17923 30725
rect 17865 30685 17877 30719
rect 17911 30685 17923 30719
rect 17865 30679 17923 30685
rect 11624 30620 13584 30648
rect 17880 30648 17908 30679
rect 17954 30676 17960 30728
rect 18012 30716 18018 30728
rect 18325 30719 18383 30725
rect 18325 30716 18337 30719
rect 18012 30688 18337 30716
rect 18012 30676 18018 30688
rect 18325 30685 18337 30688
rect 18371 30685 18383 30719
rect 18325 30679 18383 30685
rect 19245 30719 19303 30725
rect 19245 30685 19257 30719
rect 19291 30716 19303 30719
rect 19334 30716 19340 30728
rect 19291 30688 19340 30716
rect 19291 30685 19303 30688
rect 19245 30679 19303 30685
rect 19334 30676 19340 30688
rect 19392 30676 19398 30728
rect 19996 30725 20024 30824
rect 21284 30784 21312 30880
rect 22002 30852 22008 30864
rect 20272 30756 21312 30784
rect 21475 30824 22008 30852
rect 20272 30725 20300 30756
rect 19981 30719 20039 30725
rect 19981 30685 19993 30719
rect 20027 30685 20039 30719
rect 19981 30679 20039 30685
rect 20257 30719 20315 30725
rect 20257 30685 20269 30719
rect 20303 30685 20315 30719
rect 20257 30679 20315 30685
rect 20349 30719 20407 30725
rect 20349 30685 20361 30719
rect 20395 30685 20407 30719
rect 20349 30679 20407 30685
rect 18046 30648 18052 30660
rect 17880 30620 18052 30648
rect 11624 30580 11652 30620
rect 18046 30608 18052 30620
rect 18104 30608 18110 30660
rect 18138 30608 18144 30660
rect 18196 30608 18202 30660
rect 18230 30608 18236 30660
rect 18288 30608 18294 30660
rect 18810 30651 18868 30657
rect 18810 30648 18822 30651
rect 18340 30620 18822 30648
rect 4264 30552 11652 30580
rect 11793 30583 11851 30589
rect 4157 30543 4215 30549
rect 11793 30549 11805 30583
rect 11839 30580 11851 30583
rect 11974 30580 11980 30592
rect 11839 30552 11980 30580
rect 11839 30549 11851 30552
rect 11793 30543 11851 30549
rect 11974 30540 11980 30552
rect 12032 30540 12038 30592
rect 12710 30540 12716 30592
rect 12768 30580 12774 30592
rect 16850 30580 16856 30592
rect 12768 30552 16856 30580
rect 12768 30540 12774 30552
rect 16850 30540 16856 30552
rect 16908 30540 16914 30592
rect 18156 30580 18184 30608
rect 18340 30580 18368 30620
rect 18810 30617 18822 30620
rect 18856 30617 18868 30651
rect 20165 30651 20223 30657
rect 20165 30648 20177 30651
rect 18810 30611 18868 30617
rect 18984 30620 20177 30648
rect 18156 30552 18368 30580
rect 18598 30540 18604 30592
rect 18656 30540 18662 30592
rect 18690 30540 18696 30592
rect 18748 30540 18754 30592
rect 18984 30589 19012 30620
rect 20165 30617 20177 30620
rect 20211 30617 20223 30651
rect 20165 30611 20223 30617
rect 18969 30583 19027 30589
rect 18969 30549 18981 30583
rect 19015 30549 19027 30583
rect 18969 30543 19027 30549
rect 19058 30540 19064 30592
rect 19116 30580 19122 30592
rect 20364 30580 20392 30679
rect 20438 30676 20444 30728
rect 20496 30716 20502 30728
rect 20993 30719 21051 30725
rect 20993 30716 21005 30719
rect 20496 30688 21005 30716
rect 20496 30676 20502 30688
rect 20993 30685 21005 30688
rect 21039 30685 21051 30719
rect 20993 30679 21051 30685
rect 21174 30676 21180 30728
rect 21232 30716 21238 30728
rect 21475 30716 21503 30824
rect 22002 30812 22008 30824
rect 22060 30812 22066 30864
rect 22296 30852 22324 30880
rect 22204 30824 22324 30852
rect 22848 30852 22876 30880
rect 24486 30852 24492 30864
rect 22848 30824 24492 30852
rect 22204 30784 22232 30824
rect 24486 30812 24492 30824
rect 24544 30812 24550 30864
rect 24780 30793 24808 30892
rect 26053 30889 26065 30892
rect 26099 30889 26111 30923
rect 26053 30883 26111 30889
rect 24946 30812 24952 30864
rect 25004 30812 25010 30864
rect 24765 30787 24823 30793
rect 24765 30784 24777 30787
rect 21836 30756 22232 30784
rect 22848 30756 24777 30784
rect 21232 30688 21503 30716
rect 21545 30719 21603 30725
rect 21232 30676 21238 30688
rect 21545 30685 21557 30719
rect 21591 30685 21603 30719
rect 21545 30679 21603 30685
rect 20530 30608 20536 30660
rect 20588 30648 20594 30660
rect 21560 30648 21588 30679
rect 21634 30676 21640 30728
rect 21692 30716 21698 30728
rect 21836 30725 21864 30756
rect 22848 30728 22876 30756
rect 24765 30753 24777 30756
rect 24811 30753 24823 30787
rect 24964 30784 24992 30812
rect 26068 30784 26096 30883
rect 26418 30880 26424 30932
rect 26476 30920 26482 30932
rect 26694 30920 26700 30932
rect 26476 30892 26700 30920
rect 26476 30880 26482 30892
rect 26694 30880 26700 30892
rect 26752 30880 26758 30932
rect 29730 30920 29736 30932
rect 27080 30892 29736 30920
rect 26602 30784 26608 30796
rect 24964 30756 25452 30784
rect 26068 30756 26280 30784
rect 24765 30747 24823 30753
rect 21821 30719 21879 30725
rect 21692 30688 21737 30716
rect 21692 30676 21698 30688
rect 21821 30685 21833 30719
rect 21867 30685 21879 30719
rect 21821 30679 21879 30685
rect 22002 30676 22008 30728
rect 22060 30725 22066 30728
rect 22060 30719 22109 30725
rect 22060 30685 22063 30719
rect 22097 30685 22109 30719
rect 22060 30679 22109 30685
rect 22060 30676 22066 30679
rect 22830 30676 22836 30728
rect 22888 30676 22894 30728
rect 23750 30676 23756 30728
rect 23808 30676 23814 30728
rect 24670 30676 24676 30728
rect 24728 30676 24734 30728
rect 24857 30719 24915 30725
rect 24857 30685 24869 30719
rect 24903 30716 24915 30719
rect 25038 30716 25044 30728
rect 24903 30688 25044 30716
rect 24903 30685 24915 30688
rect 24857 30679 24915 30685
rect 25038 30676 25044 30688
rect 25096 30676 25102 30728
rect 25424 30725 25452 30756
rect 26252 30725 26280 30756
rect 26436 30756 26608 30784
rect 26436 30725 26464 30756
rect 26602 30744 26608 30756
rect 26660 30744 26666 30796
rect 27080 30728 27108 30892
rect 29730 30880 29736 30892
rect 29788 30880 29794 30932
rect 32217 30923 32275 30929
rect 32217 30889 32229 30923
rect 32263 30920 32275 30923
rect 32582 30920 32588 30932
rect 32263 30892 32588 30920
rect 32263 30889 32275 30892
rect 32217 30883 32275 30889
rect 32582 30880 32588 30892
rect 32640 30880 32646 30932
rect 32674 30880 32680 30932
rect 32732 30880 32738 30932
rect 37550 30920 37556 30932
rect 36832 30892 37556 30920
rect 31018 30852 31024 30864
rect 28276 30824 31024 30852
rect 28276 30793 28304 30824
rect 31018 30812 31024 30824
rect 31076 30812 31082 30864
rect 31202 30812 31208 30864
rect 31260 30852 31266 30864
rect 31662 30852 31668 30864
rect 31260 30824 31668 30852
rect 31260 30812 31266 30824
rect 31662 30812 31668 30824
rect 31720 30812 31726 30864
rect 32692 30852 32720 30880
rect 32232 30824 32720 30852
rect 28261 30787 28319 30793
rect 28261 30753 28273 30787
rect 28307 30753 28319 30787
rect 28261 30747 28319 30753
rect 28442 30744 28448 30796
rect 28500 30784 28506 30796
rect 28721 30787 28779 30793
rect 28721 30784 28733 30787
rect 28500 30756 28733 30784
rect 28500 30744 28506 30756
rect 28721 30753 28733 30756
rect 28767 30784 28779 30787
rect 28810 30784 28816 30796
rect 28767 30756 28816 30784
rect 28767 30753 28779 30756
rect 28721 30747 28779 30753
rect 28810 30744 28816 30756
rect 28868 30744 28874 30796
rect 30466 30744 30472 30796
rect 30524 30784 30530 30796
rect 31389 30787 31447 30793
rect 31389 30784 31401 30787
rect 30524 30756 31401 30784
rect 30524 30744 30530 30756
rect 31389 30753 31401 30756
rect 31435 30753 31447 30787
rect 32232 30784 32260 30824
rect 33134 30812 33140 30864
rect 33192 30852 33198 30864
rect 35989 30855 36047 30861
rect 35989 30852 36001 30855
rect 33192 30824 36001 30852
rect 33192 30812 33198 30824
rect 35989 30821 36001 30824
rect 36035 30821 36047 30855
rect 35989 30815 36047 30821
rect 31389 30747 31447 30753
rect 31588 30756 32260 30784
rect 25133 30719 25191 30725
rect 25133 30685 25145 30719
rect 25179 30685 25191 30719
rect 25133 30679 25191 30685
rect 25317 30719 25375 30725
rect 25317 30685 25329 30719
rect 25363 30685 25375 30719
rect 25317 30679 25375 30685
rect 25409 30719 25467 30725
rect 25409 30685 25421 30719
rect 25455 30685 25467 30719
rect 25409 30679 25467 30685
rect 26237 30719 26295 30725
rect 26237 30685 26249 30719
rect 26283 30685 26295 30719
rect 26237 30679 26295 30685
rect 26421 30719 26479 30725
rect 26421 30685 26433 30719
rect 26467 30685 26479 30719
rect 26421 30679 26479 30685
rect 26697 30719 26755 30725
rect 26697 30685 26709 30719
rect 26743 30716 26755 30719
rect 26786 30716 26792 30728
rect 26743 30688 26792 30716
rect 26743 30685 26755 30688
rect 26697 30679 26755 30685
rect 20588 30620 21588 30648
rect 21913 30651 21971 30657
rect 20588 30608 20594 30620
rect 21913 30617 21925 30651
rect 21959 30648 21971 30651
rect 23014 30648 23020 30660
rect 21959 30620 23020 30648
rect 21959 30617 21971 30620
rect 21913 30611 21971 30617
rect 23014 30608 23020 30620
rect 23072 30608 23078 30660
rect 23768 30648 23796 30676
rect 25148 30648 25176 30679
rect 23768 30620 25176 30648
rect 25332 30648 25360 30679
rect 25774 30648 25780 30660
rect 25332 30620 25780 30648
rect 25774 30608 25780 30620
rect 25832 30608 25838 30660
rect 25958 30608 25964 30660
rect 26016 30608 26022 30660
rect 26326 30608 26332 30660
rect 26384 30648 26390 30660
rect 26605 30651 26663 30657
rect 26605 30648 26617 30651
rect 26384 30620 26617 30648
rect 26384 30608 26390 30620
rect 26605 30617 26617 30620
rect 26651 30617 26663 30651
rect 26712 30648 26740 30679
rect 26786 30676 26792 30688
rect 26844 30676 26850 30728
rect 26881 30719 26939 30725
rect 26881 30685 26893 30719
rect 26927 30716 26939 30719
rect 27062 30716 27068 30728
rect 26927 30688 27068 30716
rect 26927 30685 26939 30688
rect 26881 30679 26939 30685
rect 27062 30676 27068 30688
rect 27120 30676 27126 30728
rect 27522 30676 27528 30728
rect 27580 30716 27586 30728
rect 28629 30719 28687 30725
rect 28629 30716 28641 30719
rect 27580 30688 28641 30716
rect 27580 30676 27586 30688
rect 28629 30685 28641 30688
rect 28675 30685 28687 30719
rect 28629 30679 28687 30685
rect 28902 30676 28908 30728
rect 28960 30676 28966 30728
rect 29822 30676 29828 30728
rect 29880 30676 29886 30728
rect 31202 30676 31208 30728
rect 31260 30676 31266 30728
rect 31297 30719 31355 30725
rect 31297 30685 31309 30719
rect 31343 30685 31355 30719
rect 31297 30679 31355 30685
rect 29840 30648 29868 30676
rect 26712 30620 29868 30648
rect 31312 30648 31340 30679
rect 31478 30676 31484 30728
rect 31536 30676 31542 30728
rect 31588 30648 31616 30756
rect 32122 30676 32128 30728
rect 32180 30676 32186 30728
rect 32232 30725 32260 30756
rect 32674 30744 32680 30796
rect 32732 30784 32738 30796
rect 34790 30784 34796 30796
rect 32732 30756 34796 30784
rect 32732 30744 32738 30756
rect 34790 30744 34796 30756
rect 34848 30744 34854 30796
rect 36722 30744 36728 30796
rect 36780 30744 36786 30796
rect 32217 30719 32275 30725
rect 32217 30685 32229 30719
rect 32263 30685 32275 30719
rect 32217 30679 32275 30685
rect 33781 30719 33839 30725
rect 33781 30685 33793 30719
rect 33827 30685 33839 30719
rect 33781 30679 33839 30685
rect 33965 30719 34023 30725
rect 33965 30685 33977 30719
rect 34011 30716 34023 30719
rect 34054 30716 34060 30728
rect 34011 30688 34060 30716
rect 34011 30685 34023 30688
rect 33965 30679 34023 30685
rect 31312 30620 31616 30648
rect 31757 30651 31815 30657
rect 26605 30611 26663 30617
rect 31757 30617 31769 30651
rect 31803 30648 31815 30651
rect 33796 30648 33824 30679
rect 34054 30676 34060 30688
rect 34112 30676 34118 30728
rect 35526 30676 35532 30728
rect 35584 30716 35590 30728
rect 35710 30716 35716 30728
rect 35584 30688 35716 30716
rect 35584 30676 35590 30688
rect 35710 30676 35716 30688
rect 35768 30676 35774 30728
rect 36832 30725 36860 30892
rect 37550 30880 37556 30892
rect 37608 30920 37614 30932
rect 38194 30920 38200 30932
rect 37608 30892 38200 30920
rect 37608 30880 37614 30892
rect 38194 30880 38200 30892
rect 38252 30880 38258 30932
rect 38746 30920 38752 30932
rect 38304 30892 38752 30920
rect 37185 30855 37243 30861
rect 37185 30821 37197 30855
rect 37231 30852 37243 30855
rect 37642 30852 37648 30864
rect 37231 30824 37648 30852
rect 37231 30821 37243 30824
rect 37185 30815 37243 30821
rect 37642 30812 37648 30824
rect 37700 30852 37706 30864
rect 37700 30824 37964 30852
rect 37700 30812 37706 30824
rect 37274 30744 37280 30796
rect 37332 30744 37338 30796
rect 37936 30784 37964 30824
rect 38304 30784 38332 30892
rect 38746 30880 38752 30892
rect 38804 30880 38810 30932
rect 39574 30880 39580 30932
rect 39632 30920 39638 30932
rect 39853 30923 39911 30929
rect 39853 30920 39865 30923
rect 39632 30892 39865 30920
rect 39632 30880 39638 30892
rect 39853 30889 39865 30892
rect 39899 30889 39911 30923
rect 39853 30883 39911 30889
rect 39485 30855 39543 30861
rect 39485 30852 39497 30855
rect 37936 30756 38332 30784
rect 38488 30824 39497 30852
rect 37936 30725 37964 30756
rect 35989 30719 36047 30725
rect 35989 30685 36001 30719
rect 36035 30685 36047 30719
rect 35989 30679 36047 30685
rect 36817 30719 36875 30725
rect 36817 30685 36829 30719
rect 36863 30685 36875 30719
rect 36817 30679 36875 30685
rect 37829 30719 37887 30725
rect 37829 30685 37841 30719
rect 37875 30685 37887 30719
rect 37829 30679 37887 30685
rect 37921 30719 37979 30725
rect 37921 30685 37933 30719
rect 37967 30685 37979 30719
rect 37921 30679 37979 30685
rect 34698 30648 34704 30660
rect 31803 30620 33456 30648
rect 33796 30620 34704 30648
rect 31803 30617 31815 30620
rect 31757 30611 31815 30617
rect 19116 30552 20392 30580
rect 19116 30540 19122 30552
rect 20898 30540 20904 30592
rect 20956 30580 20962 30592
rect 21361 30583 21419 30589
rect 21361 30580 21373 30583
rect 20956 30552 21373 30580
rect 20956 30540 20962 30552
rect 21361 30549 21373 30552
rect 21407 30549 21419 30583
rect 23032 30580 23060 30608
rect 33428 30592 33456 30620
rect 34532 30592 34560 30620
rect 34698 30608 34704 30620
rect 34756 30608 34762 30660
rect 36004 30648 36032 30679
rect 37844 30648 37872 30679
rect 38010 30676 38016 30728
rect 38068 30676 38074 30728
rect 38289 30719 38347 30725
rect 38289 30685 38301 30719
rect 38335 30716 38347 30719
rect 38378 30716 38384 30728
rect 38335 30688 38384 30716
rect 38335 30685 38347 30688
rect 38289 30679 38347 30685
rect 38378 30676 38384 30688
rect 38436 30676 38442 30728
rect 38028 30648 38056 30676
rect 38488 30648 38516 30824
rect 39485 30821 39497 30824
rect 39531 30821 39543 30855
rect 39485 30815 39543 30821
rect 38562 30744 38568 30796
rect 38620 30784 38626 30796
rect 41432 30784 41460 31096
rect 38620 30756 41460 30784
rect 38620 30744 38626 30756
rect 38838 30676 38844 30728
rect 38896 30676 38902 30728
rect 39040 30725 39068 30756
rect 39025 30719 39083 30725
rect 39025 30685 39037 30719
rect 39071 30685 39083 30719
rect 39301 30719 39359 30725
rect 39301 30716 39313 30719
rect 39025 30679 39083 30685
rect 39132 30688 39313 30716
rect 36004 30620 36952 30648
rect 37844 30620 38516 30648
rect 38565 30651 38623 30657
rect 36924 30592 36952 30620
rect 38565 30617 38577 30651
rect 38611 30648 38623 30651
rect 38930 30648 38936 30660
rect 38611 30620 38936 30648
rect 38611 30617 38623 30620
rect 38565 30611 38623 30617
rect 38930 30608 38936 30620
rect 38988 30608 38994 30660
rect 23290 30580 23296 30592
rect 23032 30552 23296 30580
rect 21361 30543 21419 30549
rect 23290 30540 23296 30552
rect 23348 30540 23354 30592
rect 25590 30540 25596 30592
rect 25648 30540 25654 30592
rect 25682 30540 25688 30592
rect 25740 30580 25746 30592
rect 26789 30583 26847 30589
rect 26789 30580 26801 30583
rect 25740 30552 26801 30580
rect 25740 30540 25746 30552
rect 26789 30549 26801 30552
rect 26835 30549 26847 30583
rect 26789 30543 26847 30549
rect 27430 30540 27436 30592
rect 27488 30580 27494 30592
rect 31021 30583 31079 30589
rect 31021 30580 31033 30583
rect 27488 30552 31033 30580
rect 27488 30540 27494 30552
rect 31021 30549 31033 30552
rect 31067 30549 31079 30583
rect 31021 30543 31079 30549
rect 32398 30540 32404 30592
rect 32456 30540 32462 30592
rect 33410 30540 33416 30592
rect 33468 30580 33474 30592
rect 33870 30580 33876 30592
rect 33468 30552 33876 30580
rect 33468 30540 33474 30552
rect 33870 30540 33876 30552
rect 33928 30540 33934 30592
rect 34514 30540 34520 30592
rect 34572 30540 34578 30592
rect 36906 30540 36912 30592
rect 36964 30580 36970 30592
rect 37553 30583 37611 30589
rect 37553 30580 37565 30583
rect 36964 30552 37565 30580
rect 36964 30540 36970 30552
rect 37553 30549 37565 30552
rect 37599 30549 37611 30583
rect 37553 30543 37611 30549
rect 38470 30540 38476 30592
rect 38528 30540 38534 30592
rect 38838 30540 38844 30592
rect 38896 30580 38902 30592
rect 39132 30580 39160 30688
rect 39301 30685 39313 30688
rect 39347 30685 39359 30719
rect 39301 30679 39359 30685
rect 40037 30719 40095 30725
rect 40037 30685 40049 30719
rect 40083 30716 40095 30719
rect 41322 30716 41328 30728
rect 40083 30688 41328 30716
rect 40083 30685 40095 30688
rect 40037 30679 40095 30685
rect 41322 30676 41328 30688
rect 41380 30676 41386 30728
rect 38896 30552 39160 30580
rect 38896 30540 38902 30552
rect 39206 30540 39212 30592
rect 39264 30540 39270 30592
rect 1104 30490 41400 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 41400 30490
rect 1104 30416 41400 30438
rect 2038 30336 2044 30388
rect 2096 30376 2102 30388
rect 2409 30379 2467 30385
rect 2409 30376 2421 30379
rect 2096 30348 2421 30376
rect 2096 30336 2102 30348
rect 2409 30345 2421 30348
rect 2455 30345 2467 30379
rect 2409 30339 2467 30345
rect 2774 30336 2780 30388
rect 2832 30336 2838 30388
rect 8938 30376 8944 30388
rect 8404 30348 8944 30376
rect 8036 30280 8248 30308
rect 4798 30200 4804 30252
rect 4856 30240 4862 30252
rect 7926 30240 7932 30252
rect 4856 30212 7932 30240
rect 4856 30200 4862 30212
rect 7926 30200 7932 30212
rect 7984 30200 7990 30252
rect 8036 30249 8064 30280
rect 8220 30252 8248 30280
rect 8021 30243 8079 30249
rect 8021 30209 8033 30243
rect 8067 30209 8079 30243
rect 8021 30203 8079 30209
rect 8114 30243 8172 30249
rect 8114 30209 8126 30243
rect 8160 30209 8172 30243
rect 8114 30203 8172 30209
rect 2866 30132 2872 30184
rect 2924 30132 2930 30184
rect 3053 30175 3111 30181
rect 3053 30141 3065 30175
rect 3099 30172 3111 30175
rect 3326 30172 3332 30184
rect 3099 30144 3332 30172
rect 3099 30141 3111 30144
rect 3053 30135 3111 30141
rect 3326 30132 3332 30144
rect 3384 30132 3390 30184
rect 7834 30132 7840 30184
rect 7892 30172 7898 30184
rect 8128 30172 8156 30203
rect 8202 30200 8208 30252
rect 8260 30200 8266 30252
rect 8404 30249 8432 30348
rect 8938 30336 8944 30348
rect 8996 30336 9002 30388
rect 18046 30336 18052 30388
rect 18104 30376 18110 30388
rect 18509 30379 18567 30385
rect 18509 30376 18521 30379
rect 18104 30348 18521 30376
rect 18104 30336 18110 30348
rect 18509 30345 18521 30348
rect 18555 30345 18567 30379
rect 18509 30339 18567 30345
rect 18877 30379 18935 30385
rect 18877 30345 18889 30379
rect 18923 30376 18935 30379
rect 19058 30376 19064 30388
rect 18923 30348 19064 30376
rect 18923 30345 18935 30348
rect 18877 30339 18935 30345
rect 9585 30311 9643 30317
rect 9585 30277 9597 30311
rect 9631 30277 9643 30311
rect 9585 30271 9643 30277
rect 9677 30311 9735 30317
rect 9677 30277 9689 30311
rect 9723 30308 9735 30311
rect 10870 30308 10876 30320
rect 9723 30280 10876 30308
rect 9723 30277 9735 30280
rect 9677 30271 9735 30277
rect 8570 30249 8576 30252
rect 8297 30243 8355 30249
rect 8297 30209 8309 30243
rect 8343 30209 8355 30243
rect 8297 30203 8355 30209
rect 8389 30243 8447 30249
rect 8389 30209 8401 30243
rect 8435 30209 8447 30243
rect 8389 30203 8447 30209
rect 8527 30243 8576 30249
rect 8527 30209 8539 30243
rect 8573 30209 8576 30243
rect 8527 30203 8576 30209
rect 7892 30144 8156 30172
rect 8312 30172 8340 30203
rect 8570 30200 8576 30203
rect 8628 30200 8634 30252
rect 9306 30200 9312 30252
rect 9364 30200 9370 30252
rect 9490 30249 9496 30252
rect 9457 30243 9496 30249
rect 9457 30209 9469 30243
rect 9457 30203 9496 30209
rect 9490 30200 9496 30203
rect 9548 30200 9554 30252
rect 9600 30240 9628 30271
rect 10870 30268 10876 30280
rect 10928 30308 10934 30320
rect 18892 30308 18920 30339
rect 19058 30336 19064 30348
rect 19116 30336 19122 30388
rect 19242 30376 19248 30388
rect 19168 30348 19248 30376
rect 10928 30280 18000 30308
rect 10928 30268 10934 30280
rect 17972 30252 18000 30280
rect 18340 30280 18920 30308
rect 9815 30243 9873 30249
rect 9600 30212 9766 30240
rect 8846 30172 8852 30184
rect 8312 30144 8852 30172
rect 7892 30132 7898 30144
rect 8846 30132 8852 30144
rect 8904 30172 8910 30184
rect 9738 30172 9766 30212
rect 9815 30209 9827 30243
rect 9861 30240 9873 30243
rect 9950 30240 9956 30252
rect 9861 30212 9956 30240
rect 9861 30209 9873 30212
rect 9815 30203 9873 30209
rect 9950 30200 9956 30212
rect 10008 30200 10014 30252
rect 17954 30200 17960 30252
rect 18012 30240 18018 30252
rect 18012 30212 18057 30240
rect 18012 30200 18018 30212
rect 18230 30200 18236 30252
rect 18288 30238 18294 30252
rect 18340 30249 18368 30280
rect 18966 30268 18972 30320
rect 19024 30308 19030 30320
rect 19168 30308 19196 30348
rect 19242 30336 19248 30348
rect 19300 30336 19306 30388
rect 19812 30348 20576 30376
rect 19812 30308 19840 30348
rect 19024 30280 19196 30308
rect 19260 30280 19840 30308
rect 19889 30311 19947 30317
rect 19024 30268 19030 30280
rect 18325 30243 18383 30249
rect 18325 30238 18337 30243
rect 18288 30210 18337 30238
rect 18288 30200 18294 30210
rect 18325 30209 18337 30210
rect 18371 30209 18383 30243
rect 18325 30203 18383 30209
rect 18693 30243 18751 30249
rect 18693 30209 18705 30243
rect 18739 30240 18751 30243
rect 18782 30240 18788 30252
rect 18739 30212 18788 30240
rect 18739 30209 18751 30212
rect 18693 30203 18751 30209
rect 18782 30200 18788 30212
rect 18840 30200 18846 30252
rect 18877 30243 18935 30249
rect 18877 30209 18889 30243
rect 18923 30209 18935 30243
rect 18877 30203 18935 30209
rect 8904 30144 9812 30172
rect 8904 30132 8910 30144
rect 9784 30116 9812 30144
rect 18598 30132 18604 30184
rect 18656 30172 18662 30184
rect 18892 30172 18920 30203
rect 19260 30184 19288 30280
rect 19889 30277 19901 30311
rect 19935 30308 19947 30311
rect 20438 30308 20444 30320
rect 19935 30280 20444 30308
rect 19935 30277 19947 30280
rect 19889 30271 19947 30277
rect 20438 30268 20444 30280
rect 20496 30268 20502 30320
rect 20548 30308 20576 30348
rect 22186 30336 22192 30388
rect 22244 30376 22250 30388
rect 22738 30376 22744 30388
rect 22244 30348 22744 30376
rect 22244 30336 22250 30348
rect 22738 30336 22744 30348
rect 22796 30376 22802 30388
rect 23750 30376 23756 30388
rect 22796 30348 23756 30376
rect 22796 30336 22802 30348
rect 23750 30336 23756 30348
rect 23808 30336 23814 30388
rect 24670 30336 24676 30388
rect 24728 30376 24734 30388
rect 26326 30376 26332 30388
rect 24728 30348 26332 30376
rect 24728 30336 24734 30348
rect 26326 30336 26332 30348
rect 26384 30376 26390 30388
rect 26384 30348 27200 30376
rect 26384 30336 26390 30348
rect 20717 30311 20775 30317
rect 20717 30308 20729 30311
rect 20548 30280 20729 30308
rect 20717 30277 20729 30280
rect 20763 30277 20775 30311
rect 20717 30271 20775 30277
rect 21174 30268 21180 30320
rect 21232 30268 21238 30320
rect 27172 30308 27200 30348
rect 27246 30336 27252 30388
rect 27304 30376 27310 30388
rect 27525 30379 27583 30385
rect 27525 30376 27537 30379
rect 27304 30348 27537 30376
rect 27304 30336 27310 30348
rect 27525 30345 27537 30348
rect 27571 30345 27583 30379
rect 27890 30376 27896 30388
rect 27525 30339 27583 30345
rect 27632 30348 27896 30376
rect 27632 30308 27660 30348
rect 27890 30336 27896 30348
rect 27948 30336 27954 30388
rect 30098 30336 30104 30388
rect 30156 30336 30162 30388
rect 31846 30336 31852 30388
rect 31904 30376 31910 30388
rect 32861 30379 32919 30385
rect 32861 30376 32873 30379
rect 31904 30348 32873 30376
rect 31904 30336 31910 30348
rect 32861 30345 32873 30348
rect 32907 30345 32919 30379
rect 32861 30339 32919 30345
rect 35636 30348 36400 30376
rect 35636 30308 35664 30348
rect 36372 30308 36400 30348
rect 38562 30336 38568 30388
rect 38620 30336 38626 30388
rect 37369 30311 37427 30317
rect 21284 30280 21680 30308
rect 27172 30280 27660 30308
rect 29380 30280 29868 30308
rect 19334 30200 19340 30252
rect 19392 30240 19398 30252
rect 20073 30243 20131 30249
rect 20073 30240 20085 30243
rect 19392 30212 20085 30240
rect 19392 30200 19398 30212
rect 20073 30209 20085 30212
rect 20119 30240 20131 30243
rect 20533 30243 20591 30249
rect 20119 30212 20392 30240
rect 20119 30209 20131 30212
rect 20073 30203 20131 30209
rect 18656 30144 18920 30172
rect 18656 30132 18662 30144
rect 4890 30064 4896 30116
rect 4948 30104 4954 30116
rect 4948 30076 6500 30104
rect 4948 30064 4954 30076
rect 6472 30048 6500 30076
rect 6546 30064 6552 30116
rect 6604 30104 6610 30116
rect 8665 30107 8723 30113
rect 8665 30104 8677 30107
rect 6604 30076 8677 30104
rect 6604 30064 6610 30076
rect 8665 30073 8677 30076
rect 8711 30073 8723 30107
rect 8665 30067 8723 30073
rect 9766 30064 9772 30116
rect 9824 30064 9830 30116
rect 18892 30104 18920 30144
rect 19242 30132 19248 30184
rect 19300 30132 19306 30184
rect 20364 30181 20392 30212
rect 20533 30209 20545 30243
rect 20579 30240 20591 30243
rect 21192 30240 21220 30268
rect 20579 30212 21220 30240
rect 20579 30209 20591 30212
rect 20533 30203 20591 30209
rect 20349 30175 20407 30181
rect 20349 30141 20361 30175
rect 20395 30172 20407 30175
rect 20622 30172 20628 30184
rect 20395 30144 20628 30172
rect 20395 30141 20407 30144
rect 20349 30135 20407 30141
rect 20622 30132 20628 30144
rect 20680 30132 20686 30184
rect 20901 30175 20959 30181
rect 20901 30141 20913 30175
rect 20947 30141 20959 30175
rect 20901 30135 20959 30141
rect 21085 30175 21143 30181
rect 21085 30141 21097 30175
rect 21131 30172 21143 30175
rect 21174 30172 21180 30184
rect 21131 30144 21180 30172
rect 21131 30141 21143 30144
rect 21085 30135 21143 30141
rect 20438 30104 20444 30116
rect 18892 30076 20444 30104
rect 20438 30064 20444 30076
rect 20496 30064 20502 30116
rect 20916 30104 20944 30135
rect 21174 30132 21180 30144
rect 21232 30172 21238 30184
rect 21284 30172 21312 30280
rect 21361 30243 21419 30249
rect 21361 30209 21373 30243
rect 21407 30240 21419 30243
rect 21542 30240 21548 30252
rect 21407 30212 21548 30240
rect 21407 30209 21419 30212
rect 21361 30203 21419 30209
rect 21542 30200 21548 30212
rect 21600 30200 21606 30252
rect 21652 30240 21680 30280
rect 29380 30252 29408 30280
rect 21652 30212 24348 30240
rect 24320 30184 24348 30212
rect 25958 30200 25964 30252
rect 26016 30240 26022 30252
rect 27522 30240 27528 30252
rect 26016 30212 27528 30240
rect 26016 30200 26022 30212
rect 27522 30200 27528 30212
rect 27580 30200 27586 30252
rect 27709 30243 27767 30249
rect 27709 30209 27721 30243
rect 27755 30240 27767 30243
rect 29362 30240 29368 30252
rect 27755 30212 29368 30240
rect 27755 30209 27767 30212
rect 27709 30203 27767 30209
rect 29362 30200 29368 30212
rect 29420 30200 29426 30252
rect 29454 30200 29460 30252
rect 29512 30200 29518 30252
rect 29638 30249 29644 30252
rect 29605 30243 29644 30249
rect 29605 30209 29617 30243
rect 29605 30203 29644 30209
rect 29638 30200 29644 30203
rect 29696 30200 29702 30252
rect 29840 30249 29868 30280
rect 32508 30280 32996 30308
rect 32508 30252 32536 30280
rect 29733 30243 29791 30249
rect 29733 30209 29745 30243
rect 29779 30209 29791 30243
rect 29733 30203 29791 30209
rect 29825 30243 29883 30249
rect 29825 30209 29837 30243
rect 29871 30209 29883 30243
rect 29825 30203 29883 30209
rect 29922 30243 29980 30249
rect 29922 30209 29934 30243
rect 29968 30240 29980 30243
rect 29968 30212 30328 30240
rect 29968 30209 29980 30212
rect 29922 30203 29980 30209
rect 21232 30144 21312 30172
rect 21637 30175 21695 30181
rect 21232 30132 21238 30144
rect 21637 30141 21649 30175
rect 21683 30172 21695 30175
rect 21910 30172 21916 30184
rect 21683 30144 21916 30172
rect 21683 30141 21695 30144
rect 21637 30135 21695 30141
rect 21910 30132 21916 30144
rect 21968 30132 21974 30184
rect 24302 30132 24308 30184
rect 24360 30132 24366 30184
rect 27985 30175 28043 30181
rect 27985 30141 27997 30175
rect 28031 30172 28043 30175
rect 28258 30172 28264 30184
rect 28031 30144 28264 30172
rect 28031 30141 28043 30144
rect 27985 30135 28043 30141
rect 28258 30132 28264 30144
rect 28316 30132 28322 30184
rect 21450 30104 21456 30116
rect 20732 30076 21456 30104
rect 5074 29996 5080 30048
rect 5132 30036 5138 30048
rect 6178 30036 6184 30048
rect 5132 30008 6184 30036
rect 5132 29996 5138 30008
rect 6178 29996 6184 30008
rect 6236 29996 6242 30048
rect 6454 29996 6460 30048
rect 6512 30036 6518 30048
rect 9953 30039 10011 30045
rect 9953 30036 9965 30039
rect 6512 30008 9965 30036
rect 6512 29996 6518 30008
rect 9953 30005 9965 30008
rect 9999 30005 10011 30039
rect 9953 29999 10011 30005
rect 11238 29996 11244 30048
rect 11296 30036 11302 30048
rect 13814 30036 13820 30048
rect 11296 30008 13820 30036
rect 11296 29996 11302 30008
rect 13814 29996 13820 30008
rect 13872 29996 13878 30048
rect 13906 29996 13912 30048
rect 13964 30036 13970 30048
rect 14826 30036 14832 30048
rect 13964 30008 14832 30036
rect 13964 29996 13970 30008
rect 14826 29996 14832 30008
rect 14884 29996 14890 30048
rect 18046 29996 18052 30048
rect 18104 29996 18110 30048
rect 20165 30039 20223 30045
rect 20165 30005 20177 30039
rect 20211 30036 20223 30039
rect 20732 30036 20760 30076
rect 21450 30064 21456 30076
rect 21508 30064 21514 30116
rect 21545 30107 21603 30113
rect 21545 30073 21557 30107
rect 21591 30073 21603 30107
rect 21545 30067 21603 30073
rect 20211 30008 20760 30036
rect 20211 30005 20223 30008
rect 20165 29999 20223 30005
rect 20806 29996 20812 30048
rect 20864 30036 20870 30048
rect 21560 30036 21588 30067
rect 21818 30064 21824 30116
rect 21876 30104 21882 30116
rect 26510 30104 26516 30116
rect 21876 30076 26516 30104
rect 21876 30064 21882 30076
rect 26510 30064 26516 30076
rect 26568 30104 26574 30116
rect 27893 30107 27951 30113
rect 27893 30104 27905 30107
rect 26568 30076 27905 30104
rect 26568 30064 26574 30076
rect 27893 30073 27905 30076
rect 27939 30073 27951 30107
rect 27893 30067 27951 30073
rect 28442 30064 28448 30116
rect 28500 30104 28506 30116
rect 29748 30104 29776 30203
rect 30300 30184 30328 30212
rect 31754 30200 31760 30252
rect 31812 30240 31818 30252
rect 32217 30243 32275 30249
rect 32217 30240 32229 30243
rect 31812 30212 32229 30240
rect 31812 30200 31818 30212
rect 32217 30209 32229 30212
rect 32263 30209 32275 30243
rect 32217 30203 32275 30209
rect 32401 30246 32459 30249
rect 32490 30246 32496 30252
rect 32401 30243 32496 30246
rect 32401 30209 32413 30243
rect 32447 30218 32496 30243
rect 32447 30209 32459 30218
rect 32401 30203 32459 30209
rect 32490 30200 32496 30218
rect 32548 30200 32554 30252
rect 32858 30200 32864 30252
rect 32916 30200 32922 30252
rect 32968 30249 32996 30280
rect 34624 30280 35664 30308
rect 35728 30280 36308 30308
rect 36372 30280 37320 30308
rect 32953 30243 33011 30249
rect 32953 30209 32965 30243
rect 32999 30209 33011 30243
rect 32953 30203 33011 30209
rect 30282 30132 30288 30184
rect 30340 30132 30346 30184
rect 31570 30132 31576 30184
rect 31628 30172 31634 30184
rect 32582 30172 32588 30184
rect 31628 30144 32588 30172
rect 31628 30132 31634 30144
rect 32582 30132 32588 30144
rect 32640 30172 32646 30184
rect 34624 30172 34652 30280
rect 35360 30249 35388 30280
rect 35728 30249 35756 30280
rect 36280 30252 36308 30280
rect 35253 30243 35311 30249
rect 35253 30209 35265 30243
rect 35299 30209 35311 30243
rect 35253 30203 35311 30209
rect 35345 30243 35403 30249
rect 35345 30209 35357 30243
rect 35391 30209 35403 30243
rect 35345 30203 35403 30209
rect 35713 30243 35771 30249
rect 35713 30209 35725 30243
rect 35759 30209 35771 30243
rect 35713 30203 35771 30209
rect 35805 30243 35863 30249
rect 35805 30209 35817 30243
rect 35851 30209 35863 30243
rect 36081 30243 36139 30249
rect 36081 30240 36093 30243
rect 35805 30203 35863 30209
rect 36004 30212 36093 30240
rect 32640 30144 34652 30172
rect 32640 30132 32646 30144
rect 34790 30132 34796 30184
rect 34848 30172 34854 30184
rect 35268 30172 35296 30203
rect 35728 30172 35756 30203
rect 34848 30144 35756 30172
rect 34848 30132 34854 30144
rect 33410 30104 33416 30116
rect 28500 30076 33416 30104
rect 28500 30064 28506 30076
rect 33410 30064 33416 30076
rect 33468 30064 33474 30116
rect 34606 30064 34612 30116
rect 34664 30104 34670 30116
rect 35437 30107 35495 30113
rect 35437 30104 35449 30107
rect 34664 30076 35449 30104
rect 34664 30064 34670 30076
rect 35437 30073 35449 30076
rect 35483 30073 35495 30107
rect 35437 30067 35495 30073
rect 35820 30048 35848 30203
rect 35894 30132 35900 30184
rect 35952 30132 35958 30184
rect 36004 30048 36032 30212
rect 36081 30209 36093 30212
rect 36127 30209 36139 30243
rect 36081 30203 36139 30209
rect 36262 30200 36268 30252
rect 36320 30200 36326 30252
rect 36354 30200 36360 30252
rect 36412 30200 36418 30252
rect 36170 30064 36176 30116
rect 36228 30104 36234 30116
rect 36357 30107 36415 30113
rect 36357 30104 36369 30107
rect 36228 30076 36369 30104
rect 36228 30064 36234 30076
rect 36357 30073 36369 30076
rect 36403 30073 36415 30107
rect 37292 30104 37320 30280
rect 37369 30277 37381 30311
rect 37415 30308 37427 30311
rect 38470 30308 38476 30320
rect 37415 30280 38476 30308
rect 37415 30277 37427 30280
rect 37369 30271 37427 30277
rect 38470 30268 38476 30280
rect 38528 30268 38534 30320
rect 38580 30249 38608 30336
rect 40034 30268 40040 30320
rect 40092 30268 40098 30320
rect 37921 30243 37979 30249
rect 37921 30209 37933 30243
rect 37967 30209 37979 30243
rect 37921 30203 37979 30209
rect 38565 30243 38623 30249
rect 38565 30209 38577 30243
rect 38611 30209 38623 30243
rect 38565 30203 38623 30209
rect 37550 30104 37556 30116
rect 37292 30076 37556 30104
rect 36357 30067 36415 30073
rect 37550 30064 37556 30076
rect 37608 30064 37614 30116
rect 37936 30104 37964 30203
rect 38746 30200 38752 30252
rect 38804 30240 38810 30252
rect 38933 30243 38991 30249
rect 38933 30240 38945 30243
rect 38804 30212 38945 30240
rect 38804 30200 38810 30212
rect 38933 30209 38945 30212
rect 38979 30209 38991 30243
rect 38933 30203 38991 30209
rect 38473 30175 38531 30181
rect 38473 30141 38485 30175
rect 38519 30172 38531 30175
rect 38519 30144 38976 30172
rect 38519 30141 38531 30144
rect 38473 30135 38531 30141
rect 38948 30116 38976 30144
rect 39022 30132 39028 30184
rect 39080 30172 39086 30184
rect 39301 30175 39359 30181
rect 39301 30172 39313 30175
rect 39080 30144 39313 30172
rect 39080 30132 39086 30144
rect 39301 30141 39313 30144
rect 39347 30141 39359 30175
rect 39301 30135 39359 30141
rect 39574 30132 39580 30184
rect 39632 30132 39638 30184
rect 38654 30104 38660 30116
rect 37936 30076 38660 30104
rect 38654 30064 38660 30076
rect 38712 30064 38718 30116
rect 38930 30064 38936 30116
rect 38988 30104 38994 30116
rect 38988 30076 39252 30104
rect 38988 30064 38994 30076
rect 21634 30036 21640 30048
rect 20864 30008 21640 30036
rect 20864 29996 20870 30008
rect 21634 29996 21640 30008
rect 21692 29996 21698 30048
rect 24762 29996 24768 30048
rect 24820 30036 24826 30048
rect 30006 30036 30012 30048
rect 24820 30008 30012 30036
rect 24820 29996 24826 30008
rect 30006 29996 30012 30008
rect 30064 29996 30070 30048
rect 32214 29996 32220 30048
rect 32272 29996 32278 30048
rect 32766 29996 32772 30048
rect 32824 30036 32830 30048
rect 33870 30036 33876 30048
rect 32824 30008 33876 30036
rect 32824 29996 32830 30008
rect 33870 29996 33876 30008
rect 33928 30036 33934 30048
rect 34698 30036 34704 30048
rect 33928 30008 34704 30036
rect 33928 29996 33934 30008
rect 34698 29996 34704 30008
rect 34756 29996 34762 30048
rect 35802 29996 35808 30048
rect 35860 29996 35866 30048
rect 35986 29996 35992 30048
rect 36044 29996 36050 30048
rect 36630 29996 36636 30048
rect 36688 30036 36694 30048
rect 38010 30036 38016 30048
rect 36688 30008 38016 30036
rect 36688 29996 36694 30008
rect 38010 29996 38016 30008
rect 38068 29996 38074 30048
rect 38838 29996 38844 30048
rect 38896 29996 38902 30048
rect 39114 29996 39120 30048
rect 39172 29996 39178 30048
rect 39224 30036 39252 30076
rect 41049 30039 41107 30045
rect 41049 30036 41061 30039
rect 39224 30008 41061 30036
rect 41049 30005 41061 30008
rect 41095 30005 41107 30039
rect 41049 29999 41107 30005
rect 1104 29946 41400 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 41400 29946
rect 1104 29872 41400 29894
rect 2866 29792 2872 29844
rect 2924 29832 2930 29844
rect 5258 29832 5264 29844
rect 2924 29804 5264 29832
rect 2924 29792 2930 29804
rect 5258 29792 5264 29804
rect 5316 29832 5322 29844
rect 5997 29835 6055 29841
rect 5997 29832 6009 29835
rect 5316 29804 6009 29832
rect 5316 29792 5322 29804
rect 5997 29801 6009 29804
rect 6043 29801 6055 29835
rect 5997 29795 6055 29801
rect 6730 29792 6736 29844
rect 6788 29792 6794 29844
rect 7374 29792 7380 29844
rect 7432 29832 7438 29844
rect 7837 29835 7895 29841
rect 7837 29832 7849 29835
rect 7432 29804 7849 29832
rect 7432 29792 7438 29804
rect 7837 29801 7849 29804
rect 7883 29801 7895 29835
rect 7837 29795 7895 29801
rect 7926 29792 7932 29844
rect 7984 29832 7990 29844
rect 8662 29832 8668 29844
rect 7984 29804 8668 29832
rect 7984 29792 7990 29804
rect 8662 29792 8668 29804
rect 8720 29792 8726 29844
rect 9784 29804 12848 29832
rect 4982 29724 4988 29776
rect 5040 29764 5046 29776
rect 5077 29767 5135 29773
rect 5077 29764 5089 29767
rect 5040 29736 5089 29764
rect 5040 29724 5046 29736
rect 5077 29733 5089 29736
rect 5123 29733 5135 29767
rect 5077 29727 5135 29733
rect 5184 29736 6592 29764
rect 2682 29588 2688 29640
rect 2740 29588 2746 29640
rect 4154 29520 4160 29572
rect 4212 29560 4218 29572
rect 4798 29560 4804 29572
rect 4212 29532 4804 29560
rect 4212 29520 4218 29532
rect 4798 29520 4804 29532
rect 4856 29520 4862 29572
rect 5184 29560 5212 29736
rect 5261 29699 5319 29705
rect 5261 29665 5273 29699
rect 5307 29696 5319 29699
rect 6564 29696 6592 29736
rect 7006 29724 7012 29776
rect 7064 29764 7070 29776
rect 9674 29764 9680 29776
rect 7064 29736 9680 29764
rect 7064 29724 7070 29736
rect 9674 29724 9680 29736
rect 9732 29724 9738 29776
rect 6730 29696 6736 29708
rect 5307 29668 6132 29696
rect 6564 29668 6736 29696
rect 5307 29665 5319 29668
rect 5261 29659 5319 29665
rect 5350 29588 5356 29640
rect 5408 29588 5414 29640
rect 5446 29631 5504 29637
rect 5446 29597 5458 29631
rect 5492 29597 5504 29631
rect 5721 29631 5779 29637
rect 5721 29628 5733 29631
rect 5446 29591 5504 29597
rect 5552 29600 5733 29628
rect 5460 29560 5488 29591
rect 5184 29532 5488 29560
rect 5460 29504 5488 29532
rect 2498 29452 2504 29504
rect 2556 29452 2562 29504
rect 5442 29452 5448 29504
rect 5500 29452 5506 29504
rect 5552 29492 5580 29600
rect 5721 29597 5733 29600
rect 5767 29597 5779 29631
rect 5721 29591 5779 29597
rect 5810 29588 5816 29640
rect 5868 29637 5874 29640
rect 6104 29637 6132 29668
rect 6730 29656 6736 29668
rect 6788 29656 6794 29708
rect 8202 29696 8208 29708
rect 8036 29668 8208 29696
rect 5868 29628 5876 29637
rect 6089 29631 6147 29637
rect 5868 29600 5913 29628
rect 5868 29591 5876 29600
rect 6089 29597 6101 29631
rect 6135 29597 6147 29631
rect 6089 29591 6147 29597
rect 5868 29588 5874 29591
rect 6178 29588 6184 29640
rect 6236 29588 6242 29640
rect 6454 29588 6460 29640
rect 6512 29588 6518 29640
rect 6595 29631 6653 29637
rect 6595 29597 6607 29631
rect 6641 29628 6653 29631
rect 7098 29628 7104 29640
rect 6641 29600 7104 29628
rect 6641 29597 6653 29600
rect 6595 29591 6653 29597
rect 7098 29588 7104 29600
rect 7156 29588 7162 29640
rect 7190 29588 7196 29640
rect 7248 29588 7254 29640
rect 7374 29637 7380 29640
rect 7341 29631 7380 29637
rect 7341 29597 7353 29631
rect 7341 29591 7380 29597
rect 7374 29588 7380 29591
rect 7432 29588 7438 29640
rect 7742 29637 7748 29640
rect 7699 29631 7748 29637
rect 7699 29597 7711 29631
rect 7745 29597 7748 29631
rect 7699 29591 7748 29597
rect 7742 29588 7748 29591
rect 7800 29588 7806 29640
rect 7926 29588 7932 29640
rect 7984 29628 7990 29640
rect 8036 29637 8064 29668
rect 8202 29656 8208 29668
rect 8260 29696 8266 29708
rect 9306 29696 9312 29708
rect 8260 29668 9312 29696
rect 8260 29656 8266 29668
rect 9306 29656 9312 29668
rect 9364 29696 9370 29708
rect 9784 29696 9812 29804
rect 12820 29776 12848 29804
rect 13814 29792 13820 29844
rect 13872 29792 13878 29844
rect 14366 29792 14372 29844
rect 14424 29832 14430 29844
rect 14737 29835 14795 29841
rect 14737 29832 14749 29835
rect 14424 29804 14749 29832
rect 14424 29792 14430 29804
rect 14737 29801 14749 29804
rect 14783 29801 14795 29835
rect 14737 29795 14795 29801
rect 15010 29792 15016 29844
rect 15068 29832 15074 29844
rect 17037 29835 17095 29841
rect 17037 29832 17049 29835
rect 15068 29804 17049 29832
rect 15068 29792 15074 29804
rect 17037 29801 17049 29804
rect 17083 29801 17095 29835
rect 17037 29795 17095 29801
rect 18506 29792 18512 29844
rect 18564 29832 18570 29844
rect 22186 29832 22192 29844
rect 18564 29804 22192 29832
rect 18564 29792 18570 29804
rect 22186 29792 22192 29804
rect 22244 29792 22250 29844
rect 22462 29792 22468 29844
rect 22520 29792 22526 29844
rect 24394 29792 24400 29844
rect 24452 29832 24458 29844
rect 24578 29832 24584 29844
rect 24452 29804 24584 29832
rect 24452 29792 24458 29804
rect 24578 29792 24584 29804
rect 24636 29832 24642 29844
rect 25777 29835 25835 29841
rect 25777 29832 25789 29835
rect 24636 29804 25789 29832
rect 24636 29792 24642 29804
rect 25777 29801 25789 29804
rect 25823 29801 25835 29835
rect 25777 29795 25835 29801
rect 26050 29792 26056 29844
rect 26108 29832 26114 29844
rect 26145 29835 26203 29841
rect 26145 29832 26157 29835
rect 26108 29804 26157 29832
rect 26108 29792 26114 29804
rect 26145 29801 26157 29804
rect 26191 29801 26203 29835
rect 26145 29795 26203 29801
rect 26510 29792 26516 29844
rect 26568 29792 26574 29844
rect 27614 29792 27620 29844
rect 27672 29832 27678 29844
rect 29549 29835 29607 29841
rect 29549 29832 29561 29835
rect 27672 29804 29561 29832
rect 27672 29792 27678 29804
rect 29549 29801 29561 29804
rect 29595 29801 29607 29835
rect 30558 29832 30564 29844
rect 29549 29795 29607 29801
rect 29656 29804 30564 29832
rect 11532 29736 12756 29764
rect 11532 29708 11560 29736
rect 9364 29668 9812 29696
rect 9364 29656 9370 29668
rect 8021 29631 8079 29637
rect 8021 29628 8033 29631
rect 7984 29600 8033 29628
rect 7984 29588 7990 29600
rect 8021 29597 8033 29600
rect 8067 29597 8079 29631
rect 8021 29591 8079 29597
rect 8110 29588 8116 29640
rect 8168 29628 8174 29640
rect 8570 29637 8576 29640
rect 8527 29631 8576 29637
rect 8168 29600 8213 29628
rect 8168 29588 8174 29600
rect 8527 29597 8539 29631
rect 8573 29597 8576 29631
rect 8527 29591 8576 29597
rect 8570 29588 8576 29591
rect 8628 29628 8634 29640
rect 8628 29600 9352 29628
rect 8628 29588 8634 29600
rect 5626 29520 5632 29572
rect 5684 29560 5690 29572
rect 6365 29563 6423 29569
rect 6365 29560 6377 29563
rect 5684 29532 6377 29560
rect 5684 29520 5690 29532
rect 6365 29529 6377 29532
rect 6411 29560 6423 29563
rect 7006 29560 7012 29572
rect 6411 29532 7012 29560
rect 6411 29529 6423 29532
rect 6365 29523 6423 29529
rect 7006 29520 7012 29532
rect 7064 29560 7070 29572
rect 7469 29563 7527 29569
rect 7469 29560 7481 29563
rect 7064 29532 7481 29560
rect 7064 29520 7070 29532
rect 7469 29529 7481 29532
rect 7515 29529 7527 29563
rect 7469 29523 7527 29529
rect 7561 29563 7619 29569
rect 7561 29529 7573 29563
rect 7607 29560 7619 29563
rect 7607 29532 7880 29560
rect 7607 29529 7619 29532
rect 7561 29523 7619 29529
rect 7852 29504 7880 29532
rect 8202 29520 8208 29572
rect 8260 29560 8266 29572
rect 8297 29563 8355 29569
rect 8297 29560 8309 29563
rect 8260 29532 8309 29560
rect 8260 29520 8266 29532
rect 8297 29529 8309 29532
rect 8343 29529 8355 29563
rect 8297 29523 8355 29529
rect 8389 29563 8447 29569
rect 8389 29529 8401 29563
rect 8435 29560 8447 29563
rect 9214 29560 9220 29572
rect 8435 29532 9220 29560
rect 8435 29529 8447 29532
rect 8389 29523 8447 29529
rect 9214 29520 9220 29532
rect 9272 29520 9278 29572
rect 6546 29492 6552 29504
rect 5552 29464 6552 29492
rect 6546 29452 6552 29464
rect 6604 29452 6610 29504
rect 7834 29452 7840 29504
rect 7892 29492 7898 29504
rect 8665 29495 8723 29501
rect 8665 29492 8677 29495
rect 7892 29464 8677 29492
rect 7892 29452 7898 29464
rect 8665 29461 8677 29464
rect 8711 29461 8723 29495
rect 9324 29492 9352 29600
rect 9398 29588 9404 29640
rect 9456 29588 9462 29640
rect 9508 29637 9536 29668
rect 11514 29656 11520 29708
rect 11572 29656 11578 29708
rect 12728 29696 12756 29736
rect 12802 29724 12808 29776
rect 12860 29764 12866 29776
rect 15841 29767 15899 29773
rect 15841 29764 15853 29767
rect 12860 29736 15853 29764
rect 12860 29724 12866 29736
rect 15841 29733 15853 29736
rect 15887 29733 15899 29767
rect 15841 29727 15899 29733
rect 16390 29724 16396 29776
rect 16448 29764 16454 29776
rect 21634 29764 21640 29776
rect 16448 29736 21640 29764
rect 16448 29724 16454 29736
rect 21634 29724 21640 29736
rect 21692 29724 21698 29776
rect 26326 29764 26332 29776
rect 25792 29736 26332 29764
rect 12728 29668 14320 29696
rect 9493 29631 9551 29637
rect 9493 29597 9505 29631
rect 9539 29597 9551 29631
rect 9493 29591 9551 29597
rect 9582 29588 9588 29640
rect 9640 29588 9646 29640
rect 9950 29628 9956 29640
rect 9692 29600 9956 29628
rect 9416 29560 9444 29588
rect 9600 29560 9628 29588
rect 9416 29532 9628 29560
rect 9692 29492 9720 29600
rect 9950 29588 9956 29600
rect 10008 29637 10014 29640
rect 10008 29631 10057 29637
rect 10008 29597 10011 29631
rect 10045 29628 10057 29631
rect 11974 29628 11980 29640
rect 10045 29600 11980 29628
rect 10045 29597 10057 29600
rect 10008 29591 10057 29597
rect 10008 29588 10014 29591
rect 11974 29588 11980 29600
rect 12032 29588 12038 29640
rect 12250 29588 12256 29640
rect 12308 29588 12314 29640
rect 13170 29588 13176 29640
rect 13228 29588 13234 29640
rect 13262 29588 13268 29640
rect 13320 29628 13326 29640
rect 13464 29637 13492 29668
rect 13449 29631 13507 29637
rect 13320 29600 13365 29628
rect 13320 29588 13326 29600
rect 13449 29597 13461 29631
rect 13495 29597 13507 29631
rect 13449 29591 13507 29597
rect 13638 29631 13696 29637
rect 13638 29597 13650 29631
rect 13684 29597 13696 29631
rect 13638 29591 13696 29597
rect 9766 29520 9772 29572
rect 9824 29520 9830 29572
rect 9858 29520 9864 29572
rect 9916 29520 9922 29572
rect 11698 29560 11704 29572
rect 9968 29532 11704 29560
rect 9324 29464 9720 29492
rect 9784 29492 9812 29520
rect 9968 29492 9996 29532
rect 11698 29520 11704 29532
rect 11756 29520 11762 29572
rect 11882 29520 11888 29572
rect 11940 29560 11946 29572
rect 12437 29563 12495 29569
rect 12437 29560 12449 29563
rect 11940 29532 12449 29560
rect 11940 29520 11946 29532
rect 12437 29529 12449 29532
rect 12483 29529 12495 29563
rect 12437 29523 12495 29529
rect 13354 29520 13360 29572
rect 13412 29560 13418 29572
rect 13541 29563 13599 29569
rect 13541 29560 13553 29563
rect 13412 29532 13553 29560
rect 13412 29520 13418 29532
rect 13541 29529 13553 29532
rect 13587 29529 13599 29563
rect 13541 29523 13599 29529
rect 13653 29560 13681 29591
rect 13906 29588 13912 29640
rect 13964 29588 13970 29640
rect 14090 29588 14096 29640
rect 14148 29588 14154 29640
rect 14186 29631 14244 29637
rect 14186 29597 14198 29631
rect 14232 29597 14244 29631
rect 14292 29628 14320 29668
rect 14366 29656 14372 29708
rect 14424 29696 14430 29708
rect 14424 29668 15240 29696
rect 14424 29656 14430 29668
rect 14599 29631 14657 29637
rect 14292 29600 14412 29628
rect 14186 29591 14244 29597
rect 13924 29560 13952 29588
rect 13653 29532 13952 29560
rect 14201 29560 14229 29591
rect 14384 29569 14412 29600
rect 14599 29597 14611 29631
rect 14645 29628 14657 29631
rect 14826 29628 14832 29640
rect 14645 29600 14832 29628
rect 14645 29597 14657 29600
rect 14599 29591 14657 29597
rect 14826 29588 14832 29600
rect 14884 29588 14890 29640
rect 14921 29631 14979 29637
rect 14921 29597 14933 29631
rect 14967 29628 14979 29631
rect 15010 29628 15016 29640
rect 14967 29600 15016 29628
rect 14967 29597 14979 29600
rect 14921 29591 14979 29597
rect 15010 29588 15016 29600
rect 15068 29588 15074 29640
rect 15212 29637 15240 29668
rect 20806 29656 20812 29708
rect 20864 29696 20870 29708
rect 21082 29696 21088 29708
rect 20864 29668 21088 29696
rect 20864 29656 20870 29668
rect 21082 29656 21088 29668
rect 21140 29656 21146 29708
rect 21726 29656 21732 29708
rect 21784 29696 21790 29708
rect 22370 29696 22376 29708
rect 21784 29668 22376 29696
rect 21784 29656 21790 29668
rect 22370 29656 22376 29668
rect 22428 29656 22434 29708
rect 23014 29656 23020 29708
rect 23072 29696 23078 29708
rect 23753 29699 23811 29705
rect 23072 29668 23612 29696
rect 23072 29656 23078 29668
rect 15197 29631 15255 29637
rect 15197 29597 15209 29631
rect 15243 29597 15255 29631
rect 15197 29591 15255 29597
rect 15289 29631 15347 29637
rect 15289 29597 15301 29631
rect 15335 29597 15347 29631
rect 15289 29591 15347 29597
rect 17773 29631 17831 29637
rect 17773 29597 17785 29631
rect 17819 29628 17831 29631
rect 18138 29628 18144 29640
rect 17819 29600 18144 29628
rect 17819 29597 17831 29600
rect 17773 29591 17831 29597
rect 14369 29563 14427 29569
rect 14201 29532 14320 29560
rect 9784 29464 9996 29492
rect 8665 29455 8723 29461
rect 10042 29452 10048 29504
rect 10100 29492 10106 29504
rect 10137 29495 10195 29501
rect 10137 29492 10149 29495
rect 10100 29464 10149 29492
rect 10100 29452 10106 29464
rect 10137 29461 10149 29464
rect 10183 29461 10195 29495
rect 10137 29455 10195 29461
rect 12342 29452 12348 29504
rect 12400 29492 12406 29504
rect 12621 29495 12679 29501
rect 12621 29492 12633 29495
rect 12400 29464 12633 29492
rect 12400 29452 12406 29464
rect 12621 29461 12633 29464
rect 12667 29461 12679 29495
rect 12621 29455 12679 29461
rect 12710 29452 12716 29504
rect 12768 29492 12774 29504
rect 13653 29492 13681 29532
rect 12768 29464 13681 29492
rect 14292 29492 14320 29532
rect 14369 29529 14381 29563
rect 14415 29529 14427 29563
rect 14369 29523 14427 29529
rect 14461 29563 14519 29569
rect 14461 29529 14473 29563
rect 14507 29560 14519 29563
rect 15102 29560 15108 29572
rect 14507 29532 15108 29560
rect 14507 29529 14519 29532
rect 14461 29523 14519 29529
rect 15102 29520 15108 29532
rect 15160 29520 15166 29572
rect 14642 29492 14648 29504
rect 14292 29464 14648 29492
rect 12768 29452 12774 29464
rect 14642 29452 14648 29464
rect 14700 29492 14706 29504
rect 15304 29492 15332 29591
rect 18138 29588 18144 29600
rect 18196 29628 18202 29640
rect 18196 29600 22784 29628
rect 18196 29588 18202 29600
rect 22756 29572 22784 29600
rect 23198 29588 23204 29640
rect 23256 29588 23262 29640
rect 23382 29588 23388 29640
rect 23440 29628 23446 29640
rect 23584 29637 23612 29668
rect 23753 29665 23765 29699
rect 23799 29696 23811 29699
rect 23842 29696 23848 29708
rect 23799 29668 23848 29696
rect 23799 29665 23811 29668
rect 23753 29659 23811 29665
rect 23842 29656 23848 29668
rect 23900 29656 23906 29708
rect 23477 29631 23535 29637
rect 23477 29628 23489 29631
rect 23440 29600 23489 29628
rect 23440 29588 23446 29600
rect 23477 29597 23489 29600
rect 23523 29597 23535 29631
rect 23477 29591 23535 29597
rect 23569 29631 23627 29637
rect 23569 29597 23581 29631
rect 23615 29628 23627 29631
rect 23615 29600 24348 29628
rect 23615 29597 23627 29600
rect 23569 29591 23627 29597
rect 24320 29572 24348 29600
rect 24670 29588 24676 29640
rect 24728 29588 24734 29640
rect 25792 29637 25820 29736
rect 26326 29724 26332 29736
rect 26384 29764 26390 29776
rect 26697 29767 26755 29773
rect 26697 29764 26709 29767
rect 26384 29736 26709 29764
rect 26384 29724 26390 29736
rect 26697 29733 26709 29736
rect 26743 29733 26755 29767
rect 29656 29764 29684 29804
rect 30558 29792 30564 29804
rect 30616 29792 30622 29844
rect 31570 29792 31576 29844
rect 31628 29792 31634 29844
rect 33134 29792 33140 29844
rect 33192 29832 33198 29844
rect 33321 29835 33379 29841
rect 33321 29832 33333 29835
rect 33192 29804 33333 29832
rect 33192 29792 33198 29804
rect 33321 29801 33333 29804
rect 33367 29832 33379 29835
rect 34974 29832 34980 29844
rect 33367 29804 34980 29832
rect 33367 29801 33379 29804
rect 33321 29795 33379 29801
rect 34974 29792 34980 29804
rect 35032 29792 35038 29844
rect 35802 29792 35808 29844
rect 35860 29832 35866 29844
rect 36630 29832 36636 29844
rect 35860 29804 36636 29832
rect 35860 29792 35866 29804
rect 36630 29792 36636 29804
rect 36688 29792 36694 29844
rect 37458 29792 37464 29844
rect 37516 29832 37522 29844
rect 38194 29832 38200 29844
rect 37516 29804 38200 29832
rect 37516 29792 37522 29804
rect 38194 29792 38200 29804
rect 38252 29792 38258 29844
rect 38841 29835 38899 29841
rect 38841 29801 38853 29835
rect 38887 29832 38899 29835
rect 38930 29832 38936 29844
rect 38887 29804 38936 29832
rect 38887 29801 38899 29804
rect 38841 29795 38899 29801
rect 38930 29792 38936 29804
rect 38988 29792 38994 29844
rect 39574 29792 39580 29844
rect 39632 29832 39638 29844
rect 39853 29835 39911 29841
rect 39853 29832 39865 29835
rect 39632 29804 39865 29832
rect 39632 29792 39638 29804
rect 39853 29801 39865 29804
rect 39899 29801 39911 29835
rect 39853 29795 39911 29801
rect 26697 29727 26755 29733
rect 29104 29736 29684 29764
rect 26510 29696 26516 29708
rect 25884 29668 26516 29696
rect 25777 29631 25835 29637
rect 25777 29597 25789 29631
rect 25823 29597 25835 29631
rect 25777 29591 25835 29597
rect 15562 29520 15568 29572
rect 15620 29560 15626 29572
rect 15657 29563 15715 29569
rect 15657 29560 15669 29563
rect 15620 29532 15669 29560
rect 15620 29520 15626 29532
rect 15657 29529 15669 29532
rect 15703 29529 15715 29563
rect 15657 29523 15715 29529
rect 16942 29520 16948 29572
rect 17000 29520 17006 29572
rect 17957 29563 18015 29569
rect 17957 29529 17969 29563
rect 18003 29560 18015 29563
rect 18230 29560 18236 29572
rect 18003 29532 18236 29560
rect 18003 29529 18015 29532
rect 17957 29523 18015 29529
rect 18230 29520 18236 29532
rect 18288 29520 18294 29572
rect 22186 29520 22192 29572
rect 22244 29560 22250 29572
rect 22281 29563 22339 29569
rect 22281 29560 22293 29563
rect 22244 29532 22293 29560
rect 22244 29520 22250 29532
rect 22281 29529 22293 29532
rect 22327 29529 22339 29563
rect 22281 29523 22339 29529
rect 22738 29520 22744 29572
rect 22796 29560 22802 29572
rect 22796 29532 23888 29560
rect 22796 29520 22802 29532
rect 14700 29464 15332 29492
rect 14700 29452 14706 29464
rect 15470 29452 15476 29504
rect 15528 29452 15534 29504
rect 17678 29452 17684 29504
rect 17736 29492 17742 29504
rect 18141 29495 18199 29501
rect 18141 29492 18153 29495
rect 17736 29464 18153 29492
rect 17736 29452 17742 29464
rect 18141 29461 18153 29464
rect 18187 29461 18199 29495
rect 18141 29455 18199 29461
rect 21082 29452 21088 29504
rect 21140 29492 21146 29504
rect 21818 29492 21824 29504
rect 21140 29464 21824 29492
rect 21140 29452 21146 29464
rect 21818 29452 21824 29464
rect 21876 29452 21882 29504
rect 22462 29452 22468 29504
rect 22520 29452 22526 29504
rect 22646 29452 22652 29504
rect 22704 29452 22710 29504
rect 23198 29452 23204 29504
rect 23256 29492 23262 29504
rect 23385 29495 23443 29501
rect 23385 29492 23397 29495
rect 23256 29464 23397 29492
rect 23256 29452 23262 29464
rect 23385 29461 23397 29464
rect 23431 29461 23443 29495
rect 23385 29455 23443 29461
rect 23658 29452 23664 29504
rect 23716 29492 23722 29504
rect 23753 29495 23811 29501
rect 23753 29492 23765 29495
rect 23716 29464 23765 29492
rect 23716 29452 23722 29464
rect 23753 29461 23765 29464
rect 23799 29461 23811 29495
rect 23860 29492 23888 29532
rect 24302 29520 24308 29572
rect 24360 29520 24366 29572
rect 24688 29560 24716 29588
rect 25884 29560 25912 29668
rect 26510 29656 26516 29668
rect 26568 29696 26574 29708
rect 26605 29699 26663 29705
rect 26605 29696 26617 29699
rect 26568 29668 26617 29696
rect 26568 29656 26574 29668
rect 26605 29665 26617 29668
rect 26651 29665 26663 29699
rect 28626 29696 28632 29708
rect 26605 29659 26663 29665
rect 26712 29668 28632 29696
rect 25961 29631 26019 29637
rect 25961 29597 25973 29631
rect 26007 29628 26019 29631
rect 26329 29631 26387 29637
rect 26007 29600 26280 29628
rect 26007 29597 26019 29600
rect 25961 29591 26019 29597
rect 24688 29532 25912 29560
rect 26252 29560 26280 29600
rect 26329 29597 26341 29631
rect 26375 29628 26387 29631
rect 26418 29628 26424 29640
rect 26375 29600 26424 29628
rect 26375 29597 26387 29600
rect 26329 29591 26387 29597
rect 26418 29588 26424 29600
rect 26476 29588 26482 29640
rect 26712 29637 26740 29668
rect 28626 29656 28632 29668
rect 28684 29656 28690 29708
rect 26697 29631 26755 29637
rect 26697 29597 26709 29631
rect 26743 29597 26755 29631
rect 26697 29591 26755 29597
rect 26786 29588 26792 29640
rect 26844 29588 26850 29640
rect 26881 29631 26939 29637
rect 26881 29597 26893 29631
rect 26927 29628 26939 29631
rect 29104 29628 29132 29736
rect 29730 29724 29736 29776
rect 29788 29764 29794 29776
rect 30282 29764 30288 29776
rect 29788 29736 30288 29764
rect 29788 29724 29794 29736
rect 30282 29724 30288 29736
rect 30340 29764 30346 29776
rect 30929 29767 30987 29773
rect 30929 29764 30941 29767
rect 30340 29736 30941 29764
rect 30340 29724 30346 29736
rect 30929 29733 30941 29736
rect 30975 29764 30987 29767
rect 31389 29767 31447 29773
rect 31389 29764 31401 29767
rect 30975 29736 31401 29764
rect 30975 29733 30987 29736
rect 30929 29727 30987 29733
rect 31389 29733 31401 29736
rect 31435 29733 31447 29767
rect 31389 29727 31447 29733
rect 29273 29699 29331 29705
rect 29273 29665 29285 29699
rect 29319 29696 29331 29699
rect 29319 29668 29868 29696
rect 29319 29665 29331 29668
rect 29273 29659 29331 29665
rect 26927 29600 29132 29628
rect 29181 29631 29239 29637
rect 26927 29597 26939 29600
rect 26881 29591 26939 29597
rect 26804 29560 26832 29588
rect 26252 29532 26832 29560
rect 27816 29504 27844 29600
rect 29181 29597 29193 29631
rect 29227 29597 29239 29631
rect 29181 29591 29239 29597
rect 29196 29560 29224 29591
rect 29362 29588 29368 29640
rect 29420 29588 29426 29640
rect 29454 29588 29460 29640
rect 29512 29588 29518 29640
rect 29840 29637 29868 29668
rect 30006 29656 30012 29708
rect 30064 29696 30070 29708
rect 30193 29699 30251 29705
rect 30193 29696 30205 29699
rect 30064 29668 30205 29696
rect 30064 29656 30070 29668
rect 30193 29665 30205 29668
rect 30239 29665 30251 29699
rect 30193 29659 30251 29665
rect 29733 29631 29791 29637
rect 29733 29597 29745 29631
rect 29779 29597 29791 29631
rect 29733 29591 29791 29597
rect 29825 29631 29883 29637
rect 29825 29597 29837 29631
rect 29871 29597 29883 29631
rect 29825 29591 29883 29597
rect 29472 29560 29500 29588
rect 29196 29532 29500 29560
rect 29748 29560 29776 29591
rect 30282 29588 30288 29640
rect 30340 29588 30346 29640
rect 30374 29588 30380 29640
rect 30432 29628 30438 29640
rect 30745 29631 30803 29637
rect 30745 29628 30757 29631
rect 30432 29600 30757 29628
rect 30432 29588 30438 29600
rect 30745 29597 30757 29600
rect 30791 29597 30803 29631
rect 30745 29591 30803 29597
rect 30837 29631 30895 29637
rect 30837 29597 30849 29631
rect 30883 29628 30895 29631
rect 30926 29628 30932 29640
rect 30883 29600 30932 29628
rect 30883 29597 30895 29600
rect 30837 29591 30895 29597
rect 30926 29588 30932 29600
rect 30984 29588 30990 29640
rect 31018 29588 31024 29640
rect 31076 29588 31082 29640
rect 31588 29637 31616 29792
rect 31846 29724 31852 29776
rect 31904 29764 31910 29776
rect 32306 29764 32312 29776
rect 31904 29736 32312 29764
rect 31904 29724 31910 29736
rect 32306 29724 32312 29736
rect 32364 29724 32370 29776
rect 33413 29767 33471 29773
rect 33413 29733 33425 29767
rect 33459 29764 33471 29767
rect 33502 29764 33508 29776
rect 33459 29736 33508 29764
rect 33459 29733 33471 29736
rect 33413 29727 33471 29733
rect 33502 29724 33508 29736
rect 33560 29724 33566 29776
rect 34330 29724 34336 29776
rect 34388 29764 34394 29776
rect 38562 29764 38568 29776
rect 34388 29736 38568 29764
rect 34388 29724 34394 29736
rect 38562 29724 38568 29736
rect 38620 29764 38626 29776
rect 39393 29767 39451 29773
rect 39393 29764 39405 29767
rect 38620 29736 39405 29764
rect 38620 29724 38626 29736
rect 39393 29733 39405 29736
rect 39439 29733 39451 29767
rect 39393 29727 39451 29733
rect 32766 29656 32772 29708
rect 32824 29656 32830 29708
rect 35986 29696 35992 29708
rect 32876 29668 35992 29696
rect 31205 29631 31263 29637
rect 31205 29597 31217 29631
rect 31251 29597 31263 29631
rect 31205 29591 31263 29597
rect 31573 29631 31631 29637
rect 31573 29597 31585 29631
rect 31619 29597 31631 29631
rect 31573 29591 31631 29597
rect 30101 29563 30159 29569
rect 29748 29532 29868 29560
rect 29840 29504 29868 29532
rect 30101 29529 30113 29563
rect 30147 29529 30159 29563
rect 30300 29560 30328 29588
rect 31220 29560 31248 29591
rect 31662 29588 31668 29640
rect 31720 29588 31726 29640
rect 30300 29532 31248 29560
rect 31389 29563 31447 29569
rect 30101 29523 30159 29529
rect 31389 29529 31401 29563
rect 31435 29560 31447 29563
rect 32784 29560 32812 29656
rect 32876 29640 32904 29668
rect 32858 29588 32864 29640
rect 32916 29588 32922 29640
rect 32953 29631 33011 29637
rect 32953 29597 32965 29631
rect 32999 29597 33011 29631
rect 32953 29591 33011 29597
rect 33045 29631 33103 29637
rect 33045 29597 33057 29631
rect 33091 29627 33103 29631
rect 33413 29631 33471 29637
rect 33152 29627 33364 29628
rect 33091 29600 33364 29627
rect 33091 29599 33180 29600
rect 33091 29597 33103 29599
rect 33045 29591 33103 29597
rect 31435 29532 32812 29560
rect 32968 29560 32996 29591
rect 33226 29560 33232 29572
rect 32968 29532 33232 29560
rect 31435 29529 31447 29532
rect 31389 29523 31447 29529
rect 27522 29492 27528 29504
rect 23860 29464 27528 29492
rect 23753 29455 23811 29461
rect 27522 29452 27528 29464
rect 27580 29452 27586 29504
rect 27798 29452 27804 29504
rect 27856 29452 27862 29504
rect 29822 29452 29828 29504
rect 29880 29452 29886 29504
rect 30116 29492 30144 29523
rect 33226 29520 33232 29532
rect 33284 29520 33290 29572
rect 33336 29560 33364 29600
rect 33413 29597 33425 29631
rect 33459 29628 33471 29631
rect 33502 29628 33508 29640
rect 33459 29600 33508 29628
rect 33459 29597 33471 29600
rect 33413 29591 33471 29597
rect 33502 29588 33508 29600
rect 33560 29588 33566 29640
rect 33796 29637 33824 29668
rect 35986 29656 35992 29668
rect 36044 29696 36050 29708
rect 36265 29699 36323 29705
rect 36265 29696 36277 29699
rect 36044 29668 36277 29696
rect 36044 29656 36050 29668
rect 36265 29665 36277 29668
rect 36311 29696 36323 29699
rect 39206 29696 39212 29708
rect 36311 29668 36768 29696
rect 36311 29665 36323 29668
rect 36265 29659 36323 29665
rect 33781 29631 33839 29637
rect 33781 29597 33793 29631
rect 33827 29597 33839 29631
rect 34330 29628 34336 29640
rect 33781 29591 33839 29597
rect 33888 29600 34336 29628
rect 33888 29560 33916 29600
rect 34330 29588 34336 29600
rect 34388 29588 34394 29640
rect 34698 29588 34704 29640
rect 34756 29628 34762 29640
rect 34882 29628 34888 29640
rect 34756 29600 34888 29628
rect 34756 29588 34762 29600
rect 34882 29588 34888 29600
rect 34940 29588 34946 29640
rect 34974 29588 34980 29640
rect 35032 29628 35038 29640
rect 35032 29600 35388 29628
rect 35032 29588 35038 29600
rect 33336 29532 33916 29560
rect 33980 29532 35020 29560
rect 30374 29492 30380 29504
rect 30116 29464 30380 29492
rect 30374 29452 30380 29464
rect 30432 29452 30438 29504
rect 30466 29452 30472 29504
rect 30524 29452 30530 29504
rect 31110 29452 31116 29504
rect 31168 29492 31174 29504
rect 32766 29492 32772 29504
rect 31168 29464 32772 29492
rect 31168 29452 31174 29464
rect 32766 29452 32772 29464
rect 32824 29492 32830 29504
rect 33137 29495 33195 29501
rect 33137 29492 33149 29495
rect 32824 29464 33149 29492
rect 32824 29452 32830 29464
rect 33137 29461 33149 29464
rect 33183 29492 33195 29495
rect 33980 29492 34008 29532
rect 34992 29504 35020 29532
rect 33183 29464 34008 29492
rect 33183 29461 33195 29464
rect 33137 29455 33195 29461
rect 34054 29452 34060 29504
rect 34112 29452 34118 29504
rect 34974 29452 34980 29504
rect 35032 29452 35038 29504
rect 35360 29492 35388 29600
rect 35526 29588 35532 29640
rect 35584 29628 35590 29640
rect 36740 29637 36768 29668
rect 37752 29668 39212 29696
rect 35621 29631 35679 29637
rect 35621 29628 35633 29631
rect 35584 29600 35633 29628
rect 35584 29588 35590 29600
rect 35621 29597 35633 29600
rect 35667 29597 35679 29631
rect 35621 29591 35679 29597
rect 36081 29631 36139 29637
rect 36081 29597 36093 29631
rect 36127 29597 36139 29631
rect 36081 29591 36139 29597
rect 36725 29631 36783 29637
rect 36725 29597 36737 29631
rect 36771 29597 36783 29631
rect 36725 29591 36783 29597
rect 36096 29560 36124 29591
rect 36906 29588 36912 29640
rect 36964 29588 36970 29640
rect 37752 29637 37780 29668
rect 39206 29656 39212 29668
rect 39264 29656 39270 29708
rect 37737 29631 37795 29637
rect 37737 29597 37749 29631
rect 37783 29597 37795 29631
rect 37737 29591 37795 29597
rect 38381 29631 38439 29637
rect 38381 29597 38393 29631
rect 38427 29597 38439 29631
rect 38381 29591 38439 29597
rect 36262 29560 36268 29572
rect 36096 29532 36268 29560
rect 36262 29520 36268 29532
rect 36320 29520 36326 29572
rect 37642 29520 37648 29572
rect 37700 29560 37706 29572
rect 38013 29563 38071 29569
rect 38013 29560 38025 29563
rect 37700 29532 38025 29560
rect 37700 29520 37706 29532
rect 38013 29529 38025 29532
rect 38059 29529 38071 29563
rect 38396 29560 38424 29591
rect 38470 29588 38476 29640
rect 38528 29588 38534 29640
rect 38746 29588 38752 29640
rect 38804 29628 38810 29640
rect 38841 29631 38899 29637
rect 38841 29628 38853 29631
rect 38804 29600 38853 29628
rect 38804 29588 38810 29600
rect 38841 29597 38853 29600
rect 38887 29628 38899 29631
rect 40037 29631 40095 29637
rect 38887 29600 39344 29628
rect 38887 29597 38899 29600
rect 38841 29591 38899 29597
rect 39209 29563 39267 29569
rect 39209 29560 39221 29563
rect 38396 29532 38884 29560
rect 38013 29523 38071 29529
rect 38856 29504 38884 29532
rect 39040 29532 39221 29560
rect 35802 29492 35808 29504
rect 35360 29464 35808 29492
rect 35802 29452 35808 29464
rect 35860 29452 35866 29504
rect 35897 29495 35955 29501
rect 35897 29461 35909 29495
rect 35943 29492 35955 29495
rect 36630 29492 36636 29504
rect 35943 29464 36636 29492
rect 35943 29461 35955 29464
rect 35897 29455 35955 29461
rect 36630 29452 36636 29464
rect 36688 29452 36694 29504
rect 36998 29452 37004 29504
rect 37056 29492 37062 29504
rect 38746 29492 38752 29504
rect 37056 29464 38752 29492
rect 37056 29452 37062 29464
rect 38746 29452 38752 29464
rect 38804 29452 38810 29504
rect 38838 29452 38844 29504
rect 38896 29452 38902 29504
rect 39040 29501 39068 29532
rect 39209 29529 39221 29532
rect 39255 29529 39267 29563
rect 39316 29560 39344 29600
rect 40037 29597 40049 29631
rect 40083 29628 40095 29631
rect 41506 29628 41512 29640
rect 40083 29600 41512 29628
rect 40083 29597 40095 29600
rect 40037 29591 40095 29597
rect 41506 29588 41512 29600
rect 41564 29588 41570 29640
rect 40678 29560 40684 29572
rect 39316 29532 40684 29560
rect 39209 29523 39267 29529
rect 40678 29520 40684 29532
rect 40736 29520 40742 29572
rect 39025 29495 39083 29501
rect 39025 29461 39037 29495
rect 39071 29461 39083 29495
rect 39025 29455 39083 29461
rect 1104 29402 41400 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 41400 29402
rect 1104 29328 41400 29350
rect 2682 29248 2688 29300
rect 2740 29288 2746 29300
rect 2961 29291 3019 29297
rect 2961 29288 2973 29291
rect 2740 29260 2973 29288
rect 2740 29248 2746 29260
rect 2961 29257 2973 29260
rect 3007 29257 3019 29291
rect 4522 29288 4528 29300
rect 2961 29251 3019 29257
rect 3252 29260 4528 29288
rect 2593 29223 2651 29229
rect 2593 29189 2605 29223
rect 2639 29220 2651 29223
rect 3252 29220 3280 29260
rect 4522 29248 4528 29260
rect 4580 29248 4586 29300
rect 4617 29291 4675 29297
rect 4617 29257 4629 29291
rect 4663 29288 4675 29291
rect 5350 29288 5356 29300
rect 4663 29260 5356 29288
rect 4663 29257 4675 29260
rect 4617 29251 4675 29257
rect 5350 29248 5356 29260
rect 5408 29248 5414 29300
rect 5534 29248 5540 29300
rect 5592 29288 5598 29300
rect 5997 29291 6055 29297
rect 5997 29288 6009 29291
rect 5592 29260 6009 29288
rect 5592 29248 5598 29260
rect 5997 29257 6009 29260
rect 6043 29257 6055 29291
rect 7098 29288 7104 29300
rect 5997 29251 6055 29257
rect 6104 29260 7104 29288
rect 2639 29192 3280 29220
rect 3329 29223 3387 29229
rect 2639 29189 2651 29192
rect 2593 29183 2651 29189
rect 3329 29189 3341 29223
rect 3375 29220 3387 29223
rect 3602 29220 3608 29232
rect 3375 29192 3608 29220
rect 3375 29189 3387 29192
rect 3329 29183 3387 29189
rect 3602 29180 3608 29192
rect 3660 29180 3666 29232
rect 4154 29180 4160 29232
rect 4212 29180 4218 29232
rect 4890 29180 4896 29232
rect 4948 29180 4954 29232
rect 4985 29223 5043 29229
rect 4985 29189 4997 29223
rect 5031 29220 5043 29223
rect 5902 29220 5908 29232
rect 5031 29192 5304 29220
rect 5031 29189 5043 29192
rect 4985 29183 5043 29189
rect 5276 29164 5304 29192
rect 5552 29192 5908 29220
rect 2041 29155 2099 29161
rect 2041 29121 2053 29155
rect 2087 29152 2099 29155
rect 2501 29155 2559 29161
rect 2087 29124 2176 29152
rect 2087 29121 2099 29124
rect 2041 29115 2099 29121
rect 2148 29025 2176 29124
rect 2501 29121 2513 29155
rect 2547 29152 2559 29155
rect 3234 29152 3240 29164
rect 2547 29124 3240 29152
rect 2547 29121 2559 29124
rect 2501 29115 2559 29121
rect 3234 29112 3240 29124
rect 3292 29112 3298 29164
rect 3418 29112 3424 29164
rect 3476 29112 3482 29164
rect 4709 29155 4767 29161
rect 4709 29121 4721 29155
rect 4755 29121 4767 29155
rect 4709 29115 4767 29121
rect 2777 29087 2835 29093
rect 2777 29053 2789 29087
rect 2823 29084 2835 29087
rect 3605 29087 3663 29093
rect 2823 29056 3372 29084
rect 2823 29053 2835 29056
rect 2777 29047 2835 29053
rect 3344 29028 3372 29056
rect 3605 29053 3617 29087
rect 3651 29053 3663 29087
rect 4724 29084 4752 29115
rect 5074 29112 5080 29164
rect 5132 29112 5138 29164
rect 5166 29112 5172 29164
rect 5224 29112 5230 29164
rect 5258 29112 5264 29164
rect 5316 29112 5322 29164
rect 5350 29112 5356 29164
rect 5408 29112 5414 29164
rect 5446 29155 5504 29161
rect 5446 29121 5458 29155
rect 5492 29152 5504 29155
rect 5552 29152 5580 29192
rect 5902 29180 5908 29192
rect 5960 29180 5966 29232
rect 5492 29124 5580 29152
rect 5492 29121 5504 29124
rect 5446 29115 5504 29121
rect 5626 29112 5632 29164
rect 5684 29112 5690 29164
rect 5721 29155 5779 29161
rect 5721 29121 5733 29155
rect 5767 29121 5779 29155
rect 5721 29115 5779 29121
rect 5184 29084 5212 29112
rect 4724 29056 5212 29084
rect 5736 29084 5764 29115
rect 5810 29112 5816 29164
rect 5868 29161 5874 29164
rect 5868 29152 5876 29161
rect 6104 29152 6132 29260
rect 7098 29248 7104 29260
rect 7156 29248 7162 29300
rect 7834 29248 7840 29300
rect 7892 29248 7898 29300
rect 8386 29288 8392 29300
rect 8092 29260 8392 29288
rect 7852 29220 7880 29248
rect 6380 29192 7328 29220
rect 5868 29124 6132 29152
rect 5868 29115 5876 29124
rect 5868 29112 5874 29115
rect 6270 29112 6276 29164
rect 6328 29152 6334 29164
rect 6380 29161 6408 29192
rect 6365 29155 6423 29161
rect 6365 29152 6377 29155
rect 6328 29124 6377 29152
rect 6328 29112 6334 29124
rect 6365 29121 6377 29124
rect 6411 29121 6423 29155
rect 6365 29115 6423 29121
rect 6546 29112 6552 29164
rect 6604 29112 6610 29164
rect 6638 29112 6644 29164
rect 6696 29112 6702 29164
rect 6730 29112 6736 29164
rect 6788 29112 6794 29164
rect 7300 29161 7328 29192
rect 7484 29192 7880 29220
rect 7285 29155 7343 29161
rect 7285 29121 7297 29155
rect 7331 29152 7343 29155
rect 7374 29152 7380 29164
rect 7331 29124 7380 29152
rect 7331 29121 7343 29124
rect 7285 29115 7343 29121
rect 7374 29112 7380 29124
rect 7432 29112 7438 29164
rect 7484 29161 7512 29192
rect 7469 29155 7527 29161
rect 7469 29121 7481 29155
rect 7515 29121 7527 29155
rect 7469 29115 7527 29121
rect 7558 29112 7564 29164
rect 7616 29112 7622 29164
rect 7650 29112 7656 29164
rect 7708 29112 7714 29164
rect 7926 29112 7932 29164
rect 7984 29112 7990 29164
rect 8092 29161 8120 29260
rect 8386 29248 8392 29260
rect 8444 29288 8450 29300
rect 8444 29260 9168 29288
rect 8444 29248 8450 29260
rect 9140 29232 9168 29260
rect 9674 29248 9680 29300
rect 9732 29288 9738 29300
rect 10597 29291 10655 29297
rect 10597 29288 10609 29291
rect 9732 29260 10609 29288
rect 9732 29248 9738 29260
rect 8202 29180 8208 29232
rect 8260 29180 8266 29232
rect 8570 29180 8576 29232
rect 8628 29180 8634 29232
rect 8662 29180 8668 29232
rect 8720 29180 8726 29232
rect 9122 29180 9128 29232
rect 9180 29180 9186 29232
rect 9968 29229 9996 29260
rect 10597 29257 10609 29260
rect 10643 29257 10655 29291
rect 10597 29251 10655 29257
rect 9493 29223 9551 29229
rect 9493 29189 9505 29223
rect 9539 29220 9551 29223
rect 9953 29223 10011 29229
rect 9539 29192 9720 29220
rect 9539 29189 9551 29192
rect 9493 29183 9551 29189
rect 8077 29155 8135 29161
rect 8077 29121 8089 29155
rect 8123 29121 8135 29155
rect 8077 29115 8135 29121
rect 8294 29112 8300 29164
rect 8352 29112 8358 29164
rect 8435 29155 8493 29161
rect 8435 29121 8447 29155
rect 8481 29152 8493 29155
rect 8588 29152 8616 29180
rect 8481 29124 8616 29152
rect 8680 29152 8708 29180
rect 9306 29152 9312 29164
rect 8680 29124 9312 29152
rect 8481 29121 8493 29124
rect 8435 29115 8493 29121
rect 9306 29112 9312 29124
rect 9364 29152 9370 29164
rect 9692 29161 9720 29192
rect 9953 29189 9965 29223
rect 9999 29189 10011 29223
rect 9953 29183 10011 29189
rect 10042 29180 10048 29232
rect 10100 29180 10106 29232
rect 10612 29220 10640 29251
rect 11698 29248 11704 29300
rect 11756 29288 11762 29300
rect 11756 29260 12480 29288
rect 11756 29248 11762 29260
rect 11514 29220 11520 29232
rect 10612 29192 11520 29220
rect 11514 29180 11520 29192
rect 11572 29220 11578 29232
rect 11572 29192 12296 29220
rect 11572 29180 11578 29192
rect 9858 29161 9864 29164
rect 9401 29155 9459 29161
rect 9401 29152 9413 29155
rect 9364 29124 9413 29152
rect 9364 29112 9370 29124
rect 9401 29121 9413 29124
rect 9447 29121 9459 29155
rect 9401 29115 9459 29121
rect 9585 29155 9643 29161
rect 9585 29121 9597 29155
rect 9631 29121 9643 29155
rect 9585 29115 9643 29121
rect 9677 29155 9735 29161
rect 9677 29121 9689 29155
rect 9723 29121 9735 29155
rect 9677 29115 9735 29121
rect 9825 29155 9864 29161
rect 9825 29121 9837 29155
rect 9825 29115 9864 29121
rect 5736 29056 8616 29084
rect 3605 29047 3663 29053
rect 2133 29019 2191 29025
rect 2133 28985 2145 29019
rect 2179 28985 2191 29019
rect 2133 28979 2191 28985
rect 3326 28976 3332 29028
rect 3384 29016 3390 29028
rect 3620 29016 3648 29047
rect 5828 29028 5856 29056
rect 3384 28988 3648 29016
rect 4525 29019 4583 29025
rect 3384 28976 3390 28988
rect 4525 28985 4537 29019
rect 4571 29016 4583 29019
rect 5261 29019 5319 29025
rect 4571 28988 5212 29016
rect 4571 28985 4583 28988
rect 4525 28979 4583 28985
rect 1854 28908 1860 28960
rect 1912 28908 1918 28960
rect 5184 28948 5212 28988
rect 5261 28985 5273 29019
rect 5307 29016 5319 29019
rect 5718 29016 5724 29028
rect 5307 28988 5724 29016
rect 5307 28985 5319 28988
rect 5261 28979 5319 28985
rect 5718 28976 5724 28988
rect 5776 28976 5782 29028
rect 5810 28976 5816 29028
rect 5868 28976 5874 29028
rect 5920 28988 6776 29016
rect 5920 28948 5948 28988
rect 5184 28920 5948 28948
rect 6748 28948 6776 28988
rect 6822 28976 6828 29028
rect 6880 29016 6886 29028
rect 6917 29019 6975 29025
rect 6917 29016 6929 29019
rect 6880 28988 6929 29016
rect 6880 28976 6886 28988
rect 6917 28985 6929 28988
rect 6963 28985 6975 29019
rect 6917 28979 6975 28985
rect 7374 28976 7380 29028
rect 7432 29016 7438 29028
rect 8294 29016 8300 29028
rect 7432 28988 8300 29016
rect 7432 28976 7438 28988
rect 8294 28976 8300 28988
rect 8352 28976 8358 29028
rect 8386 28976 8392 29028
rect 8444 28976 8450 29028
rect 8588 29025 8616 29056
rect 9030 29044 9036 29096
rect 9088 29084 9094 29096
rect 9125 29087 9183 29093
rect 9125 29084 9137 29087
rect 9088 29056 9137 29084
rect 9088 29044 9094 29056
rect 9125 29053 9137 29056
rect 9171 29053 9183 29087
rect 9600 29084 9628 29115
rect 9858 29112 9864 29115
rect 9916 29112 9922 29164
rect 10134 29112 10140 29164
rect 10192 29161 10198 29164
rect 10192 29155 10241 29161
rect 10192 29121 10195 29155
rect 10229 29152 10241 29155
rect 10597 29155 10655 29161
rect 10597 29152 10609 29155
rect 10229 29124 10609 29152
rect 10229 29121 10241 29124
rect 10192 29115 10241 29121
rect 10597 29121 10609 29124
rect 10643 29152 10655 29155
rect 11054 29152 11060 29164
rect 10643 29124 11060 29152
rect 10643 29121 10655 29124
rect 10597 29115 10655 29121
rect 10192 29112 10198 29115
rect 11054 29112 11060 29124
rect 11112 29112 11118 29164
rect 12268 29161 12296 29192
rect 12342 29180 12348 29232
rect 12400 29180 12406 29232
rect 12452 29220 12480 29260
rect 12526 29248 12532 29300
rect 12584 29288 12590 29300
rect 12621 29291 12679 29297
rect 12621 29288 12633 29291
rect 12584 29260 12633 29288
rect 12584 29248 12590 29260
rect 12621 29257 12633 29260
rect 12667 29257 12679 29291
rect 12621 29251 12679 29257
rect 13354 29248 13360 29300
rect 13412 29288 13418 29300
rect 13449 29291 13507 29297
rect 13449 29288 13461 29291
rect 13412 29260 13461 29288
rect 13412 29248 13418 29260
rect 13449 29257 13461 29260
rect 13495 29257 13507 29291
rect 13449 29251 13507 29257
rect 13538 29248 13544 29300
rect 13596 29288 13602 29300
rect 13633 29291 13691 29297
rect 13633 29288 13645 29291
rect 13596 29260 13645 29288
rect 13596 29248 13602 29260
rect 13633 29257 13645 29260
rect 13679 29257 13691 29291
rect 13633 29251 13691 29257
rect 13909 29291 13967 29297
rect 13909 29257 13921 29291
rect 13955 29288 13967 29291
rect 14090 29288 14096 29300
rect 13955 29260 14096 29288
rect 13955 29257 13967 29260
rect 13909 29251 13967 29257
rect 14090 29248 14096 29260
rect 14148 29248 14154 29300
rect 14185 29291 14243 29297
rect 14185 29257 14197 29291
rect 14231 29288 14243 29291
rect 14366 29288 14372 29300
rect 14231 29260 14372 29288
rect 14231 29257 14243 29260
rect 14185 29251 14243 29257
rect 14366 29248 14372 29260
rect 14424 29248 14430 29300
rect 14476 29260 15056 29288
rect 13081 29223 13139 29229
rect 13081 29220 13093 29223
rect 12452 29192 13093 29220
rect 13081 29189 13093 29192
rect 13127 29220 13139 29223
rect 14476 29220 14504 29260
rect 15028 29220 15056 29260
rect 15102 29248 15108 29300
rect 15160 29288 15166 29300
rect 15933 29291 15991 29297
rect 15933 29288 15945 29291
rect 15160 29260 15945 29288
rect 15160 29248 15166 29260
rect 15933 29257 15945 29260
rect 15979 29257 15991 29291
rect 15933 29251 15991 29257
rect 16942 29248 16948 29300
rect 17000 29288 17006 29300
rect 17589 29291 17647 29297
rect 17589 29288 17601 29291
rect 17000 29260 17601 29288
rect 17000 29248 17006 29260
rect 17589 29257 17601 29260
rect 17635 29257 17647 29291
rect 17589 29251 17647 29257
rect 17678 29248 17684 29300
rect 17736 29248 17742 29300
rect 20809 29291 20867 29297
rect 20809 29288 20821 29291
rect 18708 29260 20821 29288
rect 13127 29192 14504 29220
rect 14568 29192 14963 29220
rect 15028 29192 15608 29220
rect 13127 29189 13139 29192
rect 13081 29183 13139 29189
rect 11965 29155 12023 29161
rect 11965 29152 11977 29155
rect 11900 29124 11977 29152
rect 10410 29084 10416 29096
rect 9600 29056 10416 29084
rect 9125 29047 9183 29053
rect 10410 29044 10416 29056
rect 10468 29044 10474 29096
rect 8573 29019 8631 29025
rect 8573 28985 8585 29019
rect 8619 28985 8631 29019
rect 8941 29019 8999 29025
rect 8941 29016 8953 29019
rect 8573 28979 8631 28985
rect 8864 28988 8953 29016
rect 7006 28948 7012 28960
rect 6748 28920 7012 28948
rect 7006 28908 7012 28920
rect 7064 28908 7070 28960
rect 7834 28908 7840 28960
rect 7892 28908 7898 28960
rect 8202 28908 8208 28960
rect 8260 28948 8266 28960
rect 8404 28948 8432 28976
rect 8864 28960 8892 28988
rect 8941 28985 8953 28988
rect 8987 28985 8999 29019
rect 8941 28979 8999 28985
rect 11057 29019 11115 29025
rect 11057 28985 11069 29019
rect 11103 28985 11115 29019
rect 11057 28979 11115 28985
rect 8260 28920 8432 28948
rect 8260 28908 8266 28920
rect 8846 28908 8852 28960
rect 8904 28908 8910 28960
rect 10318 28908 10324 28960
rect 10376 28908 10382 28960
rect 11072 28948 11100 28979
rect 11606 28948 11612 28960
rect 11072 28920 11612 28948
rect 11606 28908 11612 28920
rect 11664 28908 11670 28960
rect 11900 28948 11928 29124
rect 11965 29121 11977 29124
rect 12011 29121 12023 29155
rect 11965 29115 12023 29121
rect 12125 29155 12183 29161
rect 12125 29121 12137 29155
rect 12171 29152 12183 29155
rect 12253 29155 12311 29161
rect 12171 29121 12204 29152
rect 12125 29115 12204 29121
rect 12253 29121 12265 29155
rect 12299 29121 12311 29155
rect 12253 29115 12311 29121
rect 12442 29155 12500 29161
rect 12442 29121 12454 29155
rect 12488 29152 12500 29155
rect 12710 29152 12716 29164
rect 12488 29124 12716 29152
rect 12488 29121 12500 29124
rect 12442 29115 12500 29121
rect 12176 29016 12204 29115
rect 12710 29112 12716 29124
rect 12768 29112 12774 29164
rect 12802 29112 12808 29164
rect 12860 29112 12866 29164
rect 12986 29161 12992 29164
rect 12953 29155 12992 29161
rect 12953 29121 12965 29155
rect 12953 29115 12992 29121
rect 12968 29112 12992 29115
rect 13044 29112 13050 29164
rect 13170 29112 13176 29164
rect 13228 29112 13234 29164
rect 13270 29155 13328 29161
rect 13270 29121 13282 29155
rect 13316 29152 13328 29155
rect 13446 29152 13452 29164
rect 13316 29124 13452 29152
rect 13316 29121 13328 29124
rect 13270 29115 13328 29121
rect 13446 29112 13452 29124
rect 13504 29112 13510 29164
rect 13541 29155 13599 29161
rect 13541 29121 13553 29155
rect 13587 29121 13599 29155
rect 13541 29115 13599 29121
rect 12802 29016 12808 29028
rect 12176 28988 12808 29016
rect 12802 28976 12808 28988
rect 12860 28976 12866 29028
rect 12968 29016 12996 29112
rect 13562 29084 13590 29115
rect 13722 29112 13728 29164
rect 13780 29112 13786 29164
rect 13817 29155 13875 29161
rect 13817 29121 13829 29155
rect 13863 29121 13875 29155
rect 13817 29115 13875 29121
rect 14001 29155 14059 29161
rect 14001 29121 14013 29155
rect 14047 29121 14059 29155
rect 14001 29115 14059 29121
rect 13832 29084 13860 29115
rect 13562 29056 13860 29084
rect 14016 29084 14044 29115
rect 14274 29112 14280 29164
rect 14332 29152 14338 29164
rect 14568 29152 14596 29192
rect 14332 29124 14596 29152
rect 14332 29112 14338 29124
rect 14826 29112 14832 29164
rect 14884 29112 14890 29164
rect 14935 29152 14963 29192
rect 15102 29152 15108 29164
rect 14935 29124 15108 29152
rect 15102 29112 15108 29124
rect 15160 29112 15166 29164
rect 15289 29155 15347 29161
rect 15289 29121 15301 29155
rect 15335 29121 15347 29155
rect 15289 29115 15347 29121
rect 14016 29056 14872 29084
rect 13354 29016 13360 29028
rect 12968 28988 13360 29016
rect 13354 28976 13360 28988
rect 13412 28976 13418 29028
rect 13562 29016 13590 29056
rect 13556 28988 13590 29016
rect 14844 29016 14872 29056
rect 15010 29044 15016 29096
rect 15068 29044 15074 29096
rect 15102 29016 15108 29028
rect 14844 28988 15108 29016
rect 13556 28960 13584 28988
rect 15102 28976 15108 28988
rect 15160 28976 15166 29028
rect 15304 29016 15332 29115
rect 15378 29112 15384 29164
rect 15436 29152 15442 29164
rect 15580 29161 15608 29192
rect 15838 29180 15844 29232
rect 15896 29220 15902 29232
rect 16025 29223 16083 29229
rect 16025 29220 16037 29223
rect 15896 29192 16037 29220
rect 15896 29180 15902 29192
rect 16025 29189 16037 29192
rect 16071 29220 16083 29223
rect 17313 29223 17371 29229
rect 16071 29192 16896 29220
rect 16071 29189 16083 29192
rect 16025 29183 16083 29189
rect 15565 29155 15623 29161
rect 15436 29124 15481 29152
rect 15436 29112 15442 29124
rect 15565 29121 15577 29155
rect 15611 29121 15623 29155
rect 15565 29115 15623 29121
rect 15580 29084 15608 29115
rect 15654 29112 15660 29164
rect 15712 29112 15718 29164
rect 15754 29155 15812 29161
rect 15754 29121 15766 29155
rect 15800 29152 15812 29155
rect 15800 29124 15884 29152
rect 15800 29121 15812 29124
rect 15754 29115 15812 29121
rect 15856 29084 15884 29124
rect 16206 29112 16212 29164
rect 16264 29112 16270 29164
rect 16393 29155 16451 29161
rect 16393 29121 16405 29155
rect 16439 29152 16451 29155
rect 16482 29152 16488 29164
rect 16439 29124 16488 29152
rect 16439 29121 16451 29124
rect 16393 29115 16451 29121
rect 16482 29112 16488 29124
rect 16540 29112 16546 29164
rect 16669 29155 16727 29161
rect 16669 29121 16681 29155
rect 16715 29121 16727 29155
rect 16868 29152 16896 29192
rect 17313 29189 17325 29223
rect 17359 29220 17371 29223
rect 17494 29220 17500 29232
rect 17359 29192 17500 29220
rect 17359 29189 17371 29192
rect 17313 29183 17371 29189
rect 17494 29180 17500 29192
rect 17552 29220 17558 29232
rect 17696 29220 17724 29248
rect 18708 29220 18736 29260
rect 20809 29257 20821 29260
rect 20855 29257 20867 29291
rect 20809 29251 20867 29257
rect 21634 29248 21640 29300
rect 21692 29288 21698 29300
rect 23109 29291 23167 29297
rect 23109 29288 23121 29291
rect 21692 29260 23121 29288
rect 21692 29248 21698 29260
rect 23109 29257 23121 29260
rect 23155 29257 23167 29291
rect 23109 29251 23167 29257
rect 20622 29220 20628 29232
rect 17552 29192 17724 29220
rect 17880 29192 18736 29220
rect 18800 29192 19472 29220
rect 17552 29180 17558 29192
rect 16942 29152 16948 29164
rect 16868 29124 16948 29152
rect 16669 29115 16727 29121
rect 15930 29084 15936 29096
rect 15580 29056 15792 29084
rect 15856 29056 15936 29084
rect 15764 29028 15792 29056
rect 15930 29044 15936 29056
rect 15988 29084 15994 29096
rect 16684 29084 16712 29115
rect 16942 29112 16948 29124
rect 17000 29112 17006 29164
rect 17218 29112 17224 29164
rect 17276 29112 17282 29164
rect 17402 29112 17408 29164
rect 17460 29152 17466 29164
rect 17880 29152 17908 29192
rect 17460 29124 17908 29152
rect 17957 29155 18015 29161
rect 17460 29112 17466 29124
rect 17957 29121 17969 29155
rect 18003 29121 18015 29155
rect 17957 29115 18015 29121
rect 18233 29155 18291 29161
rect 18233 29121 18245 29155
rect 18279 29152 18291 29155
rect 18322 29152 18328 29164
rect 18279 29124 18328 29152
rect 18279 29121 18291 29124
rect 18233 29115 18291 29121
rect 15988 29056 16344 29084
rect 16684 29056 17908 29084
rect 15988 29044 15994 29056
rect 15562 29016 15568 29028
rect 15304 28988 15568 29016
rect 15562 28976 15568 28988
rect 15620 28976 15626 29028
rect 15746 28976 15752 29028
rect 15804 28976 15810 29028
rect 16316 29025 16344 29056
rect 16301 29019 16359 29025
rect 16301 28985 16313 29019
rect 16347 29016 16359 29019
rect 16853 29019 16911 29025
rect 16853 29016 16865 29019
rect 16347 28988 16865 29016
rect 16347 28985 16359 28988
rect 16301 28979 16359 28985
rect 16853 28985 16865 28988
rect 16899 28985 16911 29019
rect 16853 28979 16911 28985
rect 16942 28976 16948 29028
rect 17000 28976 17006 29028
rect 17034 28976 17040 29028
rect 17092 28976 17098 29028
rect 17586 28976 17592 29028
rect 17644 29016 17650 29028
rect 17681 29019 17739 29025
rect 17681 29016 17693 29019
rect 17644 28988 17693 29016
rect 17644 28976 17650 28988
rect 17681 28985 17693 28988
rect 17727 28985 17739 29019
rect 17681 28979 17739 28985
rect 12526 28948 12532 28960
rect 11900 28920 12532 28948
rect 12526 28908 12532 28920
rect 12584 28908 12590 28960
rect 13538 28908 13544 28960
rect 13596 28908 13602 28960
rect 14182 28908 14188 28960
rect 14240 28948 14246 28960
rect 16393 28951 16451 28957
rect 16393 28948 16405 28951
rect 14240 28920 16405 28948
rect 14240 28908 14246 28920
rect 16393 28917 16405 28920
rect 16439 28917 16451 28951
rect 16960 28948 16988 28976
rect 17773 28951 17831 28957
rect 17773 28948 17785 28951
rect 16960 28920 17785 28948
rect 16393 28911 16451 28917
rect 17773 28917 17785 28920
rect 17819 28917 17831 28951
rect 17880 28948 17908 29056
rect 17972 29016 18000 29115
rect 18322 29112 18328 29124
rect 18380 29112 18386 29164
rect 18506 29112 18512 29164
rect 18564 29112 18570 29164
rect 18800 29161 18828 29192
rect 19444 29164 19472 29192
rect 20456 29192 20628 29220
rect 18785 29155 18843 29161
rect 18785 29121 18797 29155
rect 18831 29121 18843 29155
rect 18785 29115 18843 29121
rect 18874 29112 18880 29164
rect 18932 29152 18938 29164
rect 19245 29155 19303 29161
rect 19245 29152 19257 29155
rect 18932 29124 19257 29152
rect 18932 29112 18938 29124
rect 19245 29121 19257 29124
rect 19291 29121 19303 29155
rect 19245 29115 19303 29121
rect 18414 29016 18420 29028
rect 17972 28988 18420 29016
rect 18414 28976 18420 28988
rect 18472 28976 18478 29028
rect 18690 28976 18696 29028
rect 18748 28976 18754 29028
rect 19260 28960 19288 29115
rect 19426 29112 19432 29164
rect 19484 29112 19490 29164
rect 20456 29161 20484 29192
rect 20622 29180 20628 29192
rect 20680 29180 20686 29232
rect 22002 29220 22008 29232
rect 21836 29192 22008 29220
rect 20441 29155 20499 29161
rect 20441 29121 20453 29155
rect 20487 29121 20499 29155
rect 20441 29115 20499 29121
rect 20530 29112 20536 29164
rect 20588 29112 20594 29164
rect 21085 29155 21143 29161
rect 21085 29121 21097 29155
rect 21131 29152 21143 29155
rect 21450 29152 21456 29164
rect 21131 29124 21456 29152
rect 21131 29121 21143 29124
rect 21085 29115 21143 29121
rect 21450 29112 21456 29124
rect 21508 29112 21514 29164
rect 19518 29044 19524 29096
rect 19576 29084 19582 29096
rect 19613 29087 19671 29093
rect 19613 29084 19625 29087
rect 19576 29056 19625 29084
rect 19576 29044 19582 29056
rect 19613 29053 19625 29056
rect 19659 29084 19671 29087
rect 19659 29056 21036 29084
rect 19659 29053 19671 29056
rect 19613 29047 19671 29053
rect 19886 28976 19892 29028
rect 19944 29016 19950 29028
rect 20901 29019 20959 29025
rect 20901 29016 20913 29019
rect 19944 28988 20913 29016
rect 19944 28976 19950 28988
rect 20901 28985 20913 28988
rect 20947 28985 20959 29019
rect 21008 29016 21036 29056
rect 21266 29044 21272 29096
rect 21324 29044 21330 29096
rect 21361 29087 21419 29093
rect 21361 29053 21373 29087
rect 21407 29084 21419 29087
rect 21836 29084 21864 29192
rect 22002 29180 22008 29192
rect 22060 29180 22066 29232
rect 22738 29220 22744 29232
rect 22296 29192 22744 29220
rect 21910 29112 21916 29164
rect 21968 29152 21974 29164
rect 22296 29161 22324 29192
rect 22738 29180 22744 29192
rect 22796 29180 22802 29232
rect 23124 29220 23152 29251
rect 23474 29248 23480 29300
rect 23532 29288 23538 29300
rect 24121 29291 24179 29297
rect 24121 29288 24133 29291
rect 23532 29260 24133 29288
rect 23532 29248 23538 29260
rect 24121 29257 24133 29260
rect 24167 29257 24179 29291
rect 24121 29251 24179 29257
rect 26510 29248 26516 29300
rect 26568 29288 26574 29300
rect 30009 29291 30067 29297
rect 30009 29288 30021 29291
rect 26568 29260 30021 29288
rect 26568 29248 26574 29260
rect 30009 29257 30021 29260
rect 30055 29257 30067 29291
rect 30009 29251 30067 29257
rect 30466 29248 30472 29300
rect 30524 29288 30530 29300
rect 30926 29288 30932 29300
rect 30524 29260 30932 29288
rect 30524 29248 30530 29260
rect 30926 29248 30932 29260
rect 30984 29288 30990 29300
rect 31481 29291 31539 29297
rect 31481 29288 31493 29291
rect 30984 29260 31493 29288
rect 30984 29248 30990 29260
rect 31481 29257 31493 29260
rect 31527 29257 31539 29291
rect 31481 29251 31539 29257
rect 32950 29248 32956 29300
rect 33008 29288 33014 29300
rect 33008 29260 33364 29288
rect 33008 29248 33014 29260
rect 24946 29220 24952 29232
rect 23124 29192 23888 29220
rect 22189 29155 22247 29161
rect 22189 29152 22201 29155
rect 21968 29124 22201 29152
rect 21968 29112 21974 29124
rect 22189 29121 22201 29124
rect 22235 29121 22247 29155
rect 22189 29115 22247 29121
rect 22281 29155 22339 29161
rect 22281 29121 22293 29155
rect 22327 29121 22339 29155
rect 22281 29115 22339 29121
rect 22462 29112 22468 29164
rect 22520 29112 22526 29164
rect 23474 29112 23480 29164
rect 23532 29112 23538 29164
rect 23860 29158 23888 29192
rect 24412 29192 24952 29220
rect 23937 29158 23995 29161
rect 23860 29155 23995 29158
rect 23860 29130 23949 29155
rect 23937 29121 23949 29130
rect 23983 29121 23995 29155
rect 23937 29115 23995 29121
rect 24210 29112 24216 29164
rect 24268 29112 24274 29164
rect 21407 29056 21864 29084
rect 22373 29087 22431 29093
rect 21407 29053 21419 29056
rect 21361 29047 21419 29053
rect 22373 29053 22385 29087
rect 22419 29084 22431 29087
rect 22554 29084 22560 29096
rect 22419 29056 22560 29084
rect 22419 29053 22431 29056
rect 22373 29047 22431 29053
rect 22554 29044 22560 29056
rect 22612 29044 22618 29096
rect 23845 29087 23903 29093
rect 23845 29053 23857 29087
rect 23891 29084 23903 29087
rect 24412 29084 24440 29192
rect 24946 29180 24952 29192
rect 25004 29180 25010 29232
rect 31386 29220 31392 29232
rect 28966 29192 30880 29220
rect 24854 29112 24860 29164
rect 24912 29112 24918 29164
rect 25222 29112 25228 29164
rect 25280 29112 25286 29164
rect 25409 29155 25467 29161
rect 25409 29121 25421 29155
rect 25455 29121 25467 29155
rect 25409 29115 25467 29121
rect 23891 29056 24440 29084
rect 23891 29053 23903 29056
rect 23845 29047 23903 29053
rect 24486 29044 24492 29096
rect 24544 29084 24550 29096
rect 24765 29087 24823 29093
rect 24765 29084 24777 29087
rect 24544 29056 24777 29084
rect 24544 29044 24550 29056
rect 24765 29053 24777 29056
rect 24811 29053 24823 29087
rect 24765 29047 24823 29053
rect 22005 29019 22063 29025
rect 22005 29016 22017 29019
rect 21008 28988 22017 29016
rect 20901 28979 20959 28985
rect 22005 28985 22017 28988
rect 22051 28985 22063 29019
rect 22005 28979 22063 28985
rect 22186 28976 22192 29028
rect 22244 29016 22250 29028
rect 23382 29016 23388 29028
rect 22244 28988 23388 29016
rect 22244 28976 22250 28988
rect 23382 28976 23388 28988
rect 23440 28976 23446 29028
rect 25424 29016 25452 29115
rect 25498 29112 25504 29164
rect 25556 29152 25562 29164
rect 26970 29152 26976 29164
rect 25556 29124 26976 29152
rect 25556 29112 25562 29124
rect 26970 29112 26976 29124
rect 27028 29152 27034 29164
rect 28966 29152 28994 29192
rect 27028 29124 28994 29152
rect 29549 29155 29607 29161
rect 27028 29112 27034 29124
rect 29549 29121 29561 29155
rect 29595 29121 29607 29155
rect 29549 29115 29607 29121
rect 29564 29084 29592 29115
rect 29730 29112 29736 29164
rect 29788 29112 29794 29164
rect 29822 29112 29828 29164
rect 29880 29112 29886 29164
rect 30852 29084 30880 29192
rect 30944 29192 31392 29220
rect 30944 29161 30972 29192
rect 31386 29180 31392 29192
rect 31444 29220 31450 29232
rect 31444 29192 31892 29220
rect 31444 29180 31450 29192
rect 31864 29164 31892 29192
rect 32324 29192 33088 29220
rect 30929 29155 30987 29161
rect 30929 29121 30941 29155
rect 30975 29121 30987 29155
rect 30929 29115 30987 29121
rect 31110 29112 31116 29164
rect 31168 29112 31174 29164
rect 31202 29112 31208 29164
rect 31260 29112 31266 29164
rect 31481 29155 31539 29161
rect 31481 29121 31493 29155
rect 31527 29152 31539 29155
rect 31662 29152 31668 29164
rect 31527 29124 31668 29152
rect 31527 29121 31539 29124
rect 31481 29115 31539 29121
rect 31662 29112 31668 29124
rect 31720 29112 31726 29164
rect 31846 29112 31852 29164
rect 31904 29112 31910 29164
rect 32324 29161 32352 29192
rect 33060 29164 33088 29192
rect 33134 29180 33140 29232
rect 33192 29180 33198 29232
rect 32309 29155 32367 29161
rect 32309 29121 32321 29155
rect 32355 29121 32367 29155
rect 32490 29152 32496 29164
rect 32548 29161 32554 29164
rect 32548 29155 32589 29161
rect 32309 29115 32367 29121
rect 32416 29124 32496 29152
rect 31297 29087 31355 29093
rect 29564 29056 29776 29084
rect 30852 29056 31248 29084
rect 29748 29028 29776 29056
rect 25774 29016 25780 29028
rect 24136 28988 25780 29016
rect 18506 28948 18512 28960
rect 17880 28920 18512 28948
rect 17773 28911 17831 28917
rect 18506 28908 18512 28920
rect 18564 28908 18570 28960
rect 19242 28908 19248 28960
rect 19300 28908 19306 28960
rect 20625 28951 20683 28957
rect 20625 28917 20637 28951
rect 20671 28948 20683 28951
rect 20714 28948 20720 28960
rect 20671 28920 20720 28948
rect 20671 28917 20683 28920
rect 20625 28911 20683 28917
rect 20714 28908 20720 28920
rect 20772 28908 20778 28960
rect 23937 28951 23995 28957
rect 23937 28917 23949 28951
rect 23983 28948 23995 28951
rect 24136 28948 24164 28988
rect 25774 28976 25780 28988
rect 25832 28976 25838 29028
rect 27338 29016 27344 29028
rect 26436 28988 27344 29016
rect 26436 28960 26464 28988
rect 27338 28976 27344 28988
rect 27396 28976 27402 29028
rect 27586 28988 29685 29016
rect 23983 28920 24164 28948
rect 23983 28917 23995 28920
rect 23937 28911 23995 28917
rect 24302 28908 24308 28960
rect 24360 28948 24366 28960
rect 25958 28948 25964 28960
rect 24360 28920 25964 28948
rect 24360 28908 24366 28920
rect 25958 28908 25964 28920
rect 26016 28908 26022 28960
rect 26418 28908 26424 28960
rect 26476 28908 26482 28960
rect 26602 28908 26608 28960
rect 26660 28948 26666 28960
rect 27246 28948 27252 28960
rect 26660 28920 27252 28948
rect 26660 28908 26666 28920
rect 27246 28908 27252 28920
rect 27304 28948 27310 28960
rect 27586 28948 27614 28988
rect 27304 28920 27614 28948
rect 27304 28908 27310 28920
rect 28258 28908 28264 28960
rect 28316 28948 28322 28960
rect 29362 28948 29368 28960
rect 28316 28920 29368 28948
rect 28316 28908 28322 28920
rect 29362 28908 29368 28920
rect 29420 28908 29426 28960
rect 29454 28908 29460 28960
rect 29512 28948 29518 28960
rect 29549 28951 29607 28957
rect 29549 28948 29561 28951
rect 29512 28920 29561 28948
rect 29512 28908 29518 28920
rect 29549 28917 29561 28920
rect 29595 28917 29607 28951
rect 29657 28948 29685 28988
rect 29730 28976 29736 29028
rect 29788 29016 29794 29028
rect 30466 29016 30472 29028
rect 29788 28988 30472 29016
rect 29788 28976 29794 28988
rect 30466 28976 30472 28988
rect 30524 28976 30530 29028
rect 30558 28976 30564 29028
rect 30616 29016 30622 29028
rect 31110 29016 31116 29028
rect 30616 28988 31116 29016
rect 30616 28976 30622 28988
rect 31110 28976 31116 28988
rect 31168 28976 31174 29028
rect 31220 29016 31248 29056
rect 31297 29053 31309 29087
rect 31343 29084 31355 29087
rect 32416 29084 32444 29124
rect 32490 29112 32496 29124
rect 32577 29152 32589 29155
rect 32577 29124 32996 29152
rect 32577 29121 32589 29124
rect 32548 29115 32589 29121
rect 32548 29112 32554 29115
rect 31343 29056 32444 29084
rect 32769 29087 32827 29093
rect 31343 29053 31355 29056
rect 31297 29047 31355 29053
rect 32769 29053 32781 29087
rect 32815 29053 32827 29087
rect 32769 29047 32827 29053
rect 32784 29016 32812 29047
rect 32858 29044 32864 29096
rect 32916 29044 32922 29096
rect 32968 29084 32996 29124
rect 33042 29112 33048 29164
rect 33100 29112 33106 29164
rect 33152 29152 33180 29180
rect 33229 29155 33287 29161
rect 33229 29152 33241 29155
rect 33152 29124 33241 29152
rect 33229 29121 33241 29124
rect 33275 29121 33287 29155
rect 33336 29152 33364 29260
rect 33410 29248 33416 29300
rect 33468 29288 33474 29300
rect 35158 29288 35164 29300
rect 33468 29260 35164 29288
rect 33468 29248 33474 29260
rect 35158 29248 35164 29260
rect 35216 29248 35222 29300
rect 39114 29248 39120 29300
rect 39172 29248 39178 29300
rect 33686 29180 33692 29232
rect 33744 29180 33750 29232
rect 35894 29220 35900 29232
rect 34716 29192 35900 29220
rect 33413 29155 33471 29161
rect 33413 29152 33425 29155
rect 33336 29124 33425 29152
rect 33229 29115 33287 29121
rect 33413 29121 33425 29124
rect 33459 29121 33471 29155
rect 33413 29115 33471 29121
rect 34057 29155 34115 29161
rect 34057 29121 34069 29155
rect 34103 29121 34115 29155
rect 34057 29115 34115 29121
rect 34072 29084 34100 29115
rect 34422 29112 34428 29164
rect 34480 29112 34486 29164
rect 34716 29161 34744 29192
rect 35894 29180 35900 29192
rect 35952 29180 35958 29232
rect 34701 29155 34759 29161
rect 34701 29121 34713 29155
rect 34747 29121 34759 29155
rect 34701 29115 34759 29121
rect 34808 29124 35940 29152
rect 34808 29084 34836 29124
rect 35912 29096 35940 29124
rect 35986 29112 35992 29164
rect 36044 29152 36050 29164
rect 37277 29155 37335 29161
rect 37277 29152 37289 29155
rect 36044 29124 37289 29152
rect 36044 29112 36050 29124
rect 37277 29121 37289 29124
rect 37323 29121 37335 29155
rect 37277 29115 37335 29121
rect 37458 29112 37464 29164
rect 37516 29152 37522 29164
rect 37553 29155 37611 29161
rect 37553 29152 37565 29155
rect 37516 29124 37565 29152
rect 37516 29112 37522 29124
rect 37553 29121 37565 29124
rect 37599 29152 37611 29155
rect 37642 29152 37648 29164
rect 37599 29124 37648 29152
rect 37599 29121 37611 29124
rect 37553 29115 37611 29121
rect 37642 29112 37648 29124
rect 37700 29112 37706 29164
rect 38381 29155 38439 29161
rect 38381 29121 38393 29155
rect 38427 29152 38439 29155
rect 39132 29152 39160 29248
rect 38427 29124 39160 29152
rect 38427 29121 38439 29124
rect 38381 29115 38439 29121
rect 32968 29056 34836 29084
rect 34882 29044 34888 29096
rect 34940 29044 34946 29096
rect 35158 29044 35164 29096
rect 35216 29044 35222 29096
rect 35894 29044 35900 29096
rect 35952 29084 35958 29096
rect 37476 29084 37504 29112
rect 35952 29056 37504 29084
rect 35952 29044 35958 29056
rect 31220 28988 32812 29016
rect 34974 28976 34980 29028
rect 35032 29016 35038 29028
rect 35032 28988 37320 29016
rect 35032 28976 35038 28988
rect 29822 28948 29828 28960
rect 29657 28920 29828 28948
rect 29549 28911 29607 28917
rect 29822 28908 29828 28920
rect 29880 28908 29886 28960
rect 32030 28908 32036 28960
rect 32088 28948 32094 28960
rect 32306 28948 32312 28960
rect 32088 28920 32312 28948
rect 32088 28908 32094 28920
rect 32306 28908 32312 28920
rect 32364 28908 32370 28960
rect 32582 28908 32588 28960
rect 32640 28948 32646 28960
rect 32950 28948 32956 28960
rect 32640 28920 32956 28948
rect 32640 28908 32646 28920
rect 32950 28908 32956 28920
rect 33008 28908 33014 28960
rect 33594 28908 33600 28960
rect 33652 28948 33658 28960
rect 35250 28948 35256 28960
rect 33652 28920 35256 28948
rect 33652 28908 33658 28920
rect 35250 28908 35256 28920
rect 35308 28908 35314 28960
rect 37292 28948 37320 28988
rect 37366 28976 37372 29028
rect 37424 29016 37430 29028
rect 37553 29019 37611 29025
rect 37553 29016 37565 29019
rect 37424 28988 37565 29016
rect 37424 28976 37430 28988
rect 37553 28985 37565 28988
rect 37599 28985 37611 29019
rect 37553 28979 37611 28985
rect 38838 28976 38844 29028
rect 38896 29016 38902 29028
rect 39482 29016 39488 29028
rect 38896 28988 39488 29016
rect 38896 28976 38902 28988
rect 39482 28976 39488 28988
rect 39540 28976 39546 29028
rect 37642 28948 37648 28960
rect 37292 28920 37648 28948
rect 37642 28908 37648 28920
rect 37700 28948 37706 28960
rect 38565 28951 38623 28957
rect 38565 28948 38577 28951
rect 37700 28920 38577 28948
rect 37700 28908 37706 28920
rect 38565 28917 38577 28920
rect 38611 28917 38623 28951
rect 38565 28911 38623 28917
rect 1104 28858 41400 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 41400 28858
rect 1104 28784 41400 28806
rect 5350 28704 5356 28756
rect 5408 28744 5414 28756
rect 5445 28747 5503 28753
rect 5445 28744 5457 28747
rect 5408 28716 5457 28744
rect 5408 28704 5414 28716
rect 5445 28713 5457 28716
rect 5491 28713 5503 28747
rect 5445 28707 5503 28713
rect 5810 28704 5816 28756
rect 5868 28704 5874 28756
rect 11054 28704 11060 28756
rect 11112 28704 11118 28756
rect 12069 28747 12127 28753
rect 12069 28713 12081 28747
rect 12115 28744 12127 28747
rect 12250 28744 12256 28756
rect 12115 28716 12256 28744
rect 12115 28713 12127 28716
rect 12069 28707 12127 28713
rect 12250 28704 12256 28716
rect 12308 28704 12314 28756
rect 12710 28744 12716 28756
rect 12360 28716 12716 28744
rect 5261 28679 5319 28685
rect 5261 28645 5273 28679
rect 5307 28676 5319 28679
rect 5534 28676 5540 28688
rect 5307 28648 5540 28676
rect 5307 28645 5319 28648
rect 5261 28639 5319 28645
rect 5534 28636 5540 28648
rect 5592 28636 5598 28688
rect 1857 28611 1915 28617
rect 1857 28577 1869 28611
rect 1903 28608 1915 28611
rect 2498 28608 2504 28620
rect 1903 28580 2504 28608
rect 1903 28577 1915 28580
rect 1857 28571 1915 28577
rect 2498 28568 2504 28580
rect 2556 28568 2562 28620
rect 3050 28608 3056 28620
rect 2976 28580 3056 28608
rect 1394 28500 1400 28552
rect 1452 28540 1458 28552
rect 1581 28543 1639 28549
rect 1581 28540 1593 28543
rect 1452 28512 1593 28540
rect 1452 28500 1458 28512
rect 1581 28509 1593 28512
rect 1627 28509 1639 28543
rect 2976 28526 3004 28580
rect 3050 28568 3056 28580
rect 3108 28568 3114 28620
rect 4798 28568 4804 28620
rect 4856 28608 4862 28620
rect 4985 28611 5043 28617
rect 4985 28608 4997 28611
rect 4856 28580 4997 28608
rect 4856 28568 4862 28580
rect 4985 28577 4997 28580
rect 5031 28577 5043 28611
rect 4985 28571 5043 28577
rect 1581 28503 1639 28509
rect 5166 28500 5172 28552
rect 5224 28540 5230 28552
rect 5537 28543 5595 28549
rect 5537 28540 5549 28543
rect 5224 28512 5549 28540
rect 5224 28500 5230 28512
rect 5537 28509 5549 28512
rect 5583 28509 5595 28543
rect 5537 28503 5595 28509
rect 5721 28543 5779 28549
rect 5721 28509 5733 28543
rect 5767 28540 5779 28543
rect 5828 28540 5856 28704
rect 8294 28636 8300 28688
rect 8352 28676 8358 28688
rect 10962 28676 10968 28688
rect 8352 28648 10968 28676
rect 8352 28636 8358 28648
rect 7745 28611 7803 28617
rect 7745 28577 7757 28611
rect 7791 28608 7803 28611
rect 7834 28608 7840 28620
rect 7791 28580 7840 28608
rect 7791 28577 7803 28580
rect 7745 28571 7803 28577
rect 7834 28568 7840 28580
rect 7892 28568 7898 28620
rect 5767 28512 5856 28540
rect 5767 28509 5779 28512
rect 5721 28503 5779 28509
rect 5902 28500 5908 28552
rect 5960 28500 5966 28552
rect 6638 28500 6644 28552
rect 6696 28540 6702 28552
rect 7558 28540 7564 28552
rect 6696 28512 7564 28540
rect 6696 28500 6702 28512
rect 7558 28500 7564 28512
rect 7616 28540 7622 28552
rect 9876 28549 9904 28648
rect 10962 28636 10968 28648
rect 11020 28636 11026 28688
rect 11072 28676 11100 28704
rect 12360 28676 12388 28716
rect 12710 28704 12716 28716
rect 12768 28704 12774 28756
rect 14274 28744 14280 28756
rect 12912 28716 14280 28744
rect 12912 28676 12940 28716
rect 14274 28704 14280 28716
rect 14332 28704 14338 28756
rect 15010 28744 15016 28756
rect 14752 28716 15016 28744
rect 11072 28648 12388 28676
rect 12544 28648 12940 28676
rect 10152 28580 12112 28608
rect 9861 28543 9919 28549
rect 7616 28512 7972 28540
rect 7616 28500 7622 28512
rect 3602 28432 3608 28484
rect 3660 28432 3666 28484
rect 5258 28432 5264 28484
rect 5316 28472 5322 28484
rect 5813 28475 5871 28481
rect 5813 28472 5825 28475
rect 5316 28444 5825 28472
rect 5316 28432 5322 28444
rect 5813 28441 5825 28444
rect 5859 28472 5871 28475
rect 6656 28472 6684 28500
rect 5859 28444 6684 28472
rect 5859 28441 5871 28444
rect 5813 28435 5871 28441
rect 7374 28432 7380 28484
rect 7432 28472 7438 28484
rect 7837 28475 7895 28481
rect 7837 28472 7849 28475
rect 7432 28444 7849 28472
rect 7432 28432 7438 28444
rect 7837 28441 7849 28444
rect 7883 28441 7895 28475
rect 7944 28472 7972 28512
rect 9861 28509 9873 28543
rect 9907 28509 9919 28543
rect 9861 28503 9919 28509
rect 10042 28500 10048 28552
rect 10100 28500 10106 28552
rect 10152 28549 10180 28580
rect 10137 28543 10195 28549
rect 10137 28509 10149 28543
rect 10183 28509 10195 28543
rect 10137 28503 10195 28509
rect 10152 28472 10180 28503
rect 10226 28500 10232 28552
rect 10284 28500 10290 28552
rect 10689 28543 10747 28549
rect 10689 28509 10701 28543
rect 10735 28540 10747 28543
rect 11057 28543 11115 28549
rect 10735 28512 11008 28540
rect 10735 28509 10747 28512
rect 10689 28503 10747 28509
rect 7944 28444 10180 28472
rect 7837 28435 7895 28441
rect 10980 28416 11008 28512
rect 11057 28509 11069 28543
rect 11103 28540 11115 28543
rect 11103 28512 11192 28540
rect 11103 28509 11115 28512
rect 11057 28503 11115 28509
rect 11164 28472 11192 28512
rect 11330 28500 11336 28552
rect 11388 28540 11394 28552
rect 11517 28543 11575 28549
rect 11517 28540 11529 28543
rect 11388 28512 11529 28540
rect 11388 28500 11394 28512
rect 11517 28509 11529 28512
rect 11563 28509 11575 28543
rect 11517 28503 11575 28509
rect 11698 28500 11704 28552
rect 11756 28500 11762 28552
rect 11885 28543 11943 28549
rect 11885 28509 11897 28543
rect 11931 28540 11943 28543
rect 11974 28540 11980 28552
rect 11931 28512 11980 28540
rect 11931 28509 11943 28512
rect 11885 28503 11943 28509
rect 11974 28500 11980 28512
rect 12032 28500 12038 28552
rect 11606 28472 11612 28484
rect 11164 28444 11612 28472
rect 11164 28416 11192 28444
rect 11606 28432 11612 28444
rect 11664 28432 11670 28484
rect 11793 28475 11851 28481
rect 11793 28441 11805 28475
rect 11839 28441 11851 28475
rect 12084 28472 12112 28580
rect 12158 28500 12164 28552
rect 12216 28540 12222 28552
rect 12544 28549 12572 28648
rect 12529 28543 12587 28549
rect 12529 28540 12541 28543
rect 12216 28512 12541 28540
rect 12216 28500 12222 28512
rect 12529 28509 12541 28512
rect 12575 28509 12587 28543
rect 12529 28503 12587 28509
rect 12710 28500 12716 28552
rect 12768 28542 12774 28552
rect 12912 28549 12940 28648
rect 13446 28636 13452 28688
rect 13504 28676 13510 28688
rect 14752 28676 14780 28716
rect 15010 28704 15016 28716
rect 15068 28704 15074 28756
rect 15562 28704 15568 28756
rect 15620 28704 15626 28756
rect 15746 28704 15752 28756
rect 15804 28744 15810 28756
rect 15841 28747 15899 28753
rect 15841 28744 15853 28747
rect 15804 28716 15853 28744
rect 15804 28704 15810 28716
rect 15841 28713 15853 28716
rect 15887 28713 15899 28747
rect 15841 28707 15899 28713
rect 16206 28704 16212 28756
rect 16264 28744 16270 28756
rect 16301 28747 16359 28753
rect 16301 28744 16313 28747
rect 16264 28716 16313 28744
rect 16264 28704 16270 28716
rect 16301 28713 16313 28716
rect 16347 28713 16359 28747
rect 16301 28707 16359 28713
rect 17034 28704 17040 28756
rect 17092 28744 17098 28756
rect 17678 28744 17684 28756
rect 17092 28716 17684 28744
rect 17092 28704 17098 28716
rect 17678 28704 17684 28716
rect 17736 28704 17742 28756
rect 18141 28747 18199 28753
rect 18141 28713 18153 28747
rect 18187 28713 18199 28747
rect 18141 28707 18199 28713
rect 13504 28648 14780 28676
rect 13504 28636 13510 28648
rect 12805 28543 12863 28549
rect 12805 28542 12817 28543
rect 12768 28514 12817 28542
rect 12768 28500 12774 28514
rect 12805 28509 12817 28514
rect 12851 28509 12863 28543
rect 12805 28503 12863 28509
rect 12897 28543 12955 28549
rect 12897 28509 12909 28543
rect 12943 28509 12955 28543
rect 12897 28503 12955 28509
rect 13078 28500 13084 28552
rect 13136 28500 13142 28552
rect 13265 28543 13323 28549
rect 13265 28509 13277 28543
rect 13311 28540 13323 28543
rect 14090 28540 14096 28552
rect 13311 28512 14096 28540
rect 13311 28509 13323 28512
rect 13265 28503 13323 28509
rect 14090 28500 14096 28512
rect 14148 28500 14154 28552
rect 14366 28500 14372 28552
rect 14424 28500 14430 28552
rect 14752 28549 14780 28648
rect 14826 28636 14832 28688
rect 14884 28676 14890 28688
rect 18156 28676 18184 28707
rect 19426 28704 19432 28756
rect 19484 28704 19490 28756
rect 19794 28744 19800 28756
rect 19536 28716 19800 28744
rect 14884 28648 18184 28676
rect 14884 28636 14890 28648
rect 14921 28611 14979 28617
rect 14921 28577 14933 28611
rect 14967 28608 14979 28611
rect 15197 28611 15255 28617
rect 15197 28608 15209 28611
rect 14967 28580 15209 28608
rect 14967 28577 14979 28580
rect 14921 28571 14979 28577
rect 15197 28577 15209 28580
rect 15243 28577 15255 28611
rect 15197 28571 15255 28577
rect 15749 28611 15807 28617
rect 15749 28577 15761 28611
rect 15795 28608 15807 28611
rect 19536 28608 19564 28716
rect 19794 28704 19800 28716
rect 19852 28704 19858 28756
rect 20441 28747 20499 28753
rect 20441 28713 20453 28747
rect 20487 28744 20499 28747
rect 20717 28747 20775 28753
rect 20717 28744 20729 28747
rect 20487 28716 20729 28744
rect 20487 28713 20499 28716
rect 20441 28707 20499 28713
rect 20717 28713 20729 28716
rect 20763 28713 20775 28747
rect 20717 28707 20775 28713
rect 21266 28704 21272 28756
rect 21324 28744 21330 28756
rect 21542 28744 21548 28756
rect 21324 28716 21548 28744
rect 21324 28704 21330 28716
rect 21542 28704 21548 28716
rect 21600 28704 21606 28756
rect 21637 28747 21695 28753
rect 21637 28713 21649 28747
rect 21683 28744 21695 28747
rect 21726 28744 21732 28756
rect 21683 28716 21732 28744
rect 21683 28713 21695 28716
rect 21637 28707 21695 28713
rect 21726 28704 21732 28716
rect 21784 28704 21790 28756
rect 21818 28704 21824 28756
rect 21876 28704 21882 28756
rect 22094 28704 22100 28756
rect 22152 28744 22158 28756
rect 22833 28747 22891 28753
rect 22833 28744 22845 28747
rect 22152 28716 22845 28744
rect 22152 28704 22158 28716
rect 22833 28713 22845 28716
rect 22879 28713 22891 28747
rect 22833 28707 22891 28713
rect 23014 28704 23020 28756
rect 23072 28704 23078 28756
rect 23293 28747 23351 28753
rect 23293 28713 23305 28747
rect 23339 28744 23351 28747
rect 24026 28744 24032 28756
rect 23339 28716 24032 28744
rect 23339 28713 23351 28716
rect 23293 28707 23351 28713
rect 24026 28704 24032 28716
rect 24084 28704 24090 28756
rect 24394 28704 24400 28756
rect 24452 28704 24458 28756
rect 24946 28704 24952 28756
rect 25004 28704 25010 28756
rect 25314 28704 25320 28756
rect 25372 28744 25378 28756
rect 25869 28747 25927 28753
rect 25869 28744 25881 28747
rect 25372 28716 25881 28744
rect 25372 28704 25378 28716
rect 25869 28713 25881 28716
rect 25915 28713 25927 28747
rect 25869 28707 25927 28713
rect 25958 28704 25964 28756
rect 26016 28744 26022 28756
rect 26053 28747 26111 28753
rect 26053 28744 26065 28747
rect 26016 28716 26065 28744
rect 26016 28704 26022 28716
rect 26053 28713 26065 28716
rect 26099 28713 26111 28747
rect 26053 28707 26111 28713
rect 26786 28704 26792 28756
rect 26844 28744 26850 28756
rect 27706 28744 27712 28756
rect 26844 28716 27712 28744
rect 26844 28704 26850 28716
rect 27706 28704 27712 28716
rect 27764 28704 27770 28756
rect 27893 28747 27951 28753
rect 27893 28713 27905 28747
rect 27939 28744 27951 28747
rect 28166 28744 28172 28756
rect 27939 28716 28172 28744
rect 27939 28713 27951 28716
rect 27893 28707 27951 28713
rect 28166 28704 28172 28716
rect 28224 28704 28230 28756
rect 28445 28747 28503 28753
rect 28445 28744 28457 28747
rect 28276 28716 28457 28744
rect 19613 28679 19671 28685
rect 19613 28645 19625 28679
rect 19659 28645 19671 28679
rect 19613 28639 19671 28645
rect 15795 28580 19564 28608
rect 15795 28577 15807 28580
rect 15749 28571 15807 28577
rect 14645 28543 14703 28549
rect 14645 28509 14657 28543
rect 14691 28509 14703 28543
rect 14645 28503 14703 28509
rect 14737 28543 14795 28549
rect 14737 28509 14749 28543
rect 14783 28509 14795 28543
rect 14737 28503 14795 28509
rect 13173 28475 13231 28481
rect 13173 28472 13185 28475
rect 12084 28444 13185 28472
rect 11793 28435 11851 28441
rect 13173 28441 13185 28444
rect 13219 28472 13231 28475
rect 14384 28472 14412 28500
rect 13219 28444 14412 28472
rect 14660 28472 14688 28503
rect 15010 28500 15016 28552
rect 15068 28500 15074 28552
rect 15102 28500 15108 28552
rect 15160 28500 15166 28552
rect 15289 28543 15347 28549
rect 15289 28509 15301 28543
rect 15335 28540 15347 28543
rect 15378 28540 15384 28552
rect 15335 28512 15384 28540
rect 15335 28509 15347 28512
rect 15289 28503 15347 28509
rect 15378 28500 15384 28512
rect 15436 28500 15442 28552
rect 15470 28500 15476 28552
rect 15528 28500 15534 28552
rect 15930 28500 15936 28552
rect 15988 28500 15994 28552
rect 16224 28549 16252 28580
rect 16209 28543 16267 28549
rect 16209 28509 16221 28543
rect 16255 28509 16267 28543
rect 16209 28503 16267 28509
rect 16393 28543 16451 28549
rect 16393 28509 16405 28543
rect 16439 28540 16451 28543
rect 17221 28543 17279 28549
rect 16439 28512 17172 28540
rect 16439 28509 16451 28512
rect 16393 28503 16451 28509
rect 15488 28472 15516 28500
rect 14660 28444 15516 28472
rect 13219 28441 13231 28444
rect 13173 28435 13231 28441
rect 5902 28364 5908 28416
rect 5960 28404 5966 28416
rect 6089 28407 6147 28413
rect 6089 28404 6101 28407
rect 5960 28376 6101 28404
rect 5960 28364 5966 28376
rect 6089 28373 6101 28376
rect 6135 28373 6147 28407
rect 6089 28367 6147 28373
rect 6178 28364 6184 28416
rect 6236 28404 6242 28416
rect 7267 28407 7325 28413
rect 7267 28404 7279 28407
rect 6236 28376 7279 28404
rect 6236 28364 6242 28376
rect 7267 28373 7279 28376
rect 7313 28373 7325 28407
rect 7267 28367 7325 28373
rect 7742 28364 7748 28416
rect 7800 28404 7806 28416
rect 8846 28404 8852 28416
rect 7800 28376 8852 28404
rect 7800 28364 7806 28376
rect 8846 28364 8852 28376
rect 8904 28364 8910 28416
rect 9858 28364 9864 28416
rect 9916 28404 9922 28416
rect 10226 28404 10232 28416
rect 9916 28376 10232 28404
rect 9916 28364 9922 28376
rect 10226 28364 10232 28376
rect 10284 28364 10290 28416
rect 10413 28407 10471 28413
rect 10413 28373 10425 28407
rect 10459 28404 10471 28407
rect 10502 28404 10508 28416
rect 10459 28376 10508 28404
rect 10459 28373 10471 28376
rect 10413 28367 10471 28373
rect 10502 28364 10508 28376
rect 10560 28364 10566 28416
rect 10962 28364 10968 28416
rect 11020 28364 11026 28416
rect 11146 28364 11152 28416
rect 11204 28364 11210 28416
rect 11238 28364 11244 28416
rect 11296 28364 11302 28416
rect 11514 28364 11520 28416
rect 11572 28404 11578 28416
rect 11808 28404 11836 28435
rect 15562 28432 15568 28484
rect 15620 28472 15626 28484
rect 15838 28472 15844 28484
rect 15620 28444 15844 28472
rect 15620 28432 15626 28444
rect 15838 28432 15844 28444
rect 15896 28432 15902 28484
rect 17037 28475 17095 28481
rect 17037 28441 17049 28475
rect 17083 28441 17095 28475
rect 17037 28435 17095 28441
rect 11572 28376 11836 28404
rect 11572 28364 11578 28376
rect 11974 28364 11980 28416
rect 12032 28404 12038 28416
rect 12345 28407 12403 28413
rect 12345 28404 12357 28407
rect 12032 28376 12357 28404
rect 12032 28364 12038 28376
rect 12345 28373 12357 28376
rect 12391 28373 12403 28407
rect 12345 28367 12403 28373
rect 12618 28364 12624 28416
rect 12676 28404 12682 28416
rect 12713 28407 12771 28413
rect 12713 28404 12725 28407
rect 12676 28376 12725 28404
rect 12676 28364 12682 28376
rect 12713 28373 12725 28376
rect 12759 28373 12771 28407
rect 12713 28367 12771 28373
rect 13262 28364 13268 28416
rect 13320 28404 13326 28416
rect 13449 28407 13507 28413
rect 13449 28404 13461 28407
rect 13320 28376 13461 28404
rect 13320 28364 13326 28376
rect 13449 28373 13461 28376
rect 13495 28373 13507 28407
rect 13449 28367 13507 28373
rect 14461 28407 14519 28413
rect 14461 28373 14473 28407
rect 14507 28404 14519 28407
rect 14826 28404 14832 28416
rect 14507 28376 14832 28404
rect 14507 28373 14519 28376
rect 14461 28367 14519 28373
rect 14826 28364 14832 28376
rect 14884 28364 14890 28416
rect 14918 28364 14924 28416
rect 14976 28404 14982 28416
rect 17052 28404 17080 28435
rect 14976 28376 17080 28404
rect 17144 28404 17172 28512
rect 17221 28509 17233 28543
rect 17267 28540 17279 28543
rect 17402 28540 17408 28552
rect 17267 28512 17408 28540
rect 17267 28509 17279 28512
rect 17221 28503 17279 28509
rect 17402 28500 17408 28512
rect 17460 28500 17466 28552
rect 18138 28500 18144 28552
rect 18196 28500 18202 28552
rect 18230 28500 18236 28552
rect 18288 28540 18294 28552
rect 18325 28543 18383 28549
rect 18325 28540 18337 28543
rect 18288 28512 18337 28540
rect 18288 28500 18294 28512
rect 18325 28509 18337 28512
rect 18371 28509 18383 28543
rect 18325 28503 18383 28509
rect 17494 28432 17500 28484
rect 17552 28432 17558 28484
rect 17678 28432 17684 28484
rect 17736 28432 17742 28484
rect 18340 28472 18368 28503
rect 18506 28500 18512 28552
rect 18564 28540 18570 28552
rect 19628 28540 19656 28639
rect 19886 28636 19892 28688
rect 19944 28636 19950 28688
rect 19981 28679 20039 28685
rect 19981 28645 19993 28679
rect 20027 28676 20039 28679
rect 21836 28676 21864 28704
rect 22554 28676 22560 28688
rect 20027 28648 21864 28676
rect 22020 28648 22560 28676
rect 20027 28645 20039 28648
rect 19981 28639 20039 28645
rect 19904 28549 19932 28636
rect 20165 28611 20223 28617
rect 20165 28577 20177 28611
rect 20211 28608 20223 28611
rect 20211 28580 20392 28608
rect 20211 28577 20223 28580
rect 20165 28571 20223 28577
rect 20364 28552 20392 28580
rect 21174 28568 21180 28620
rect 21232 28617 21238 28620
rect 21232 28597 21241 28617
rect 22020 28608 22048 28648
rect 22554 28636 22560 28648
rect 22612 28636 22618 28688
rect 23032 28676 23060 28704
rect 23032 28648 23152 28676
rect 21284 28597 22048 28608
rect 21232 28580 22048 28597
rect 21232 28569 21312 28580
rect 21232 28568 21238 28569
rect 18564 28512 19656 28540
rect 19889 28543 19947 28549
rect 18564 28500 18570 28512
rect 19889 28509 19901 28543
rect 19935 28540 19947 28543
rect 20257 28543 20315 28549
rect 20257 28540 20269 28543
rect 19935 28512 20269 28540
rect 19935 28509 19947 28512
rect 19889 28503 19947 28509
rect 20257 28509 20269 28512
rect 20303 28509 20315 28543
rect 20257 28503 20315 28509
rect 20346 28500 20352 28552
rect 20404 28500 20410 28552
rect 20441 28543 20499 28549
rect 20441 28509 20453 28543
rect 20487 28509 20499 28543
rect 20441 28503 20499 28509
rect 20901 28543 20959 28549
rect 20901 28509 20913 28543
rect 20947 28542 20959 28543
rect 20990 28542 20996 28552
rect 20947 28514 20996 28542
rect 20947 28509 20959 28514
rect 20901 28503 20959 28509
rect 19150 28472 19156 28484
rect 18340 28444 19156 28472
rect 19150 28432 19156 28444
rect 19208 28432 19214 28484
rect 19242 28432 19248 28484
rect 19300 28432 19306 28484
rect 19518 28481 19524 28484
rect 19461 28475 19524 28481
rect 19461 28441 19473 28475
rect 19507 28441 19524 28475
rect 19461 28435 19524 28441
rect 19518 28432 19524 28435
rect 19576 28432 19582 28484
rect 19794 28432 19800 28484
rect 19852 28472 19858 28484
rect 20456 28472 20484 28503
rect 20990 28500 20996 28514
rect 21048 28500 21054 28552
rect 21082 28500 21088 28552
rect 21140 28500 21146 28552
rect 21450 28500 21456 28552
rect 21508 28500 21514 28552
rect 21542 28500 21548 28552
rect 21600 28540 21606 28552
rect 22020 28549 22048 28580
rect 22094 28568 22100 28620
rect 22152 28608 22158 28620
rect 22189 28611 22247 28617
rect 22189 28608 22201 28611
rect 22152 28580 22201 28608
rect 22152 28568 22158 28580
rect 22189 28577 22201 28580
rect 22235 28608 22247 28611
rect 22462 28608 22468 28620
rect 22235 28580 22468 28608
rect 22235 28577 22247 28580
rect 22189 28571 22247 28577
rect 22462 28568 22468 28580
rect 22520 28568 22526 28620
rect 21729 28543 21787 28549
rect 21729 28540 21741 28543
rect 21600 28512 21741 28540
rect 21600 28500 21606 28512
rect 21729 28509 21741 28512
rect 21775 28509 21787 28543
rect 21729 28503 21787 28509
rect 22005 28543 22063 28549
rect 22005 28509 22017 28543
rect 22051 28509 22063 28543
rect 22005 28503 22063 28509
rect 22281 28543 22339 28549
rect 22281 28509 22293 28543
rect 22327 28509 22339 28543
rect 22281 28503 22339 28509
rect 19852 28444 20484 28472
rect 19852 28432 19858 28444
rect 21266 28432 21272 28484
rect 21324 28432 21330 28484
rect 21468 28472 21496 28500
rect 22186 28472 22192 28484
rect 21468 28444 22192 28472
rect 22186 28432 22192 28444
rect 22244 28472 22250 28484
rect 22296 28472 22324 28503
rect 22554 28500 22560 28552
rect 22612 28540 22618 28552
rect 22833 28543 22891 28549
rect 22833 28540 22845 28543
rect 22612 28512 22845 28540
rect 22612 28500 22618 28512
rect 22833 28509 22845 28512
rect 22879 28509 22891 28543
rect 22833 28503 22891 28509
rect 23014 28500 23020 28552
rect 23072 28500 23078 28552
rect 23124 28549 23152 28648
rect 23566 28636 23572 28688
rect 23624 28636 23630 28688
rect 24412 28676 24440 28704
rect 23952 28648 24440 28676
rect 23109 28543 23167 28549
rect 23109 28509 23121 28543
rect 23155 28509 23167 28543
rect 23109 28503 23167 28509
rect 23382 28500 23388 28552
rect 23440 28500 23446 28552
rect 23474 28500 23480 28552
rect 23532 28500 23538 28552
rect 23658 28500 23664 28552
rect 23716 28500 23722 28552
rect 23750 28500 23756 28552
rect 23808 28500 23814 28552
rect 23845 28543 23903 28549
rect 23845 28509 23857 28543
rect 23891 28540 23903 28543
rect 23952 28540 23980 28648
rect 24486 28636 24492 28688
rect 24544 28676 24550 28688
rect 28276 28676 28304 28716
rect 28445 28713 28457 28716
rect 28491 28713 28503 28747
rect 28445 28707 28503 28713
rect 28718 28704 28724 28756
rect 28776 28744 28782 28756
rect 28813 28747 28871 28753
rect 28813 28744 28825 28747
rect 28776 28716 28825 28744
rect 28776 28704 28782 28716
rect 28813 28713 28825 28716
rect 28859 28713 28871 28747
rect 29178 28744 29184 28756
rect 28813 28707 28871 28713
rect 29012 28716 29184 28744
rect 29012 28676 29040 28716
rect 29178 28704 29184 28716
rect 29236 28704 29242 28756
rect 29454 28704 29460 28756
rect 29512 28744 29518 28756
rect 30006 28744 30012 28756
rect 29512 28716 30012 28744
rect 29512 28704 29518 28716
rect 30006 28704 30012 28716
rect 30064 28744 30070 28756
rect 31018 28744 31024 28756
rect 30064 28716 31024 28744
rect 30064 28704 30070 28716
rect 31018 28704 31024 28716
rect 31076 28704 31082 28756
rect 36262 28704 36268 28756
rect 36320 28744 36326 28756
rect 36722 28744 36728 28756
rect 36320 28716 36728 28744
rect 36320 28704 36326 28716
rect 36722 28704 36728 28716
rect 36780 28744 36786 28756
rect 36909 28747 36967 28753
rect 36909 28744 36921 28747
rect 36780 28716 36921 28744
rect 36780 28704 36786 28716
rect 36909 28713 36921 28716
rect 36955 28713 36967 28747
rect 36909 28707 36967 28713
rect 24544 28648 28304 28676
rect 28645 28648 29040 28676
rect 24544 28636 24550 28648
rect 26878 28608 26884 28620
rect 26160 28580 26740 28608
rect 24397 28543 24455 28549
rect 23891 28512 23980 28540
rect 24029 28537 24087 28543
rect 23891 28509 23903 28512
rect 23845 28503 23903 28509
rect 24029 28503 24041 28537
rect 24075 28503 24087 28537
rect 24397 28509 24409 28543
rect 24443 28509 24455 28543
rect 24397 28503 24455 28509
rect 24765 28543 24823 28549
rect 24765 28509 24777 28543
rect 24811 28540 24823 28543
rect 24854 28540 24860 28552
rect 24811 28512 24860 28540
rect 24811 28509 24823 28512
rect 24765 28503 24823 28509
rect 22244 28444 22784 28472
rect 22244 28432 22250 28444
rect 22756 28416 22784 28444
rect 17402 28404 17408 28416
rect 17144 28376 17408 28404
rect 14976 28364 14982 28376
rect 17402 28364 17408 28376
rect 17460 28404 17466 28416
rect 17773 28407 17831 28413
rect 17773 28404 17785 28407
rect 17460 28376 17785 28404
rect 17460 28364 17466 28376
rect 17773 28373 17785 28376
rect 17819 28373 17831 28407
rect 17773 28367 17831 28373
rect 18506 28364 18512 28416
rect 18564 28404 18570 28416
rect 20165 28407 20223 28413
rect 20165 28404 20177 28407
rect 18564 28376 20177 28404
rect 18564 28364 18570 28376
rect 20165 28373 20177 28376
rect 20211 28373 20223 28407
rect 20165 28367 20223 28373
rect 20625 28407 20683 28413
rect 20625 28373 20637 28407
rect 20671 28404 20683 28407
rect 20714 28404 20720 28416
rect 20671 28376 20720 28404
rect 20671 28373 20683 28376
rect 20625 28367 20683 28373
rect 20714 28364 20720 28376
rect 20772 28364 20778 28416
rect 22738 28364 22744 28416
rect 22796 28364 22802 28416
rect 23492 28404 23520 28500
rect 24029 28497 24087 28503
rect 23937 28475 23995 28481
rect 23937 28472 23949 28475
rect 23768 28444 23949 28472
rect 23768 28404 23796 28444
rect 23937 28441 23949 28444
rect 23983 28441 23995 28475
rect 23937 28435 23995 28441
rect 24044 28416 24072 28497
rect 23492 28376 23796 28404
rect 24026 28364 24032 28416
rect 24084 28364 24090 28416
rect 24412 28404 24440 28503
rect 24854 28500 24860 28512
rect 24912 28500 24918 28552
rect 25038 28500 25044 28552
rect 25096 28500 25102 28552
rect 25314 28500 25320 28552
rect 25372 28540 25378 28552
rect 25409 28543 25467 28549
rect 25409 28540 25421 28543
rect 25372 28512 25421 28540
rect 25372 28500 25378 28512
rect 25409 28509 25421 28512
rect 25455 28509 25467 28543
rect 25409 28503 25467 28509
rect 25498 28500 25504 28552
rect 25556 28500 25562 28552
rect 26160 28549 26188 28580
rect 26712 28552 26740 28580
rect 26804 28580 26884 28608
rect 25593 28543 25651 28549
rect 25593 28509 25605 28543
rect 25639 28540 25651 28543
rect 26145 28543 26203 28549
rect 25639 28512 25820 28540
rect 25639 28509 25651 28512
rect 25593 28503 25651 28509
rect 24486 28432 24492 28484
rect 24544 28472 24550 28484
rect 24581 28475 24639 28481
rect 24581 28472 24593 28475
rect 24544 28444 24593 28472
rect 24544 28432 24550 28444
rect 24581 28441 24593 28444
rect 24627 28441 24639 28475
rect 24581 28435 24639 28441
rect 24673 28475 24731 28481
rect 24673 28441 24685 28475
rect 24719 28472 24731 28475
rect 24946 28472 24952 28484
rect 24719 28444 24952 28472
rect 24719 28441 24731 28444
rect 24673 28435 24731 28441
rect 24946 28432 24952 28444
rect 25004 28432 25010 28484
rect 25056 28472 25084 28500
rect 25608 28472 25636 28503
rect 25056 28444 25636 28472
rect 25685 28475 25743 28481
rect 25685 28441 25697 28475
rect 25731 28441 25743 28475
rect 25792 28472 25820 28512
rect 26145 28509 26157 28543
rect 26191 28509 26203 28543
rect 26145 28503 26203 28509
rect 26418 28500 26424 28552
rect 26476 28500 26482 28552
rect 26513 28543 26571 28549
rect 26513 28509 26525 28543
rect 26559 28540 26571 28543
rect 26602 28540 26608 28552
rect 26559 28512 26608 28540
rect 26559 28509 26571 28512
rect 26513 28503 26571 28509
rect 26602 28500 26608 28512
rect 26660 28500 26666 28552
rect 26694 28500 26700 28552
rect 26752 28500 26758 28552
rect 26804 28549 26832 28580
rect 26878 28568 26884 28580
rect 26936 28568 26942 28620
rect 27985 28611 28043 28617
rect 27985 28608 27997 28611
rect 27080 28580 27292 28608
rect 27080 28549 27108 28580
rect 27264 28552 27292 28580
rect 27356 28580 27997 28608
rect 26789 28543 26847 28549
rect 26789 28509 26801 28543
rect 26835 28509 26847 28543
rect 26973 28543 27031 28549
rect 26973 28534 26985 28543
rect 26896 28518 26985 28534
rect 26789 28503 26847 28509
rect 25792 28444 26004 28472
rect 25685 28435 25743 28441
rect 24762 28404 24768 28416
rect 24412 28376 24768 28404
rect 24762 28364 24768 28376
rect 24820 28364 24826 28416
rect 25222 28364 25228 28416
rect 25280 28404 25286 28416
rect 25700 28404 25728 28435
rect 25280 28376 25728 28404
rect 25280 28364 25286 28376
rect 25866 28364 25872 28416
rect 25924 28413 25930 28416
rect 25924 28407 25943 28413
rect 25931 28373 25943 28407
rect 25976 28404 26004 28444
rect 26234 28432 26240 28484
rect 26292 28472 26298 28484
rect 26329 28475 26387 28481
rect 26329 28472 26341 28475
rect 26292 28444 26341 28472
rect 26292 28432 26298 28444
rect 26329 28441 26341 28444
rect 26375 28441 26387 28475
rect 26878 28466 26884 28518
rect 26936 28509 26985 28518
rect 27019 28509 27031 28543
rect 26936 28506 27031 28509
rect 26936 28466 26942 28506
rect 26973 28503 27031 28506
rect 27065 28543 27123 28549
rect 27065 28509 27077 28543
rect 27111 28509 27123 28543
rect 27065 28503 27123 28509
rect 27154 28500 27160 28552
rect 27212 28500 27218 28552
rect 27246 28500 27252 28552
rect 27304 28500 27310 28552
rect 27356 28472 27384 28580
rect 27985 28577 27997 28580
rect 28031 28577 28043 28611
rect 28645 28608 28673 28648
rect 27985 28571 28043 28577
rect 28552 28580 28673 28608
rect 27430 28500 27436 28552
rect 27488 28500 27494 28552
rect 27522 28500 27528 28552
rect 27580 28500 27586 28552
rect 27709 28543 27767 28549
rect 27709 28509 27721 28543
rect 27755 28509 27767 28543
rect 27709 28503 27767 28509
rect 26329 28435 26387 28441
rect 27176 28444 27384 28472
rect 27448 28472 27476 28500
rect 27724 28472 27752 28503
rect 27448 28444 27752 28472
rect 26697 28407 26755 28413
rect 26697 28404 26709 28407
rect 25976 28376 26709 28404
rect 25924 28367 25943 28373
rect 26697 28373 26709 28376
rect 26743 28373 26755 28407
rect 26697 28367 26755 28373
rect 25924 28364 25930 28367
rect 26878 28364 26884 28416
rect 26936 28404 26942 28416
rect 27176 28404 27204 28444
rect 26936 28376 27204 28404
rect 26936 28364 26942 28376
rect 27246 28364 27252 28416
rect 27304 28404 27310 28416
rect 27341 28407 27399 28413
rect 27341 28404 27353 28407
rect 27304 28376 27353 28404
rect 27304 28364 27310 28376
rect 27341 28373 27353 28376
rect 27387 28373 27399 28407
rect 27341 28367 27399 28373
rect 27522 28364 27528 28416
rect 27580 28404 27586 28416
rect 27706 28404 27712 28416
rect 27580 28376 27712 28404
rect 27580 28364 27586 28376
rect 27706 28364 27712 28376
rect 27764 28364 27770 28416
rect 28000 28404 28028 28571
rect 28099 28556 28157 28562
rect 28099 28553 28111 28556
rect 28092 28522 28111 28553
rect 28145 28542 28157 28556
rect 28350 28542 28356 28552
rect 28145 28522 28356 28542
rect 28092 28514 28356 28522
rect 28350 28500 28356 28514
rect 28408 28500 28414 28552
rect 28445 28543 28503 28549
rect 28445 28509 28457 28543
rect 28491 28540 28503 28543
rect 28552 28540 28580 28580
rect 28491 28512 28580 28540
rect 28629 28543 28687 28549
rect 28491 28509 28503 28512
rect 28445 28503 28503 28509
rect 28629 28509 28641 28543
rect 28675 28509 28687 28543
rect 28629 28503 28687 28509
rect 28166 28432 28172 28484
rect 28224 28432 28230 28484
rect 28184 28404 28212 28432
rect 28000 28376 28212 28404
rect 28258 28364 28264 28416
rect 28316 28364 28322 28416
rect 28350 28364 28356 28416
rect 28408 28404 28414 28416
rect 28645 28404 28673 28503
rect 28902 28500 28908 28552
rect 28960 28540 28966 28552
rect 29012 28540 29040 28648
rect 29086 28636 29092 28688
rect 29144 28676 29150 28688
rect 32309 28679 32367 28685
rect 32309 28676 32321 28679
rect 29144 28648 32321 28676
rect 29144 28636 29150 28648
rect 32309 28645 32321 28648
rect 32355 28645 32367 28679
rect 34330 28676 34336 28688
rect 32309 28639 32367 28645
rect 33796 28648 34336 28676
rect 29362 28568 29368 28620
rect 29420 28608 29426 28620
rect 33686 28608 33692 28620
rect 29420 28580 33692 28608
rect 29420 28568 29426 28580
rect 33686 28568 33692 28580
rect 33744 28568 33750 28620
rect 28960 28512 29040 28540
rect 28960 28500 28966 28512
rect 29178 28500 29184 28552
rect 29236 28549 29242 28552
rect 29236 28503 29244 28549
rect 29236 28500 29242 28503
rect 29822 28500 29828 28552
rect 29880 28540 29886 28552
rect 31021 28543 31079 28549
rect 31021 28540 31033 28543
rect 29880 28512 31033 28540
rect 29880 28500 29886 28512
rect 31021 28509 31033 28512
rect 31067 28540 31079 28543
rect 31202 28540 31208 28552
rect 31067 28512 31208 28540
rect 31067 28509 31079 28512
rect 31021 28503 31079 28509
rect 31202 28500 31208 28512
rect 31260 28500 31266 28552
rect 31386 28500 31392 28552
rect 31444 28540 31450 28552
rect 31481 28543 31539 28549
rect 31481 28540 31493 28543
rect 31444 28512 31493 28540
rect 31444 28500 31450 28512
rect 31481 28509 31493 28512
rect 31527 28509 31539 28543
rect 31481 28503 31539 28509
rect 31665 28543 31723 28549
rect 31665 28509 31677 28543
rect 31711 28540 31723 28543
rect 32030 28540 32036 28552
rect 31711 28512 32036 28540
rect 31711 28509 31723 28512
rect 31665 28503 31723 28509
rect 32030 28500 32036 28512
rect 32088 28500 32094 28552
rect 32585 28543 32643 28549
rect 32585 28509 32597 28543
rect 32631 28540 32643 28543
rect 32766 28540 32772 28552
rect 32631 28512 32772 28540
rect 32631 28509 32643 28512
rect 32585 28503 32643 28509
rect 32766 28500 32772 28512
rect 32824 28500 32830 28552
rect 33796 28549 33824 28648
rect 34330 28636 34336 28648
rect 34388 28636 34394 28688
rect 34698 28636 34704 28688
rect 34756 28636 34762 28688
rect 37826 28676 37832 28688
rect 35728 28648 37832 28676
rect 34514 28608 34520 28620
rect 34164 28580 34520 28608
rect 34164 28552 34192 28580
rect 34514 28568 34520 28580
rect 34572 28608 34578 28620
rect 35253 28611 35311 28617
rect 34572 28580 35112 28608
rect 34572 28568 34578 28580
rect 33505 28543 33563 28549
rect 33505 28509 33517 28543
rect 33551 28509 33563 28543
rect 33505 28503 33563 28509
rect 33781 28543 33839 28549
rect 33781 28509 33793 28543
rect 33827 28509 33839 28543
rect 33781 28503 33839 28509
rect 28813 28475 28871 28481
rect 28813 28441 28825 28475
rect 28859 28441 28871 28475
rect 28813 28435 28871 28441
rect 28408 28376 28673 28404
rect 28828 28404 28856 28435
rect 28994 28432 29000 28484
rect 29052 28432 29058 28484
rect 29089 28475 29147 28481
rect 29089 28441 29101 28475
rect 29135 28472 29147 28475
rect 29638 28472 29644 28484
rect 29135 28444 29644 28472
rect 29135 28441 29147 28444
rect 29089 28435 29147 28441
rect 29638 28432 29644 28444
rect 29696 28432 29702 28484
rect 31036 28444 31616 28472
rect 31036 28416 31064 28444
rect 29178 28404 29184 28416
rect 28828 28376 29184 28404
rect 28408 28364 28414 28376
rect 29178 28364 29184 28376
rect 29236 28364 29242 28416
rect 31018 28364 31024 28416
rect 31076 28364 31082 28416
rect 31297 28407 31355 28413
rect 31297 28373 31309 28407
rect 31343 28404 31355 28407
rect 31386 28404 31392 28416
rect 31343 28376 31392 28404
rect 31343 28373 31355 28376
rect 31297 28367 31355 28373
rect 31386 28364 31392 28376
rect 31444 28364 31450 28416
rect 31588 28413 31616 28444
rect 32122 28432 32128 28484
rect 32180 28432 32186 28484
rect 32309 28475 32367 28481
rect 32309 28441 32321 28475
rect 32355 28472 32367 28475
rect 33520 28472 33548 28503
rect 34146 28500 34152 28552
rect 34204 28500 34210 28552
rect 34790 28500 34796 28552
rect 34848 28540 34854 28552
rect 34885 28543 34943 28549
rect 34885 28540 34897 28543
rect 34848 28512 34897 28540
rect 34848 28500 34854 28512
rect 34885 28509 34897 28512
rect 34931 28509 34943 28543
rect 34885 28503 34943 28509
rect 34974 28500 34980 28552
rect 35032 28500 35038 28552
rect 35084 28540 35112 28580
rect 35253 28577 35265 28611
rect 35299 28608 35311 28611
rect 35342 28608 35348 28620
rect 35299 28580 35348 28608
rect 35299 28577 35311 28580
rect 35253 28571 35311 28577
rect 35342 28568 35348 28580
rect 35400 28568 35406 28620
rect 35084 28512 35388 28540
rect 35360 28481 35388 28512
rect 35526 28500 35532 28552
rect 35584 28540 35590 28552
rect 35728 28549 35756 28648
rect 37826 28636 37832 28648
rect 37884 28636 37890 28688
rect 35820 28580 36952 28608
rect 35820 28552 35848 28580
rect 35713 28543 35771 28549
rect 35713 28540 35725 28543
rect 35584 28512 35725 28540
rect 35584 28500 35590 28512
rect 35713 28509 35725 28512
rect 35759 28509 35771 28543
rect 35713 28503 35771 28509
rect 35802 28500 35808 28552
rect 35860 28500 35866 28552
rect 36924 28549 36952 28580
rect 35897 28543 35955 28549
rect 35897 28509 35909 28543
rect 35943 28509 35955 28543
rect 35897 28503 35955 28509
rect 36909 28543 36967 28549
rect 36909 28509 36921 28543
rect 36955 28509 36967 28543
rect 36909 28503 36967 28509
rect 37093 28543 37151 28549
rect 37093 28509 37105 28543
rect 37139 28540 37151 28543
rect 37550 28540 37556 28552
rect 37139 28512 37556 28540
rect 37139 28509 37151 28512
rect 37093 28503 37151 28509
rect 35345 28475 35403 28481
rect 32355 28444 35296 28472
rect 32355 28441 32367 28444
rect 32309 28435 32367 28441
rect 31573 28407 31631 28413
rect 31573 28373 31585 28407
rect 31619 28373 31631 28407
rect 32140 28404 32168 28432
rect 32493 28407 32551 28413
rect 32493 28404 32505 28407
rect 32140 28376 32505 28404
rect 31573 28367 31631 28373
rect 32493 28373 32505 28376
rect 32539 28373 32551 28407
rect 32493 28367 32551 28373
rect 32582 28364 32588 28416
rect 32640 28404 32646 28416
rect 33597 28407 33655 28413
rect 33597 28404 33609 28407
rect 32640 28376 33609 28404
rect 32640 28364 32646 28376
rect 33597 28373 33609 28376
rect 33643 28373 33655 28407
rect 33597 28367 33655 28373
rect 33962 28364 33968 28416
rect 34020 28404 34026 28416
rect 34974 28404 34980 28416
rect 34020 28376 34980 28404
rect 34020 28364 34026 28376
rect 34974 28364 34980 28376
rect 35032 28364 35038 28416
rect 35268 28404 35296 28444
rect 35345 28441 35357 28475
rect 35391 28441 35403 28475
rect 35345 28435 35403 28441
rect 35618 28404 35624 28416
rect 35268 28376 35624 28404
rect 35618 28364 35624 28376
rect 35676 28404 35682 28416
rect 35912 28404 35940 28503
rect 37550 28500 37556 28512
rect 37608 28540 37614 28552
rect 37826 28540 37832 28552
rect 37608 28512 37832 28540
rect 37608 28500 37614 28512
rect 37826 28500 37832 28512
rect 37884 28500 37890 28552
rect 36081 28475 36139 28481
rect 36081 28441 36093 28475
rect 36127 28472 36139 28475
rect 36814 28472 36820 28484
rect 36127 28444 36820 28472
rect 36127 28441 36139 28444
rect 36081 28435 36139 28441
rect 36814 28432 36820 28444
rect 36872 28432 36878 28484
rect 35676 28376 35940 28404
rect 35676 28364 35682 28376
rect 1104 28314 41400 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 41400 28314
rect 1104 28240 41400 28262
rect 1854 28160 1860 28212
rect 1912 28160 1918 28212
rect 5442 28160 5448 28212
rect 5500 28200 5506 28212
rect 6178 28200 6184 28212
rect 5500 28172 6184 28200
rect 5500 28160 5506 28172
rect 6178 28160 6184 28172
rect 6236 28160 6242 28212
rect 9306 28160 9312 28212
rect 9364 28200 9370 28212
rect 10965 28203 11023 28209
rect 10965 28200 10977 28203
rect 9364 28172 10977 28200
rect 9364 28160 9370 28172
rect 1673 28135 1731 28141
rect 1673 28101 1685 28135
rect 1719 28132 1731 28135
rect 1872 28132 1900 28160
rect 3050 28132 3056 28144
rect 1719 28104 1900 28132
rect 2898 28104 3056 28132
rect 1719 28101 1731 28104
rect 1673 28095 1731 28101
rect 3050 28092 3056 28104
rect 3108 28092 3114 28144
rect 5718 28092 5724 28144
rect 5776 28092 5782 28144
rect 5905 28135 5963 28141
rect 5905 28101 5917 28135
rect 5951 28132 5963 28135
rect 5951 28104 8340 28132
rect 5951 28101 5963 28104
rect 5905 28095 5963 28101
rect 1394 28024 1400 28076
rect 1452 28024 1458 28076
rect 4982 28024 4988 28076
rect 5040 28064 5046 28076
rect 5350 28064 5356 28076
rect 5040 28036 5356 28064
rect 5040 28024 5046 28036
rect 5350 28024 5356 28036
rect 5408 28064 5414 28076
rect 5920 28064 5948 28095
rect 5408 28036 5948 28064
rect 5408 28024 5414 28036
rect 3326 27956 3332 28008
rect 3384 27996 3390 28008
rect 3421 27999 3479 28005
rect 3421 27996 3433 27999
rect 3384 27968 3433 27996
rect 3384 27956 3390 27968
rect 3421 27965 3433 27968
rect 3467 27965 3479 27999
rect 3421 27959 3479 27965
rect 5997 27999 6055 28005
rect 5997 27965 6009 27999
rect 6043 27996 6055 27999
rect 6086 27996 6092 28008
rect 6043 27968 6092 27996
rect 6043 27965 6055 27968
rect 5997 27959 6055 27965
rect 6086 27956 6092 27968
rect 6144 27956 6150 28008
rect 8312 27872 8340 28104
rect 10796 27996 10824 28172
rect 10965 28169 10977 28172
rect 11011 28169 11023 28203
rect 10965 28163 11023 28169
rect 11238 28160 11244 28212
rect 11296 28160 11302 28212
rect 12526 28160 12532 28212
rect 12584 28200 12590 28212
rect 12621 28203 12679 28209
rect 12621 28200 12633 28203
rect 12584 28172 12633 28200
rect 12584 28160 12590 28172
rect 12621 28169 12633 28172
rect 12667 28169 12679 28203
rect 12621 28163 12679 28169
rect 12710 28160 12716 28212
rect 12768 28200 12774 28212
rect 13446 28200 13452 28212
rect 12768 28172 13452 28200
rect 12768 28160 12774 28172
rect 13446 28160 13452 28172
rect 13504 28160 13510 28212
rect 14182 28160 14188 28212
rect 14240 28160 14246 28212
rect 20990 28160 20996 28212
rect 21048 28200 21054 28212
rect 21174 28200 21180 28212
rect 21048 28172 21180 28200
rect 21048 28160 21054 28172
rect 21174 28160 21180 28172
rect 21232 28160 21238 28212
rect 22278 28160 22284 28212
rect 22336 28200 22342 28212
rect 22336 28172 23336 28200
rect 22336 28160 22342 28172
rect 10873 28135 10931 28141
rect 10873 28101 10885 28135
rect 10919 28132 10931 28135
rect 11256 28132 11284 28160
rect 10919 28104 11284 28132
rect 10919 28101 10931 28104
rect 10873 28095 10931 28101
rect 11882 28092 11888 28144
rect 11940 28132 11946 28144
rect 14200 28132 14228 28160
rect 11940 28104 14228 28132
rect 11940 28092 11946 28104
rect 12158 28024 12164 28076
rect 12216 28024 12222 28076
rect 12250 28024 12256 28076
rect 12308 28064 12314 28076
rect 12452 28073 12480 28104
rect 14458 28092 14464 28144
rect 14516 28132 14522 28144
rect 15562 28132 15568 28144
rect 14516 28104 15568 28132
rect 14516 28092 14522 28104
rect 15562 28092 15568 28104
rect 15620 28092 15626 28144
rect 19058 28092 19064 28144
rect 19116 28132 19122 28144
rect 19242 28132 19248 28144
rect 19116 28104 19248 28132
rect 19116 28092 19122 28104
rect 19242 28092 19248 28104
rect 19300 28092 19306 28144
rect 21266 28132 21272 28144
rect 21008 28104 21272 28132
rect 12345 28067 12403 28073
rect 12345 28064 12357 28067
rect 12308 28036 12357 28064
rect 12308 28024 12314 28036
rect 12345 28033 12357 28036
rect 12391 28033 12403 28067
rect 12345 28027 12403 28033
rect 12437 28067 12495 28073
rect 12437 28033 12449 28067
rect 12483 28033 12495 28067
rect 12437 28027 12495 28033
rect 12529 28067 12587 28073
rect 12529 28033 12541 28067
rect 12575 28033 12587 28067
rect 12529 28027 12587 28033
rect 12544 27996 12572 28027
rect 12618 28024 12624 28076
rect 12676 28064 12682 28076
rect 12713 28067 12771 28073
rect 12713 28064 12725 28067
rect 12676 28036 12725 28064
rect 12676 28024 12682 28036
rect 12713 28033 12725 28036
rect 12759 28033 12771 28067
rect 12713 28027 12771 28033
rect 14182 28024 14188 28076
rect 14240 28064 14246 28076
rect 15378 28064 15384 28076
rect 14240 28036 15384 28064
rect 14240 28024 14246 28036
rect 15378 28024 15384 28036
rect 15436 28024 15442 28076
rect 15838 28024 15844 28076
rect 15896 28064 15902 28076
rect 18046 28064 18052 28076
rect 15896 28036 18052 28064
rect 15896 28024 15902 28036
rect 18046 28024 18052 28036
rect 18104 28024 18110 28076
rect 20806 28024 20812 28076
rect 20864 28024 20870 28076
rect 21008 28073 21036 28104
rect 21266 28092 21272 28104
rect 21324 28092 21330 28144
rect 22830 28092 22836 28144
rect 22888 28132 22894 28144
rect 23014 28132 23020 28144
rect 22888 28104 23020 28132
rect 22888 28092 22894 28104
rect 23014 28092 23020 28104
rect 23072 28092 23078 28144
rect 23308 28132 23336 28172
rect 23382 28160 23388 28212
rect 23440 28200 23446 28212
rect 23842 28200 23848 28212
rect 23440 28172 23848 28200
rect 23440 28160 23446 28172
rect 23842 28160 23848 28172
rect 23900 28200 23906 28212
rect 24946 28200 24952 28212
rect 23900 28172 24952 28200
rect 23900 28160 23906 28172
rect 24946 28160 24952 28172
rect 25004 28160 25010 28212
rect 25866 28160 25872 28212
rect 25924 28200 25930 28212
rect 26418 28200 26424 28212
rect 25924 28172 26424 28200
rect 25924 28160 25930 28172
rect 26418 28160 26424 28172
rect 26476 28160 26482 28212
rect 27246 28160 27252 28212
rect 27304 28160 27310 28212
rect 27448 28172 28307 28200
rect 23750 28132 23756 28144
rect 23308 28104 23756 28132
rect 23750 28092 23756 28104
rect 23808 28092 23814 28144
rect 25314 28092 25320 28144
rect 25372 28132 25378 28144
rect 27264 28132 27292 28160
rect 25372 28104 27292 28132
rect 25372 28092 25378 28104
rect 20993 28067 21051 28073
rect 20993 28033 21005 28067
rect 21039 28033 21051 28067
rect 20993 28027 21051 28033
rect 21085 28067 21143 28073
rect 21085 28033 21097 28067
rect 21131 28064 21143 28067
rect 21818 28064 21824 28076
rect 21131 28036 21824 28064
rect 21131 28033 21143 28036
rect 21085 28027 21143 28033
rect 13538 27996 13544 28008
rect 10796 27968 13544 27996
rect 13538 27956 13544 27968
rect 13596 27956 13602 28008
rect 17678 27956 17684 28008
rect 17736 27996 17742 28008
rect 19334 27996 19340 28008
rect 17736 27968 19340 27996
rect 17736 27956 17742 27968
rect 19334 27956 19340 27968
rect 19392 27996 19398 28008
rect 20346 27996 20352 28008
rect 19392 27968 20352 27996
rect 19392 27956 19398 27968
rect 20346 27956 20352 27968
rect 20404 27996 20410 28008
rect 21100 27996 21128 28027
rect 21818 28024 21824 28036
rect 21876 28024 21882 28076
rect 22554 28024 22560 28076
rect 22612 28064 22618 28076
rect 24026 28064 24032 28076
rect 22612 28036 24032 28064
rect 22612 28024 22618 28036
rect 24026 28024 24032 28036
rect 24084 28024 24090 28076
rect 26252 28073 26280 28104
rect 26237 28067 26295 28073
rect 26237 28033 26249 28067
rect 26283 28033 26295 28067
rect 26237 28027 26295 28033
rect 26418 28024 26424 28076
rect 26476 28024 26482 28076
rect 26973 28067 27031 28073
rect 26973 28064 26985 28067
rect 26712 28036 26985 28064
rect 26712 28008 26740 28036
rect 26973 28033 26985 28036
rect 27019 28033 27031 28067
rect 26973 28027 27031 28033
rect 27157 28067 27215 28073
rect 27157 28033 27169 28067
rect 27203 28064 27215 28067
rect 27246 28064 27252 28076
rect 27203 28036 27252 28064
rect 27203 28033 27215 28036
rect 27157 28027 27215 28033
rect 20404 27968 21128 27996
rect 20404 27956 20410 27968
rect 22738 27956 22744 28008
rect 22796 27996 22802 28008
rect 23474 27996 23480 28008
rect 22796 27968 23480 27996
rect 22796 27956 22802 27968
rect 23474 27956 23480 27968
rect 23532 27956 23538 28008
rect 23658 27956 23664 28008
rect 23716 27996 23722 28008
rect 24854 27996 24860 28008
rect 23716 27968 24860 27996
rect 23716 27956 23722 27968
rect 24854 27956 24860 27968
rect 24912 27956 24918 28008
rect 26694 27956 26700 28008
rect 26752 27956 26758 28008
rect 26988 27996 27016 28027
rect 27246 28024 27252 28036
rect 27304 28064 27310 28076
rect 27448 28064 27476 28172
rect 27522 28092 27528 28144
rect 27580 28132 27586 28144
rect 28077 28135 28135 28141
rect 28077 28132 28089 28135
rect 27580 28104 28089 28132
rect 27580 28092 27586 28104
rect 28077 28101 28089 28104
rect 28123 28101 28135 28135
rect 28077 28095 28135 28101
rect 27304 28036 27476 28064
rect 27801 28067 27859 28073
rect 27304 28024 27310 28036
rect 27801 28033 27813 28067
rect 27847 28064 27859 28067
rect 27847 28036 27946 28064
rect 27847 28033 27859 28036
rect 27801 28027 27859 28033
rect 27614 27996 27620 28008
rect 26988 27968 27620 27996
rect 27614 27956 27620 27968
rect 27672 27956 27678 28008
rect 8662 27888 8668 27940
rect 8720 27928 8726 27940
rect 13630 27928 13636 27940
rect 8720 27900 13636 27928
rect 8720 27888 8726 27900
rect 13630 27888 13636 27900
rect 13688 27888 13694 27940
rect 14274 27888 14280 27940
rect 14332 27928 14338 27940
rect 15010 27928 15016 27940
rect 14332 27900 15016 27928
rect 14332 27888 14338 27900
rect 15010 27888 15016 27900
rect 15068 27928 15074 27940
rect 17218 27928 17224 27940
rect 15068 27900 17224 27928
rect 15068 27888 15074 27900
rect 17218 27888 17224 27900
rect 17276 27928 17282 27940
rect 20901 27931 20959 27937
rect 17276 27900 20760 27928
rect 17276 27888 17282 27900
rect 4706 27820 4712 27872
rect 4764 27860 4770 27872
rect 5445 27863 5503 27869
rect 5445 27860 5457 27863
rect 4764 27832 5457 27860
rect 4764 27820 4770 27832
rect 5445 27829 5457 27832
rect 5491 27829 5503 27863
rect 5445 27823 5503 27829
rect 8294 27820 8300 27872
rect 8352 27820 8358 27872
rect 10042 27820 10048 27872
rect 10100 27860 10106 27872
rect 10318 27860 10324 27872
rect 10100 27832 10324 27860
rect 10100 27820 10106 27832
rect 10318 27820 10324 27832
rect 10376 27820 10382 27872
rect 11977 27863 12035 27869
rect 11977 27829 11989 27863
rect 12023 27860 12035 27863
rect 12158 27860 12164 27872
rect 12023 27832 12164 27860
rect 12023 27829 12035 27832
rect 11977 27823 12035 27829
rect 12158 27820 12164 27832
rect 12216 27820 12222 27872
rect 19518 27820 19524 27872
rect 19576 27860 19582 27872
rect 20625 27863 20683 27869
rect 20625 27860 20637 27863
rect 19576 27832 20637 27860
rect 19576 27820 19582 27832
rect 20625 27829 20637 27832
rect 20671 27829 20683 27863
rect 20732 27860 20760 27900
rect 20901 27897 20913 27931
rect 20947 27928 20959 27931
rect 25038 27928 25044 27940
rect 20947 27900 25044 27928
rect 20947 27897 20959 27900
rect 20901 27891 20959 27897
rect 25038 27888 25044 27900
rect 25096 27888 25102 27940
rect 25130 27888 25136 27940
rect 25188 27928 25194 27940
rect 27522 27928 27528 27940
rect 25188 27900 27528 27928
rect 25188 27888 25194 27900
rect 27522 27888 27528 27900
rect 27580 27888 27586 27940
rect 27918 27928 27946 28036
rect 27982 28024 27988 28076
rect 28040 28024 28046 28076
rect 28166 28024 28172 28076
rect 28224 28024 28230 28076
rect 28279 28064 28307 28172
rect 28350 28160 28356 28212
rect 28408 28160 28414 28212
rect 28534 28160 28540 28212
rect 28592 28160 28598 28212
rect 28828 28172 28994 28200
rect 28445 28135 28503 28141
rect 28445 28101 28457 28135
rect 28491 28132 28503 28135
rect 28552 28132 28580 28160
rect 28828 28132 28856 28172
rect 28491 28104 28580 28132
rect 28644 28104 28856 28132
rect 28966 28132 28994 28172
rect 29086 28160 29092 28212
rect 29144 28160 29150 28212
rect 32306 28160 32312 28212
rect 32364 28200 32370 28212
rect 32582 28200 32588 28212
rect 32364 28172 32588 28200
rect 32364 28160 32370 28172
rect 32582 28160 32588 28172
rect 32640 28160 32646 28212
rect 34330 28200 34336 28212
rect 33796 28172 34336 28200
rect 29104 28132 29132 28160
rect 28966 28104 29132 28132
rect 28491 28101 28503 28104
rect 28445 28095 28503 28101
rect 28644 28064 28672 28104
rect 31754 28092 31760 28144
rect 31812 28132 31818 28144
rect 32766 28132 32772 28144
rect 31812 28104 32772 28132
rect 31812 28092 31818 28104
rect 32766 28092 32772 28104
rect 32824 28092 32830 28144
rect 33796 28141 33824 28172
rect 34330 28160 34336 28172
rect 34388 28160 34394 28212
rect 34698 28160 34704 28212
rect 34756 28160 34762 28212
rect 37458 28160 37464 28212
rect 37516 28200 37522 28212
rect 37645 28203 37703 28209
rect 37645 28200 37657 28203
rect 37516 28172 37657 28200
rect 37516 28160 37522 28172
rect 37645 28169 37657 28172
rect 37691 28169 37703 28203
rect 37645 28163 37703 28169
rect 38289 28203 38347 28209
rect 38289 28169 38301 28203
rect 38335 28200 38347 28203
rect 38378 28200 38384 28212
rect 38335 28172 38384 28200
rect 38335 28169 38347 28172
rect 38289 28163 38347 28169
rect 38378 28160 38384 28172
rect 38436 28160 38442 28212
rect 33781 28135 33839 28141
rect 33781 28101 33793 28135
rect 33827 28101 33839 28135
rect 34716 28132 34744 28160
rect 33781 28095 33839 28101
rect 34072 28104 34744 28132
rect 28279 28036 28672 28064
rect 28813 28067 28871 28073
rect 28813 28033 28825 28067
rect 28859 28033 28871 28067
rect 28813 28027 28871 28033
rect 28074 27956 28080 28008
rect 28132 27996 28138 28008
rect 28534 27996 28540 28008
rect 28132 27968 28540 27996
rect 28132 27956 28138 27968
rect 28534 27956 28540 27968
rect 28592 27956 28598 28008
rect 28828 27996 28856 28027
rect 28902 28024 28908 28076
rect 28960 28024 28966 28076
rect 29270 28024 29276 28076
rect 29328 28024 29334 28076
rect 31570 28024 31576 28076
rect 31628 28064 31634 28076
rect 34072 28073 34100 28104
rect 35710 28092 35716 28144
rect 35768 28132 35774 28144
rect 35768 28104 38654 28132
rect 35768 28092 35774 28104
rect 34057 28067 34115 28073
rect 31628 28036 32996 28064
rect 31628 28024 31634 28036
rect 29288 27996 29316 28024
rect 28828 27968 29316 27996
rect 27918 27900 28304 27928
rect 21266 27860 21272 27872
rect 20732 27832 21272 27860
rect 20625 27823 20683 27829
rect 21266 27820 21272 27832
rect 21324 27820 21330 27872
rect 22278 27820 22284 27872
rect 22336 27860 22342 27872
rect 25958 27860 25964 27872
rect 22336 27832 25964 27860
rect 22336 27820 22342 27832
rect 25958 27820 25964 27832
rect 26016 27820 26022 27872
rect 26142 27820 26148 27872
rect 26200 27860 26206 27872
rect 26237 27863 26295 27869
rect 26237 27860 26249 27863
rect 26200 27832 26249 27860
rect 26200 27820 26206 27832
rect 26237 27829 26249 27832
rect 26283 27829 26295 27863
rect 26237 27823 26295 27829
rect 26878 27820 26884 27872
rect 26936 27860 26942 27872
rect 27341 27863 27399 27869
rect 27341 27860 27353 27863
rect 26936 27832 27353 27860
rect 26936 27820 26942 27832
rect 27341 27829 27353 27832
rect 27387 27829 27399 27863
rect 27341 27823 27399 27829
rect 27706 27820 27712 27872
rect 27764 27860 27770 27872
rect 27918 27860 27946 27900
rect 28276 27872 28304 27900
rect 28350 27888 28356 27940
rect 28408 27928 28414 27940
rect 28408 27900 28856 27928
rect 28408 27888 28414 27900
rect 27764 27832 27946 27860
rect 27764 27820 27770 27832
rect 28258 27820 28264 27872
rect 28316 27820 28322 27872
rect 28718 27820 28724 27872
rect 28776 27820 28782 27872
rect 28828 27860 28856 27900
rect 29086 27888 29092 27940
rect 29144 27888 29150 27940
rect 32968 27928 32996 28036
rect 34057 28033 34069 28067
rect 34103 28033 34115 28067
rect 34057 28027 34115 28033
rect 34514 28024 34520 28076
rect 34572 28064 34578 28076
rect 34885 28067 34943 28073
rect 34885 28064 34897 28067
rect 34572 28036 34897 28064
rect 34572 28024 34578 28036
rect 34885 28033 34897 28036
rect 34931 28033 34943 28067
rect 34885 28027 34943 28033
rect 35894 28024 35900 28076
rect 35952 28024 35958 28076
rect 35989 28067 36047 28073
rect 35989 28033 36001 28067
rect 36035 28064 36047 28067
rect 36906 28064 36912 28076
rect 36035 28036 36912 28064
rect 36035 28033 36047 28036
rect 35989 28027 36047 28033
rect 36906 28024 36912 28036
rect 36964 28064 36970 28076
rect 37921 28067 37979 28073
rect 37921 28064 37933 28067
rect 36964 28036 37933 28064
rect 36964 28024 36970 28036
rect 37921 28033 37933 28036
rect 37967 28033 37979 28067
rect 37921 28027 37979 28033
rect 38010 28024 38016 28076
rect 38068 28024 38074 28076
rect 38286 28024 38292 28076
rect 38344 28024 38350 28076
rect 38473 28067 38531 28073
rect 38473 28033 38485 28067
rect 38519 28033 38531 28067
rect 38626 28064 38654 28104
rect 40034 28092 40040 28144
rect 40092 28092 40098 28144
rect 40678 28092 40684 28144
rect 40736 28132 40742 28144
rect 41049 28135 41107 28141
rect 41049 28132 41061 28135
rect 40736 28104 41061 28132
rect 40736 28092 40742 28104
rect 41049 28101 41061 28104
rect 41095 28101 41107 28135
rect 41049 28095 41107 28101
rect 39022 28064 39028 28076
rect 39080 28073 39086 28076
rect 38626 28036 39028 28064
rect 38473 28027 38531 28033
rect 33962 27956 33968 28008
rect 34020 27956 34026 28008
rect 35526 27956 35532 28008
rect 35584 27956 35590 28008
rect 35912 27996 35940 28024
rect 36081 27999 36139 28005
rect 36081 27996 36093 27999
rect 35912 27968 36093 27996
rect 36081 27965 36093 27968
rect 36127 27965 36139 27999
rect 36081 27959 36139 27965
rect 36357 27999 36415 28005
rect 36357 27965 36369 27999
rect 36403 27996 36415 27999
rect 36446 27996 36452 28008
rect 36403 27968 36452 27996
rect 36403 27965 36415 27968
rect 36357 27959 36415 27965
rect 36446 27956 36452 27968
rect 36504 27956 36510 28008
rect 36538 27956 36544 28008
rect 36596 27956 36602 28008
rect 36725 27999 36783 28005
rect 36725 27965 36737 27999
rect 36771 27965 36783 27999
rect 36725 27959 36783 27965
rect 34241 27931 34299 27937
rect 34241 27928 34253 27931
rect 32968 27900 34253 27928
rect 34241 27897 34253 27900
rect 34287 27897 34299 27931
rect 34241 27891 34299 27897
rect 31018 27860 31024 27872
rect 28828 27832 31024 27860
rect 31018 27820 31024 27832
rect 31076 27820 31082 27872
rect 31294 27820 31300 27872
rect 31352 27860 31358 27872
rect 31846 27860 31852 27872
rect 31352 27832 31852 27860
rect 31352 27820 31358 27832
rect 31846 27820 31852 27832
rect 31904 27860 31910 27872
rect 32582 27860 32588 27872
rect 31904 27832 32588 27860
rect 31904 27820 31910 27832
rect 32582 27820 32588 27832
rect 32640 27820 32646 27872
rect 33778 27820 33784 27872
rect 33836 27820 33842 27872
rect 34698 27820 34704 27872
rect 34756 27860 34762 27872
rect 35544 27860 35572 27956
rect 35986 27888 35992 27940
rect 36044 27928 36050 27940
rect 36740 27928 36768 27959
rect 37366 27956 37372 28008
rect 37424 27996 37430 28008
rect 37461 27999 37519 28005
rect 37461 27996 37473 27999
rect 37424 27968 37473 27996
rect 37424 27956 37430 27968
rect 37461 27965 37473 27968
rect 37507 27965 37519 27999
rect 37461 27959 37519 27965
rect 37553 27999 37611 28005
rect 37553 27965 37565 27999
rect 37599 27965 37611 27999
rect 37553 27959 37611 27965
rect 37829 27999 37887 28005
rect 37829 27965 37841 27999
rect 37875 27965 37887 27999
rect 38028 27996 38056 28024
rect 38488 27996 38516 28027
rect 39022 28024 39028 28036
rect 39080 28027 39090 28073
rect 39080 28024 39086 28027
rect 38028 27968 38516 27996
rect 37829 27959 37887 27965
rect 37568 27928 37596 27959
rect 36044 27900 36768 27928
rect 37200 27900 37596 27928
rect 36044 27888 36050 27900
rect 34756 27832 35572 27860
rect 34756 27820 34762 27832
rect 36354 27820 36360 27872
rect 36412 27860 36418 27872
rect 37200 27860 37228 27900
rect 36412 27832 37228 27860
rect 36412 27820 36418 27832
rect 37274 27820 37280 27872
rect 37332 27820 37338 27872
rect 37550 27820 37556 27872
rect 37608 27860 37614 27872
rect 37844 27860 37872 27959
rect 39298 27956 39304 28008
rect 39356 27956 39362 28008
rect 37608 27832 37872 27860
rect 37608 27820 37614 27832
rect 1104 27770 41400 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 41400 27770
rect 1104 27696 41400 27718
rect 8205 27659 8263 27665
rect 8205 27656 8217 27659
rect 6012 27628 8217 27656
rect 6012 27600 6040 27628
rect 8205 27625 8217 27628
rect 8251 27625 8263 27659
rect 8205 27619 8263 27625
rect 8294 27616 8300 27668
rect 8352 27656 8358 27668
rect 9493 27659 9551 27665
rect 9493 27656 9505 27659
rect 8352 27628 9505 27656
rect 8352 27616 8358 27628
rect 9493 27625 9505 27628
rect 9539 27625 9551 27659
rect 9493 27619 9551 27625
rect 10410 27616 10416 27668
rect 10468 27656 10474 27668
rect 10505 27659 10563 27665
rect 10505 27656 10517 27659
rect 10468 27628 10517 27656
rect 10468 27616 10474 27628
rect 10505 27625 10517 27628
rect 10551 27656 10563 27659
rect 10962 27656 10968 27668
rect 10551 27628 10968 27656
rect 10551 27625 10563 27628
rect 10505 27619 10563 27625
rect 10962 27616 10968 27628
rect 11020 27616 11026 27668
rect 12342 27616 12348 27668
rect 12400 27656 12406 27668
rect 12618 27656 12624 27668
rect 12400 27628 12624 27656
rect 12400 27616 12406 27628
rect 12618 27616 12624 27628
rect 12676 27616 12682 27668
rect 13541 27659 13599 27665
rect 13541 27625 13553 27659
rect 13587 27656 13599 27659
rect 13814 27656 13820 27668
rect 13587 27628 13820 27656
rect 13587 27625 13599 27628
rect 13541 27619 13599 27625
rect 13814 27616 13820 27628
rect 13872 27616 13878 27668
rect 15838 27656 15844 27668
rect 13924 27628 15844 27656
rect 4614 27548 4620 27600
rect 4672 27588 4678 27600
rect 4893 27591 4951 27597
rect 4893 27588 4905 27591
rect 4672 27560 4905 27588
rect 4672 27548 4678 27560
rect 4893 27557 4905 27560
rect 4939 27588 4951 27591
rect 4939 27560 5304 27588
rect 4939 27557 4951 27560
rect 4893 27551 4951 27557
rect 4890 27344 4896 27396
rect 4948 27384 4954 27396
rect 5074 27384 5080 27396
rect 4948 27356 5080 27384
rect 4948 27344 4954 27356
rect 5074 27344 5080 27356
rect 5132 27384 5138 27396
rect 5169 27387 5227 27393
rect 5169 27384 5181 27387
rect 5132 27356 5181 27384
rect 5132 27344 5138 27356
rect 5169 27353 5181 27356
rect 5215 27353 5227 27387
rect 5169 27347 5227 27353
rect 5276 27316 5304 27560
rect 5994 27548 6000 27600
rect 6052 27548 6058 27600
rect 8846 27588 8852 27600
rect 6656 27560 8852 27588
rect 6656 27529 6684 27560
rect 8846 27548 8852 27560
rect 8904 27548 8910 27600
rect 13924 27588 13952 27628
rect 15838 27616 15844 27628
rect 15896 27616 15902 27668
rect 15930 27616 15936 27668
rect 15988 27656 15994 27668
rect 16577 27659 16635 27665
rect 16577 27656 16589 27659
rect 15988 27628 16589 27656
rect 15988 27616 15994 27628
rect 16577 27625 16589 27628
rect 16623 27625 16635 27659
rect 19518 27656 19524 27668
rect 16577 27619 16635 27625
rect 19352 27628 19524 27656
rect 9789 27560 13952 27588
rect 6641 27523 6699 27529
rect 6641 27489 6653 27523
rect 6687 27489 6699 27523
rect 6641 27483 6699 27489
rect 7760 27492 9536 27520
rect 7760 27464 7788 27492
rect 5626 27412 5632 27464
rect 5684 27452 5690 27464
rect 5810 27452 5816 27464
rect 5684 27424 5816 27452
rect 5684 27412 5690 27424
rect 5810 27412 5816 27424
rect 5868 27452 5874 27464
rect 5905 27455 5963 27461
rect 5905 27452 5917 27455
rect 5868 27424 5917 27452
rect 5868 27412 5874 27424
rect 5905 27421 5917 27424
rect 5951 27421 5963 27455
rect 5905 27415 5963 27421
rect 5994 27412 6000 27464
rect 6052 27461 6058 27464
rect 6052 27455 6081 27461
rect 6069 27421 6081 27455
rect 6052 27415 6081 27421
rect 6181 27455 6239 27461
rect 6181 27421 6193 27455
rect 6227 27452 6239 27455
rect 6227 27424 6408 27452
rect 6227 27421 6239 27424
rect 6181 27415 6239 27421
rect 6052 27412 6058 27415
rect 6380 27396 6408 27424
rect 7742 27412 7748 27464
rect 7800 27412 7806 27464
rect 7837 27455 7895 27461
rect 7837 27421 7849 27455
rect 7883 27421 7895 27455
rect 7837 27415 7895 27421
rect 8021 27455 8079 27461
rect 8021 27421 8033 27455
rect 8067 27421 8079 27455
rect 8021 27415 8079 27421
rect 8113 27455 8171 27461
rect 8113 27421 8125 27455
rect 8159 27452 8171 27455
rect 8294 27452 8300 27464
rect 8159 27424 8300 27452
rect 8159 27421 8171 27424
rect 8113 27415 8171 27421
rect 5350 27344 5356 27396
rect 5408 27344 5414 27396
rect 5445 27387 5503 27393
rect 5445 27353 5457 27387
rect 5491 27384 5503 27387
rect 6362 27384 6368 27396
rect 5491 27356 6368 27384
rect 5491 27353 5503 27356
rect 5445 27347 5503 27353
rect 6362 27344 6368 27356
rect 6420 27344 6426 27396
rect 7006 27344 7012 27396
rect 7064 27384 7070 27396
rect 7561 27387 7619 27393
rect 7561 27384 7573 27387
rect 7064 27356 7573 27384
rect 7064 27344 7070 27356
rect 7561 27353 7573 27356
rect 7607 27353 7619 27387
rect 7561 27347 7619 27353
rect 6270 27316 6276 27328
rect 5276 27288 6276 27316
rect 6270 27276 6276 27288
rect 6328 27276 6334 27328
rect 7852 27316 7880 27415
rect 7926 27344 7932 27396
rect 7984 27384 7990 27396
rect 8036 27384 8064 27415
rect 8294 27412 8300 27424
rect 8352 27412 8358 27464
rect 8404 27461 8432 27492
rect 8588 27464 8616 27492
rect 8389 27455 8447 27461
rect 8389 27421 8401 27455
rect 8435 27421 8447 27455
rect 8389 27415 8447 27421
rect 8478 27412 8484 27464
rect 8536 27412 8542 27464
rect 8570 27412 8576 27464
rect 8628 27412 8634 27464
rect 8665 27455 8723 27461
rect 8665 27421 8677 27455
rect 8711 27421 8723 27455
rect 8665 27415 8723 27421
rect 8680 27384 8708 27415
rect 8754 27412 8760 27464
rect 8812 27412 8818 27464
rect 9508 27448 9536 27492
rect 9789 27464 9817 27560
rect 15102 27548 15108 27600
rect 15160 27588 15166 27600
rect 15749 27591 15807 27597
rect 15749 27588 15761 27591
rect 15160 27560 15761 27588
rect 15160 27548 15166 27560
rect 15749 27557 15761 27560
rect 15795 27557 15807 27591
rect 15749 27551 15807 27557
rect 19245 27591 19303 27597
rect 19245 27557 19257 27591
rect 19291 27557 19303 27591
rect 19245 27551 19303 27557
rect 9968 27492 10180 27520
rect 9677 27455 9735 27461
rect 9508 27442 9628 27448
rect 9677 27442 9689 27455
rect 9508 27421 9689 27442
rect 9723 27421 9735 27455
rect 9508 27420 9735 27421
rect 9600 27415 9735 27420
rect 9600 27414 9720 27415
rect 9766 27412 9772 27464
rect 9824 27412 9830 27464
rect 9968 27461 9996 27492
rect 9953 27455 10011 27461
rect 9953 27452 9965 27455
rect 9876 27424 9965 27452
rect 7984 27356 8985 27384
rect 7984 27344 7990 27356
rect 8386 27316 8392 27328
rect 7852 27288 8392 27316
rect 8386 27276 8392 27288
rect 8444 27276 8450 27328
rect 8957 27316 8985 27356
rect 9876 27316 9904 27424
rect 9953 27421 9965 27424
rect 9999 27421 10011 27455
rect 9953 27415 10011 27421
rect 10045 27455 10103 27461
rect 10045 27421 10057 27455
rect 10091 27421 10103 27455
rect 10152 27452 10180 27492
rect 10318 27480 10324 27532
rect 10376 27520 10382 27532
rect 10505 27523 10563 27529
rect 10505 27520 10517 27523
rect 10376 27492 10517 27520
rect 10376 27480 10382 27492
rect 10505 27489 10517 27492
rect 10551 27489 10563 27523
rect 10505 27483 10563 27489
rect 13538 27480 13544 27532
rect 13596 27520 13602 27532
rect 15289 27523 15347 27529
rect 15289 27520 15301 27523
rect 13596 27492 15301 27520
rect 13596 27480 13602 27492
rect 15289 27489 15301 27492
rect 15335 27489 15347 27523
rect 15289 27483 15347 27489
rect 15841 27523 15899 27529
rect 15841 27489 15853 27523
rect 15887 27520 15899 27523
rect 19260 27520 19288 27551
rect 15887 27492 16620 27520
rect 15887 27489 15899 27492
rect 15841 27483 15899 27489
rect 16592 27464 16620 27492
rect 16776 27492 19288 27520
rect 16776 27464 16804 27492
rect 10413 27455 10471 27461
rect 10413 27452 10425 27455
rect 10152 27424 10425 27452
rect 10045 27415 10103 27421
rect 10413 27421 10425 27424
rect 10459 27452 10471 27455
rect 12434 27452 12440 27464
rect 10459 27424 12440 27452
rect 10459 27421 10471 27424
rect 10413 27415 10471 27421
rect 10061 27328 10089 27415
rect 12434 27412 12440 27424
rect 12492 27412 12498 27464
rect 13449 27455 13507 27461
rect 13449 27421 13461 27455
rect 13495 27421 13507 27455
rect 13449 27415 13507 27421
rect 13633 27455 13691 27461
rect 13633 27421 13645 27455
rect 13679 27452 13691 27455
rect 15657 27455 15715 27461
rect 13679 27424 13952 27452
rect 13679 27421 13691 27424
rect 13633 27415 13691 27421
rect 10137 27387 10195 27393
rect 10137 27353 10149 27387
rect 10183 27384 10195 27387
rect 10318 27384 10324 27396
rect 10183 27356 10324 27384
rect 10183 27353 10195 27356
rect 10137 27347 10195 27353
rect 10318 27344 10324 27356
rect 10376 27384 10382 27396
rect 13464 27384 13492 27415
rect 13924 27396 13952 27424
rect 15657 27421 15669 27455
rect 15703 27452 15715 27455
rect 15746 27452 15752 27464
rect 15703 27424 15752 27452
rect 15703 27421 15715 27424
rect 15657 27415 15715 27421
rect 15746 27412 15752 27424
rect 15804 27412 15810 27464
rect 16206 27412 16212 27464
rect 16264 27412 16270 27464
rect 16485 27455 16543 27461
rect 16485 27421 16497 27455
rect 16531 27421 16543 27455
rect 16485 27415 16543 27421
rect 13722 27384 13728 27396
rect 10376 27356 12848 27384
rect 13464 27356 13728 27384
rect 10376 27344 10382 27356
rect 12820 27328 12848 27356
rect 13722 27344 13728 27356
rect 13780 27344 13786 27396
rect 13906 27344 13912 27396
rect 13964 27344 13970 27396
rect 15105 27387 15163 27393
rect 15105 27353 15117 27387
rect 15151 27384 15163 27387
rect 15562 27384 15568 27396
rect 15151 27356 15568 27384
rect 15151 27353 15163 27356
rect 15105 27347 15163 27353
rect 15562 27344 15568 27356
rect 15620 27384 15626 27396
rect 15930 27384 15936 27396
rect 15620 27356 15936 27384
rect 15620 27344 15626 27356
rect 15930 27344 15936 27356
rect 15988 27344 15994 27396
rect 16500 27384 16528 27415
rect 16574 27412 16580 27464
rect 16632 27412 16638 27464
rect 16758 27412 16764 27464
rect 16816 27412 16822 27464
rect 17586 27412 17592 27464
rect 17644 27412 17650 27464
rect 17773 27455 17831 27461
rect 17773 27421 17785 27455
rect 17819 27452 17831 27455
rect 17954 27452 17960 27464
rect 17819 27424 17960 27452
rect 17819 27421 17831 27424
rect 17773 27415 17831 27421
rect 17954 27412 17960 27424
rect 18012 27452 18018 27464
rect 18417 27455 18475 27461
rect 18417 27452 18429 27455
rect 18012 27424 18429 27452
rect 18012 27412 18018 27424
rect 18417 27421 18429 27424
rect 18463 27421 18475 27455
rect 19352 27452 19380 27628
rect 19518 27616 19524 27628
rect 19576 27616 19582 27668
rect 25958 27656 25964 27668
rect 21560 27628 25964 27656
rect 19429 27591 19487 27597
rect 19429 27557 19441 27591
rect 19475 27588 19487 27591
rect 19610 27588 19616 27600
rect 19475 27560 19616 27588
rect 19475 27557 19487 27560
rect 19429 27551 19487 27557
rect 19610 27548 19616 27560
rect 19668 27588 19674 27600
rect 21560 27588 21588 27628
rect 25958 27616 25964 27628
rect 26016 27616 26022 27668
rect 26418 27616 26424 27668
rect 26476 27656 26482 27668
rect 26881 27659 26939 27665
rect 26881 27656 26893 27659
rect 26476 27628 26893 27656
rect 26476 27616 26482 27628
rect 26881 27625 26893 27628
rect 26927 27625 26939 27659
rect 26881 27619 26939 27625
rect 27246 27616 27252 27668
rect 27304 27616 27310 27668
rect 27338 27616 27344 27668
rect 27396 27656 27402 27668
rect 27396 27628 28994 27656
rect 27396 27616 27402 27628
rect 19668 27560 21588 27588
rect 22741 27591 22799 27597
rect 19668 27548 19674 27560
rect 22741 27557 22753 27591
rect 22787 27588 22799 27591
rect 23106 27588 23112 27600
rect 22787 27560 23112 27588
rect 22787 27557 22799 27560
rect 22741 27551 22799 27557
rect 23106 27548 23112 27560
rect 23164 27548 23170 27600
rect 23198 27548 23204 27600
rect 23256 27548 23262 27600
rect 23382 27548 23388 27600
rect 23440 27588 23446 27600
rect 24949 27591 25007 27597
rect 24949 27588 24961 27591
rect 23440 27560 24961 27588
rect 23440 27548 23446 27560
rect 24949 27557 24961 27560
rect 24995 27588 25007 27591
rect 26326 27588 26332 27600
rect 24995 27560 26332 27588
rect 24995 27557 25007 27560
rect 24949 27551 25007 27557
rect 26326 27548 26332 27560
rect 26384 27548 26390 27600
rect 26602 27548 26608 27600
rect 26660 27548 26666 27600
rect 27798 27588 27804 27600
rect 27264 27560 27804 27588
rect 22370 27520 22376 27532
rect 22296 27492 22376 27520
rect 18417 27415 18475 27421
rect 18800 27424 19380 27452
rect 19613 27455 19671 27461
rect 18049 27387 18107 27393
rect 16500 27356 17632 27384
rect 8957 27288 9904 27316
rect 10042 27276 10048 27328
rect 10100 27276 10106 27328
rect 10229 27319 10287 27325
rect 10229 27285 10241 27319
rect 10275 27316 10287 27319
rect 10410 27316 10416 27328
rect 10275 27288 10416 27316
rect 10275 27285 10287 27288
rect 10229 27279 10287 27285
rect 10410 27276 10416 27288
rect 10468 27316 10474 27328
rect 10778 27316 10784 27328
rect 10468 27288 10784 27316
rect 10468 27276 10474 27288
rect 10778 27276 10784 27288
rect 10836 27276 10842 27328
rect 12802 27276 12808 27328
rect 12860 27316 12866 27328
rect 14366 27316 14372 27328
rect 12860 27288 14372 27316
rect 12860 27276 12866 27288
rect 14366 27276 14372 27288
rect 14424 27316 14430 27328
rect 16500 27316 16528 27356
rect 17604 27325 17632 27356
rect 18049 27353 18061 27387
rect 18095 27384 18107 27387
rect 18138 27384 18144 27396
rect 18095 27356 18144 27384
rect 18095 27353 18107 27356
rect 18049 27347 18107 27353
rect 18138 27344 18144 27356
rect 18196 27344 18202 27396
rect 18233 27387 18291 27393
rect 18233 27353 18245 27387
rect 18279 27384 18291 27387
rect 18322 27384 18328 27396
rect 18279 27356 18328 27384
rect 18279 27353 18291 27356
rect 18233 27347 18291 27353
rect 18322 27344 18328 27356
rect 18380 27384 18386 27396
rect 18800 27384 18828 27424
rect 19613 27421 19625 27455
rect 19659 27452 19671 27455
rect 19978 27452 19984 27464
rect 19659 27424 19984 27452
rect 19659 27421 19671 27424
rect 19613 27415 19671 27421
rect 19978 27412 19984 27424
rect 20036 27452 20042 27464
rect 20530 27452 20536 27464
rect 20036 27424 20536 27452
rect 20036 27412 20042 27424
rect 20530 27412 20536 27424
rect 20588 27412 20594 27464
rect 22296 27461 22324 27492
rect 22370 27480 22376 27492
rect 22428 27520 22434 27532
rect 23216 27520 23244 27548
rect 27264 27532 27292 27560
rect 27798 27548 27804 27560
rect 27856 27548 27862 27600
rect 22428 27492 23244 27520
rect 22428 27480 22434 27492
rect 23842 27480 23848 27532
rect 23900 27520 23906 27532
rect 24394 27520 24400 27532
rect 23900 27492 24400 27520
rect 23900 27480 23906 27492
rect 24394 27480 24400 27492
rect 24452 27480 24458 27532
rect 25038 27480 25044 27532
rect 25096 27520 25102 27532
rect 25590 27520 25596 27532
rect 25096 27492 25596 27520
rect 25096 27480 25102 27492
rect 25590 27480 25596 27492
rect 25648 27480 25654 27532
rect 25866 27520 25872 27532
rect 25716 27492 25872 27520
rect 22281 27455 22339 27461
rect 22281 27421 22293 27455
rect 22327 27421 22339 27455
rect 22281 27415 22339 27421
rect 22649 27455 22707 27461
rect 22649 27421 22661 27455
rect 22695 27452 22707 27455
rect 22833 27455 22891 27461
rect 22695 27424 22784 27452
rect 22695 27421 22707 27424
rect 22649 27415 22707 27421
rect 18380 27356 18828 27384
rect 18380 27344 18386 27356
rect 19242 27344 19248 27396
rect 19300 27384 19306 27396
rect 22554 27384 22560 27396
rect 19300 27356 22560 27384
rect 19300 27344 19306 27356
rect 22554 27344 22560 27356
rect 22612 27344 22618 27396
rect 22756 27328 22784 27424
rect 22833 27421 22845 27455
rect 22879 27452 22891 27455
rect 22879 27424 23060 27452
rect 22879 27421 22891 27424
rect 22833 27415 22891 27421
rect 23032 27328 23060 27424
rect 24762 27412 24768 27464
rect 24820 27412 24826 27464
rect 25133 27455 25191 27461
rect 25133 27421 25145 27455
rect 25179 27421 25191 27455
rect 25133 27415 25191 27421
rect 24581 27387 24639 27393
rect 24581 27353 24593 27387
rect 24627 27384 24639 27387
rect 25148 27384 25176 27415
rect 25222 27412 25228 27464
rect 25280 27452 25286 27464
rect 25716 27452 25744 27492
rect 25866 27480 25872 27492
rect 25924 27520 25930 27532
rect 25924 27492 27108 27520
rect 25924 27480 25930 27492
rect 25280 27424 25744 27452
rect 25777 27455 25835 27461
rect 25280 27412 25286 27424
rect 25777 27421 25789 27455
rect 25823 27452 25835 27455
rect 26050 27452 26056 27464
rect 25823 27424 26056 27452
rect 25823 27421 25835 27424
rect 25777 27415 25835 27421
rect 26050 27412 26056 27424
rect 26108 27412 26114 27464
rect 26145 27455 26203 27461
rect 26145 27421 26157 27455
rect 26191 27452 26203 27455
rect 26191 27424 26280 27452
rect 26191 27421 26203 27424
rect 26145 27415 26203 27421
rect 24627 27356 25176 27384
rect 24627 27353 24639 27356
rect 24581 27347 24639 27353
rect 14424 27288 16528 27316
rect 17589 27319 17647 27325
rect 14424 27276 14430 27288
rect 17589 27285 17601 27319
rect 17635 27285 17647 27319
rect 17589 27279 17647 27285
rect 18874 27276 18880 27328
rect 18932 27316 18938 27328
rect 19610 27316 19616 27328
rect 18932 27288 19616 27316
rect 18932 27276 18938 27288
rect 19610 27276 19616 27288
rect 19668 27276 19674 27328
rect 22094 27276 22100 27328
rect 22152 27276 22158 27328
rect 22738 27276 22744 27328
rect 22796 27276 22802 27328
rect 23014 27276 23020 27328
rect 23072 27276 23078 27328
rect 26252 27316 26280 27424
rect 26510 27412 26516 27464
rect 26568 27412 26574 27464
rect 27080 27461 27108 27492
rect 27246 27480 27252 27532
rect 27304 27480 27310 27532
rect 27341 27523 27399 27529
rect 27341 27489 27353 27523
rect 27387 27520 27399 27523
rect 28166 27520 28172 27532
rect 27387 27492 28172 27520
rect 27387 27489 27399 27492
rect 27341 27483 27399 27489
rect 28166 27480 28172 27492
rect 28224 27480 28230 27532
rect 28966 27520 28994 27628
rect 29178 27616 29184 27668
rect 29236 27656 29242 27668
rect 30098 27656 30104 27668
rect 29236 27628 30104 27656
rect 29236 27616 29242 27628
rect 30098 27616 30104 27628
rect 30156 27616 30162 27668
rect 30282 27616 30288 27668
rect 30340 27656 30346 27668
rect 30653 27659 30711 27665
rect 30653 27656 30665 27659
rect 30340 27628 30665 27656
rect 30340 27616 30346 27628
rect 30653 27625 30665 27628
rect 30699 27625 30711 27659
rect 30653 27619 30711 27625
rect 31018 27616 31024 27668
rect 31076 27656 31082 27668
rect 36078 27656 36084 27668
rect 31076 27628 36084 27656
rect 31076 27616 31082 27628
rect 36078 27616 36084 27628
rect 36136 27616 36142 27668
rect 37185 27659 37243 27665
rect 37185 27625 37197 27659
rect 37231 27625 37243 27659
rect 37185 27619 37243 27625
rect 30926 27548 30932 27600
rect 30984 27548 30990 27600
rect 31662 27548 31668 27600
rect 31720 27548 31726 27600
rect 31757 27591 31815 27597
rect 31757 27557 31769 27591
rect 31803 27588 31815 27591
rect 32398 27588 32404 27600
rect 31803 27560 32404 27588
rect 31803 27557 31815 27560
rect 31757 27551 31815 27557
rect 32398 27548 32404 27560
rect 32456 27548 32462 27600
rect 32766 27548 32772 27600
rect 32824 27588 32830 27600
rect 37200 27588 37228 27619
rect 37642 27616 37648 27668
rect 37700 27616 37706 27668
rect 39298 27616 39304 27668
rect 39356 27656 39362 27668
rect 39853 27659 39911 27665
rect 39853 27656 39865 27659
rect 39356 27628 39865 27656
rect 39356 27616 39362 27628
rect 39853 27625 39865 27628
rect 39899 27625 39911 27659
rect 39853 27619 39911 27625
rect 38289 27591 38347 27597
rect 38289 27588 38301 27591
rect 32824 27560 37228 27588
rect 37936 27560 38301 27588
rect 32824 27548 32830 27560
rect 29638 27520 29644 27532
rect 28966 27492 29644 27520
rect 29638 27480 29644 27492
rect 29696 27520 29702 27532
rect 30282 27520 30288 27532
rect 29696 27492 30288 27520
rect 29696 27480 29702 27492
rect 30282 27480 30288 27492
rect 30340 27480 30346 27532
rect 31113 27523 31171 27529
rect 31113 27489 31125 27523
rect 31159 27520 31171 27523
rect 31478 27520 31484 27532
rect 31159 27492 31484 27520
rect 31159 27489 31171 27492
rect 31113 27483 31171 27489
rect 31478 27480 31484 27492
rect 31536 27480 31542 27532
rect 31680 27520 31708 27548
rect 37366 27520 37372 27532
rect 31680 27492 31984 27520
rect 27065 27455 27123 27461
rect 27065 27421 27077 27455
rect 27111 27452 27123 27455
rect 27430 27452 27436 27464
rect 27111 27424 27436 27452
rect 27111 27421 27123 27424
rect 27065 27415 27123 27421
rect 27430 27412 27436 27424
rect 27488 27412 27494 27464
rect 28534 27412 28540 27464
rect 28592 27452 28598 27464
rect 30834 27452 30840 27464
rect 28592 27424 30840 27452
rect 28592 27412 28598 27424
rect 30834 27412 30840 27424
rect 30892 27412 30898 27464
rect 31018 27412 31024 27464
rect 31076 27412 31082 27464
rect 31202 27412 31208 27464
rect 31260 27412 31266 27464
rect 31389 27455 31447 27461
rect 31389 27421 31401 27455
rect 31435 27452 31447 27455
rect 31570 27452 31576 27464
rect 31435 27424 31576 27452
rect 31435 27421 31447 27424
rect 31389 27415 31447 27421
rect 31570 27412 31576 27424
rect 31628 27462 31634 27464
rect 31628 27461 31708 27462
rect 31628 27455 31723 27461
rect 31628 27434 31677 27455
rect 31628 27412 31634 27434
rect 31665 27421 31677 27434
rect 31711 27421 31723 27455
rect 31665 27415 31723 27421
rect 31846 27412 31852 27464
rect 31904 27412 31910 27464
rect 31956 27461 31984 27492
rect 34164 27492 37372 27520
rect 31941 27455 31999 27461
rect 31941 27421 31953 27455
rect 31987 27421 31999 27455
rect 31941 27415 31999 27421
rect 32125 27455 32183 27461
rect 32125 27421 32137 27455
rect 32171 27421 32183 27455
rect 32125 27415 32183 27421
rect 32309 27455 32367 27461
rect 32309 27421 32321 27455
rect 32355 27452 32367 27455
rect 32490 27452 32496 27464
rect 32355 27424 32496 27452
rect 32355 27421 32367 27424
rect 32309 27415 32367 27421
rect 26326 27344 26332 27396
rect 26384 27384 26390 27396
rect 31110 27384 31116 27396
rect 26384 27356 31116 27384
rect 26384 27344 26390 27356
rect 31110 27344 31116 27356
rect 31168 27344 31174 27396
rect 32140 27384 32168 27415
rect 32490 27412 32496 27424
rect 32548 27412 32554 27464
rect 33318 27412 33324 27464
rect 33376 27412 33382 27464
rect 33410 27412 33416 27464
rect 33468 27412 33474 27464
rect 33597 27455 33655 27461
rect 33597 27421 33609 27455
rect 33643 27452 33655 27455
rect 33965 27455 34023 27461
rect 33643 27424 33732 27452
rect 33643 27421 33655 27424
rect 33597 27415 33655 27421
rect 32582 27384 32588 27396
rect 32140 27356 32588 27384
rect 32582 27344 32588 27356
rect 32640 27384 32646 27396
rect 33428 27384 33456 27412
rect 32640 27356 33456 27384
rect 32640 27344 32646 27356
rect 33704 27328 33732 27424
rect 33965 27421 33977 27455
rect 34011 27421 34023 27455
rect 33965 27415 34023 27421
rect 33980 27384 34008 27415
rect 34054 27412 34060 27464
rect 34112 27452 34118 27464
rect 34164 27461 34192 27492
rect 37366 27480 37372 27492
rect 37424 27480 37430 27532
rect 37936 27529 37964 27560
rect 38289 27557 38301 27560
rect 38335 27557 38347 27591
rect 38289 27551 38347 27557
rect 37921 27523 37979 27529
rect 37921 27489 37933 27523
rect 37967 27489 37979 27523
rect 37921 27483 37979 27489
rect 38028 27492 38884 27520
rect 34149 27455 34207 27461
rect 34149 27452 34161 27455
rect 34112 27424 34161 27452
rect 34112 27412 34118 27424
rect 34149 27421 34161 27424
rect 34195 27421 34207 27455
rect 34698 27452 34704 27464
rect 34149 27415 34207 27421
rect 34256 27424 34704 27452
rect 34256 27384 34284 27424
rect 34698 27412 34704 27424
rect 34756 27412 34762 27464
rect 34885 27455 34943 27461
rect 34885 27421 34897 27455
rect 34931 27452 34943 27455
rect 34974 27452 34980 27464
rect 34931 27424 34980 27452
rect 34931 27421 34943 27424
rect 34885 27415 34943 27421
rect 34974 27412 34980 27424
rect 35032 27412 35038 27464
rect 35437 27455 35495 27461
rect 35437 27421 35449 27455
rect 35483 27421 35495 27455
rect 35437 27415 35495 27421
rect 35621 27455 35679 27461
rect 35621 27421 35633 27455
rect 35667 27452 35679 27455
rect 36354 27452 36360 27464
rect 35667 27424 36360 27452
rect 35667 27421 35679 27424
rect 35621 27415 35679 27421
rect 33980 27356 34284 27384
rect 34422 27344 34428 27396
rect 34480 27344 34486 27396
rect 35066 27344 35072 27396
rect 35124 27384 35130 27396
rect 35452 27384 35480 27415
rect 36354 27412 36360 27424
rect 36412 27412 36418 27464
rect 36630 27412 36636 27464
rect 36688 27412 36694 27464
rect 37274 27412 37280 27464
rect 37332 27452 37338 27464
rect 38028 27461 38056 27492
rect 38856 27464 38884 27492
rect 37553 27455 37611 27461
rect 37553 27452 37565 27455
rect 37332 27424 37565 27452
rect 37332 27412 37338 27424
rect 37553 27421 37565 27424
rect 37599 27421 37611 27455
rect 37553 27415 37611 27421
rect 38013 27455 38071 27461
rect 38013 27421 38025 27455
rect 38059 27421 38071 27455
rect 38013 27415 38071 27421
rect 38194 27412 38200 27464
rect 38252 27452 38258 27464
rect 38252 27424 38424 27452
rect 38252 27412 38258 27424
rect 36648 27384 36676 27412
rect 35124 27356 36676 27384
rect 37093 27387 37151 27393
rect 35124 27344 35130 27356
rect 37093 27353 37105 27387
rect 37139 27384 37151 27387
rect 37139 27356 38240 27384
rect 37139 27353 37151 27356
rect 37093 27347 37151 27353
rect 31481 27319 31539 27325
rect 31481 27316 31493 27319
rect 26252 27288 31493 27316
rect 31481 27285 31493 27288
rect 31527 27285 31539 27319
rect 31481 27279 31539 27285
rect 32122 27276 32128 27328
rect 32180 27316 32186 27328
rect 32217 27319 32275 27325
rect 32217 27316 32229 27319
rect 32180 27288 32229 27316
rect 32180 27276 32186 27288
rect 32217 27285 32229 27288
rect 32263 27285 32275 27319
rect 32217 27279 32275 27285
rect 33226 27276 33232 27328
rect 33284 27316 33290 27328
rect 33502 27316 33508 27328
rect 33284 27288 33508 27316
rect 33284 27276 33290 27288
rect 33502 27276 33508 27288
rect 33560 27276 33566 27328
rect 33686 27276 33692 27328
rect 33744 27276 33750 27328
rect 33962 27276 33968 27328
rect 34020 27316 34026 27328
rect 34698 27316 34704 27328
rect 34020 27288 34704 27316
rect 34020 27276 34026 27288
rect 34698 27276 34704 27288
rect 34756 27276 34762 27328
rect 34790 27276 34796 27328
rect 34848 27276 34854 27328
rect 35526 27276 35532 27328
rect 35584 27276 35590 27328
rect 38212 27325 38240 27356
rect 38286 27344 38292 27396
rect 38344 27344 38350 27396
rect 38197 27319 38255 27325
rect 38197 27285 38209 27319
rect 38243 27285 38255 27319
rect 38396 27316 38424 27424
rect 38470 27412 38476 27464
rect 38528 27452 38534 27464
rect 38565 27455 38623 27461
rect 38565 27452 38577 27455
rect 38528 27424 38577 27452
rect 38528 27412 38534 27424
rect 38565 27421 38577 27424
rect 38611 27421 38623 27455
rect 38565 27415 38623 27421
rect 38838 27412 38844 27464
rect 38896 27412 38902 27464
rect 39577 27455 39635 27461
rect 39577 27421 39589 27455
rect 39623 27452 39635 27455
rect 39850 27452 39856 27464
rect 39623 27424 39856 27452
rect 39623 27421 39635 27424
rect 39577 27415 39635 27421
rect 39850 27412 39856 27424
rect 39908 27412 39914 27464
rect 40037 27455 40095 27461
rect 40037 27421 40049 27455
rect 40083 27452 40095 27455
rect 41690 27452 41696 27464
rect 40083 27424 41696 27452
rect 40083 27421 40095 27424
rect 40037 27415 40095 27421
rect 41690 27412 41696 27424
rect 41748 27412 41754 27464
rect 38473 27319 38531 27325
rect 38473 27316 38485 27319
rect 38396 27288 38485 27316
rect 38197 27279 38255 27285
rect 38473 27285 38485 27288
rect 38519 27285 38531 27319
rect 38473 27279 38531 27285
rect 39390 27276 39396 27328
rect 39448 27276 39454 27328
rect 1104 27226 41400 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 41400 27226
rect 1104 27152 41400 27174
rect 5534 27072 5540 27124
rect 5592 27112 5598 27124
rect 5994 27112 6000 27124
rect 5592 27084 6000 27112
rect 5592 27072 5598 27084
rect 5994 27072 6000 27084
rect 6052 27072 6058 27124
rect 6917 27115 6975 27121
rect 6917 27081 6929 27115
rect 6963 27112 6975 27115
rect 7006 27112 7012 27124
rect 6963 27084 7012 27112
rect 6963 27081 6975 27084
rect 6917 27075 6975 27081
rect 7006 27072 7012 27084
rect 7064 27072 7070 27124
rect 7742 27112 7748 27124
rect 7484 27084 7748 27112
rect 3050 27044 3056 27056
rect 2990 27016 3056 27044
rect 3050 27004 3056 27016
rect 3108 27044 3114 27056
rect 3878 27044 3884 27056
rect 3108 27016 3884 27044
rect 3108 27004 3114 27016
rect 3878 27004 3884 27016
rect 3936 27004 3942 27056
rect 5813 27047 5871 27053
rect 5813 27013 5825 27047
rect 5859 27044 5871 27047
rect 5902 27044 5908 27056
rect 5859 27016 5908 27044
rect 5859 27013 5871 27016
rect 5813 27007 5871 27013
rect 5902 27004 5908 27016
rect 5960 27004 5966 27056
rect 6733 27047 6791 27053
rect 6733 27013 6745 27047
rect 6779 27044 6791 27047
rect 6822 27044 6828 27056
rect 6779 27016 6828 27044
rect 6779 27013 6791 27016
rect 6733 27007 6791 27013
rect 6822 27004 6828 27016
rect 6880 27004 6886 27056
rect 7484 26985 7512 27084
rect 7742 27072 7748 27084
rect 7800 27072 7806 27124
rect 7926 27072 7932 27124
rect 7984 27072 7990 27124
rect 8294 27072 8300 27124
rect 8352 27112 8358 27124
rect 8665 27115 8723 27121
rect 8665 27112 8677 27115
rect 8352 27084 8677 27112
rect 8352 27072 8358 27084
rect 8665 27081 8677 27084
rect 8711 27081 8723 27115
rect 8665 27075 8723 27081
rect 8938 27072 8944 27124
rect 8996 27112 9002 27124
rect 9033 27115 9091 27121
rect 9033 27112 9045 27115
rect 8996 27084 9045 27112
rect 8996 27072 9002 27084
rect 9033 27081 9045 27084
rect 9079 27112 9091 27115
rect 9122 27112 9128 27124
rect 9079 27084 9128 27112
rect 9079 27081 9091 27084
rect 9033 27075 9091 27081
rect 9122 27072 9128 27084
rect 9180 27072 9186 27124
rect 9766 27112 9772 27124
rect 9600 27084 9772 27112
rect 7944 27044 7972 27072
rect 9600 27053 9628 27084
rect 9766 27072 9772 27084
rect 9824 27072 9830 27124
rect 9858 27072 9864 27124
rect 9916 27072 9922 27124
rect 10042 27072 10048 27124
rect 10100 27112 10106 27124
rect 10597 27115 10655 27121
rect 10597 27112 10609 27115
rect 10100 27084 10609 27112
rect 10100 27072 10106 27084
rect 10597 27081 10609 27084
rect 10643 27081 10655 27115
rect 10597 27075 10655 27081
rect 12342 27072 12348 27124
rect 12400 27072 12406 27124
rect 12526 27072 12532 27124
rect 12584 27112 12590 27124
rect 12621 27115 12679 27121
rect 12621 27112 12633 27115
rect 12584 27084 12633 27112
rect 12584 27072 12590 27084
rect 12621 27081 12633 27084
rect 12667 27081 12679 27115
rect 12621 27075 12679 27081
rect 12802 27072 12808 27124
rect 12860 27072 12866 27124
rect 12986 27072 12992 27124
rect 13044 27112 13050 27124
rect 13044 27084 13308 27112
rect 13044 27072 13050 27084
rect 7760 27016 7972 27044
rect 8205 27047 8263 27053
rect 7760 26985 7788 27016
rect 8205 27013 8217 27047
rect 8251 27044 8263 27047
rect 9585 27047 9643 27053
rect 8251 27016 9536 27044
rect 8251 27013 8263 27016
rect 8205 27007 8263 27013
rect 7469 26979 7527 26985
rect 7469 26945 7481 26979
rect 7515 26945 7527 26979
rect 7469 26939 7527 26945
rect 7561 26979 7619 26985
rect 7561 26945 7573 26979
rect 7607 26945 7619 26979
rect 7561 26939 7619 26945
rect 7745 26979 7803 26985
rect 7745 26945 7757 26979
rect 7791 26945 7803 26979
rect 7745 26939 7803 26945
rect 7837 26979 7895 26985
rect 7837 26945 7849 26979
rect 7883 26945 7895 26979
rect 7837 26939 7895 26945
rect 1394 26868 1400 26920
rect 1452 26908 1458 26920
rect 1489 26911 1547 26917
rect 1489 26908 1501 26911
rect 1452 26880 1501 26908
rect 1452 26868 1458 26880
rect 1489 26877 1501 26880
rect 1535 26908 1547 26911
rect 1535 26880 1624 26908
rect 1535 26877 1547 26880
rect 1489 26871 1547 26877
rect 1596 26772 1624 26880
rect 1762 26868 1768 26920
rect 1820 26868 1826 26920
rect 6086 26868 6092 26920
rect 6144 26908 6150 26920
rect 7009 26911 7067 26917
rect 7009 26908 7021 26911
rect 6144 26880 7021 26908
rect 6144 26868 6150 26880
rect 7009 26877 7021 26880
rect 7055 26908 7067 26911
rect 7374 26908 7380 26920
rect 7055 26880 7380 26908
rect 7055 26877 7067 26880
rect 7009 26871 7067 26877
rect 7374 26868 7380 26880
rect 7432 26868 7438 26920
rect 2866 26800 2872 26852
rect 2924 26840 2930 26852
rect 5537 26843 5595 26849
rect 5537 26840 5549 26843
rect 2924 26812 5549 26840
rect 2924 26800 2930 26812
rect 5537 26809 5549 26812
rect 5583 26809 5595 26843
rect 7576 26840 7604 26939
rect 7852 26908 7880 26939
rect 7926 26936 7932 26988
rect 7984 26936 7990 26988
rect 8110 26985 8116 26988
rect 8077 26979 8116 26985
rect 8077 26945 8089 26979
rect 8077 26939 8116 26945
rect 8110 26936 8116 26939
rect 8168 26936 8174 26988
rect 8294 26936 8300 26988
rect 8352 26936 8358 26988
rect 8435 26979 8493 26985
rect 8435 26945 8447 26979
rect 8481 26976 8493 26979
rect 8570 26976 8576 26988
rect 8481 26948 8576 26976
rect 8481 26945 8493 26948
rect 8435 26939 8493 26945
rect 8570 26936 8576 26948
rect 8628 26936 8634 26988
rect 8846 26936 8852 26988
rect 8904 26936 8910 26988
rect 9398 26985 9404 26988
rect 9125 26979 9183 26985
rect 9125 26945 9137 26979
rect 9171 26945 9183 26979
rect 9125 26939 9183 26945
rect 9217 26979 9275 26985
rect 9217 26945 9229 26979
rect 9263 26945 9275 26979
rect 9217 26939 9275 26945
rect 9365 26979 9404 26985
rect 9365 26945 9377 26979
rect 9365 26939 9404 26945
rect 7852 26880 8616 26908
rect 8588 26849 8616 26880
rect 8573 26843 8631 26849
rect 7576 26812 7972 26840
rect 5537 26803 5595 26809
rect 2406 26772 2412 26784
rect 1596 26744 2412 26772
rect 2406 26732 2412 26744
rect 2464 26732 2470 26784
rect 3234 26732 3240 26784
rect 3292 26732 3298 26784
rect 3510 26732 3516 26784
rect 3568 26772 3574 26784
rect 4798 26772 4804 26784
rect 3568 26744 4804 26772
rect 3568 26732 3574 26744
rect 4798 26732 4804 26744
rect 4856 26772 4862 26784
rect 6457 26775 6515 26781
rect 6457 26772 6469 26775
rect 4856 26744 6469 26772
rect 4856 26732 4862 26744
rect 6457 26741 6469 26744
rect 6503 26741 6515 26775
rect 6457 26735 6515 26741
rect 7285 26775 7343 26781
rect 7285 26741 7297 26775
rect 7331 26772 7343 26775
rect 7834 26772 7840 26784
rect 7331 26744 7840 26772
rect 7331 26741 7343 26744
rect 7285 26735 7343 26741
rect 7834 26732 7840 26744
rect 7892 26732 7898 26784
rect 7944 26772 7972 26812
rect 8573 26809 8585 26843
rect 8619 26809 8631 26843
rect 8573 26803 8631 26809
rect 8662 26772 8668 26784
rect 7944 26744 8668 26772
rect 8662 26732 8668 26744
rect 8720 26732 8726 26784
rect 9030 26732 9036 26784
rect 9088 26772 9094 26784
rect 9140 26772 9168 26939
rect 9232 26840 9260 26939
rect 9398 26936 9404 26939
rect 9456 26936 9462 26988
rect 9508 26985 9536 27016
rect 9585 27013 9597 27047
rect 9631 27013 9643 27047
rect 9585 27007 9643 27013
rect 10229 27047 10287 27053
rect 10229 27013 10241 27047
rect 10275 27044 10287 27047
rect 10686 27044 10692 27056
rect 10275 27016 10692 27044
rect 10275 27013 10287 27016
rect 10229 27007 10287 27013
rect 10686 27004 10692 27016
rect 10744 27044 10750 27056
rect 11790 27044 11796 27056
rect 10744 27016 11796 27044
rect 10744 27004 10750 27016
rect 11790 27004 11796 27016
rect 11848 27044 11854 27056
rect 12066 27044 12072 27056
rect 11848 27016 12072 27044
rect 11848 27004 11854 27016
rect 12066 27004 12072 27016
rect 12124 27004 12130 27056
rect 9493 26979 9551 26985
rect 9493 26945 9505 26979
rect 9539 26945 9551 26979
rect 9493 26939 9551 26945
rect 9721 26979 9779 26985
rect 9721 26945 9733 26979
rect 9767 26976 9779 26979
rect 9767 26948 9868 26976
rect 9767 26945 9779 26948
rect 9721 26939 9779 26945
rect 9508 26908 9536 26939
rect 9508 26880 9628 26908
rect 9490 26840 9496 26852
rect 9232 26812 9496 26840
rect 9490 26800 9496 26812
rect 9548 26800 9554 26852
rect 9600 26840 9628 26880
rect 9674 26840 9680 26852
rect 9600 26812 9680 26840
rect 9674 26800 9680 26812
rect 9732 26800 9738 26852
rect 9840 26772 9868 26948
rect 9950 26936 9956 26988
rect 10008 26936 10014 26988
rect 10042 26936 10048 26988
rect 10100 26936 10106 26988
rect 10318 26936 10324 26988
rect 10376 26936 10382 26988
rect 10418 26979 10476 26985
rect 10418 26945 10430 26979
rect 10464 26945 10476 26979
rect 10418 26939 10476 26945
rect 12437 26979 12495 26985
rect 12437 26945 12449 26979
rect 12483 26976 12495 26979
rect 12526 26976 12532 26988
rect 12483 26948 12532 26976
rect 12483 26945 12495 26948
rect 12437 26939 12495 26945
rect 10433 26772 10461 26939
rect 12526 26936 12532 26948
rect 12584 26936 12590 26988
rect 12713 26979 12771 26985
rect 12713 26945 12725 26979
rect 12759 26976 12771 26979
rect 12820 26976 12848 27072
rect 13280 27053 13308 27084
rect 13998 27072 14004 27124
rect 14056 27112 14062 27124
rect 14369 27115 14427 27121
rect 14369 27112 14381 27115
rect 14056 27084 14381 27112
rect 14056 27072 14062 27084
rect 14369 27081 14381 27084
rect 14415 27112 14427 27115
rect 14550 27112 14556 27124
rect 14415 27084 14556 27112
rect 14415 27081 14427 27084
rect 14369 27075 14427 27081
rect 14550 27072 14556 27084
rect 14608 27072 14614 27124
rect 14918 27072 14924 27124
rect 14976 27072 14982 27124
rect 15746 27072 15752 27124
rect 15804 27072 15810 27124
rect 15930 27072 15936 27124
rect 15988 27112 15994 27124
rect 15988 27084 16444 27112
rect 15988 27072 15994 27084
rect 13265 27047 13323 27053
rect 13265 27013 13277 27047
rect 13311 27013 13323 27047
rect 13265 27007 13323 27013
rect 13722 27004 13728 27056
rect 13780 27044 13786 27056
rect 14737 27047 14795 27053
rect 14737 27044 14749 27047
rect 13780 27016 14749 27044
rect 13780 27004 13786 27016
rect 14737 27013 14749 27016
rect 14783 27013 14795 27047
rect 14737 27007 14795 27013
rect 15028 27016 16068 27044
rect 12759 26948 12848 26976
rect 12897 26979 12955 26985
rect 12897 26966 12909 26979
rect 12759 26945 12771 26948
rect 12713 26939 12771 26945
rect 12876 26945 12909 26966
rect 12943 26945 12955 26979
rect 12876 26939 12955 26945
rect 13045 26979 13103 26985
rect 13045 26945 13057 26979
rect 13091 26945 13103 26979
rect 13045 26939 13103 26945
rect 12876 26938 12940 26939
rect 11882 26868 11888 26920
rect 11940 26868 11946 26920
rect 12253 26843 12311 26849
rect 12253 26809 12265 26843
rect 12299 26840 12311 26843
rect 12434 26840 12440 26852
rect 12299 26812 12440 26840
rect 12299 26809 12311 26812
rect 12253 26803 12311 26809
rect 12434 26800 12440 26812
rect 12492 26800 12498 26852
rect 12876 26840 12904 26938
rect 13060 26908 13088 26939
rect 13170 26936 13176 26988
rect 13228 26936 13234 26988
rect 13403 26979 13461 26985
rect 13403 26945 13415 26979
rect 13449 26976 13461 26979
rect 13538 26976 13544 26988
rect 13449 26948 13544 26976
rect 13449 26945 13481 26948
rect 13403 26939 13481 26945
rect 13060 26880 13400 26908
rect 13372 26852 13400 26880
rect 13170 26840 13176 26852
rect 12876 26812 13176 26840
rect 13170 26800 13176 26812
rect 13228 26800 13234 26852
rect 13354 26800 13360 26852
rect 13412 26800 13418 26852
rect 10778 26772 10784 26784
rect 9088 26744 10784 26772
rect 9088 26732 9094 26744
rect 10778 26732 10784 26744
rect 10836 26772 10842 26784
rect 13453 26772 13481 26939
rect 13538 26936 13544 26948
rect 13596 26936 13602 26988
rect 13814 26936 13820 26988
rect 13872 26976 13878 26988
rect 13909 26979 13967 26985
rect 13909 26976 13921 26979
rect 13872 26948 13921 26976
rect 13872 26936 13878 26948
rect 13909 26945 13921 26948
rect 13955 26945 13967 26979
rect 13909 26939 13967 26945
rect 14182 26936 14188 26988
rect 14240 26936 14246 26988
rect 14277 26979 14335 26985
rect 14277 26945 14289 26979
rect 14323 26976 14335 26979
rect 14366 26976 14372 26988
rect 14323 26948 14372 26976
rect 14323 26945 14335 26948
rect 14277 26939 14335 26945
rect 14366 26936 14372 26948
rect 14424 26936 14430 26988
rect 14550 26936 14556 26988
rect 14608 26976 14614 26988
rect 15028 26985 15056 27016
rect 14829 26979 14887 26985
rect 14829 26976 14841 26979
rect 14608 26948 14841 26976
rect 14608 26936 14614 26948
rect 14829 26945 14841 26948
rect 14875 26945 14887 26979
rect 15013 26979 15071 26985
rect 15013 26976 15025 26979
rect 14829 26939 14887 26945
rect 14936 26948 15025 26976
rect 14645 26911 14703 26917
rect 14645 26908 14657 26911
rect 13832 26880 14657 26908
rect 13541 26843 13599 26849
rect 13541 26809 13553 26843
rect 13587 26840 13599 26843
rect 13832 26840 13860 26880
rect 14645 26877 14657 26880
rect 14691 26877 14703 26911
rect 14645 26871 14703 26877
rect 13587 26812 13860 26840
rect 13587 26809 13599 26812
rect 13541 26803 13599 26809
rect 14090 26800 14096 26852
rect 14148 26800 14154 26852
rect 14936 26840 14964 26948
rect 15013 26945 15025 26948
rect 15059 26945 15071 26979
rect 15013 26939 15071 26945
rect 15102 26936 15108 26988
rect 15160 26936 15166 26988
rect 15286 26985 15292 26988
rect 15253 26979 15292 26985
rect 15253 26945 15265 26979
rect 15253 26939 15292 26945
rect 15286 26936 15292 26939
rect 15344 26936 15350 26988
rect 15378 26936 15384 26988
rect 15436 26936 15442 26988
rect 15470 26936 15476 26988
rect 15528 26936 15534 26988
rect 15562 26936 15568 26988
rect 15620 26985 15626 26988
rect 16040 26985 16068 27016
rect 16416 26985 16444 27084
rect 16574 27072 16580 27124
rect 16632 27112 16638 27124
rect 16853 27115 16911 27121
rect 16853 27112 16865 27115
rect 16632 27084 16865 27112
rect 16632 27072 16638 27084
rect 16853 27081 16865 27084
rect 16899 27081 16911 27115
rect 16853 27075 16911 27081
rect 17954 27072 17960 27124
rect 18012 27112 18018 27124
rect 18233 27115 18291 27121
rect 18233 27112 18245 27115
rect 18012 27084 18245 27112
rect 18012 27072 18018 27084
rect 18233 27081 18245 27084
rect 18279 27081 18291 27115
rect 18233 27075 18291 27081
rect 19061 27115 19119 27121
rect 19061 27081 19073 27115
rect 19107 27081 19119 27115
rect 19061 27075 19119 27081
rect 18350 27047 18408 27053
rect 16500 27016 17724 27044
rect 15620 26976 15628 26985
rect 16025 26979 16083 26985
rect 15620 26948 15665 26976
rect 15620 26939 15628 26948
rect 16025 26945 16037 26979
rect 16071 26945 16083 26979
rect 16025 26939 16083 26945
rect 16393 26979 16451 26985
rect 16393 26945 16405 26979
rect 16439 26945 16451 26979
rect 16393 26939 16451 26945
rect 15620 26936 15626 26939
rect 15841 26911 15899 26917
rect 15841 26908 15853 26911
rect 15028 26880 15853 26908
rect 15028 26852 15056 26880
rect 15841 26877 15853 26880
rect 15887 26877 15899 26911
rect 16500 26908 16528 27016
rect 16669 26979 16727 26985
rect 16669 26945 16681 26979
rect 16715 26945 16727 26979
rect 16669 26939 16727 26945
rect 17497 26979 17555 26985
rect 17497 26945 17509 26979
rect 17543 26976 17555 26979
rect 17586 26976 17592 26988
rect 17543 26948 17592 26976
rect 17543 26945 17555 26948
rect 17497 26939 17555 26945
rect 15841 26871 15899 26877
rect 15948 26880 16528 26908
rect 14384 26812 14964 26840
rect 10836 26744 13481 26772
rect 10836 26732 10842 26744
rect 13722 26732 13728 26784
rect 13780 26732 13786 26784
rect 13906 26732 13912 26784
rect 13964 26772 13970 26784
rect 14384 26772 14412 26812
rect 15010 26800 15016 26852
rect 15068 26800 15074 26852
rect 15378 26800 15384 26852
rect 15436 26840 15442 26852
rect 15948 26840 15976 26880
rect 15436 26812 15976 26840
rect 15436 26800 15442 26812
rect 16298 26800 16304 26852
rect 16356 26800 16362 26852
rect 16684 26840 16712 26939
rect 17586 26936 17592 26948
rect 17644 26936 17650 26988
rect 17696 26985 17724 27016
rect 18350 27013 18362 27047
rect 18396 27044 18408 27047
rect 19076 27044 19104 27075
rect 19242 27072 19248 27124
rect 19300 27072 19306 27124
rect 22094 27072 22100 27124
rect 22152 27072 22158 27124
rect 22922 27072 22928 27124
rect 22980 27112 22986 27124
rect 23109 27115 23167 27121
rect 23109 27112 23121 27115
rect 22980 27084 23121 27112
rect 22980 27072 22986 27084
rect 23109 27081 23121 27084
rect 23155 27081 23167 27115
rect 23109 27075 23167 27081
rect 23382 27072 23388 27124
rect 23440 27072 23446 27124
rect 23566 27072 23572 27124
rect 23624 27112 23630 27124
rect 23624 27084 24716 27112
rect 23624 27072 23630 27084
rect 18396 27016 19104 27044
rect 18396 27013 18408 27016
rect 18350 27007 18408 27013
rect 17681 26979 17739 26985
rect 17681 26945 17693 26979
rect 17727 26976 17739 26979
rect 17865 26979 17923 26985
rect 17865 26976 17877 26979
rect 17727 26948 17877 26976
rect 17727 26945 17739 26948
rect 17681 26939 17739 26945
rect 17865 26945 17877 26948
rect 17911 26945 17923 26979
rect 17865 26939 17923 26945
rect 18064 26948 18368 26976
rect 17313 26911 17371 26917
rect 17313 26877 17325 26911
rect 17359 26908 17371 26911
rect 18064 26908 18092 26948
rect 18340 26920 18368 26948
rect 18690 26936 18696 26988
rect 18748 26976 18754 26988
rect 19260 26976 19288 27072
rect 19978 27004 19984 27056
rect 20036 27044 20042 27056
rect 20990 27044 20996 27056
rect 20036 27016 20996 27044
rect 20036 27004 20042 27016
rect 20990 27004 20996 27016
rect 21048 27004 21054 27056
rect 18748 26948 19288 26976
rect 18748 26936 18754 26948
rect 19334 26936 19340 26988
rect 19392 26936 19398 26988
rect 19705 26979 19763 26985
rect 19705 26976 19717 26979
rect 19536 26948 19717 26976
rect 17359 26880 18092 26908
rect 18141 26911 18199 26917
rect 17359 26877 17371 26880
rect 17313 26871 17371 26877
rect 18141 26877 18153 26911
rect 18187 26877 18199 26911
rect 18141 26871 18199 26877
rect 18156 26840 18184 26871
rect 18322 26868 18328 26920
rect 18380 26868 18386 26920
rect 18785 26911 18843 26917
rect 18785 26877 18797 26911
rect 18831 26908 18843 26911
rect 19536 26908 19564 26948
rect 19705 26945 19717 26948
rect 19751 26976 19763 26979
rect 22002 26976 22008 26988
rect 19751 26948 22008 26976
rect 19751 26945 19763 26948
rect 19705 26939 19763 26945
rect 22002 26936 22008 26948
rect 22060 26936 22066 26988
rect 22112 26976 22140 27072
rect 22281 26979 22339 26985
rect 22281 26976 22293 26979
rect 22112 26948 22293 26976
rect 22281 26945 22293 26948
rect 22327 26945 22339 26979
rect 22281 26939 22339 26945
rect 22649 26979 22707 26985
rect 22649 26945 22661 26979
rect 22695 26976 22707 26979
rect 22830 26976 22836 26988
rect 22695 26948 22836 26976
rect 22695 26945 22707 26948
rect 22649 26939 22707 26945
rect 22830 26936 22836 26948
rect 22888 26936 22894 26988
rect 22925 26979 22983 26985
rect 22925 26945 22937 26979
rect 22971 26945 22983 26979
rect 22925 26939 22983 26945
rect 23201 26979 23259 26985
rect 23201 26945 23213 26979
rect 23247 26976 23259 26979
rect 23400 26976 23428 27072
rect 23247 26948 23428 26976
rect 23584 26976 23612 27072
rect 24688 27044 24716 27084
rect 28626 27072 28632 27124
rect 28684 27112 28690 27124
rect 30834 27112 30840 27124
rect 28684 27084 30840 27112
rect 28684 27072 28690 27084
rect 25409 27047 25467 27053
rect 25409 27044 25421 27047
rect 24688 27016 25421 27044
rect 25409 27013 25421 27016
rect 25455 27013 25467 27047
rect 25409 27007 25467 27013
rect 26602 27004 26608 27056
rect 26660 27044 26666 27056
rect 29086 27044 29092 27056
rect 26660 27016 29092 27044
rect 26660 27004 26666 27016
rect 29086 27004 29092 27016
rect 29144 27004 29150 27056
rect 23845 26979 23903 26985
rect 23845 26976 23857 26979
rect 23584 26948 23857 26976
rect 23247 26945 23259 26948
rect 23201 26939 23259 26945
rect 23845 26945 23857 26948
rect 23891 26945 23903 26979
rect 23845 26939 23903 26945
rect 24305 26979 24363 26985
rect 24305 26945 24317 26979
rect 24351 26976 24363 26979
rect 25038 26976 25044 26988
rect 24351 26948 25044 26976
rect 24351 26945 24363 26948
rect 24305 26939 24363 26945
rect 18831 26880 19564 26908
rect 18831 26877 18843 26880
rect 18785 26871 18843 26877
rect 19610 26868 19616 26920
rect 19668 26908 19674 26920
rect 21082 26908 21088 26920
rect 19668 26880 21088 26908
rect 19668 26868 19674 26880
rect 21082 26868 21088 26880
rect 21140 26868 21146 26920
rect 21821 26911 21879 26917
rect 21821 26877 21833 26911
rect 21867 26908 21879 26911
rect 22741 26911 22799 26917
rect 21867 26880 22094 26908
rect 21867 26877 21879 26880
rect 21821 26871 21879 26877
rect 19153 26843 19211 26849
rect 19153 26840 19165 26843
rect 16684 26812 17816 26840
rect 18156 26812 19165 26840
rect 13964 26744 14412 26772
rect 13964 26732 13970 26744
rect 14458 26732 14464 26784
rect 14516 26772 14522 26784
rect 14553 26775 14611 26781
rect 14553 26772 14565 26775
rect 14516 26744 14565 26772
rect 14516 26732 14522 26744
rect 14553 26741 14565 26744
rect 14599 26772 14611 26775
rect 16574 26772 16580 26784
rect 14599 26744 16580 26772
rect 14599 26741 14611 26744
rect 14553 26735 14611 26741
rect 16574 26732 16580 26744
rect 16632 26732 16638 26784
rect 17788 26772 17816 26812
rect 19153 26809 19165 26812
rect 19199 26809 19211 26843
rect 19153 26803 19211 26809
rect 19242 26800 19248 26852
rect 19300 26840 19306 26852
rect 21913 26843 21971 26849
rect 21913 26840 21925 26843
rect 19300 26812 21925 26840
rect 19300 26800 19306 26812
rect 21913 26809 21925 26812
rect 21959 26809 21971 26843
rect 21913 26803 21971 26809
rect 22066 26784 22094 26880
rect 22741 26877 22753 26911
rect 22787 26877 22799 26911
rect 22940 26908 22968 26939
rect 25038 26936 25044 26948
rect 25096 26936 25102 26988
rect 25130 26936 25136 26988
rect 25188 26976 25194 26988
rect 25593 26979 25651 26985
rect 25593 26976 25605 26979
rect 25188 26948 25605 26976
rect 25188 26936 25194 26948
rect 25593 26945 25605 26948
rect 25639 26945 25651 26979
rect 25593 26939 25651 26945
rect 25869 26979 25927 26985
rect 25869 26945 25881 26979
rect 25915 26976 25927 26979
rect 26418 26976 26424 26988
rect 25915 26948 26424 26976
rect 25915 26945 25927 26948
rect 25869 26939 25927 26945
rect 26418 26936 26424 26948
rect 26476 26936 26482 26988
rect 28166 26976 28172 26988
rect 26528 26948 28172 26976
rect 23477 26911 23535 26917
rect 22940 26880 23428 26908
rect 22741 26871 22799 26877
rect 22756 26784 22784 26871
rect 23400 26849 23428 26880
rect 23477 26877 23489 26911
rect 23523 26877 23535 26911
rect 23477 26871 23535 26877
rect 23385 26843 23443 26849
rect 23385 26809 23397 26843
rect 23431 26809 23443 26843
rect 23492 26840 23520 26871
rect 23566 26868 23572 26920
rect 23624 26908 23630 26920
rect 23661 26911 23719 26917
rect 23661 26908 23673 26911
rect 23624 26880 23673 26908
rect 23624 26868 23630 26880
rect 23661 26877 23673 26880
rect 23707 26908 23719 26911
rect 24026 26908 24032 26920
rect 23707 26880 24032 26908
rect 23707 26877 23719 26880
rect 23661 26871 23719 26877
rect 24026 26868 24032 26880
rect 24084 26868 24090 26920
rect 24581 26911 24639 26917
rect 24581 26877 24593 26911
rect 24627 26908 24639 26911
rect 24762 26908 24768 26920
rect 24627 26880 24768 26908
rect 24627 26877 24639 26880
rect 24581 26871 24639 26877
rect 24596 26840 24624 26871
rect 24762 26868 24768 26880
rect 24820 26908 24826 26920
rect 26528 26908 26556 26948
rect 28166 26936 28172 26948
rect 28224 26976 28230 26988
rect 28534 26976 28540 26988
rect 28224 26948 28540 26976
rect 28224 26936 28230 26948
rect 28534 26936 28540 26948
rect 28592 26936 28598 26988
rect 29472 26985 29500 27084
rect 30834 27072 30840 27084
rect 30892 27072 30898 27124
rect 31110 27072 31116 27124
rect 31168 27072 31174 27124
rect 31573 27115 31631 27121
rect 31573 27081 31585 27115
rect 31619 27112 31631 27115
rect 31754 27112 31760 27124
rect 31619 27084 31760 27112
rect 31619 27081 31631 27084
rect 31573 27075 31631 27081
rect 31754 27072 31760 27084
rect 31812 27072 31818 27124
rect 33410 27072 33416 27124
rect 33468 27072 33474 27124
rect 33689 27115 33747 27121
rect 33689 27081 33701 27115
rect 33735 27112 33747 27115
rect 33778 27112 33784 27124
rect 33735 27084 33784 27112
rect 33735 27081 33747 27084
rect 33689 27075 33747 27081
rect 33778 27072 33784 27084
rect 33836 27072 33842 27124
rect 34882 27112 34888 27124
rect 34164 27084 34888 27112
rect 33428 27044 33456 27072
rect 34164 27044 34192 27084
rect 34882 27072 34888 27084
rect 34940 27112 34946 27124
rect 39390 27112 39396 27124
rect 34940 27084 37044 27112
rect 34940 27072 34946 27084
rect 34974 27044 34980 27056
rect 29840 27016 33456 27044
rect 33520 27016 34192 27044
rect 29457 26979 29515 26985
rect 29457 26945 29469 26979
rect 29503 26945 29515 26979
rect 29457 26939 29515 26945
rect 29840 26920 29868 27016
rect 31202 26936 31208 26988
rect 31260 26976 31266 26988
rect 31389 26979 31447 26985
rect 31389 26976 31401 26979
rect 31260 26948 31401 26976
rect 31260 26936 31266 26948
rect 31389 26945 31401 26948
rect 31435 26945 31447 26979
rect 31389 26939 31447 26945
rect 32030 26936 32036 26988
rect 32088 26976 32094 26988
rect 32398 26976 32404 26988
rect 32088 26948 32404 26976
rect 32088 26936 32094 26948
rect 32398 26936 32404 26948
rect 32456 26976 32462 26988
rect 32456 26948 32720 26976
rect 32456 26936 32462 26948
rect 24820 26880 26556 26908
rect 26973 26911 27031 26917
rect 24820 26868 24826 26880
rect 26973 26877 26985 26911
rect 27019 26908 27031 26911
rect 27154 26908 27160 26920
rect 27019 26880 27160 26908
rect 27019 26877 27031 26880
rect 26973 26871 27031 26877
rect 27154 26868 27160 26880
rect 27212 26908 27218 26920
rect 28074 26908 28080 26920
rect 27212 26880 28080 26908
rect 27212 26868 27218 26880
rect 28074 26868 28080 26880
rect 28132 26868 28138 26920
rect 29733 26911 29791 26917
rect 29733 26877 29745 26911
rect 29779 26908 29791 26911
rect 29822 26908 29828 26920
rect 29779 26880 29828 26908
rect 29779 26877 29791 26880
rect 29733 26871 29791 26877
rect 29822 26868 29828 26880
rect 29880 26868 29886 26920
rect 30282 26868 30288 26920
rect 30340 26908 30346 26920
rect 31297 26911 31355 26917
rect 31297 26908 31309 26911
rect 30340 26880 31309 26908
rect 30340 26868 30346 26880
rect 31297 26877 31309 26880
rect 31343 26877 31355 26911
rect 31297 26871 31355 26877
rect 31662 26868 31668 26920
rect 31720 26868 31726 26920
rect 31757 26911 31815 26917
rect 31757 26877 31769 26911
rect 31803 26908 31815 26911
rect 32582 26908 32588 26920
rect 31803 26880 32588 26908
rect 31803 26877 31815 26880
rect 31757 26871 31815 26877
rect 32582 26868 32588 26880
rect 32640 26868 32646 26920
rect 32692 26908 32720 26948
rect 33318 26936 33324 26988
rect 33376 26976 33382 26988
rect 33520 26976 33548 27016
rect 33376 26948 33548 26976
rect 33376 26936 33382 26948
rect 33870 26936 33876 26988
rect 33928 26936 33934 26988
rect 34164 26985 34192 27016
rect 34808 27016 34980 27044
rect 34149 26979 34207 26985
rect 34149 26945 34161 26979
rect 34195 26945 34207 26979
rect 34149 26939 34207 26945
rect 34238 26936 34244 26988
rect 34296 26976 34302 26988
rect 34808 26985 34836 27016
rect 34974 27004 34980 27016
rect 35032 27044 35038 27056
rect 35032 27016 35848 27044
rect 35032 27004 35038 27016
rect 35820 26988 35848 27016
rect 36078 27004 36084 27056
rect 36136 27044 36142 27056
rect 36630 27044 36636 27056
rect 36136 27016 36636 27044
rect 36136 27004 36142 27016
rect 36630 27004 36636 27016
rect 36688 27004 36694 27056
rect 37016 26988 37044 27084
rect 39316 27084 39396 27112
rect 38286 27044 38292 27056
rect 37568 27016 38292 27044
rect 34425 26979 34483 26985
rect 34425 26976 34437 26979
rect 34296 26948 34437 26976
rect 34296 26936 34302 26948
rect 34425 26945 34437 26948
rect 34471 26945 34483 26979
rect 34425 26939 34483 26945
rect 34609 26979 34667 26985
rect 34609 26945 34621 26979
rect 34655 26976 34667 26979
rect 34793 26979 34851 26985
rect 34793 26976 34805 26979
rect 34655 26948 34805 26976
rect 34655 26945 34667 26948
rect 34609 26939 34667 26945
rect 34793 26945 34805 26948
rect 34839 26945 34851 26979
rect 34793 26939 34851 26945
rect 34885 26979 34943 26985
rect 34885 26945 34897 26979
rect 34931 26945 34943 26979
rect 34885 26939 34943 26945
rect 33686 26908 33692 26920
rect 32692 26880 33692 26908
rect 33686 26868 33692 26880
rect 33744 26908 33750 26920
rect 34900 26908 34928 26939
rect 35802 26936 35808 26988
rect 35860 26936 35866 26988
rect 36446 26936 36452 26988
rect 36504 26936 36510 26988
rect 36998 26936 37004 26988
rect 37056 26936 37062 26988
rect 37366 26936 37372 26988
rect 37424 26976 37430 26988
rect 37568 26985 37596 27016
rect 37553 26979 37611 26985
rect 37553 26976 37565 26979
rect 37424 26948 37565 26976
rect 37424 26936 37430 26948
rect 37553 26945 37565 26948
rect 37599 26945 37611 26979
rect 37553 26939 37611 26945
rect 37737 26979 37795 26985
rect 37737 26945 37749 26979
rect 37783 26976 37795 26979
rect 37826 26976 37832 26988
rect 37783 26948 37832 26976
rect 37783 26945 37795 26948
rect 37737 26939 37795 26945
rect 37826 26936 37832 26948
rect 37884 26936 37890 26988
rect 38028 26985 38056 27016
rect 38286 27004 38292 27016
rect 38344 27004 38350 27056
rect 39316 27053 39344 27084
rect 39390 27072 39396 27084
rect 39448 27072 39454 27124
rect 39482 27072 39488 27124
rect 39540 27112 39546 27124
rect 40773 27115 40831 27121
rect 40773 27112 40785 27115
rect 39540 27084 40785 27112
rect 39540 27072 39546 27084
rect 40773 27081 40785 27084
rect 40819 27081 40831 27115
rect 40773 27075 40831 27081
rect 39301 27047 39359 27053
rect 39301 27013 39313 27047
rect 39347 27013 39359 27047
rect 39301 27007 39359 27013
rect 40034 27004 40040 27056
rect 40092 27004 40098 27056
rect 38013 26979 38071 26985
rect 38013 26945 38025 26979
rect 38059 26945 38071 26979
rect 38013 26939 38071 26945
rect 38102 26936 38108 26988
rect 38160 26976 38166 26988
rect 38197 26979 38255 26985
rect 38197 26976 38209 26979
rect 38160 26948 38209 26976
rect 38160 26936 38166 26948
rect 38197 26945 38209 26948
rect 38243 26945 38255 26979
rect 38197 26939 38255 26945
rect 36464 26908 36492 26936
rect 33744 26880 36492 26908
rect 39025 26911 39083 26917
rect 33744 26868 33750 26880
rect 39025 26877 39037 26911
rect 39071 26877 39083 26911
rect 39025 26871 39083 26877
rect 27338 26840 27344 26852
rect 23492 26812 24624 26840
rect 25516 26812 27344 26840
rect 23385 26803 23443 26809
rect 18509 26775 18567 26781
rect 18509 26772 18521 26775
rect 17788 26744 18521 26772
rect 18509 26741 18521 26744
rect 18555 26741 18567 26775
rect 18509 26735 18567 26741
rect 18874 26732 18880 26784
rect 18932 26732 18938 26784
rect 19521 26775 19579 26781
rect 19521 26741 19533 26775
rect 19567 26772 19579 26775
rect 20162 26772 20168 26784
rect 19567 26744 20168 26772
rect 19567 26741 19579 26744
rect 19521 26735 19579 26741
rect 20162 26732 20168 26744
rect 20220 26732 20226 26784
rect 22066 26744 22100 26784
rect 22094 26732 22100 26744
rect 22152 26732 22158 26784
rect 22738 26732 22744 26784
rect 22796 26732 22802 26784
rect 23198 26732 23204 26784
rect 23256 26772 23262 26784
rect 23293 26775 23351 26781
rect 23293 26772 23305 26775
rect 23256 26744 23305 26772
rect 23256 26732 23262 26744
rect 23293 26741 23305 26744
rect 23339 26741 23351 26775
rect 23293 26735 23351 26741
rect 24026 26732 24032 26784
rect 24084 26732 24090 26784
rect 24210 26732 24216 26784
rect 24268 26772 24274 26784
rect 24397 26775 24455 26781
rect 24397 26772 24409 26775
rect 24268 26744 24409 26772
rect 24268 26732 24274 26744
rect 24397 26741 24409 26744
rect 24443 26741 24455 26775
rect 24397 26735 24455 26741
rect 24489 26775 24547 26781
rect 24489 26741 24501 26775
rect 24535 26772 24547 26775
rect 24578 26772 24584 26784
rect 24535 26744 24584 26772
rect 24535 26741 24547 26744
rect 24489 26735 24547 26741
rect 24578 26732 24584 26744
rect 24636 26732 24642 26784
rect 25130 26732 25136 26784
rect 25188 26772 25194 26784
rect 25516 26772 25544 26812
rect 27338 26800 27344 26812
rect 27396 26800 27402 26852
rect 34164 26812 34560 26840
rect 25188 26744 25544 26772
rect 25777 26775 25835 26781
rect 25188 26732 25194 26744
rect 25777 26741 25789 26775
rect 25823 26772 25835 26775
rect 26050 26772 26056 26784
rect 25823 26744 26056 26772
rect 25823 26741 25835 26744
rect 25777 26735 25835 26741
rect 26050 26732 26056 26744
rect 26108 26772 26114 26784
rect 27433 26775 27491 26781
rect 27433 26772 27445 26775
rect 26108 26744 27445 26772
rect 26108 26732 26114 26744
rect 27433 26741 27445 26744
rect 27479 26741 27491 26775
rect 27433 26735 27491 26741
rect 29270 26732 29276 26784
rect 29328 26732 29334 26784
rect 29454 26732 29460 26784
rect 29512 26772 29518 26784
rect 29641 26775 29699 26781
rect 29641 26772 29653 26775
rect 29512 26744 29653 26772
rect 29512 26732 29518 26744
rect 29641 26741 29653 26744
rect 29687 26772 29699 26775
rect 34164 26772 34192 26812
rect 29687 26744 34192 26772
rect 29687 26741 29699 26744
rect 29641 26735 29699 26741
rect 34422 26732 34428 26784
rect 34480 26732 34486 26784
rect 34532 26772 34560 26812
rect 34698 26800 34704 26852
rect 34756 26840 34762 26852
rect 34977 26843 35035 26849
rect 34977 26840 34989 26843
rect 34756 26812 34989 26840
rect 34756 26800 34762 26812
rect 34977 26809 34989 26812
rect 35023 26809 35035 26843
rect 34977 26803 35035 26809
rect 36538 26772 36544 26784
rect 34532 26744 36544 26772
rect 36538 26732 36544 26744
rect 36596 26732 36602 26784
rect 37553 26775 37611 26781
rect 37553 26741 37565 26775
rect 37599 26772 37611 26775
rect 37642 26772 37648 26784
rect 37599 26744 37648 26772
rect 37599 26741 37611 26744
rect 37553 26735 37611 26741
rect 37642 26732 37648 26744
rect 37700 26732 37706 26784
rect 38013 26775 38071 26781
rect 38013 26741 38025 26775
rect 38059 26772 38071 26775
rect 38838 26772 38844 26784
rect 38059 26744 38844 26772
rect 38059 26741 38071 26744
rect 38013 26735 38071 26741
rect 38838 26732 38844 26744
rect 38896 26732 38902 26784
rect 39040 26772 39068 26871
rect 39298 26772 39304 26784
rect 39040 26744 39304 26772
rect 39298 26732 39304 26744
rect 39356 26732 39362 26784
rect 1104 26682 41400 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 41400 26682
rect 1104 26608 41400 26630
rect 1762 26528 1768 26580
rect 1820 26568 1826 26580
rect 2133 26571 2191 26577
rect 2133 26568 2145 26571
rect 1820 26540 2145 26568
rect 1820 26528 1826 26540
rect 2133 26537 2145 26540
rect 2179 26537 2191 26571
rect 2133 26531 2191 26537
rect 5534 26528 5540 26580
rect 5592 26568 5598 26580
rect 8481 26571 8539 26577
rect 5592 26540 8340 26568
rect 5592 26528 5598 26540
rect 8312 26512 8340 26540
rect 8481 26537 8493 26571
rect 8527 26568 8539 26571
rect 8846 26568 8852 26580
rect 8527 26540 8852 26568
rect 8527 26537 8539 26540
rect 8481 26531 8539 26537
rect 8846 26528 8852 26540
rect 8904 26528 8910 26580
rect 9585 26571 9643 26577
rect 9585 26537 9597 26571
rect 9631 26537 9643 26571
rect 9585 26531 9643 26537
rect 2869 26503 2927 26509
rect 2869 26500 2881 26503
rect 2746 26472 2881 26500
rect 2317 26367 2375 26373
rect 2317 26333 2329 26367
rect 2363 26364 2375 26367
rect 2746 26364 2774 26472
rect 2869 26469 2881 26472
rect 2915 26469 2927 26503
rect 2869 26463 2927 26469
rect 5813 26503 5871 26509
rect 5813 26469 5825 26503
rect 5859 26500 5871 26503
rect 6546 26500 6552 26512
rect 5859 26472 6552 26500
rect 5859 26469 5871 26472
rect 5813 26463 5871 26469
rect 6546 26460 6552 26472
rect 6604 26460 6610 26512
rect 8294 26460 8300 26512
rect 8352 26460 8358 26512
rect 8754 26460 8760 26512
rect 8812 26500 8818 26512
rect 9600 26500 9628 26531
rect 9674 26528 9680 26580
rect 9732 26568 9738 26580
rect 10686 26568 10692 26580
rect 9732 26540 10692 26568
rect 9732 26528 9738 26540
rect 8812 26472 9628 26500
rect 8812 26460 8818 26472
rect 3418 26392 3424 26444
rect 3476 26392 3482 26444
rect 4614 26432 4620 26444
rect 3712 26404 4620 26432
rect 2363 26336 2774 26364
rect 2363 26333 2375 26336
rect 2317 26327 2375 26333
rect 3234 26324 3240 26376
rect 3292 26364 3298 26376
rect 3329 26367 3387 26373
rect 3329 26364 3341 26367
rect 3292 26336 3341 26364
rect 3292 26324 3298 26336
rect 3329 26333 3341 26336
rect 3375 26364 3387 26367
rect 3712 26364 3740 26404
rect 4614 26392 4620 26404
rect 4672 26432 4678 26444
rect 4672 26404 8248 26432
rect 4672 26392 4678 26404
rect 3375 26336 3740 26364
rect 3375 26333 3387 26336
rect 3329 26327 3387 26333
rect 3786 26324 3792 26376
rect 3844 26324 3850 26376
rect 8018 26373 8024 26376
rect 7837 26367 7895 26373
rect 6288 26336 7052 26364
rect 3510 26296 3516 26308
rect 3344 26268 3516 26296
rect 3237 26231 3295 26237
rect 3237 26197 3249 26231
rect 3283 26228 3295 26231
rect 3344 26228 3372 26268
rect 3510 26256 3516 26268
rect 3568 26256 3574 26308
rect 3970 26256 3976 26308
rect 4028 26296 4034 26308
rect 4065 26299 4123 26305
rect 4065 26296 4077 26299
rect 4028 26268 4077 26296
rect 4028 26256 4034 26268
rect 4065 26265 4077 26268
rect 4111 26265 4123 26299
rect 4065 26259 4123 26265
rect 4172 26268 4554 26296
rect 3283 26200 3372 26228
rect 3283 26197 3295 26200
rect 3237 26191 3295 26197
rect 3878 26188 3884 26240
rect 3936 26228 3942 26240
rect 4172 26228 4200 26268
rect 3936 26200 4200 26228
rect 4448 26228 4476 26268
rect 5810 26256 5816 26308
rect 5868 26296 5874 26308
rect 6288 26305 6316 26336
rect 7024 26308 7052 26336
rect 7837 26333 7849 26367
rect 7883 26333 7895 26367
rect 7837 26327 7895 26333
rect 7985 26367 8024 26373
rect 7985 26333 7997 26367
rect 7985 26327 8024 26333
rect 6089 26299 6147 26305
rect 6089 26296 6101 26299
rect 5868 26268 6101 26296
rect 5868 26256 5874 26268
rect 6089 26265 6101 26268
rect 6135 26265 6147 26299
rect 6089 26259 6147 26265
rect 6273 26299 6331 26305
rect 6273 26265 6285 26299
rect 6319 26265 6331 26299
rect 6273 26259 6331 26265
rect 6362 26256 6368 26308
rect 6420 26296 6426 26308
rect 6822 26296 6828 26308
rect 6420 26268 6828 26296
rect 6420 26256 6426 26268
rect 6822 26256 6828 26268
rect 6880 26256 6886 26308
rect 7006 26256 7012 26308
rect 7064 26256 7070 26308
rect 7852 26296 7880 26327
rect 8018 26324 8024 26327
rect 8076 26324 8082 26376
rect 8220 26373 8248 26404
rect 8864 26404 9260 26432
rect 8205 26367 8263 26373
rect 8205 26333 8217 26367
rect 8251 26333 8263 26367
rect 8205 26327 8263 26333
rect 8343 26367 8401 26373
rect 8343 26333 8355 26367
rect 8389 26364 8401 26367
rect 8570 26364 8576 26376
rect 8389 26336 8576 26364
rect 8389 26333 8401 26336
rect 8343 26327 8401 26333
rect 8570 26324 8576 26336
rect 8628 26324 8634 26376
rect 8113 26299 8171 26305
rect 7852 26268 8064 26296
rect 7098 26228 7104 26240
rect 4448 26200 7104 26228
rect 3936 26188 3942 26200
rect 7098 26188 7104 26200
rect 7156 26188 7162 26240
rect 8036 26228 8064 26268
rect 8113 26265 8125 26299
rect 8159 26296 8171 26299
rect 8864 26296 8892 26404
rect 8938 26324 8944 26376
rect 8996 26324 9002 26376
rect 9122 26373 9128 26376
rect 9089 26367 9128 26373
rect 9089 26333 9101 26367
rect 9089 26327 9128 26333
rect 9122 26324 9128 26327
rect 9180 26324 9186 26376
rect 9232 26364 9260 26404
rect 9447 26367 9505 26373
rect 9447 26364 9459 26367
rect 9232 26336 9459 26364
rect 9447 26333 9459 26336
rect 9493 26364 9505 26367
rect 9784 26364 9812 26540
rect 10686 26528 10692 26540
rect 10744 26528 10750 26580
rect 11330 26528 11336 26580
rect 11388 26568 11394 26580
rect 11388 26540 11652 26568
rect 11388 26528 11394 26540
rect 9493 26336 9812 26364
rect 9968 26472 11560 26500
rect 9493 26333 9505 26336
rect 9447 26327 9505 26333
rect 8159 26268 8892 26296
rect 9217 26299 9275 26305
rect 8159 26265 8171 26268
rect 8113 26259 8171 26265
rect 9217 26265 9229 26299
rect 9263 26265 9275 26299
rect 9217 26259 9275 26265
rect 9232 26228 9260 26259
rect 9306 26256 9312 26308
rect 9364 26256 9370 26308
rect 9968 26296 9996 26472
rect 10962 26432 10968 26444
rect 10520 26404 10968 26432
rect 10520 26373 10548 26404
rect 10962 26392 10968 26404
rect 11020 26392 11026 26444
rect 11532 26376 11560 26472
rect 10505 26367 10563 26373
rect 10505 26333 10517 26367
rect 10551 26333 10563 26367
rect 10505 26327 10563 26333
rect 10689 26367 10747 26373
rect 10689 26333 10701 26367
rect 10735 26364 10747 26367
rect 10735 26336 11009 26364
rect 10735 26333 10747 26336
rect 10689 26327 10747 26333
rect 9416 26268 9996 26296
rect 9416 26240 9444 26268
rect 10042 26256 10048 26308
rect 10100 26296 10106 26308
rect 10410 26296 10416 26308
rect 10100 26268 10416 26296
rect 10100 26256 10106 26268
rect 10410 26256 10416 26268
rect 10468 26256 10474 26308
rect 9398 26228 9404 26240
rect 8036 26200 9404 26228
rect 9398 26188 9404 26200
rect 9456 26188 9462 26240
rect 10686 26188 10692 26240
rect 10744 26188 10750 26240
rect 10981 26228 11009 26336
rect 11238 26324 11244 26376
rect 11296 26324 11302 26376
rect 11422 26373 11428 26376
rect 11389 26367 11428 26373
rect 11389 26333 11401 26367
rect 11389 26327 11428 26333
rect 11422 26324 11428 26327
rect 11480 26324 11486 26376
rect 11514 26324 11520 26376
rect 11572 26324 11578 26376
rect 11624 26373 11652 26540
rect 11882 26528 11888 26580
rect 11940 26528 11946 26580
rect 12434 26528 12440 26580
rect 12492 26528 12498 26580
rect 13541 26571 13599 26577
rect 13541 26537 13553 26571
rect 13587 26568 13599 26571
rect 13630 26568 13636 26580
rect 13587 26540 13636 26568
rect 13587 26537 13599 26540
rect 13541 26531 13599 26537
rect 13630 26528 13636 26540
rect 13688 26528 13694 26580
rect 14458 26528 14464 26580
rect 14516 26528 14522 26580
rect 16482 26528 16488 26580
rect 16540 26528 16546 26580
rect 16666 26528 16672 26580
rect 16724 26528 16730 26580
rect 16758 26528 16764 26580
rect 16816 26528 16822 26580
rect 18785 26571 18843 26577
rect 18785 26537 18797 26571
rect 18831 26568 18843 26571
rect 18874 26568 18880 26580
rect 18831 26540 18880 26568
rect 18831 26537 18843 26540
rect 18785 26531 18843 26537
rect 18874 26528 18880 26540
rect 18932 26528 18938 26580
rect 19334 26528 19340 26580
rect 19392 26528 19398 26580
rect 19426 26528 19432 26580
rect 19484 26568 19490 26580
rect 19484 26540 19932 26568
rect 19484 26528 19490 26540
rect 11790 26373 11796 26376
rect 11609 26367 11667 26373
rect 11609 26333 11621 26367
rect 11655 26333 11667 26367
rect 11609 26327 11667 26333
rect 11747 26367 11796 26373
rect 11747 26333 11759 26367
rect 11793 26333 11796 26367
rect 11747 26327 11796 26333
rect 11790 26324 11796 26327
rect 11848 26324 11854 26376
rect 11900 26364 11928 26528
rect 12452 26373 12480 26528
rect 12526 26460 12532 26512
rect 12584 26500 12590 26512
rect 14476 26500 14504 26528
rect 16500 26500 16528 26528
rect 12584 26472 14504 26500
rect 16408 26472 16528 26500
rect 12584 26460 12590 26472
rect 14274 26392 14280 26444
rect 14332 26392 14338 26444
rect 12069 26367 12127 26373
rect 12069 26364 12081 26367
rect 11900 26336 12081 26364
rect 12069 26333 12081 26336
rect 12115 26333 12127 26367
rect 12069 26327 12127 26333
rect 12253 26367 12311 26373
rect 12253 26333 12265 26367
rect 12299 26364 12311 26367
rect 12437 26367 12495 26373
rect 12299 26336 12408 26364
rect 12299 26333 12311 26336
rect 12253 26327 12311 26333
rect 12380 26240 12408 26336
rect 12437 26333 12449 26367
rect 12483 26333 12495 26367
rect 12437 26327 12495 26333
rect 12618 26324 12624 26376
rect 12676 26364 12682 26376
rect 12676 26336 12848 26364
rect 12676 26324 12682 26336
rect 12526 26256 12532 26308
rect 12584 26296 12590 26308
rect 12713 26299 12771 26305
rect 12713 26296 12725 26299
rect 12584 26268 12725 26296
rect 12584 26256 12590 26268
rect 12713 26265 12725 26268
rect 12759 26265 12771 26299
rect 12820 26296 12848 26336
rect 13262 26324 13268 26376
rect 13320 26324 13326 26376
rect 13357 26367 13415 26373
rect 13357 26333 13369 26367
rect 13403 26364 13415 26367
rect 13446 26364 13452 26376
rect 13403 26336 13452 26364
rect 13403 26333 13415 26336
rect 13357 26327 13415 26333
rect 13446 26324 13452 26336
rect 13504 26324 13510 26376
rect 13538 26324 13544 26376
rect 13596 26364 13602 26376
rect 13633 26367 13691 26373
rect 13633 26364 13645 26367
rect 13596 26336 13645 26364
rect 13596 26324 13602 26336
rect 13633 26333 13645 26336
rect 13679 26364 13691 26367
rect 14292 26364 14320 26392
rect 13679 26336 14320 26364
rect 16117 26367 16175 26373
rect 13679 26333 13691 26336
rect 13633 26327 13691 26333
rect 16117 26333 16129 26367
rect 16163 26364 16175 26367
rect 16206 26364 16212 26376
rect 16163 26336 16212 26364
rect 16163 26333 16175 26336
rect 16117 26327 16175 26333
rect 16206 26324 16212 26336
rect 16264 26324 16270 26376
rect 16408 26373 16436 26472
rect 16393 26367 16451 26373
rect 16393 26333 16405 26367
rect 16439 26333 16451 26367
rect 16393 26327 16451 26333
rect 16485 26367 16543 26373
rect 16485 26333 16497 26367
rect 16531 26364 16543 26367
rect 16776 26364 16804 26528
rect 17034 26460 17040 26512
rect 17092 26500 17098 26512
rect 18969 26503 19027 26509
rect 18969 26500 18981 26503
rect 17092 26472 18981 26500
rect 17092 26460 17098 26472
rect 18969 26469 18981 26472
rect 19015 26469 19027 26503
rect 18969 26463 19027 26469
rect 19150 26460 19156 26512
rect 19208 26500 19214 26512
rect 19610 26500 19616 26512
rect 19208 26472 19616 26500
rect 19208 26460 19214 26472
rect 19610 26460 19616 26472
rect 19668 26460 19674 26512
rect 19797 26503 19855 26509
rect 19797 26469 19809 26503
rect 19843 26469 19855 26503
rect 19904 26500 19932 26540
rect 20070 26528 20076 26580
rect 20128 26568 20134 26580
rect 20346 26568 20352 26580
rect 20128 26540 20352 26568
rect 20128 26528 20134 26540
rect 20346 26528 20352 26540
rect 20404 26528 20410 26580
rect 20622 26528 20628 26580
rect 20680 26568 20686 26580
rect 20717 26571 20775 26577
rect 20717 26568 20729 26571
rect 20680 26540 20729 26568
rect 20680 26528 20686 26540
rect 20717 26537 20729 26540
rect 20763 26537 20775 26571
rect 22649 26571 22707 26577
rect 22649 26568 22661 26571
rect 20717 26531 20775 26537
rect 21836 26540 22661 26568
rect 21545 26503 21603 26509
rect 21545 26500 21557 26503
rect 19904 26472 21557 26500
rect 19797 26463 19855 26469
rect 21545 26469 21557 26472
rect 21591 26469 21603 26503
rect 21545 26463 21603 26469
rect 19812 26432 19840 26463
rect 18248 26404 19840 26432
rect 17773 26367 17831 26373
rect 17773 26364 17785 26367
rect 16531 26336 16804 26364
rect 16868 26336 17785 26364
rect 16531 26333 16543 26336
rect 16485 26327 16543 26333
rect 13081 26299 13139 26305
rect 13081 26296 13093 26299
rect 12820 26268 13093 26296
rect 12713 26259 12771 26265
rect 13081 26265 13093 26268
rect 13127 26265 13139 26299
rect 13081 26259 13139 26265
rect 13906 26256 13912 26308
rect 13964 26256 13970 26308
rect 14642 26256 14648 26308
rect 14700 26296 14706 26308
rect 16301 26299 16359 26305
rect 16301 26296 16313 26299
rect 14700 26268 16313 26296
rect 14700 26256 14706 26268
rect 16301 26265 16313 26268
rect 16347 26296 16359 26299
rect 16868 26296 16896 26336
rect 17773 26333 17785 26336
rect 17819 26333 17831 26367
rect 17773 26327 17831 26333
rect 18138 26324 18144 26376
rect 18196 26364 18202 26376
rect 18248 26364 18276 26404
rect 20438 26392 20444 26444
rect 20496 26392 20502 26444
rect 20622 26392 20628 26444
rect 20680 26432 20686 26444
rect 20680 26404 20944 26432
rect 20680 26392 20686 26404
rect 18196 26336 18276 26364
rect 18196 26324 18202 26336
rect 18322 26324 18328 26376
rect 18380 26324 18386 26376
rect 18690 26364 18696 26376
rect 18524 26336 18696 26364
rect 16347 26268 16896 26296
rect 16347 26265 16359 26268
rect 16301 26259 16359 26265
rect 17586 26256 17592 26308
rect 17644 26296 17650 26308
rect 17681 26299 17739 26305
rect 17681 26296 17693 26299
rect 17644 26268 17693 26296
rect 17644 26256 17650 26268
rect 17681 26265 17693 26268
rect 17727 26296 17739 26299
rect 17727 26268 18184 26296
rect 17727 26265 17739 26268
rect 17681 26259 17739 26265
rect 12342 26228 12348 26240
rect 10981 26200 12348 26228
rect 12342 26188 12348 26200
rect 12400 26228 12408 26240
rect 13924 26228 13952 26256
rect 12400 26200 13952 26228
rect 12400 26188 12406 26200
rect 14918 26188 14924 26240
rect 14976 26228 14982 26240
rect 15194 26228 15200 26240
rect 14976 26200 15200 26228
rect 14976 26188 14982 26200
rect 15194 26188 15200 26200
rect 15252 26188 15258 26240
rect 18156 26228 18184 26268
rect 18230 26256 18236 26308
rect 18288 26256 18294 26308
rect 18524 26296 18552 26336
rect 18690 26324 18696 26336
rect 18748 26324 18754 26376
rect 18874 26324 18880 26376
rect 18932 26364 18938 26376
rect 19245 26367 19303 26373
rect 19245 26364 19257 26367
rect 18932 26336 19257 26364
rect 18932 26324 18938 26336
rect 19245 26333 19257 26336
rect 19291 26333 19303 26367
rect 19245 26327 19303 26333
rect 19426 26324 19432 26376
rect 19484 26364 19490 26376
rect 19613 26367 19671 26373
rect 19613 26364 19625 26367
rect 19484 26336 19625 26364
rect 19484 26324 19490 26336
rect 19613 26333 19625 26336
rect 19659 26364 19671 26367
rect 20456 26364 20484 26392
rect 20916 26373 20944 26404
rect 19659 26336 20484 26364
rect 20717 26367 20775 26373
rect 19659 26333 19671 26336
rect 19613 26327 19671 26333
rect 20717 26333 20729 26367
rect 20763 26333 20775 26367
rect 20717 26327 20775 26333
rect 20901 26367 20959 26373
rect 20901 26333 20913 26367
rect 20947 26364 20959 26367
rect 21542 26364 21548 26376
rect 20947 26336 21548 26364
rect 20947 26333 20959 26336
rect 20901 26327 20959 26333
rect 18340 26268 18552 26296
rect 18601 26299 18659 26305
rect 18340 26228 18368 26268
rect 18601 26265 18613 26299
rect 18647 26265 18659 26299
rect 18708 26296 18736 26324
rect 18785 26299 18843 26305
rect 18785 26296 18797 26299
rect 18708 26268 18797 26296
rect 18601 26259 18659 26265
rect 18785 26265 18797 26268
rect 18831 26265 18843 26299
rect 20732 26296 20760 26327
rect 21542 26324 21548 26336
rect 21600 26324 21606 26376
rect 21726 26324 21732 26376
rect 21784 26324 21790 26376
rect 21836 26373 21864 26540
rect 22649 26537 22661 26540
rect 22695 26568 22707 26571
rect 22738 26568 22744 26580
rect 22695 26540 22744 26568
rect 22695 26537 22707 26540
rect 22649 26531 22707 26537
rect 22738 26528 22744 26540
rect 22796 26528 22802 26580
rect 23658 26568 23664 26580
rect 23216 26540 23664 26568
rect 22094 26460 22100 26512
rect 22152 26460 22158 26512
rect 23216 26500 23244 26540
rect 23658 26528 23664 26540
rect 23716 26528 23722 26580
rect 23750 26528 23756 26580
rect 23808 26528 23814 26580
rect 23937 26571 23995 26577
rect 23937 26537 23949 26571
rect 23983 26568 23995 26571
rect 24026 26568 24032 26580
rect 23983 26540 24032 26568
rect 23983 26537 23995 26540
rect 23937 26531 23995 26537
rect 24026 26528 24032 26540
rect 24084 26568 24090 26580
rect 24394 26568 24400 26580
rect 24084 26540 24400 26568
rect 24084 26528 24090 26540
rect 24394 26528 24400 26540
rect 24452 26528 24458 26580
rect 24578 26528 24584 26580
rect 24636 26568 24642 26580
rect 25038 26568 25044 26580
rect 24636 26540 25044 26568
rect 24636 26528 24642 26540
rect 25038 26528 25044 26540
rect 25096 26528 25102 26580
rect 25314 26528 25320 26580
rect 25372 26528 25378 26580
rect 26418 26528 26424 26580
rect 26476 26568 26482 26580
rect 27798 26568 27804 26580
rect 26476 26540 27804 26568
rect 26476 26528 26482 26540
rect 27798 26528 27804 26540
rect 27856 26568 27862 26580
rect 28810 26568 28816 26580
rect 27856 26540 28816 26568
rect 27856 26528 27862 26540
rect 28810 26528 28816 26540
rect 28868 26528 28874 26580
rect 29362 26528 29368 26580
rect 29420 26568 29426 26580
rect 29549 26571 29607 26577
rect 29549 26568 29561 26571
rect 29420 26540 29561 26568
rect 29420 26528 29426 26540
rect 29549 26537 29561 26540
rect 29595 26537 29607 26571
rect 29549 26531 29607 26537
rect 30006 26528 30012 26580
rect 30064 26528 30070 26580
rect 31662 26528 31668 26580
rect 31720 26568 31726 26580
rect 31849 26571 31907 26577
rect 31849 26568 31861 26571
rect 31720 26540 31861 26568
rect 31720 26528 31726 26540
rect 31849 26537 31861 26540
rect 31895 26537 31907 26571
rect 31849 26531 31907 26537
rect 22572 26472 23244 26500
rect 23293 26503 23351 26509
rect 22112 26432 22140 26460
rect 22112 26404 22508 26432
rect 22112 26373 22140 26404
rect 21821 26367 21879 26373
rect 21821 26333 21833 26367
rect 21867 26333 21879 26367
rect 21821 26327 21879 26333
rect 22097 26367 22155 26373
rect 22097 26333 22109 26367
rect 22143 26333 22155 26367
rect 22097 26327 22155 26333
rect 22186 26324 22192 26376
rect 22244 26324 22250 26376
rect 21913 26299 21971 26305
rect 20732 26268 21864 26296
rect 18785 26259 18843 26265
rect 18156 26200 18368 26228
rect 18616 26228 18644 26259
rect 18874 26228 18880 26240
rect 18616 26200 18880 26228
rect 18874 26188 18880 26200
rect 18932 26228 18938 26240
rect 19058 26228 19064 26240
rect 18932 26200 19064 26228
rect 18932 26188 18938 26200
rect 19058 26188 19064 26200
rect 19116 26188 19122 26240
rect 20898 26188 20904 26240
rect 20956 26228 20962 26240
rect 21726 26228 21732 26240
rect 20956 26200 21732 26228
rect 20956 26188 20962 26200
rect 21726 26188 21732 26200
rect 21784 26188 21790 26240
rect 21836 26228 21864 26268
rect 21913 26265 21925 26299
rect 21959 26296 21971 26299
rect 22480 26296 22508 26404
rect 22572 26373 22600 26472
rect 23293 26469 23305 26503
rect 23339 26469 23351 26503
rect 23768 26500 23796 26528
rect 24121 26503 24179 26509
rect 24121 26500 24133 26503
rect 23768 26472 24133 26500
rect 23293 26463 23351 26469
rect 24121 26469 24133 26472
rect 24167 26469 24179 26503
rect 24121 26463 24179 26469
rect 23308 26432 23336 26463
rect 24210 26460 24216 26512
rect 24268 26500 24274 26512
rect 25501 26503 25559 26509
rect 25501 26500 25513 26503
rect 24268 26472 25513 26500
rect 24268 26460 24274 26472
rect 25501 26469 25513 26472
rect 25547 26469 25559 26503
rect 30193 26503 30251 26509
rect 30193 26500 30205 26503
rect 25501 26463 25559 26469
rect 29196 26472 30205 26500
rect 22664 26404 23336 26432
rect 22557 26367 22615 26373
rect 22557 26333 22569 26367
rect 22603 26333 22615 26367
rect 22557 26327 22615 26333
rect 22664 26296 22692 26404
rect 23382 26392 23388 26444
rect 23440 26432 23446 26444
rect 23845 26435 23903 26441
rect 23845 26432 23857 26435
rect 23440 26404 23857 26432
rect 23440 26392 23446 26404
rect 23845 26401 23857 26404
rect 23891 26432 23903 26435
rect 25777 26435 25835 26441
rect 23891 26404 25360 26432
rect 23891 26401 23903 26404
rect 23845 26395 23903 26401
rect 22738 26324 22744 26376
rect 22796 26324 22802 26376
rect 23569 26367 23627 26373
rect 23569 26333 23581 26367
rect 23615 26364 23627 26367
rect 23658 26364 23664 26376
rect 23615 26336 23664 26364
rect 23615 26333 23627 26336
rect 23569 26327 23627 26333
rect 23658 26324 23664 26336
rect 23716 26324 23722 26376
rect 23750 26324 23756 26376
rect 23808 26324 23814 26376
rect 24302 26324 24308 26376
rect 24360 26364 24366 26376
rect 24397 26367 24455 26373
rect 24397 26364 24409 26367
rect 24360 26336 24409 26364
rect 24360 26324 24366 26336
rect 24397 26333 24409 26336
rect 24443 26333 24455 26367
rect 24397 26327 24455 26333
rect 24762 26324 24768 26376
rect 24820 26324 24826 26376
rect 24857 26367 24915 26373
rect 24857 26333 24869 26367
rect 24903 26364 24915 26367
rect 24946 26364 24952 26376
rect 24903 26336 24952 26364
rect 24903 26333 24915 26336
rect 24857 26327 24915 26333
rect 24946 26324 24952 26336
rect 25004 26324 25010 26376
rect 25130 26324 25136 26376
rect 25188 26324 25194 26376
rect 25222 26324 25228 26376
rect 25280 26324 25286 26376
rect 25332 26364 25360 26404
rect 25777 26401 25789 26435
rect 25823 26432 25835 26435
rect 26142 26432 26148 26444
rect 25823 26404 26148 26432
rect 25823 26401 25835 26404
rect 25777 26395 25835 26401
rect 26142 26392 26148 26404
rect 26200 26392 26206 26444
rect 28902 26432 28908 26444
rect 26896 26404 28908 26432
rect 25961 26367 26019 26373
rect 25961 26364 25973 26367
rect 25332 26336 25973 26364
rect 25961 26333 25973 26336
rect 26007 26333 26019 26367
rect 25961 26327 26019 26333
rect 26326 26324 26332 26376
rect 26384 26324 26390 26376
rect 26694 26324 26700 26376
rect 26752 26364 26758 26376
rect 26896 26364 26924 26404
rect 28902 26392 28908 26404
rect 28960 26392 28966 26444
rect 26752 26336 26924 26364
rect 26752 26324 26758 26336
rect 26970 26324 26976 26376
rect 27028 26324 27034 26376
rect 27522 26324 27528 26376
rect 27580 26324 27586 26376
rect 27617 26367 27675 26373
rect 27617 26333 27629 26367
rect 27663 26333 27675 26367
rect 27617 26327 27675 26333
rect 21959 26268 22232 26296
rect 22480 26268 22692 26296
rect 23293 26299 23351 26305
rect 21959 26265 21971 26268
rect 21913 26259 21971 26265
rect 22094 26228 22100 26240
rect 21836 26200 22100 26228
rect 22094 26188 22100 26200
rect 22152 26188 22158 26240
rect 22204 26228 22232 26268
rect 23293 26265 23305 26299
rect 23339 26296 23351 26299
rect 25041 26299 25099 26305
rect 25041 26296 25053 26299
rect 23339 26268 25053 26296
rect 23339 26265 23351 26268
rect 23293 26259 23351 26265
rect 25041 26265 25053 26268
rect 25087 26265 25099 26299
rect 25041 26259 25099 26265
rect 22370 26228 22376 26240
rect 22204 26200 22376 26228
rect 22370 26188 22376 26200
rect 22428 26188 22434 26240
rect 23477 26231 23535 26237
rect 23477 26197 23489 26231
rect 23523 26228 23535 26231
rect 23934 26228 23940 26240
rect 23523 26200 23940 26228
rect 23523 26197 23535 26200
rect 23477 26191 23535 26197
rect 23934 26188 23940 26200
rect 23992 26228 23998 26240
rect 24578 26228 24584 26240
rect 23992 26200 24584 26228
rect 23992 26188 23998 26200
rect 24578 26188 24584 26200
rect 24636 26188 24642 26240
rect 24762 26188 24768 26240
rect 24820 26228 24826 26240
rect 25240 26228 25268 26324
rect 25590 26256 25596 26308
rect 25648 26296 25654 26308
rect 26513 26299 26571 26305
rect 26513 26296 26525 26299
rect 25648 26268 26525 26296
rect 25648 26256 25654 26268
rect 26513 26265 26525 26268
rect 26559 26265 26571 26299
rect 26988 26296 27016 26324
rect 27632 26296 27660 26327
rect 27798 26324 27804 26376
rect 27856 26324 27862 26376
rect 27893 26367 27951 26373
rect 27893 26333 27905 26367
rect 27939 26333 27951 26367
rect 27893 26327 27951 26333
rect 28997 26367 29055 26373
rect 28997 26333 29009 26367
rect 29043 26364 29055 26367
rect 29196 26364 29224 26472
rect 30193 26469 30205 26472
rect 30239 26469 30251 26503
rect 30193 26463 30251 26469
rect 30469 26503 30527 26509
rect 30469 26469 30481 26503
rect 30515 26500 30527 26503
rect 30742 26500 30748 26512
rect 30515 26472 30748 26500
rect 30515 26469 30527 26472
rect 30469 26463 30527 26469
rect 30742 26460 30748 26472
rect 30800 26460 30806 26512
rect 31864 26500 31892 26531
rect 32030 26528 32036 26580
rect 32088 26528 32094 26580
rect 33042 26528 33048 26580
rect 33100 26568 33106 26580
rect 33100 26540 34192 26568
rect 33100 26528 33106 26540
rect 31864 26472 33456 26500
rect 29270 26392 29276 26444
rect 29328 26392 29334 26444
rect 29638 26392 29644 26444
rect 29696 26392 29702 26444
rect 32122 26432 32128 26444
rect 30576 26404 32128 26432
rect 29043 26336 29224 26364
rect 29288 26364 29316 26392
rect 29825 26367 29883 26373
rect 29825 26364 29837 26367
rect 29288 26336 29837 26364
rect 29043 26333 29055 26336
rect 28997 26327 29055 26333
rect 29825 26333 29837 26336
rect 29871 26333 29883 26367
rect 29825 26327 29883 26333
rect 30377 26367 30435 26373
rect 30377 26333 30389 26367
rect 30423 26333 30435 26367
rect 30377 26327 30435 26333
rect 26988 26268 27660 26296
rect 26513 26259 26571 26265
rect 27632 26240 27660 26268
rect 27908 26240 27936 26327
rect 28626 26256 28632 26308
rect 28684 26296 28690 26308
rect 29181 26299 29239 26305
rect 29181 26296 29193 26299
rect 28684 26268 29193 26296
rect 28684 26256 28690 26268
rect 29181 26265 29193 26268
rect 29227 26265 29239 26299
rect 29181 26259 29239 26265
rect 29362 26256 29368 26308
rect 29420 26296 29426 26308
rect 29549 26299 29607 26305
rect 29549 26296 29561 26299
rect 29420 26268 29561 26296
rect 29420 26256 29426 26268
rect 29549 26265 29561 26268
rect 29595 26265 29607 26299
rect 29549 26259 29607 26265
rect 30392 26296 30420 26327
rect 30466 26324 30472 26376
rect 30524 26364 30530 26376
rect 30576 26373 30604 26404
rect 32122 26392 32128 26404
rect 32180 26392 32186 26444
rect 30561 26367 30619 26373
rect 30561 26364 30573 26367
rect 30524 26336 30573 26364
rect 30524 26324 30530 26336
rect 30561 26333 30573 26336
rect 30607 26333 30619 26367
rect 30561 26327 30619 26333
rect 30653 26367 30711 26373
rect 30653 26333 30665 26367
rect 30699 26364 30711 26367
rect 30834 26364 30840 26376
rect 30699 26336 30840 26364
rect 30699 26333 30711 26336
rect 30653 26327 30711 26333
rect 30834 26324 30840 26336
rect 30892 26324 30898 26376
rect 31018 26324 31024 26376
rect 31076 26324 31082 26376
rect 32030 26364 32036 26376
rect 31880 26336 32036 26364
rect 31036 26296 31064 26324
rect 31880 26305 31908 26336
rect 32030 26324 32036 26336
rect 32088 26364 32094 26376
rect 32217 26367 32275 26373
rect 32217 26364 32229 26367
rect 32088 26336 32229 26364
rect 32088 26324 32094 26336
rect 32217 26333 32229 26336
rect 32263 26364 32275 26367
rect 32582 26364 32588 26376
rect 32263 26336 32588 26364
rect 32263 26333 32275 26336
rect 32217 26327 32275 26333
rect 32582 26324 32588 26336
rect 32640 26324 32646 26376
rect 32692 26373 32720 26472
rect 33428 26432 33456 26472
rect 33502 26460 33508 26512
rect 33560 26460 33566 26512
rect 33428 26404 33548 26432
rect 33520 26376 33548 26404
rect 32677 26367 32735 26373
rect 32677 26333 32689 26367
rect 32723 26333 32735 26367
rect 32677 26327 32735 26333
rect 32766 26324 32772 26376
rect 32824 26364 32830 26376
rect 32861 26367 32919 26373
rect 32861 26364 32873 26367
rect 32824 26336 32873 26364
rect 32824 26324 32830 26336
rect 32861 26333 32873 26336
rect 32907 26333 32919 26367
rect 32861 26327 32919 26333
rect 33226 26324 33232 26376
rect 33284 26324 33290 26376
rect 33502 26324 33508 26376
rect 33560 26324 33566 26376
rect 33965 26367 34023 26373
rect 33965 26333 33977 26367
rect 34011 26364 34023 26367
rect 34054 26364 34060 26376
rect 34011 26336 34060 26364
rect 34011 26333 34023 26336
rect 33965 26327 34023 26333
rect 34054 26324 34060 26336
rect 34112 26324 34118 26376
rect 34164 26373 34192 26540
rect 37366 26528 37372 26580
rect 37424 26568 37430 26580
rect 37550 26568 37556 26580
rect 37424 26540 37556 26568
rect 37424 26528 37430 26540
rect 37550 26528 37556 26540
rect 37608 26528 37614 26580
rect 38286 26528 38292 26580
rect 38344 26568 38350 26580
rect 38933 26571 38991 26577
rect 38933 26568 38945 26571
rect 38344 26540 38945 26568
rect 38344 26528 38350 26540
rect 38933 26537 38945 26540
rect 38979 26537 38991 26571
rect 38933 26531 38991 26537
rect 35897 26503 35955 26509
rect 35897 26469 35909 26503
rect 35943 26500 35955 26503
rect 36538 26500 36544 26512
rect 35943 26472 36544 26500
rect 35943 26469 35955 26472
rect 35897 26463 35955 26469
rect 36538 26460 36544 26472
rect 36596 26460 36602 26512
rect 34238 26392 34244 26444
rect 34296 26432 34302 26444
rect 34296 26404 36400 26432
rect 34296 26392 34302 26404
rect 35912 26373 35940 26404
rect 34149 26367 34207 26373
rect 34149 26333 34161 26367
rect 34195 26333 34207 26367
rect 34149 26327 34207 26333
rect 35897 26367 35955 26373
rect 35897 26333 35909 26367
rect 35943 26333 35955 26367
rect 35897 26327 35955 26333
rect 35986 26324 35992 26376
rect 36044 26324 36050 26376
rect 36078 26324 36084 26376
rect 36136 26324 36142 26376
rect 36372 26373 36400 26404
rect 36173 26367 36231 26373
rect 36173 26333 36185 26367
rect 36219 26333 36231 26367
rect 36173 26327 36231 26333
rect 36357 26367 36415 26373
rect 36357 26333 36369 26367
rect 36403 26333 36415 26367
rect 36357 26327 36415 26333
rect 38841 26367 38899 26373
rect 38841 26333 38853 26367
rect 38887 26364 38899 26367
rect 39669 26367 39727 26373
rect 39669 26364 39681 26367
rect 38887 26336 39681 26364
rect 38887 26333 38899 26336
rect 38841 26327 38899 26333
rect 39669 26333 39681 26336
rect 39715 26333 39727 26367
rect 39669 26327 39727 26333
rect 30392 26268 31064 26296
rect 31665 26299 31723 26305
rect 24820 26200 25268 26228
rect 24820 26188 24826 26200
rect 25958 26188 25964 26240
rect 26016 26188 26022 26240
rect 26881 26231 26939 26237
rect 26881 26197 26893 26231
rect 26927 26228 26939 26231
rect 27062 26228 27068 26240
rect 26927 26200 27068 26228
rect 26927 26197 26939 26200
rect 26881 26191 26939 26197
rect 27062 26188 27068 26200
rect 27120 26188 27126 26240
rect 27338 26188 27344 26240
rect 27396 26188 27402 26240
rect 27614 26188 27620 26240
rect 27672 26188 27678 26240
rect 27890 26188 27896 26240
rect 27948 26188 27954 26240
rect 27982 26188 27988 26240
rect 28040 26228 28046 26240
rect 28442 26228 28448 26240
rect 28040 26200 28448 26228
rect 28040 26188 28046 26200
rect 28442 26188 28448 26200
rect 28500 26188 28506 26240
rect 29270 26188 29276 26240
rect 29328 26228 29334 26240
rect 30392 26228 30420 26268
rect 31665 26265 31677 26299
rect 31711 26265 31723 26299
rect 31665 26259 31723 26265
rect 31865 26299 31923 26305
rect 31865 26265 31877 26299
rect 31911 26265 31923 26299
rect 32784 26296 32812 26324
rect 36004 26296 36032 26324
rect 36188 26296 36216 26327
rect 37090 26296 37096 26308
rect 31865 26259 31923 26265
rect 31956 26268 32812 26296
rect 32876 26268 33916 26296
rect 36004 26268 37096 26296
rect 29328 26200 30420 26228
rect 31680 26228 31708 26259
rect 31754 26228 31760 26240
rect 31680 26200 31760 26228
rect 29328 26188 29334 26200
rect 31754 26188 31760 26200
rect 31812 26228 31818 26240
rect 31956 26228 31984 26268
rect 31812 26200 31984 26228
rect 31812 26188 31818 26200
rect 32122 26188 32128 26240
rect 32180 26228 32186 26240
rect 32876 26228 32904 26268
rect 32180 26200 32904 26228
rect 32180 26188 32186 26200
rect 33686 26188 33692 26240
rect 33744 26228 33750 26240
rect 33781 26231 33839 26237
rect 33781 26228 33793 26231
rect 33744 26200 33793 26228
rect 33744 26188 33750 26200
rect 33781 26197 33793 26200
rect 33827 26197 33839 26231
rect 33888 26228 33916 26268
rect 37090 26256 37096 26268
rect 37148 26256 37154 26308
rect 39301 26299 39359 26305
rect 39301 26265 39313 26299
rect 39347 26265 39359 26299
rect 39301 26259 39359 26265
rect 39485 26299 39543 26305
rect 39485 26265 39497 26299
rect 39531 26296 39543 26299
rect 39758 26296 39764 26308
rect 39531 26268 39764 26296
rect 39531 26265 39543 26268
rect 39485 26259 39543 26265
rect 36265 26231 36323 26237
rect 36265 26228 36277 26231
rect 33888 26200 36277 26228
rect 33781 26191 33839 26197
rect 36265 26197 36277 26200
rect 36311 26197 36323 26231
rect 36265 26191 36323 26197
rect 39206 26188 39212 26240
rect 39264 26228 39270 26240
rect 39316 26228 39344 26259
rect 39758 26256 39764 26268
rect 39816 26256 39822 26308
rect 39942 26256 39948 26308
rect 40000 26256 40006 26308
rect 40678 26256 40684 26308
rect 40736 26256 40742 26308
rect 39960 26228 39988 26256
rect 39264 26200 39988 26228
rect 39264 26188 39270 26200
rect 40494 26188 40500 26240
rect 40552 26228 40558 26240
rect 40773 26231 40831 26237
rect 40773 26228 40785 26231
rect 40552 26200 40785 26228
rect 40552 26188 40558 26200
rect 40773 26197 40785 26200
rect 40819 26197 40831 26231
rect 40773 26191 40831 26197
rect 1104 26138 41400 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 41400 26138
rect 1104 26064 41400 26086
rect 4617 26027 4675 26033
rect 4617 25993 4629 26027
rect 4663 26024 4675 26027
rect 5534 26024 5540 26036
rect 4663 25996 5540 26024
rect 4663 25993 4675 25996
rect 4617 25987 4675 25993
rect 5534 25984 5540 25996
rect 5592 25984 5598 26036
rect 8389 26027 8447 26033
rect 8389 25993 8401 26027
rect 8435 26024 8447 26027
rect 8938 26024 8944 26036
rect 8435 25996 8944 26024
rect 8435 25993 8447 25996
rect 8389 25987 8447 25993
rect 8938 25984 8944 25996
rect 8996 25984 9002 26036
rect 10965 26027 11023 26033
rect 10965 25993 10977 26027
rect 11011 26024 11023 26027
rect 11238 26024 11244 26036
rect 11011 25996 11244 26024
rect 11011 25993 11023 25996
rect 10965 25987 11023 25993
rect 11238 25984 11244 25996
rect 11296 25984 11302 26036
rect 11514 25984 11520 26036
rect 11572 26024 11578 26036
rect 12802 26024 12808 26036
rect 11572 25996 12808 26024
rect 11572 25984 11578 25996
rect 12802 25984 12808 25996
rect 12860 25984 12866 26036
rect 20438 26024 20444 26036
rect 20272 25996 20444 26024
rect 20272 25968 20300 25996
rect 20438 25984 20444 25996
rect 20496 26024 20502 26036
rect 21361 26027 21419 26033
rect 20496 25996 21312 26024
rect 20496 25984 20502 25996
rect 2406 25916 2412 25968
rect 2464 25956 2470 25968
rect 3786 25956 3792 25968
rect 2464 25928 3792 25956
rect 2464 25916 2470 25928
rect 3786 25916 3792 25928
rect 3844 25956 3850 25968
rect 3844 25928 6408 25956
rect 3844 25916 3850 25928
rect 2958 25848 2964 25900
rect 3016 25848 3022 25900
rect 4525 25891 4583 25897
rect 4525 25857 4537 25891
rect 4571 25888 4583 25891
rect 5442 25888 5448 25900
rect 4571 25860 5448 25888
rect 4571 25857 4583 25860
rect 4525 25851 4583 25857
rect 5442 25848 5448 25860
rect 5500 25848 5506 25900
rect 6380 25832 6408 25928
rect 9306 25916 9312 25968
rect 9364 25956 9370 25968
rect 9582 25956 9588 25968
rect 9364 25928 9588 25956
rect 9364 25916 9370 25928
rect 9582 25916 9588 25928
rect 9640 25916 9646 25968
rect 10689 25959 10747 25965
rect 10689 25925 10701 25959
rect 10735 25956 10747 25959
rect 10735 25928 11652 25956
rect 10735 25925 10747 25928
rect 10689 25919 10747 25925
rect 11624 25900 11652 25928
rect 13170 25916 13176 25968
rect 13228 25956 13234 25968
rect 14090 25956 14096 25968
rect 13228 25928 14096 25956
rect 13228 25916 13234 25928
rect 14090 25916 14096 25928
rect 14148 25916 14154 25968
rect 18230 25916 18236 25968
rect 18288 25956 18294 25968
rect 18785 25959 18843 25965
rect 18785 25956 18797 25959
rect 18288 25928 18797 25956
rect 18288 25916 18294 25928
rect 18785 25925 18797 25928
rect 18831 25956 18843 25959
rect 19150 25956 19156 25968
rect 18831 25928 19156 25956
rect 18831 25925 18843 25928
rect 18785 25919 18843 25925
rect 19150 25916 19156 25928
rect 19208 25956 19214 25968
rect 19337 25959 19395 25965
rect 19337 25956 19349 25959
rect 19208 25928 19349 25956
rect 19208 25916 19214 25928
rect 19337 25925 19349 25928
rect 19383 25925 19395 25959
rect 19337 25919 19395 25925
rect 20254 25916 20260 25968
rect 20312 25916 20318 25968
rect 20732 25928 21220 25956
rect 6914 25848 6920 25900
rect 6972 25888 6978 25900
rect 7837 25891 7895 25897
rect 7837 25888 7849 25891
rect 6972 25860 7849 25888
rect 6972 25848 6978 25860
rect 7837 25857 7849 25860
rect 7883 25857 7895 25891
rect 7837 25851 7895 25857
rect 8021 25891 8079 25897
rect 8021 25857 8033 25891
rect 8067 25857 8079 25891
rect 8021 25851 8079 25857
rect 4801 25823 4859 25829
rect 4801 25789 4813 25823
rect 4847 25789 4859 25823
rect 4801 25783 4859 25789
rect 3418 25712 3424 25764
rect 3476 25752 3482 25764
rect 3878 25752 3884 25764
rect 3476 25724 3884 25752
rect 3476 25712 3482 25724
rect 3878 25712 3884 25724
rect 3936 25752 3942 25764
rect 4816 25752 4844 25783
rect 6362 25780 6368 25832
rect 6420 25780 6426 25832
rect 7098 25780 7104 25832
rect 7156 25820 7162 25832
rect 7558 25820 7564 25832
rect 7156 25792 7564 25820
rect 7156 25780 7162 25792
rect 7558 25780 7564 25792
rect 7616 25780 7622 25832
rect 8036 25820 8064 25851
rect 8110 25848 8116 25900
rect 8168 25848 8174 25900
rect 8205 25891 8263 25897
rect 8205 25857 8217 25891
rect 8251 25888 8263 25891
rect 9030 25888 9036 25900
rect 8251 25860 9036 25888
rect 8251 25857 8263 25860
rect 8205 25851 8263 25857
rect 9030 25848 9036 25860
rect 9088 25848 9094 25900
rect 10410 25848 10416 25900
rect 10468 25848 10474 25900
rect 10597 25891 10655 25897
rect 10597 25857 10609 25891
rect 10643 25857 10655 25891
rect 10597 25851 10655 25857
rect 8570 25820 8576 25832
rect 8036 25792 8576 25820
rect 8570 25780 8576 25792
rect 8628 25820 8634 25832
rect 9582 25820 9588 25832
rect 8628 25792 9588 25820
rect 8628 25780 8634 25792
rect 9582 25780 9588 25792
rect 9640 25820 9646 25832
rect 10612 25820 10640 25851
rect 10778 25848 10784 25900
rect 10836 25848 10842 25900
rect 11606 25848 11612 25900
rect 11664 25848 11670 25900
rect 13630 25848 13636 25900
rect 13688 25848 13694 25900
rect 15194 25848 15200 25900
rect 15252 25848 15258 25900
rect 16942 25848 16948 25900
rect 17000 25848 17006 25900
rect 17405 25891 17463 25897
rect 17405 25857 17417 25891
rect 17451 25888 17463 25891
rect 17586 25888 17592 25900
rect 17451 25860 17592 25888
rect 17451 25857 17463 25860
rect 17405 25851 17463 25857
rect 17586 25848 17592 25860
rect 17644 25848 17650 25900
rect 19245 25891 19303 25897
rect 19245 25857 19257 25891
rect 19291 25857 19303 25891
rect 19245 25851 19303 25857
rect 13648 25820 13676 25848
rect 9640 25792 13676 25820
rect 19260 25820 19288 25851
rect 19426 25848 19432 25900
rect 19484 25848 19490 25900
rect 20070 25848 20076 25900
rect 20128 25848 20134 25900
rect 19334 25820 19340 25832
rect 19260 25792 19340 25820
rect 9640 25780 9646 25792
rect 19334 25780 19340 25792
rect 19392 25820 19398 25832
rect 20088 25820 20116 25848
rect 19392 25792 20116 25820
rect 19392 25780 19398 25792
rect 3936 25724 7236 25752
rect 3936 25712 3942 25724
rect 7208 25696 7236 25724
rect 9214 25712 9220 25764
rect 9272 25752 9278 25764
rect 9272 25724 11836 25752
rect 9272 25712 9278 25724
rect 11808 25696 11836 25724
rect 20732 25696 20760 25928
rect 20809 25891 20867 25897
rect 20809 25857 20821 25891
rect 20855 25888 20867 25891
rect 20898 25888 20904 25900
rect 20855 25860 20904 25888
rect 20855 25857 20867 25860
rect 20809 25851 20867 25857
rect 20898 25848 20904 25860
rect 20956 25848 20962 25900
rect 21192 25897 21220 25928
rect 20993 25891 21051 25897
rect 20993 25857 21005 25891
rect 21039 25857 21051 25891
rect 20993 25851 21051 25857
rect 21085 25891 21143 25897
rect 21085 25857 21097 25891
rect 21131 25857 21143 25891
rect 21085 25851 21143 25857
rect 21177 25891 21235 25897
rect 21177 25857 21189 25891
rect 21223 25857 21235 25891
rect 21284 25888 21312 25996
rect 21361 25993 21373 26027
rect 21407 26024 21419 26027
rect 22002 26024 22008 26036
rect 21407 25996 22008 26024
rect 21407 25993 21419 25996
rect 21361 25987 21419 25993
rect 22002 25984 22008 25996
rect 22060 25984 22066 26036
rect 22094 25984 22100 26036
rect 22152 26024 22158 26036
rect 23566 26024 23572 26036
rect 22152 25996 23572 26024
rect 22152 25984 22158 25996
rect 23566 25984 23572 25996
rect 23624 25984 23630 26036
rect 23750 25984 23756 26036
rect 23808 26024 23814 26036
rect 25041 26027 25099 26033
rect 25041 26024 25053 26027
rect 23808 25996 25053 26024
rect 23808 25984 23814 25996
rect 25041 25993 25053 25996
rect 25087 25993 25099 26027
rect 25041 25987 25099 25993
rect 25148 25996 26280 26024
rect 22278 25916 22284 25968
rect 22336 25916 22342 25968
rect 21361 25891 21419 25897
rect 21361 25888 21373 25891
rect 21284 25860 21373 25888
rect 21177 25851 21235 25857
rect 21361 25857 21373 25860
rect 21407 25857 21419 25891
rect 21361 25851 21419 25857
rect 21008 25752 21036 25851
rect 21100 25820 21128 25851
rect 22002 25820 22008 25832
rect 21100 25792 22008 25820
rect 22002 25780 22008 25792
rect 22060 25820 22066 25832
rect 22296 25820 22324 25916
rect 22060 25792 22324 25820
rect 25148 25820 25176 25996
rect 25240 25928 26096 25956
rect 25240 25897 25268 25928
rect 26068 25900 26096 25928
rect 26252 25900 26280 25996
rect 27430 25984 27436 26036
rect 27488 26024 27494 26036
rect 28077 26027 28135 26033
rect 28077 26024 28089 26027
rect 27488 25996 28089 26024
rect 27488 25984 27494 25996
rect 28077 25993 28089 25996
rect 28123 25993 28135 26027
rect 28077 25987 28135 25993
rect 28626 25984 28632 26036
rect 28684 25984 28690 26036
rect 28718 25984 28724 26036
rect 28776 26024 28782 26036
rect 28776 25996 28994 26024
rect 28776 25984 28782 25996
rect 26602 25916 26608 25968
rect 26660 25956 26666 25968
rect 27246 25956 27252 25968
rect 26660 25928 27252 25956
rect 26660 25916 26666 25928
rect 25225 25891 25283 25897
rect 25225 25857 25237 25891
rect 25271 25857 25283 25891
rect 25225 25851 25283 25857
rect 25317 25891 25375 25897
rect 25317 25857 25329 25891
rect 25363 25857 25375 25891
rect 25317 25851 25375 25857
rect 25332 25820 25360 25851
rect 25406 25848 25412 25900
rect 25464 25848 25470 25900
rect 25547 25891 25605 25897
rect 25547 25857 25559 25891
rect 25593 25888 25605 25891
rect 25958 25888 25964 25900
rect 25593 25860 25964 25888
rect 25593 25857 25605 25860
rect 25547 25851 25605 25857
rect 25958 25848 25964 25860
rect 26016 25848 26022 25900
rect 26050 25848 26056 25900
rect 26108 25848 26114 25900
rect 26234 25848 26240 25900
rect 26292 25848 26298 25900
rect 26329 25891 26387 25897
rect 26329 25857 26341 25891
rect 26375 25888 26387 25891
rect 26878 25888 26884 25900
rect 26375 25860 26884 25888
rect 26375 25857 26387 25860
rect 26329 25851 26387 25857
rect 26878 25848 26884 25860
rect 26936 25848 26942 25900
rect 26988 25897 27016 25928
rect 27246 25916 27252 25928
rect 27304 25916 27310 25968
rect 28644 25956 28672 25984
rect 27908 25928 28672 25956
rect 28966 25956 28994 25996
rect 32030 25984 32036 26036
rect 32088 26024 32094 26036
rect 34238 26024 34244 26036
rect 32088 25996 34244 26024
rect 32088 25984 32094 25996
rect 34238 25984 34244 25996
rect 34296 25984 34302 26036
rect 34330 25984 34336 26036
rect 34388 25984 34394 26036
rect 35526 26024 35532 26036
rect 35268 25996 35532 26024
rect 34348 25956 34376 25984
rect 28966 25928 34376 25956
rect 26973 25891 27031 25897
rect 26973 25857 26985 25891
rect 27019 25857 27031 25891
rect 26973 25851 27031 25857
rect 27062 25848 27068 25900
rect 27120 25888 27126 25900
rect 27157 25891 27215 25897
rect 27157 25888 27169 25891
rect 27120 25860 27169 25888
rect 27120 25848 27126 25860
rect 27157 25857 27169 25860
rect 27203 25857 27215 25891
rect 27157 25851 27215 25857
rect 27338 25848 27344 25900
rect 27396 25888 27402 25900
rect 27908 25897 27936 25928
rect 35066 25916 35072 25968
rect 35124 25956 35130 25968
rect 35268 25965 35296 25996
rect 35526 25984 35532 25996
rect 35584 25984 35590 26036
rect 37458 25984 37464 26036
rect 37516 25984 37522 26036
rect 37553 26027 37611 26033
rect 37553 25993 37565 26027
rect 37599 26024 37611 26027
rect 37734 26024 37740 26036
rect 37599 25996 37740 26024
rect 37599 25993 37611 25996
rect 37553 25987 37611 25993
rect 37734 25984 37740 25996
rect 37792 25984 37798 26036
rect 39758 25984 39764 26036
rect 39816 26024 39822 26036
rect 41049 26027 41107 26033
rect 41049 26024 41061 26027
rect 39816 25996 41061 26024
rect 39816 25984 39822 25996
rect 41049 25993 41061 25996
rect 41095 25993 41107 26027
rect 41049 25987 41107 25993
rect 35253 25959 35311 25965
rect 35253 25956 35265 25959
rect 35124 25928 35265 25956
rect 35124 25916 35130 25928
rect 35253 25925 35265 25928
rect 35299 25925 35311 25959
rect 37476 25956 37504 25984
rect 38565 25959 38623 25965
rect 37476 25928 37780 25956
rect 35253 25919 35311 25925
rect 27709 25891 27767 25897
rect 27709 25888 27721 25891
rect 27396 25860 27721 25888
rect 27396 25848 27402 25860
rect 27709 25857 27721 25860
rect 27755 25857 27767 25891
rect 27709 25851 27767 25857
rect 27893 25891 27951 25897
rect 27893 25857 27905 25891
rect 27939 25857 27951 25891
rect 27893 25851 27951 25857
rect 28169 25891 28227 25897
rect 28169 25857 28181 25891
rect 28215 25888 28227 25891
rect 28215 25860 28396 25888
rect 28215 25857 28227 25860
rect 28169 25851 28227 25857
rect 25148 25792 25360 25820
rect 25685 25823 25743 25829
rect 22060 25780 22066 25792
rect 25685 25789 25697 25823
rect 25731 25820 25743 25823
rect 25866 25820 25872 25832
rect 25731 25792 25872 25820
rect 25731 25789 25743 25792
rect 25685 25783 25743 25789
rect 23014 25752 23020 25764
rect 21008 25724 23020 25752
rect 21008 25696 21036 25724
rect 23014 25712 23020 25724
rect 23072 25712 23078 25764
rect 24946 25712 24952 25764
rect 25004 25752 25010 25764
rect 25700 25752 25728 25783
rect 25866 25780 25872 25792
rect 25924 25780 25930 25832
rect 25976 25792 27384 25820
rect 25004 25724 25728 25752
rect 25004 25712 25010 25724
rect 4062 25644 4068 25696
rect 4120 25684 4126 25696
rect 4157 25687 4215 25693
rect 4157 25684 4169 25687
rect 4120 25656 4169 25684
rect 4120 25644 4126 25656
rect 4157 25653 4169 25656
rect 4203 25653 4215 25687
rect 4157 25647 4215 25653
rect 7190 25644 7196 25696
rect 7248 25684 7254 25696
rect 9858 25684 9864 25696
rect 7248 25656 9864 25684
rect 7248 25644 7254 25656
rect 9858 25644 9864 25656
rect 9916 25644 9922 25696
rect 11790 25644 11796 25696
rect 11848 25644 11854 25696
rect 15010 25644 15016 25696
rect 15068 25644 15074 25696
rect 15746 25644 15752 25696
rect 15804 25684 15810 25696
rect 16761 25687 16819 25693
rect 16761 25684 16773 25687
rect 15804 25656 16773 25684
rect 15804 25644 15810 25656
rect 16761 25653 16773 25656
rect 16807 25653 16819 25687
rect 16761 25647 16819 25653
rect 18874 25644 18880 25696
rect 18932 25684 18938 25696
rect 19061 25687 19119 25693
rect 19061 25684 19073 25687
rect 18932 25656 19073 25684
rect 18932 25644 18938 25656
rect 19061 25653 19073 25656
rect 19107 25684 19119 25687
rect 19334 25684 19340 25696
rect 19107 25656 19340 25684
rect 19107 25653 19119 25656
rect 19061 25647 19119 25653
rect 19334 25644 19340 25656
rect 19392 25644 19398 25696
rect 20625 25687 20683 25693
rect 20625 25653 20637 25687
rect 20671 25684 20683 25687
rect 20714 25684 20720 25696
rect 20671 25656 20720 25684
rect 20671 25653 20683 25656
rect 20625 25647 20683 25653
rect 20714 25644 20720 25656
rect 20772 25644 20778 25696
rect 20990 25644 20996 25696
rect 21048 25644 21054 25696
rect 21542 25644 21548 25696
rect 21600 25684 21606 25696
rect 25976 25684 26004 25792
rect 26050 25712 26056 25764
rect 26108 25752 26114 25764
rect 27249 25755 27307 25761
rect 27249 25752 27261 25755
rect 26108 25724 27261 25752
rect 26108 25712 26114 25724
rect 27249 25721 27261 25724
rect 27295 25721 27307 25755
rect 27356 25752 27384 25792
rect 27614 25780 27620 25832
rect 27672 25820 27678 25832
rect 28261 25823 28319 25829
rect 28261 25820 28273 25823
rect 27672 25792 28273 25820
rect 27672 25780 27678 25792
rect 28261 25789 28273 25792
rect 28307 25789 28319 25823
rect 28368 25820 28396 25860
rect 28442 25848 28448 25900
rect 28500 25848 28506 25900
rect 29362 25848 29368 25900
rect 29420 25848 29426 25900
rect 29914 25848 29920 25900
rect 29972 25848 29978 25900
rect 30190 25848 30196 25900
rect 30248 25848 30254 25900
rect 30558 25888 30564 25900
rect 30300 25860 30564 25888
rect 30300 25820 30328 25860
rect 30558 25848 30564 25860
rect 30616 25848 30622 25900
rect 30745 25891 30803 25897
rect 30745 25857 30757 25891
rect 30791 25888 30803 25891
rect 31110 25888 31116 25900
rect 30791 25860 31116 25888
rect 30791 25857 30803 25860
rect 30745 25851 30803 25857
rect 31110 25848 31116 25860
rect 31168 25848 31174 25900
rect 32030 25848 32036 25900
rect 32088 25888 32094 25900
rect 33410 25888 33416 25900
rect 32088 25860 33416 25888
rect 32088 25848 32094 25860
rect 33410 25848 33416 25860
rect 33468 25848 33474 25900
rect 35437 25891 35495 25897
rect 35437 25857 35449 25891
rect 35483 25857 35495 25891
rect 35437 25851 35495 25857
rect 35529 25891 35587 25897
rect 35529 25857 35541 25891
rect 35575 25857 35587 25891
rect 35529 25851 35587 25857
rect 28368 25792 30328 25820
rect 28261 25783 28319 25789
rect 30374 25780 30380 25832
rect 30432 25780 30438 25832
rect 33226 25780 33232 25832
rect 33284 25820 33290 25832
rect 34790 25820 34796 25832
rect 33284 25792 34796 25820
rect 33284 25780 33290 25792
rect 34790 25780 34796 25792
rect 34848 25780 34854 25832
rect 35342 25780 35348 25832
rect 35400 25820 35406 25832
rect 35452 25820 35480 25851
rect 35400 25792 35480 25820
rect 35400 25780 35406 25792
rect 34885 25755 34943 25761
rect 34885 25752 34897 25755
rect 27356 25724 34897 25752
rect 27249 25715 27307 25721
rect 34808 25696 34836 25724
rect 34885 25721 34897 25724
rect 34931 25752 34943 25755
rect 35544 25752 35572 25851
rect 35802 25848 35808 25900
rect 35860 25888 35866 25900
rect 37277 25891 37335 25897
rect 37277 25888 37289 25891
rect 35860 25860 37289 25888
rect 35860 25848 35866 25860
rect 37277 25857 37289 25860
rect 37323 25888 37335 25891
rect 37458 25888 37464 25900
rect 37323 25860 37464 25888
rect 37323 25857 37335 25860
rect 37277 25851 37335 25857
rect 37458 25848 37464 25860
rect 37516 25848 37522 25900
rect 37752 25897 37780 25928
rect 38565 25925 38577 25959
rect 38611 25956 38623 25959
rect 39206 25956 39212 25968
rect 38611 25928 39212 25956
rect 38611 25925 38623 25928
rect 38565 25919 38623 25925
rect 39206 25916 39212 25928
rect 39264 25916 39270 25968
rect 40034 25916 40040 25968
rect 40092 25916 40098 25968
rect 37737 25891 37795 25897
rect 37737 25857 37749 25891
rect 37783 25888 37795 25891
rect 37826 25888 37832 25900
rect 37783 25860 37832 25888
rect 37783 25857 37795 25860
rect 37737 25851 37795 25857
rect 37826 25848 37832 25860
rect 37884 25848 37890 25900
rect 38105 25891 38163 25897
rect 38105 25857 38117 25891
rect 38151 25888 38163 25891
rect 38286 25888 38292 25900
rect 38151 25860 38292 25888
rect 38151 25857 38163 25860
rect 38105 25851 38163 25857
rect 38286 25848 38292 25860
rect 38344 25848 38350 25900
rect 36078 25780 36084 25832
rect 36136 25820 36142 25832
rect 38841 25823 38899 25829
rect 38841 25820 38853 25823
rect 36136 25792 38853 25820
rect 36136 25780 36142 25792
rect 38841 25789 38853 25792
rect 38887 25789 38899 25823
rect 38841 25783 38899 25789
rect 39298 25780 39304 25832
rect 39356 25780 39362 25832
rect 39574 25780 39580 25832
rect 39632 25780 39638 25832
rect 35802 25752 35808 25764
rect 34931 25724 35808 25752
rect 34931 25721 34943 25724
rect 34885 25715 34943 25721
rect 35802 25712 35808 25724
rect 35860 25712 35866 25764
rect 21600 25656 26004 25684
rect 21600 25644 21606 25656
rect 27430 25644 27436 25696
rect 27488 25644 27494 25696
rect 27798 25644 27804 25696
rect 27856 25644 27862 25696
rect 34790 25644 34796 25696
rect 34848 25644 34854 25696
rect 35529 25687 35587 25693
rect 35529 25653 35541 25687
rect 35575 25684 35587 25687
rect 36078 25684 36084 25696
rect 35575 25656 36084 25684
rect 35575 25653 35587 25656
rect 35529 25647 35587 25653
rect 36078 25644 36084 25656
rect 36136 25644 36142 25696
rect 38286 25644 38292 25696
rect 38344 25644 38350 25696
rect 1104 25594 41400 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 41400 25594
rect 1104 25520 41400 25542
rect 3789 25483 3847 25489
rect 3789 25449 3801 25483
rect 3835 25480 3847 25483
rect 3970 25480 3976 25492
rect 3835 25452 3976 25480
rect 3835 25449 3847 25452
rect 3789 25443 3847 25449
rect 3970 25440 3976 25452
rect 4028 25440 4034 25492
rect 4062 25440 4068 25492
rect 4120 25440 4126 25492
rect 5718 25440 5724 25492
rect 5776 25480 5782 25492
rect 5776 25452 7328 25480
rect 5776 25440 5782 25452
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25344 1455 25347
rect 2406 25344 2412 25356
rect 1443 25316 2412 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 2406 25304 2412 25316
rect 2464 25304 2470 25356
rect 3050 25276 3056 25288
rect 2806 25248 3056 25276
rect 3050 25236 3056 25248
rect 3108 25236 3114 25288
rect 3973 25279 4031 25285
rect 3973 25245 3985 25279
rect 4019 25276 4031 25279
rect 4080 25276 4108 25440
rect 7300 25412 7328 25452
rect 7374 25440 7380 25492
rect 7432 25480 7438 25492
rect 9769 25483 9827 25489
rect 7432 25452 7880 25480
rect 7432 25440 7438 25452
rect 7300 25384 7420 25412
rect 7190 25304 7196 25356
rect 7248 25304 7254 25356
rect 7392 25344 7420 25384
rect 7558 25372 7564 25424
rect 7616 25412 7622 25424
rect 7745 25415 7803 25421
rect 7745 25412 7757 25415
rect 7616 25384 7757 25412
rect 7616 25372 7622 25384
rect 7745 25381 7757 25384
rect 7791 25381 7803 25415
rect 7852 25412 7880 25452
rect 9769 25449 9781 25483
rect 9815 25480 9827 25483
rect 9950 25480 9956 25492
rect 9815 25452 9956 25480
rect 9815 25449 9827 25452
rect 9769 25443 9827 25449
rect 9950 25440 9956 25452
rect 10008 25440 10014 25492
rect 11882 25480 11888 25492
rect 10658 25452 11888 25480
rect 10658 25412 10686 25452
rect 11882 25440 11888 25452
rect 11940 25480 11946 25492
rect 13446 25480 13452 25492
rect 11940 25452 13452 25480
rect 11940 25440 11946 25452
rect 13446 25440 13452 25452
rect 13504 25480 13510 25492
rect 14277 25483 14335 25489
rect 14277 25480 14289 25483
rect 13504 25452 14289 25480
rect 13504 25440 13510 25452
rect 14277 25449 14289 25452
rect 14323 25449 14335 25483
rect 14277 25443 14335 25449
rect 20254 25440 20260 25492
rect 20312 25480 20318 25492
rect 20806 25480 20812 25492
rect 20312 25452 20812 25480
rect 20312 25440 20318 25452
rect 20806 25440 20812 25452
rect 20864 25440 20870 25492
rect 20898 25440 20904 25492
rect 20956 25480 20962 25492
rect 25409 25483 25467 25489
rect 20956 25452 25084 25480
rect 20956 25440 20962 25452
rect 7852 25384 10686 25412
rect 7745 25375 7803 25381
rect 10658 25344 10686 25384
rect 11790 25372 11796 25424
rect 11848 25372 11854 25424
rect 13725 25415 13783 25421
rect 13725 25381 13737 25415
rect 13771 25412 13783 25415
rect 13906 25412 13912 25424
rect 13771 25384 13912 25412
rect 13771 25381 13783 25384
rect 13725 25375 13783 25381
rect 13906 25372 13912 25384
rect 13964 25412 13970 25424
rect 14090 25412 14096 25424
rect 13964 25384 14096 25412
rect 13964 25372 13970 25384
rect 14090 25372 14096 25384
rect 14148 25372 14154 25424
rect 20456 25384 21220 25412
rect 20456 25356 20484 25384
rect 7392 25316 9536 25344
rect 7466 25276 7472 25288
rect 4019 25248 4108 25276
rect 7024 25248 7472 25276
rect 4019 25245 4031 25248
rect 3973 25239 4031 25245
rect 1670 25168 1676 25220
rect 1728 25168 1734 25220
rect 7024 25217 7052 25248
rect 7466 25236 7472 25248
rect 7524 25276 7530 25288
rect 7524 25248 8340 25276
rect 7524 25236 7530 25248
rect 7009 25211 7067 25217
rect 7009 25177 7021 25211
rect 7055 25177 7067 25211
rect 7009 25171 7067 25177
rect 7282 25168 7288 25220
rect 7340 25208 7346 25220
rect 7561 25211 7619 25217
rect 7561 25208 7573 25211
rect 7340 25180 7573 25208
rect 7340 25168 7346 25180
rect 7561 25177 7573 25180
rect 7607 25177 7619 25211
rect 7561 25171 7619 25177
rect 3142 25100 3148 25152
rect 3200 25140 3206 25152
rect 4062 25140 4068 25152
rect 3200 25112 4068 25140
rect 3200 25100 3206 25112
rect 4062 25100 4068 25112
rect 4120 25100 4126 25152
rect 6638 25100 6644 25152
rect 6696 25100 6702 25152
rect 7101 25143 7159 25149
rect 7101 25109 7113 25143
rect 7147 25140 7159 25143
rect 7466 25140 7472 25152
rect 7147 25112 7472 25140
rect 7147 25109 7159 25112
rect 7101 25103 7159 25109
rect 7466 25100 7472 25112
rect 7524 25100 7530 25152
rect 8312 25140 8340 25248
rect 9214 25236 9220 25288
rect 9272 25236 9278 25288
rect 9398 25236 9404 25288
rect 9456 25236 9462 25288
rect 9508 25285 9536 25316
rect 10612 25316 10686 25344
rect 9493 25279 9551 25285
rect 9493 25245 9505 25279
rect 9539 25245 9551 25279
rect 9493 25239 9551 25245
rect 9582 25236 9588 25288
rect 9640 25236 9646 25288
rect 9766 25236 9772 25288
rect 9824 25236 9830 25288
rect 10502 25236 10508 25288
rect 10560 25236 10566 25288
rect 10612 25285 10640 25316
rect 10778 25304 10784 25356
rect 10836 25304 10842 25356
rect 10873 25347 10931 25353
rect 10873 25313 10885 25347
rect 10919 25344 10931 25347
rect 11146 25344 11152 25356
rect 10919 25316 11152 25344
rect 10919 25313 10931 25316
rect 10873 25307 10931 25313
rect 11146 25304 11152 25316
rect 11204 25344 11210 25356
rect 12253 25347 12311 25353
rect 12253 25344 12265 25347
rect 11204 25316 12265 25344
rect 11204 25304 11210 25316
rect 12253 25313 12265 25316
rect 12299 25344 12311 25347
rect 13357 25347 13415 25353
rect 13357 25344 13369 25347
rect 12299 25316 13369 25344
rect 12299 25313 12311 25316
rect 12253 25307 12311 25313
rect 13357 25313 13369 25316
rect 13403 25344 13415 25347
rect 13538 25344 13544 25356
rect 13403 25316 13544 25344
rect 13403 25313 13415 25316
rect 13357 25307 13415 25313
rect 13538 25304 13544 25316
rect 13596 25304 13602 25356
rect 14734 25304 14740 25356
rect 14792 25304 14798 25356
rect 15010 25304 15016 25356
rect 15068 25304 15074 25356
rect 19058 25344 19064 25356
rect 17972 25316 19064 25344
rect 10597 25279 10655 25285
rect 10597 25245 10609 25279
rect 10643 25245 10655 25279
rect 10796 25276 10824 25304
rect 11241 25279 11299 25285
rect 11241 25276 11253 25279
rect 10796 25248 11253 25276
rect 10597 25239 10655 25245
rect 11241 25245 11253 25248
rect 11287 25245 11299 25279
rect 11241 25239 11299 25245
rect 11425 25279 11483 25285
rect 11425 25245 11437 25279
rect 11471 25245 11483 25279
rect 11425 25239 11483 25245
rect 11517 25279 11575 25285
rect 11517 25245 11529 25279
rect 11563 25245 11575 25279
rect 11517 25239 11575 25245
rect 9030 25168 9036 25220
rect 9088 25208 9094 25220
rect 9416 25208 9444 25236
rect 9088 25180 9444 25208
rect 9784 25208 9812 25236
rect 10226 25208 10232 25220
rect 9784 25180 10232 25208
rect 9088 25168 9094 25180
rect 10226 25168 10232 25180
rect 10284 25208 10290 25220
rect 11440 25208 11468 25239
rect 10284 25180 11468 25208
rect 11532 25208 11560 25239
rect 11882 25236 11888 25288
rect 11940 25276 11946 25288
rect 11977 25279 12035 25285
rect 11977 25276 11989 25279
rect 11940 25248 11989 25276
rect 11940 25236 11946 25248
rect 11977 25245 11989 25248
rect 12023 25245 12035 25279
rect 11977 25239 12035 25245
rect 12066 25236 12072 25288
rect 12124 25236 12130 25288
rect 12158 25236 12164 25288
rect 12216 25236 12222 25288
rect 12342 25236 12348 25288
rect 12400 25236 12406 25288
rect 12437 25279 12495 25285
rect 12437 25245 12449 25279
rect 12483 25276 12495 25279
rect 12526 25276 12532 25288
rect 12483 25248 12532 25276
rect 12483 25245 12495 25248
rect 12437 25239 12495 25245
rect 12526 25236 12532 25248
rect 12584 25276 12590 25288
rect 17037 25279 17095 25285
rect 17037 25276 17049 25279
rect 12584 25248 13584 25276
rect 16146 25248 17049 25276
rect 12584 25236 12590 25248
rect 12360 25208 12388 25236
rect 11532 25180 12388 25208
rect 10284 25168 10290 25180
rect 13556 25152 13584 25248
rect 17037 25245 17049 25248
rect 17083 25276 17095 25279
rect 17126 25276 17132 25288
rect 17083 25248 17132 25276
rect 17083 25245 17095 25248
rect 17037 25239 17095 25245
rect 17126 25236 17132 25248
rect 17184 25236 17190 25288
rect 17972 25285 18000 25316
rect 19058 25304 19064 25316
rect 19116 25304 19122 25356
rect 20438 25304 20444 25356
rect 20496 25304 20502 25356
rect 20533 25347 20591 25353
rect 20533 25313 20545 25347
rect 20579 25344 20591 25347
rect 20898 25344 20904 25356
rect 20579 25316 20904 25344
rect 20579 25313 20591 25316
rect 20533 25307 20591 25313
rect 20898 25304 20904 25316
rect 20956 25304 20962 25356
rect 21192 25353 21220 25384
rect 21836 25356 21864 25452
rect 22554 25372 22560 25424
rect 22612 25412 22618 25424
rect 24949 25415 25007 25421
rect 24949 25412 24961 25415
rect 22612 25384 24961 25412
rect 22612 25372 22618 25384
rect 24949 25381 24961 25384
rect 24995 25381 25007 25415
rect 25056 25412 25084 25452
rect 25409 25449 25421 25483
rect 25455 25480 25467 25483
rect 25498 25480 25504 25492
rect 25455 25452 25504 25480
rect 25455 25449 25467 25452
rect 25409 25443 25467 25449
rect 25498 25440 25504 25452
rect 25556 25440 25562 25492
rect 27798 25440 27804 25492
rect 27856 25480 27862 25492
rect 27893 25483 27951 25489
rect 27893 25480 27905 25483
rect 27856 25452 27905 25480
rect 27856 25440 27862 25452
rect 27893 25449 27905 25452
rect 27939 25449 27951 25483
rect 27893 25443 27951 25449
rect 29549 25483 29607 25489
rect 29549 25449 29561 25483
rect 29595 25480 29607 25483
rect 29638 25480 29644 25492
rect 29595 25452 29644 25480
rect 29595 25449 29607 25452
rect 29549 25443 29607 25449
rect 29638 25440 29644 25452
rect 29696 25440 29702 25492
rect 29914 25440 29920 25492
rect 29972 25480 29978 25492
rect 30285 25483 30343 25489
rect 30285 25480 30297 25483
rect 29972 25452 30297 25480
rect 29972 25440 29978 25452
rect 30285 25449 30297 25452
rect 30331 25449 30343 25483
rect 30285 25443 30343 25449
rect 31113 25483 31171 25489
rect 31113 25449 31125 25483
rect 31159 25449 31171 25483
rect 31113 25443 31171 25449
rect 31128 25412 31156 25443
rect 31478 25440 31484 25492
rect 31536 25440 31542 25492
rect 32122 25480 32128 25492
rect 31648 25452 32128 25480
rect 31648 25412 31676 25452
rect 32122 25440 32128 25452
rect 32180 25440 32186 25492
rect 32766 25440 32772 25492
rect 32824 25440 32830 25492
rect 33781 25483 33839 25489
rect 33781 25480 33793 25483
rect 33060 25452 33793 25480
rect 31941 25415 31999 25421
rect 31941 25412 31953 25415
rect 25056 25384 28764 25412
rect 24949 25375 25007 25381
rect 28736 25356 28764 25384
rect 29748 25384 31676 25412
rect 31726 25384 31953 25412
rect 21177 25347 21235 25353
rect 21177 25313 21189 25347
rect 21223 25344 21235 25347
rect 21223 25316 21772 25344
rect 21223 25313 21235 25316
rect 21177 25307 21235 25313
rect 17957 25279 18015 25285
rect 17957 25245 17969 25279
rect 18003 25245 18015 25279
rect 17957 25239 18015 25245
rect 18046 25236 18052 25288
rect 18104 25276 18110 25288
rect 19242 25276 19248 25288
rect 18104 25248 19248 25276
rect 18104 25236 18110 25248
rect 19242 25236 19248 25248
rect 19300 25236 19306 25288
rect 19978 25236 19984 25288
rect 20036 25276 20042 25288
rect 20165 25279 20223 25285
rect 20036 25248 20116 25276
rect 20036 25236 20042 25248
rect 14185 25211 14243 25217
rect 14185 25208 14197 25211
rect 13832 25180 14197 25208
rect 10321 25143 10379 25149
rect 10321 25140 10333 25143
rect 8312 25112 10333 25140
rect 10321 25109 10333 25112
rect 10367 25109 10379 25143
rect 10321 25103 10379 25109
rect 11057 25143 11115 25149
rect 11057 25109 11069 25143
rect 11103 25140 11115 25143
rect 11514 25140 11520 25152
rect 11103 25112 11520 25140
rect 11103 25109 11115 25112
rect 11057 25103 11115 25109
rect 11514 25100 11520 25112
rect 11572 25100 11578 25152
rect 13538 25100 13544 25152
rect 13596 25100 13602 25152
rect 13832 25149 13860 25180
rect 14185 25177 14197 25180
rect 14231 25177 14243 25211
rect 14185 25171 14243 25177
rect 16666 25168 16672 25220
rect 16724 25168 16730 25220
rect 18233 25211 18291 25217
rect 18233 25177 18245 25211
rect 18279 25208 18291 25211
rect 18506 25208 18512 25220
rect 18279 25180 18512 25208
rect 18279 25177 18291 25180
rect 18233 25171 18291 25177
rect 18506 25168 18512 25180
rect 18564 25168 18570 25220
rect 20088 25208 20116 25248
rect 20165 25245 20177 25279
rect 20211 25276 20223 25279
rect 20990 25276 20996 25288
rect 20211 25248 20996 25276
rect 20211 25245 20223 25248
rect 20165 25239 20223 25245
rect 20990 25236 20996 25248
rect 21048 25276 21054 25288
rect 21269 25279 21327 25285
rect 21269 25276 21281 25279
rect 21048 25248 21281 25276
rect 21048 25236 21054 25248
rect 21269 25245 21281 25248
rect 21315 25245 21327 25279
rect 21269 25239 21327 25245
rect 21637 25279 21695 25285
rect 21637 25245 21649 25279
rect 21683 25245 21695 25279
rect 21744 25276 21772 25316
rect 21818 25304 21824 25356
rect 21876 25304 21882 25356
rect 27522 25344 27528 25356
rect 25056 25316 27292 25344
rect 22094 25276 22100 25288
rect 21744 25248 22100 25276
rect 21637 25239 21695 25245
rect 20625 25211 20683 25217
rect 20088 25180 20300 25208
rect 13817 25143 13875 25149
rect 13817 25109 13829 25143
rect 13863 25109 13875 25143
rect 13817 25103 13875 25109
rect 15654 25100 15660 25152
rect 15712 25140 15718 25152
rect 16485 25143 16543 25149
rect 16485 25140 16497 25143
rect 15712 25112 16497 25140
rect 15712 25100 15718 25112
rect 16485 25109 16497 25112
rect 16531 25109 16543 25143
rect 16485 25103 16543 25109
rect 17957 25143 18015 25149
rect 17957 25109 17969 25143
rect 18003 25140 18015 25143
rect 18138 25140 18144 25152
rect 18003 25112 18144 25140
rect 18003 25109 18015 25112
rect 17957 25103 18015 25109
rect 18138 25100 18144 25112
rect 18196 25100 18202 25152
rect 20070 25100 20076 25152
rect 20128 25140 20134 25152
rect 20165 25143 20223 25149
rect 20165 25140 20177 25143
rect 20128 25112 20177 25140
rect 20128 25100 20134 25112
rect 20165 25109 20177 25112
rect 20211 25109 20223 25143
rect 20272 25140 20300 25180
rect 20625 25177 20637 25211
rect 20671 25208 20683 25211
rect 21542 25208 21548 25220
rect 20671 25180 21548 25208
rect 20671 25177 20683 25180
rect 20625 25171 20683 25177
rect 21542 25168 21548 25180
rect 21600 25168 21606 25220
rect 21652 25208 21680 25239
rect 22094 25236 22100 25248
rect 22152 25236 22158 25288
rect 22738 25236 22744 25288
rect 22796 25276 22802 25288
rect 25056 25276 25084 25316
rect 22796 25248 25084 25276
rect 22796 25236 22802 25248
rect 25130 25236 25136 25288
rect 25188 25236 25194 25288
rect 25225 25279 25283 25285
rect 25225 25245 25237 25279
rect 25271 25245 25283 25279
rect 25225 25239 25283 25245
rect 22002 25208 22008 25220
rect 21652 25180 22008 25208
rect 21652 25140 21680 25180
rect 22002 25168 22008 25180
rect 22060 25168 22066 25220
rect 23382 25168 23388 25220
rect 23440 25208 23446 25220
rect 24486 25208 24492 25220
rect 23440 25180 24492 25208
rect 23440 25168 23446 25180
rect 24486 25168 24492 25180
rect 24544 25168 24550 25220
rect 20272 25112 21680 25140
rect 20165 25103 20223 25109
rect 22186 25100 22192 25152
rect 22244 25140 22250 25152
rect 24946 25140 24952 25152
rect 22244 25112 24952 25140
rect 22244 25100 22250 25112
rect 24946 25100 24952 25112
rect 25004 25100 25010 25152
rect 25240 25140 25268 25239
rect 25314 25236 25320 25288
rect 25372 25276 25378 25288
rect 25501 25279 25559 25285
rect 25501 25276 25513 25279
rect 25372 25248 25513 25276
rect 25372 25236 25378 25248
rect 25501 25245 25513 25248
rect 25547 25276 25559 25279
rect 25547 25248 27228 25276
rect 25547 25245 25559 25248
rect 25501 25239 25559 25245
rect 26970 25140 26976 25152
rect 25240 25112 26976 25140
rect 26970 25100 26976 25112
rect 27028 25100 27034 25152
rect 27200 25140 27228 25248
rect 27264 25208 27292 25316
rect 27356 25316 27528 25344
rect 27356 25285 27384 25316
rect 27522 25304 27528 25316
rect 27580 25304 27586 25356
rect 28718 25304 28724 25356
rect 28776 25304 28782 25356
rect 27341 25279 27399 25285
rect 27341 25245 27353 25279
rect 27387 25245 27399 25279
rect 27341 25239 27399 25245
rect 27614 25236 27620 25288
rect 27672 25236 27678 25288
rect 27709 25279 27767 25285
rect 27709 25245 27721 25279
rect 27755 25276 27767 25279
rect 28902 25276 28908 25288
rect 27755 25248 28908 25276
rect 27755 25245 27767 25248
rect 27709 25239 27767 25245
rect 28902 25236 28908 25248
rect 28960 25236 28966 25288
rect 29638 25236 29644 25288
rect 29696 25276 29702 25288
rect 29748 25285 29776 25384
rect 30561 25347 30619 25353
rect 30561 25313 30573 25347
rect 30607 25344 30619 25347
rect 31205 25347 31263 25353
rect 31205 25344 31217 25347
rect 30607 25316 31217 25344
rect 30607 25313 30619 25316
rect 30561 25307 30619 25313
rect 31205 25313 31217 25316
rect 31251 25344 31263 25347
rect 31726 25344 31754 25384
rect 31941 25381 31953 25384
rect 31987 25381 31999 25415
rect 31941 25375 31999 25381
rect 32490 25372 32496 25424
rect 32548 25412 32554 25424
rect 33060 25412 33088 25452
rect 33781 25449 33793 25452
rect 33827 25449 33839 25483
rect 33781 25443 33839 25449
rect 34790 25440 34796 25492
rect 34848 25480 34854 25492
rect 34977 25483 35035 25489
rect 34977 25480 34989 25483
rect 34848 25452 34989 25480
rect 34848 25440 34854 25452
rect 34977 25449 34989 25452
rect 35023 25449 35035 25483
rect 36722 25480 36728 25492
rect 34977 25443 35035 25449
rect 35452 25452 36728 25480
rect 32548 25384 33088 25412
rect 33137 25415 33195 25421
rect 32548 25372 32554 25384
rect 33137 25381 33149 25415
rect 33183 25412 33195 25415
rect 33962 25412 33968 25424
rect 33183 25384 33968 25412
rect 33183 25381 33195 25384
rect 33137 25375 33195 25381
rect 33152 25344 33180 25375
rect 33962 25372 33968 25384
rect 34020 25372 34026 25424
rect 33594 25344 33600 25356
rect 31251 25316 31754 25344
rect 31956 25316 33180 25344
rect 33336 25316 33600 25344
rect 31251 25313 31263 25316
rect 31205 25307 31263 25313
rect 29733 25279 29791 25285
rect 29733 25276 29745 25279
rect 29696 25248 29745 25276
rect 29696 25236 29702 25248
rect 29733 25245 29745 25248
rect 29779 25245 29791 25279
rect 29733 25239 29791 25245
rect 29825 25279 29883 25285
rect 29825 25245 29837 25279
rect 29871 25245 29883 25279
rect 29825 25239 29883 25245
rect 27525 25211 27583 25217
rect 27525 25208 27537 25211
rect 27264 25180 27537 25208
rect 27525 25177 27537 25180
rect 27571 25208 27583 25211
rect 27890 25208 27896 25220
rect 27571 25180 27896 25208
rect 27571 25177 27583 25180
rect 27525 25171 27583 25177
rect 27890 25168 27896 25180
rect 27948 25168 27954 25220
rect 29840 25208 29868 25239
rect 29914 25236 29920 25288
rect 29972 25236 29978 25288
rect 30006 25236 30012 25288
rect 30064 25236 30070 25288
rect 30374 25236 30380 25288
rect 30432 25276 30438 25288
rect 30469 25279 30527 25285
rect 30469 25276 30481 25279
rect 30432 25248 30481 25276
rect 30432 25236 30438 25248
rect 30469 25245 30481 25248
rect 30515 25245 30527 25279
rect 30469 25239 30527 25245
rect 30650 25236 30656 25288
rect 30708 25236 30714 25288
rect 30745 25279 30803 25285
rect 30745 25245 30757 25279
rect 30791 25276 30803 25279
rect 30834 25276 30840 25288
rect 30791 25248 30840 25276
rect 30791 25245 30803 25248
rect 30745 25239 30803 25245
rect 30834 25236 30840 25248
rect 30892 25236 30898 25288
rect 31956 25285 31984 25316
rect 33336 25288 33364 25316
rect 33594 25304 33600 25316
rect 33652 25344 33658 25356
rect 34057 25347 34115 25353
rect 34057 25344 34069 25347
rect 33652 25316 34069 25344
rect 33652 25304 33658 25316
rect 34057 25313 34069 25316
rect 34103 25313 34115 25347
rect 34057 25307 34115 25313
rect 34238 25304 34244 25356
rect 34296 25344 34302 25356
rect 35345 25347 35403 25353
rect 35345 25344 35357 25347
rect 34296 25316 35357 25344
rect 34296 25304 34302 25316
rect 35345 25313 35357 25316
rect 35391 25313 35403 25347
rect 35345 25307 35403 25313
rect 31113 25279 31171 25285
rect 31113 25245 31125 25279
rect 31159 25245 31171 25279
rect 31113 25239 31171 25245
rect 31941 25279 31999 25285
rect 31941 25245 31953 25279
rect 31987 25245 31999 25279
rect 31941 25239 31999 25245
rect 30282 25208 30288 25220
rect 29840 25180 30288 25208
rect 30282 25168 30288 25180
rect 30340 25208 30346 25220
rect 31128 25208 31156 25239
rect 32030 25236 32036 25288
rect 32088 25276 32094 25288
rect 32217 25279 32275 25285
rect 32217 25276 32229 25279
rect 32088 25248 32229 25276
rect 32088 25236 32094 25248
rect 32217 25245 32229 25248
rect 32263 25245 32275 25279
rect 32217 25239 32275 25245
rect 32398 25236 32404 25288
rect 32456 25236 32462 25288
rect 32674 25236 32680 25288
rect 32732 25236 32738 25288
rect 32950 25236 32956 25288
rect 33008 25236 33014 25288
rect 33045 25279 33103 25285
rect 33045 25245 33057 25279
rect 33091 25245 33103 25279
rect 33045 25239 33103 25245
rect 33229 25279 33287 25285
rect 33229 25245 33241 25279
rect 33275 25245 33287 25279
rect 33229 25239 33287 25245
rect 30340 25180 31156 25208
rect 30340 25168 30346 25180
rect 27798 25140 27804 25152
rect 27200 25112 27804 25140
rect 27798 25100 27804 25112
rect 27856 25100 27862 25152
rect 31128 25140 31156 25180
rect 31754 25168 31760 25220
rect 31812 25208 31818 25220
rect 32048 25208 32076 25236
rect 31812 25180 32076 25208
rect 32125 25211 32183 25217
rect 31812 25168 31818 25180
rect 32125 25177 32137 25211
rect 32171 25208 32183 25211
rect 32416 25208 32444 25236
rect 32171 25180 32444 25208
rect 32692 25208 32720 25236
rect 33060 25208 33088 25239
rect 32692 25180 33088 25208
rect 32171 25177 32183 25180
rect 32125 25171 32183 25177
rect 32490 25140 32496 25152
rect 31128 25112 32496 25140
rect 32490 25100 32496 25112
rect 32548 25100 32554 25152
rect 32950 25100 32956 25152
rect 33008 25140 33014 25152
rect 33244 25140 33272 25239
rect 33318 25236 33324 25288
rect 33376 25236 33382 25288
rect 33413 25279 33471 25285
rect 33413 25245 33425 25279
rect 33459 25245 33471 25279
rect 33413 25239 33471 25245
rect 33008 25112 33272 25140
rect 33428 25140 33456 25239
rect 34146 25236 34152 25288
rect 34204 25276 34210 25288
rect 35452 25276 35480 25452
rect 36722 25440 36728 25452
rect 36780 25480 36786 25492
rect 36780 25452 37780 25480
rect 36780 25440 36786 25452
rect 37550 25412 37556 25424
rect 35728 25384 37556 25412
rect 35728 25285 35756 25384
rect 37550 25372 37556 25384
rect 37608 25412 37614 25424
rect 37645 25415 37703 25421
rect 37645 25412 37657 25415
rect 37608 25384 37657 25412
rect 37608 25372 37614 25384
rect 37645 25381 37657 25384
rect 37691 25381 37703 25415
rect 37752 25412 37780 25452
rect 37826 25440 37832 25492
rect 37884 25440 37890 25492
rect 39574 25440 39580 25492
rect 39632 25480 39638 25492
rect 39853 25483 39911 25489
rect 39853 25480 39865 25483
rect 39632 25452 39865 25480
rect 39632 25440 39638 25452
rect 39853 25449 39865 25452
rect 39899 25449 39911 25483
rect 39853 25443 39911 25449
rect 40126 25440 40132 25492
rect 40184 25480 40190 25492
rect 40773 25483 40831 25489
rect 40773 25480 40785 25483
rect 40184 25452 40785 25480
rect 40184 25440 40190 25452
rect 40773 25449 40785 25452
rect 40819 25449 40831 25483
rect 40773 25443 40831 25449
rect 38933 25415 38991 25421
rect 38933 25412 38945 25415
rect 37752 25384 38945 25412
rect 37645 25375 37703 25381
rect 38933 25381 38945 25384
rect 38979 25381 38991 25415
rect 38933 25375 38991 25381
rect 35802 25304 35808 25356
rect 35860 25304 35866 25356
rect 37829 25347 37887 25353
rect 37829 25344 37841 25347
rect 37476 25316 37841 25344
rect 36078 25285 36084 25288
rect 34204 25248 35480 25276
rect 35529 25279 35587 25285
rect 34204 25236 34210 25248
rect 35529 25245 35541 25279
rect 35575 25245 35587 25279
rect 35529 25239 35587 25245
rect 35713 25279 35771 25285
rect 35713 25245 35725 25279
rect 35759 25245 35771 25279
rect 35713 25239 35771 25245
rect 35915 25279 35973 25285
rect 35915 25245 35927 25279
rect 35961 25276 35973 25279
rect 35961 25248 36032 25276
rect 35961 25245 35973 25248
rect 35915 25239 35973 25245
rect 33594 25168 33600 25220
rect 33652 25208 33658 25220
rect 33689 25211 33747 25217
rect 33689 25208 33701 25211
rect 33652 25180 33701 25208
rect 33652 25168 33658 25180
rect 33689 25177 33701 25180
rect 33735 25208 33747 25211
rect 35544 25208 35572 25239
rect 33735 25180 35572 25208
rect 36004 25208 36032 25248
rect 36075 25239 36084 25285
rect 36136 25276 36142 25288
rect 36136 25248 36175 25276
rect 36078 25236 36084 25239
rect 36136 25236 36142 25248
rect 36998 25236 37004 25288
rect 37056 25236 37062 25288
rect 37090 25236 37096 25288
rect 37148 25276 37154 25288
rect 37185 25279 37243 25285
rect 37185 25276 37197 25279
rect 37148 25248 37197 25276
rect 37148 25236 37154 25248
rect 37185 25245 37197 25248
rect 37231 25245 37243 25279
rect 37185 25239 37243 25245
rect 37277 25279 37335 25285
rect 37277 25245 37289 25279
rect 37323 25276 37335 25279
rect 37366 25276 37372 25288
rect 37323 25248 37372 25276
rect 37323 25245 37335 25248
rect 37277 25239 37335 25245
rect 37366 25236 37372 25248
rect 37424 25236 37430 25288
rect 37476 25285 37504 25316
rect 37829 25313 37841 25316
rect 37875 25344 37887 25347
rect 38286 25344 38292 25356
rect 37875 25316 38292 25344
rect 37875 25313 37887 25316
rect 37829 25307 37887 25313
rect 38286 25304 38292 25316
rect 38344 25304 38350 25356
rect 37461 25279 37519 25285
rect 37461 25245 37473 25279
rect 37507 25245 37519 25279
rect 37461 25239 37519 25245
rect 37737 25279 37795 25285
rect 37737 25245 37749 25279
rect 37783 25245 37795 25279
rect 37737 25239 37795 25245
rect 38749 25279 38807 25285
rect 38749 25245 38761 25279
rect 38795 25276 38807 25279
rect 39758 25276 39764 25288
rect 38795 25248 39764 25276
rect 38795 25245 38807 25248
rect 38749 25239 38807 25245
rect 36004 25180 36216 25208
rect 33735 25177 33747 25180
rect 33689 25171 33747 25177
rect 36188 25152 36216 25180
rect 37752 25152 37780 25239
rect 39758 25236 39764 25248
rect 39816 25236 39822 25288
rect 40034 25236 40040 25288
rect 40092 25236 40098 25288
rect 40494 25168 40500 25220
rect 40552 25208 40558 25220
rect 40681 25211 40739 25217
rect 40681 25208 40693 25211
rect 40552 25180 40693 25208
rect 40552 25168 40558 25180
rect 40681 25177 40693 25180
rect 40727 25177 40739 25211
rect 40681 25171 40739 25177
rect 34333 25143 34391 25149
rect 34333 25140 34345 25143
rect 33428 25112 34345 25140
rect 33008 25100 33014 25112
rect 34333 25109 34345 25112
rect 34379 25109 34391 25143
rect 34333 25103 34391 25109
rect 36170 25100 36176 25152
rect 36228 25100 36234 25152
rect 37090 25100 37096 25152
rect 37148 25100 37154 25152
rect 37734 25100 37740 25152
rect 37792 25100 37798 25152
rect 38102 25100 38108 25152
rect 38160 25100 38166 25152
rect 1104 25050 41400 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 41400 25050
rect 1104 24976 41400 24998
rect 1670 24896 1676 24948
rect 1728 24936 1734 24948
rect 1857 24939 1915 24945
rect 1857 24936 1869 24939
rect 1728 24908 1869 24936
rect 1728 24896 1734 24908
rect 1857 24905 1869 24908
rect 1903 24905 1915 24939
rect 1857 24899 1915 24905
rect 2866 24896 2872 24948
rect 2924 24896 2930 24948
rect 2961 24939 3019 24945
rect 2961 24905 2973 24939
rect 3007 24936 3019 24939
rect 3142 24936 3148 24948
rect 3007 24908 3148 24936
rect 3007 24905 3019 24908
rect 2961 24899 3019 24905
rect 3142 24896 3148 24908
rect 3200 24896 3206 24948
rect 5074 24936 5080 24948
rect 4632 24908 5080 24936
rect 2041 24803 2099 24809
rect 2041 24769 2053 24803
rect 2087 24800 2099 24803
rect 2087 24772 2544 24800
rect 2087 24769 2099 24772
rect 2041 24763 2099 24769
rect 2516 24673 2544 24772
rect 3970 24760 3976 24812
rect 4028 24800 4034 24812
rect 4632 24809 4660 24908
rect 5074 24896 5080 24908
rect 5132 24896 5138 24948
rect 5169 24939 5227 24945
rect 5169 24905 5181 24939
rect 5215 24936 5227 24939
rect 5626 24936 5632 24948
rect 5215 24908 5632 24936
rect 5215 24905 5227 24908
rect 5169 24899 5227 24905
rect 5626 24896 5632 24908
rect 5684 24896 5690 24948
rect 5810 24896 5816 24948
rect 5868 24896 5874 24948
rect 6638 24896 6644 24948
rect 6696 24896 6702 24948
rect 7466 24896 7472 24948
rect 7524 24936 7530 24948
rect 8110 24936 8116 24948
rect 7524 24908 8116 24936
rect 7524 24896 7530 24908
rect 8110 24896 8116 24908
rect 8168 24896 8174 24948
rect 9674 24936 9680 24948
rect 8450 24908 9680 24936
rect 6656 24868 6684 24896
rect 4816 24840 5764 24868
rect 4341 24803 4399 24809
rect 4341 24800 4353 24803
rect 4028 24772 4353 24800
rect 4028 24760 4034 24772
rect 4341 24769 4353 24772
rect 4387 24769 4399 24803
rect 4341 24763 4399 24769
rect 4525 24803 4583 24809
rect 4525 24769 4537 24803
rect 4571 24769 4583 24803
rect 4525 24763 4583 24769
rect 4617 24803 4675 24809
rect 4617 24769 4629 24803
rect 4663 24769 4675 24803
rect 4617 24763 4675 24769
rect 3145 24735 3203 24741
rect 3145 24701 3157 24735
rect 3191 24732 3203 24735
rect 3878 24732 3884 24744
rect 3191 24704 3884 24732
rect 3191 24701 3203 24704
rect 3145 24695 3203 24701
rect 3878 24692 3884 24704
rect 3936 24692 3942 24744
rect 2501 24667 2559 24673
rect 2501 24633 2513 24667
rect 2547 24633 2559 24667
rect 4540 24664 4568 24763
rect 4709 24735 4767 24741
rect 4709 24701 4721 24735
rect 4755 24732 4767 24735
rect 4816 24732 4844 24840
rect 4893 24803 4951 24809
rect 4893 24769 4905 24803
rect 4939 24800 4951 24803
rect 5074 24800 5080 24812
rect 4939 24772 5080 24800
rect 4939 24769 4951 24772
rect 4893 24763 4951 24769
rect 5074 24760 5080 24772
rect 5132 24760 5138 24812
rect 5166 24760 5172 24812
rect 5224 24806 5230 24812
rect 5353 24806 5411 24809
rect 5224 24803 5411 24806
rect 5224 24778 5365 24803
rect 5224 24760 5230 24778
rect 5353 24769 5365 24778
rect 5399 24769 5411 24803
rect 5353 24763 5411 24769
rect 5534 24760 5540 24812
rect 5592 24760 5598 24812
rect 4755 24704 4844 24732
rect 4755 24701 4767 24704
rect 4709 24695 4767 24701
rect 5258 24692 5264 24744
rect 5316 24692 5322 24744
rect 5626 24692 5632 24744
rect 5684 24732 5690 24744
rect 5736 24732 5764 24840
rect 6196 24840 6684 24868
rect 6196 24809 6224 24840
rect 7098 24828 7104 24880
rect 7156 24828 7162 24880
rect 8018 24828 8024 24880
rect 8076 24868 8082 24880
rect 8450 24868 8478 24908
rect 9674 24896 9680 24908
rect 9732 24896 9738 24948
rect 9766 24896 9772 24948
rect 9824 24896 9830 24948
rect 10965 24939 11023 24945
rect 10965 24905 10977 24939
rect 11011 24905 11023 24939
rect 10965 24899 11023 24905
rect 11241 24939 11299 24945
rect 11241 24905 11253 24939
rect 11287 24936 11299 24939
rect 12066 24936 12072 24948
rect 11287 24908 12072 24936
rect 11287 24905 11299 24908
rect 11241 24899 11299 24905
rect 10980 24868 11008 24899
rect 12066 24896 12072 24908
rect 12124 24896 12130 24948
rect 12250 24896 12256 24948
rect 12308 24936 12314 24948
rect 13906 24936 13912 24948
rect 12308 24908 13912 24936
rect 12308 24896 12314 24908
rect 13906 24896 13912 24908
rect 13964 24936 13970 24948
rect 14001 24939 14059 24945
rect 14001 24936 14013 24939
rect 13964 24908 14013 24936
rect 13964 24896 13970 24908
rect 14001 24905 14013 24908
rect 14047 24905 14059 24939
rect 14001 24899 14059 24905
rect 14826 24896 14832 24948
rect 14884 24896 14890 24948
rect 15105 24939 15163 24945
rect 15105 24905 15117 24939
rect 15151 24936 15163 24939
rect 15194 24936 15200 24948
rect 15151 24908 15200 24936
rect 15151 24905 15163 24908
rect 15105 24899 15163 24905
rect 15194 24896 15200 24908
rect 15252 24896 15258 24948
rect 18417 24939 18475 24945
rect 18417 24936 18429 24939
rect 17420 24908 18429 24936
rect 12342 24868 12348 24880
rect 8076 24840 8478 24868
rect 9646 24840 12348 24868
rect 8076 24828 8082 24840
rect 6181 24803 6239 24809
rect 6181 24769 6193 24803
rect 6227 24769 6239 24803
rect 6181 24763 6239 24769
rect 6362 24760 6368 24812
rect 6420 24760 6426 24812
rect 8202 24760 8208 24812
rect 8260 24760 8266 24812
rect 8294 24760 8300 24812
rect 8352 24800 8358 24812
rect 8573 24803 8631 24809
rect 8573 24800 8585 24803
rect 8352 24772 8585 24800
rect 8352 24760 8358 24772
rect 8573 24769 8585 24772
rect 8619 24769 8631 24803
rect 8573 24763 8631 24769
rect 8665 24803 8723 24809
rect 8665 24769 8677 24803
rect 8711 24800 8723 24803
rect 8754 24800 8760 24812
rect 8711 24772 8760 24800
rect 8711 24769 8723 24772
rect 8665 24763 8723 24769
rect 8754 24760 8760 24772
rect 8812 24760 8818 24812
rect 9493 24803 9551 24809
rect 9493 24800 9505 24803
rect 8864 24772 9505 24800
rect 5684 24704 5764 24732
rect 5684 24692 5690 24704
rect 5902 24692 5908 24744
rect 5960 24692 5966 24744
rect 6641 24735 6699 24741
rect 6641 24732 6653 24735
rect 6012 24704 6653 24732
rect 4614 24664 4620 24676
rect 4540 24636 4620 24664
rect 2501 24627 2559 24633
rect 4614 24624 4620 24636
rect 4672 24624 4678 24676
rect 5166 24624 5172 24676
rect 5224 24624 5230 24676
rect 6012 24673 6040 24704
rect 6641 24701 6653 24704
rect 6687 24701 6699 24735
rect 6641 24695 6699 24701
rect 5997 24667 6055 24673
rect 5997 24633 6009 24667
rect 6043 24633 6055 24667
rect 8225 24664 8253 24760
rect 8864 24664 8892 24772
rect 9493 24769 9505 24772
rect 9539 24800 9551 24803
rect 9646 24800 9674 24840
rect 12342 24828 12348 24840
rect 12400 24828 12406 24880
rect 12802 24828 12808 24880
rect 12860 24868 12866 24880
rect 13630 24868 13636 24880
rect 12860 24840 13216 24868
rect 12860 24828 12866 24840
rect 9539 24772 9674 24800
rect 9539 24769 9551 24772
rect 9493 24763 9551 24769
rect 10226 24760 10232 24812
rect 10284 24800 10290 24812
rect 10781 24803 10839 24809
rect 10781 24800 10793 24803
rect 10284 24772 10793 24800
rect 10284 24760 10290 24772
rect 10781 24769 10793 24772
rect 10827 24769 10839 24803
rect 10781 24763 10839 24769
rect 10873 24803 10931 24809
rect 10873 24769 10885 24803
rect 10919 24800 10931 24803
rect 11146 24800 11152 24812
rect 10919 24772 11152 24800
rect 10919 24769 10931 24772
rect 10873 24763 10931 24769
rect 11146 24760 11152 24772
rect 11204 24760 11210 24812
rect 13188 24809 13216 24840
rect 13418 24840 13636 24868
rect 11241 24803 11299 24809
rect 11241 24769 11253 24803
rect 11287 24800 11299 24803
rect 12161 24803 12219 24809
rect 12161 24800 12173 24803
rect 11287 24772 12173 24800
rect 11287 24769 11299 24772
rect 11241 24763 11299 24769
rect 12161 24769 12173 24772
rect 12207 24800 12219 24803
rect 12989 24803 13047 24809
rect 12989 24800 13001 24803
rect 12207 24772 12848 24800
rect 12207 24769 12219 24772
rect 12161 24763 12219 24769
rect 9306 24692 9312 24744
rect 9364 24692 9370 24744
rect 9861 24735 9919 24741
rect 9861 24701 9873 24735
rect 9907 24701 9919 24735
rect 9861 24695 9919 24701
rect 8225 24636 8892 24664
rect 5997 24627 6055 24633
rect 9214 24624 9220 24676
rect 9272 24664 9278 24676
rect 9876 24664 9904 24695
rect 12345 24667 12403 24673
rect 12345 24664 12357 24667
rect 9272 24636 12357 24664
rect 9272 24624 9278 24636
rect 12345 24633 12357 24636
rect 12391 24633 12403 24667
rect 12345 24627 12403 24633
rect 4341 24599 4399 24605
rect 4341 24565 4353 24599
rect 4387 24596 4399 24599
rect 5184 24596 5212 24624
rect 12820 24608 12848 24772
rect 12912 24772 13001 24800
rect 4387 24568 5212 24596
rect 4387 24565 4399 24568
rect 4341 24559 4399 24565
rect 8846 24556 8852 24608
rect 8904 24556 8910 24608
rect 11149 24599 11207 24605
rect 11149 24565 11161 24599
rect 11195 24596 11207 24599
rect 11974 24596 11980 24608
rect 11195 24568 11980 24596
rect 11195 24565 11207 24568
rect 11149 24559 11207 24565
rect 11974 24556 11980 24568
rect 12032 24556 12038 24608
rect 12802 24556 12808 24608
rect 12860 24556 12866 24608
rect 12912 24596 12940 24772
rect 12989 24769 13001 24772
rect 13035 24769 13047 24803
rect 12989 24763 13047 24769
rect 13173 24803 13231 24809
rect 13173 24769 13185 24803
rect 13219 24769 13231 24803
rect 13173 24763 13231 24769
rect 13188 24732 13216 24763
rect 13262 24760 13268 24812
rect 13320 24760 13326 24812
rect 13418 24809 13446 24840
rect 13630 24828 13636 24840
rect 13688 24828 13694 24880
rect 14274 24868 14280 24880
rect 13740 24840 14280 24868
rect 13740 24809 13768 24840
rect 14274 24828 14280 24840
rect 14332 24828 14338 24880
rect 14366 24828 14372 24880
rect 14424 24868 14430 24880
rect 14844 24868 14872 24896
rect 15473 24871 15531 24877
rect 15473 24868 15485 24871
rect 14424 24840 15485 24868
rect 14424 24828 14430 24840
rect 15473 24837 15485 24840
rect 15519 24837 15531 24871
rect 15473 24831 15531 24837
rect 15565 24871 15623 24877
rect 15565 24837 15577 24871
rect 15611 24868 15623 24871
rect 15654 24868 15660 24880
rect 15611 24840 15660 24868
rect 15611 24837 15623 24840
rect 15565 24831 15623 24837
rect 15654 24828 15660 24840
rect 15712 24828 15718 24880
rect 13403 24803 13461 24809
rect 13403 24769 13415 24803
rect 13449 24769 13461 24803
rect 13403 24763 13461 24769
rect 13725 24803 13783 24809
rect 13725 24769 13737 24803
rect 13771 24769 13783 24803
rect 13725 24763 13783 24769
rect 13814 24760 13820 24812
rect 13872 24760 13878 24812
rect 14458 24760 14464 24812
rect 14516 24760 14522 24812
rect 14642 24760 14648 24812
rect 14700 24760 14706 24812
rect 14734 24760 14740 24812
rect 14792 24760 14798 24812
rect 14829 24803 14887 24809
rect 14829 24769 14841 24803
rect 14875 24800 14887 24803
rect 17034 24800 17040 24812
rect 14875 24772 17040 24800
rect 14875 24769 14887 24772
rect 14829 24763 14887 24769
rect 14660 24732 14688 24760
rect 13188 24704 14688 24732
rect 13170 24624 13176 24676
rect 13228 24664 13234 24676
rect 13228 24636 13584 24664
rect 13228 24624 13234 24636
rect 13262 24596 13268 24608
rect 12912 24568 13268 24596
rect 13262 24556 13268 24568
rect 13320 24556 13326 24608
rect 13556 24605 13584 24636
rect 13630 24624 13636 24676
rect 13688 24664 13694 24676
rect 14844 24664 14872 24763
rect 17034 24760 17040 24772
rect 17092 24760 17098 24812
rect 17313 24803 17371 24809
rect 17313 24769 17325 24803
rect 17359 24800 17371 24803
rect 17420 24800 17448 24908
rect 18417 24905 18429 24908
rect 18463 24936 18475 24939
rect 19058 24936 19064 24948
rect 18463 24908 19064 24936
rect 18463 24905 18475 24908
rect 18417 24899 18475 24905
rect 19058 24896 19064 24908
rect 19116 24896 19122 24948
rect 19242 24896 19248 24948
rect 19300 24936 19306 24948
rect 19889 24939 19947 24945
rect 19889 24936 19901 24939
rect 19300 24908 19901 24936
rect 19300 24896 19306 24908
rect 19889 24905 19901 24908
rect 19935 24905 19947 24939
rect 19889 24899 19947 24905
rect 22002 24896 22008 24948
rect 22060 24896 22066 24948
rect 22296 24908 23244 24936
rect 18046 24868 18052 24880
rect 17696 24840 18052 24868
rect 17359 24772 17448 24800
rect 17497 24803 17555 24809
rect 17359 24769 17371 24772
rect 17313 24763 17371 24769
rect 17497 24769 17509 24803
rect 17543 24800 17555 24803
rect 17696 24800 17724 24840
rect 18046 24828 18052 24840
rect 18104 24828 18110 24880
rect 19521 24871 19579 24877
rect 19168 24840 19380 24868
rect 17543 24772 17724 24800
rect 17773 24803 17831 24809
rect 17543 24769 17555 24772
rect 17497 24763 17555 24769
rect 17773 24769 17785 24803
rect 17819 24800 17831 24803
rect 19061 24803 19119 24809
rect 17819 24772 18092 24800
rect 17819 24769 17831 24772
rect 17773 24763 17831 24769
rect 15562 24692 15568 24744
rect 15620 24732 15626 24744
rect 15746 24732 15752 24744
rect 15620 24704 15752 24732
rect 15620 24692 15626 24704
rect 15746 24692 15752 24704
rect 15804 24692 15810 24744
rect 17589 24735 17647 24741
rect 17589 24701 17601 24735
rect 17635 24701 17647 24735
rect 17589 24695 17647 24701
rect 13688 24636 14872 24664
rect 13688 24624 13694 24636
rect 13541 24599 13599 24605
rect 13541 24565 13553 24599
rect 13587 24565 13599 24599
rect 13541 24559 13599 24565
rect 15013 24599 15071 24605
rect 15013 24565 15025 24599
rect 15059 24596 15071 24599
rect 15102 24596 15108 24608
rect 15059 24568 15108 24596
rect 15059 24565 15071 24568
rect 15013 24559 15071 24565
rect 15102 24556 15108 24568
rect 15160 24556 15166 24608
rect 15470 24556 15476 24608
rect 15528 24596 15534 24608
rect 17034 24596 17040 24608
rect 15528 24568 17040 24596
rect 15528 24556 15534 24568
rect 17034 24556 17040 24568
rect 17092 24556 17098 24608
rect 17310 24556 17316 24608
rect 17368 24556 17374 24608
rect 17604 24596 17632 24695
rect 17770 24624 17776 24676
rect 17828 24664 17834 24676
rect 18064 24673 18092 24772
rect 19061 24769 19073 24803
rect 19107 24800 19119 24803
rect 19168 24800 19196 24840
rect 19107 24772 19196 24800
rect 19107 24769 19119 24772
rect 19061 24763 19119 24769
rect 19242 24760 19248 24812
rect 19300 24760 19306 24812
rect 19352 24800 19380 24840
rect 19521 24837 19533 24871
rect 19567 24868 19579 24871
rect 19610 24868 19616 24880
rect 19567 24840 19616 24868
rect 19567 24837 19579 24840
rect 19521 24831 19579 24837
rect 19610 24828 19616 24840
rect 19668 24828 19674 24880
rect 19726 24871 19784 24877
rect 19726 24868 19738 24871
rect 19720 24837 19738 24868
rect 19772 24837 19784 24871
rect 19720 24831 19784 24837
rect 20916 24840 21220 24868
rect 19720 24800 19748 24831
rect 20254 24800 20260 24812
rect 19352 24772 20260 24800
rect 20254 24760 20260 24772
rect 20312 24760 20318 24812
rect 20625 24803 20683 24809
rect 20625 24769 20637 24803
rect 20671 24800 20683 24803
rect 20806 24800 20812 24812
rect 20671 24772 20812 24800
rect 20671 24769 20683 24772
rect 20625 24763 20683 24769
rect 20806 24760 20812 24772
rect 20864 24760 20870 24812
rect 19153 24735 19211 24741
rect 19153 24701 19165 24735
rect 19199 24701 19211 24735
rect 19153 24695 19211 24701
rect 19337 24735 19395 24741
rect 19337 24701 19349 24735
rect 19383 24732 19395 24735
rect 20916 24732 20944 24840
rect 20993 24803 21051 24809
rect 20993 24769 21005 24803
rect 21039 24800 21051 24803
rect 21039 24772 21128 24800
rect 21039 24769 21051 24772
rect 20993 24763 21051 24769
rect 19383 24704 20944 24732
rect 19383 24701 19395 24704
rect 19337 24695 19395 24701
rect 17957 24667 18015 24673
rect 17957 24664 17969 24667
rect 17828 24636 17969 24664
rect 17828 24624 17834 24636
rect 17957 24633 17969 24636
rect 18003 24633 18015 24667
rect 17957 24627 18015 24633
rect 18049 24667 18107 24673
rect 18049 24633 18061 24667
rect 18095 24664 18107 24667
rect 18877 24667 18935 24673
rect 18877 24664 18889 24667
rect 18095 24636 18889 24664
rect 18095 24633 18107 24636
rect 18049 24627 18107 24633
rect 18877 24633 18889 24636
rect 18923 24633 18935 24667
rect 18877 24627 18935 24633
rect 18417 24599 18475 24605
rect 18417 24596 18429 24599
rect 17604 24568 18429 24596
rect 18417 24565 18429 24568
rect 18463 24596 18475 24599
rect 18506 24596 18512 24608
rect 18463 24568 18512 24596
rect 18463 24565 18475 24568
rect 18417 24559 18475 24565
rect 18506 24556 18512 24568
rect 18564 24556 18570 24608
rect 18598 24556 18604 24608
rect 18656 24556 18662 24608
rect 19168 24596 19196 24695
rect 19705 24599 19763 24605
rect 19705 24596 19717 24599
rect 19168 24568 19717 24596
rect 19705 24565 19717 24568
rect 19751 24596 19763 24599
rect 19794 24596 19800 24608
rect 19751 24568 19800 24596
rect 19751 24565 19763 24568
rect 19705 24559 19763 24565
rect 19794 24556 19800 24568
rect 19852 24556 19858 24608
rect 21100 24596 21128 24772
rect 21192 24732 21220 24840
rect 21818 24828 21824 24880
rect 21876 24828 21882 24880
rect 22094 24828 22100 24880
rect 22152 24828 22158 24880
rect 22186 24828 22192 24880
rect 22244 24828 22250 24880
rect 21361 24803 21419 24809
rect 21361 24769 21373 24803
rect 21407 24800 21419 24803
rect 21542 24800 21548 24812
rect 21407 24772 21548 24800
rect 21407 24769 21419 24772
rect 21361 24763 21419 24769
rect 21542 24760 21548 24772
rect 21600 24800 21606 24812
rect 22296 24800 22324 24908
rect 22833 24871 22891 24877
rect 22833 24837 22845 24871
rect 22879 24837 22891 24871
rect 23216 24868 23244 24908
rect 23658 24896 23664 24948
rect 23716 24936 23722 24948
rect 25498 24936 25504 24948
rect 23716 24908 25504 24936
rect 23716 24896 23722 24908
rect 25498 24896 25504 24908
rect 25556 24896 25562 24948
rect 26970 24896 26976 24948
rect 27028 24896 27034 24948
rect 27614 24896 27620 24948
rect 27672 24936 27678 24948
rect 27672 24908 28396 24936
rect 27672 24896 27678 24908
rect 27249 24871 27307 24877
rect 23216 24840 26556 24868
rect 22833 24831 22891 24837
rect 21600 24772 22324 24800
rect 21600 24760 21606 24772
rect 22554 24760 22560 24812
rect 22612 24760 22618 24812
rect 22650 24803 22708 24809
rect 22650 24769 22662 24803
rect 22696 24769 22708 24803
rect 22650 24763 22708 24769
rect 22373 24735 22431 24741
rect 22373 24732 22385 24735
rect 21192 24704 22385 24732
rect 22373 24701 22385 24704
rect 22419 24701 22431 24735
rect 22373 24695 22431 24701
rect 22462 24692 22468 24744
rect 22520 24732 22526 24744
rect 22665 24732 22693 24763
rect 22520 24704 22693 24732
rect 22848 24732 22876 24831
rect 26528 24812 26556 24840
rect 27249 24837 27261 24871
rect 27295 24868 27307 24871
rect 27338 24868 27344 24880
rect 27295 24840 27344 24868
rect 27295 24837 27307 24840
rect 27249 24831 27307 24837
rect 27338 24828 27344 24840
rect 27396 24828 27402 24880
rect 27430 24828 27436 24880
rect 27488 24828 27494 24880
rect 28092 24840 28304 24868
rect 22922 24760 22928 24812
rect 22980 24760 22986 24812
rect 23014 24760 23020 24812
rect 23072 24809 23078 24812
rect 23072 24800 23080 24809
rect 23072 24772 23117 24800
rect 23072 24763 23080 24772
rect 23072 24760 23078 24763
rect 26510 24760 26516 24812
rect 26568 24760 26574 24812
rect 26973 24803 27031 24809
rect 26973 24769 26985 24803
rect 27019 24800 27031 24803
rect 27448 24800 27476 24828
rect 28092 24812 28120 24840
rect 27019 24772 27476 24800
rect 27019 24769 27031 24772
rect 26973 24763 27031 24769
rect 28074 24760 28080 24812
rect 28132 24760 28138 24812
rect 28276 24809 28304 24840
rect 28169 24803 28227 24809
rect 28169 24769 28181 24803
rect 28215 24769 28227 24803
rect 28169 24763 28227 24769
rect 28261 24803 28319 24809
rect 28261 24769 28273 24803
rect 28307 24769 28319 24803
rect 28261 24763 28319 24769
rect 24670 24732 24676 24744
rect 22848 24704 24676 24732
rect 22520 24692 22526 24704
rect 24670 24692 24676 24704
rect 24728 24692 24734 24744
rect 27985 24735 28043 24741
rect 27985 24732 27997 24735
rect 24780 24704 27997 24732
rect 21266 24624 21272 24676
rect 21324 24624 21330 24676
rect 24780 24664 24808 24704
rect 27985 24701 27997 24704
rect 28031 24701 28043 24735
rect 28184 24732 28212 24763
rect 28368 24732 28396 24908
rect 28902 24896 28908 24948
rect 28960 24936 28966 24948
rect 33321 24939 33379 24945
rect 33321 24936 33333 24939
rect 28960 24908 33333 24936
rect 28960 24896 28966 24908
rect 33321 24905 33333 24908
rect 33367 24936 33379 24939
rect 33367 24908 34376 24936
rect 33367 24905 33379 24908
rect 33321 24899 33379 24905
rect 34348 24880 34376 24908
rect 35342 24896 35348 24948
rect 35400 24936 35406 24948
rect 35400 24908 35572 24936
rect 35400 24896 35406 24908
rect 28460 24840 28672 24868
rect 28460 24809 28488 24840
rect 28644 24812 28672 24840
rect 29638 24828 29644 24880
rect 29696 24868 29702 24880
rect 30006 24868 30012 24880
rect 29696 24840 30012 24868
rect 29696 24828 29702 24840
rect 30006 24828 30012 24840
rect 30064 24828 30070 24880
rect 32398 24868 32404 24880
rect 32140 24840 32404 24868
rect 28445 24803 28503 24809
rect 28445 24769 28457 24803
rect 28491 24769 28503 24803
rect 28445 24763 28503 24769
rect 28534 24760 28540 24812
rect 28592 24760 28598 24812
rect 28626 24760 28632 24812
rect 28684 24760 28690 24812
rect 28718 24760 28724 24812
rect 28776 24800 28782 24812
rect 30926 24800 30932 24812
rect 28776 24772 30932 24800
rect 28776 24760 28782 24772
rect 30926 24760 30932 24772
rect 30984 24760 30990 24812
rect 32140 24809 32168 24840
rect 32398 24828 32404 24840
rect 32456 24828 32462 24880
rect 33962 24868 33968 24880
rect 32600 24840 33968 24868
rect 32600 24809 32628 24840
rect 33962 24828 33968 24840
rect 34020 24828 34026 24880
rect 34330 24828 34336 24880
rect 34388 24828 34394 24880
rect 32125 24803 32183 24809
rect 32125 24769 32137 24803
rect 32171 24769 32183 24803
rect 32125 24763 32183 24769
rect 32309 24803 32367 24809
rect 32309 24769 32321 24803
rect 32355 24800 32367 24803
rect 32585 24803 32643 24809
rect 32585 24800 32597 24803
rect 32355 24772 32597 24800
rect 32355 24769 32367 24772
rect 32309 24763 32367 24769
rect 32585 24769 32597 24772
rect 32631 24769 32643 24803
rect 32585 24763 32643 24769
rect 32858 24760 32864 24812
rect 32916 24800 32922 24812
rect 33045 24803 33103 24809
rect 33045 24800 33057 24803
rect 32916 24772 33057 24800
rect 32916 24760 32922 24772
rect 33045 24769 33057 24772
rect 33091 24769 33103 24803
rect 33045 24763 33103 24769
rect 33134 24760 33140 24812
rect 33192 24800 33198 24812
rect 33229 24803 33287 24809
rect 33229 24800 33241 24803
rect 33192 24772 33241 24800
rect 33192 24760 33198 24772
rect 33229 24769 33241 24772
rect 33275 24769 33287 24803
rect 33229 24763 33287 24769
rect 34054 24760 34060 24812
rect 34112 24800 34118 24812
rect 35342 24809 35348 24812
rect 34149 24803 34207 24809
rect 34149 24800 34161 24803
rect 34112 24772 34161 24800
rect 34112 24760 34118 24772
rect 34149 24769 34161 24772
rect 34195 24800 34207 24803
rect 35335 24803 35348 24809
rect 35335 24800 35347 24803
rect 34195 24772 34284 24800
rect 35303 24772 35347 24800
rect 34195 24769 34207 24772
rect 34149 24763 34207 24769
rect 34256 24744 34284 24772
rect 35335 24769 35347 24772
rect 35335 24763 35348 24769
rect 35342 24760 35348 24763
rect 35400 24760 35406 24812
rect 35544 24809 35572 24908
rect 40126 24828 40132 24880
rect 40184 24828 40190 24880
rect 35529 24803 35587 24809
rect 35529 24769 35541 24803
rect 35575 24800 35587 24803
rect 35618 24800 35624 24812
rect 35575 24772 35624 24800
rect 35575 24769 35587 24772
rect 35529 24763 35587 24769
rect 35618 24760 35624 24772
rect 35676 24760 35682 24812
rect 36538 24800 36544 24812
rect 35820 24772 36544 24800
rect 30650 24732 30656 24744
rect 28184 24704 28304 24732
rect 28368 24704 30656 24732
rect 27985 24695 28043 24701
rect 21376 24636 24808 24664
rect 27065 24667 27123 24673
rect 21376 24596 21404 24636
rect 27065 24633 27077 24667
rect 27111 24664 27123 24667
rect 27111 24636 27292 24664
rect 27111 24633 27123 24636
rect 27065 24627 27123 24633
rect 27264 24608 27292 24636
rect 28276 24608 28304 24704
rect 30650 24692 30656 24704
rect 30708 24732 30714 24744
rect 31202 24732 31208 24744
rect 30708 24704 31208 24732
rect 30708 24692 30714 24704
rect 31202 24692 31208 24704
rect 31260 24692 31266 24744
rect 32030 24692 32036 24744
rect 32088 24732 32094 24744
rect 32677 24735 32735 24741
rect 32677 24732 32689 24735
rect 32088 24704 32689 24732
rect 32088 24692 32094 24704
rect 32677 24701 32689 24704
rect 32723 24701 32735 24735
rect 32677 24695 32735 24701
rect 33410 24692 33416 24744
rect 33468 24732 33474 24744
rect 33965 24735 34023 24741
rect 33965 24732 33977 24735
rect 33468 24704 33977 24732
rect 33468 24692 33474 24704
rect 33965 24701 33977 24704
rect 34011 24701 34023 24735
rect 33965 24695 34023 24701
rect 34238 24692 34244 24744
rect 34296 24692 34302 24744
rect 28442 24624 28448 24676
rect 28500 24664 28506 24676
rect 35820 24664 35848 24772
rect 36538 24760 36544 24772
rect 36596 24800 36602 24812
rect 39022 24800 39028 24812
rect 36596 24772 39028 24800
rect 36596 24760 36602 24772
rect 39022 24760 39028 24772
rect 39080 24760 39086 24812
rect 36446 24692 36452 24744
rect 36504 24732 36510 24744
rect 39298 24732 39304 24744
rect 36504 24704 39304 24732
rect 36504 24692 36510 24704
rect 39298 24692 39304 24704
rect 39356 24692 39362 24744
rect 39574 24692 39580 24744
rect 39632 24692 39638 24744
rect 39942 24692 39948 24744
rect 40000 24732 40006 24744
rect 41049 24735 41107 24741
rect 41049 24732 41061 24735
rect 40000 24704 41061 24732
rect 40000 24692 40006 24704
rect 41049 24701 41061 24704
rect 41095 24701 41107 24735
rect 41049 24695 41107 24701
rect 28500 24636 35848 24664
rect 28500 24624 28506 24636
rect 21100 24568 21404 24596
rect 21910 24556 21916 24608
rect 21968 24596 21974 24608
rect 23014 24596 23020 24608
rect 21968 24568 23020 24596
rect 21968 24556 21974 24568
rect 23014 24556 23020 24568
rect 23072 24556 23078 24608
rect 23201 24599 23259 24605
rect 23201 24565 23213 24599
rect 23247 24596 23259 24599
rect 23842 24596 23848 24608
rect 23247 24568 23848 24596
rect 23247 24565 23259 24568
rect 23201 24559 23259 24565
rect 23842 24556 23848 24568
rect 23900 24556 23906 24608
rect 24486 24556 24492 24608
rect 24544 24596 24550 24608
rect 25958 24596 25964 24608
rect 24544 24568 25964 24596
rect 24544 24556 24550 24568
rect 25958 24556 25964 24568
rect 26016 24556 26022 24608
rect 27246 24556 27252 24608
rect 27304 24556 27310 24608
rect 28258 24556 28264 24608
rect 28316 24556 28322 24608
rect 29638 24556 29644 24608
rect 29696 24596 29702 24608
rect 30834 24596 30840 24608
rect 29696 24568 30840 24596
rect 29696 24556 29702 24568
rect 30834 24556 30840 24568
rect 30892 24556 30898 24608
rect 31294 24556 31300 24608
rect 31352 24596 31358 24608
rect 32030 24596 32036 24608
rect 31352 24568 32036 24596
rect 31352 24556 31358 24568
rect 32030 24556 32036 24568
rect 32088 24556 32094 24608
rect 32122 24556 32128 24608
rect 32180 24556 32186 24608
rect 32582 24556 32588 24608
rect 32640 24556 32646 24608
rect 32858 24556 32864 24608
rect 32916 24596 32922 24608
rect 32953 24599 33011 24605
rect 32953 24596 32965 24599
rect 32916 24568 32965 24596
rect 32916 24556 32922 24568
rect 32953 24565 32965 24568
rect 32999 24565 33011 24599
rect 32953 24559 33011 24565
rect 33594 24556 33600 24608
rect 33652 24596 33658 24608
rect 34333 24599 34391 24605
rect 34333 24596 34345 24599
rect 33652 24568 34345 24596
rect 33652 24556 33658 24568
rect 34333 24565 34345 24568
rect 34379 24565 34391 24599
rect 34333 24559 34391 24565
rect 35437 24599 35495 24605
rect 35437 24565 35449 24599
rect 35483 24596 35495 24599
rect 36170 24596 36176 24608
rect 35483 24568 36176 24596
rect 35483 24565 35495 24568
rect 35437 24559 35495 24565
rect 36170 24556 36176 24568
rect 36228 24556 36234 24608
rect 1104 24506 41400 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 41400 24506
rect 1104 24432 41400 24454
rect 4890 24352 4896 24404
rect 4948 24352 4954 24404
rect 4982 24352 4988 24404
rect 5040 24352 5046 24404
rect 5074 24352 5080 24404
rect 5132 24352 5138 24404
rect 5626 24352 5632 24404
rect 5684 24352 5690 24404
rect 6822 24352 6828 24404
rect 6880 24392 6886 24404
rect 8297 24395 8355 24401
rect 6880 24364 7972 24392
rect 6880 24352 6886 24364
rect 3789 24327 3847 24333
rect 3789 24293 3801 24327
rect 3835 24293 3847 24327
rect 3789 24287 3847 24293
rect 2961 24191 3019 24197
rect 2961 24157 2973 24191
rect 3007 24188 3019 24191
rect 3804 24188 3832 24287
rect 3878 24216 3884 24268
rect 3936 24256 3942 24268
rect 4341 24259 4399 24265
rect 4341 24256 4353 24259
rect 3936 24228 4353 24256
rect 3936 24216 3942 24228
rect 4341 24225 4353 24228
rect 4387 24225 4399 24259
rect 4341 24219 4399 24225
rect 3007 24160 3832 24188
rect 4157 24191 4215 24197
rect 3007 24157 3019 24160
rect 2961 24151 3019 24157
rect 4157 24157 4169 24191
rect 4203 24188 4215 24191
rect 4706 24188 4712 24200
rect 4203 24160 4712 24188
rect 4203 24157 4215 24160
rect 4157 24151 4215 24157
rect 4706 24148 4712 24160
rect 4764 24148 4770 24200
rect 4893 24191 4951 24197
rect 4893 24157 4905 24191
rect 4939 24188 4951 24191
rect 5000 24188 5028 24352
rect 5092 24197 5120 24352
rect 5261 24327 5319 24333
rect 5261 24293 5273 24327
rect 5307 24293 5319 24327
rect 5261 24287 5319 24293
rect 7377 24327 7435 24333
rect 7377 24293 7389 24327
rect 7423 24324 7435 24327
rect 7742 24324 7748 24336
rect 7423 24296 7748 24324
rect 7423 24293 7435 24296
rect 7377 24287 7435 24293
rect 4939 24160 5028 24188
rect 5077 24191 5135 24197
rect 4939 24157 4951 24160
rect 4893 24151 4951 24157
rect 5077 24157 5089 24191
rect 5123 24157 5135 24191
rect 5077 24151 5135 24157
rect 5169 24191 5227 24197
rect 5169 24157 5181 24191
rect 5215 24188 5227 24191
rect 5276 24188 5304 24287
rect 7742 24284 7748 24296
rect 7800 24284 7806 24336
rect 7944 24324 7972 24364
rect 8297 24361 8309 24395
rect 8343 24392 8355 24395
rect 9306 24392 9312 24404
rect 8343 24364 9312 24392
rect 8343 24361 8355 24364
rect 8297 24355 8355 24361
rect 9306 24352 9312 24364
rect 9364 24352 9370 24404
rect 9490 24352 9496 24404
rect 9548 24352 9554 24404
rect 9646 24364 12112 24392
rect 9646 24324 9674 24364
rect 7944 24296 9674 24324
rect 7009 24259 7067 24265
rect 5920 24228 6960 24256
rect 5215 24160 5304 24188
rect 5215 24157 5227 24160
rect 5169 24151 5227 24157
rect 5350 24148 5356 24200
rect 5408 24188 5414 24200
rect 5920 24197 5948 24228
rect 5537 24191 5595 24197
rect 5537 24188 5549 24191
rect 5408 24160 5549 24188
rect 5408 24148 5414 24160
rect 5537 24157 5549 24160
rect 5583 24188 5595 24191
rect 5905 24191 5963 24197
rect 5905 24188 5917 24191
rect 5583 24160 5917 24188
rect 5583 24157 5595 24160
rect 5537 24151 5595 24157
rect 5905 24157 5917 24160
rect 5951 24157 5963 24191
rect 5905 24151 5963 24157
rect 6454 24148 6460 24200
rect 6512 24188 6518 24200
rect 6733 24191 6791 24197
rect 6733 24188 6745 24191
rect 6512 24160 6745 24188
rect 6512 24148 6518 24160
rect 6733 24157 6745 24160
rect 6779 24157 6791 24191
rect 6932 24188 6960 24228
rect 7009 24225 7021 24259
rect 7055 24256 7067 24259
rect 7190 24256 7196 24268
rect 7055 24228 7196 24256
rect 7055 24225 7067 24228
rect 7009 24219 7067 24225
rect 7190 24216 7196 24228
rect 7248 24216 7254 24268
rect 7944 24265 7972 24296
rect 11146 24284 11152 24336
rect 11204 24324 11210 24336
rect 12084 24324 12112 24364
rect 12250 24352 12256 24404
rect 12308 24392 12314 24404
rect 13998 24392 14004 24404
rect 12308 24364 14004 24392
rect 12308 24352 12314 24364
rect 13998 24352 14004 24364
rect 14056 24352 14062 24404
rect 14458 24352 14464 24404
rect 14516 24392 14522 24404
rect 14553 24395 14611 24401
rect 14553 24392 14565 24395
rect 14516 24364 14565 24392
rect 14516 24352 14522 24364
rect 14553 24361 14565 24364
rect 14599 24361 14611 24395
rect 14553 24355 14611 24361
rect 17310 24352 17316 24404
rect 17368 24352 17374 24404
rect 17770 24352 17776 24404
rect 17828 24352 17834 24404
rect 19334 24352 19340 24404
rect 19392 24392 19398 24404
rect 19702 24392 19708 24404
rect 19392 24364 19708 24392
rect 19392 24352 19398 24364
rect 19702 24352 19708 24364
rect 19760 24352 19766 24404
rect 21266 24352 21272 24404
rect 21324 24392 21330 24404
rect 21910 24392 21916 24404
rect 21324 24364 21916 24392
rect 21324 24352 21330 24364
rect 21910 24352 21916 24364
rect 21968 24352 21974 24404
rect 22373 24395 22431 24401
rect 22373 24361 22385 24395
rect 22419 24392 22431 24395
rect 22554 24392 22560 24404
rect 22419 24364 22560 24392
rect 22419 24361 22431 24364
rect 22373 24355 22431 24361
rect 22554 24352 22560 24364
rect 22612 24352 22618 24404
rect 23290 24352 23296 24404
rect 23348 24352 23354 24404
rect 23845 24395 23903 24401
rect 23845 24361 23857 24395
rect 23891 24392 23903 24395
rect 23891 24364 24348 24392
rect 23891 24361 23903 24364
rect 23845 24355 23903 24361
rect 12526 24324 12532 24336
rect 11204 24296 12020 24324
rect 12084 24296 12532 24324
rect 11204 24284 11210 24296
rect 7929 24259 7987 24265
rect 7929 24225 7941 24259
rect 7975 24225 7987 24259
rect 7929 24219 7987 24225
rect 8496 24228 9260 24256
rect 6932 24160 8064 24188
rect 6733 24151 6791 24157
rect 5258 24080 5264 24132
rect 5316 24080 5322 24132
rect 5626 24080 5632 24132
rect 5684 24080 5690 24132
rect 5718 24080 5724 24132
rect 5776 24080 5782 24132
rect 6914 24080 6920 24132
rect 6972 24080 6978 24132
rect 7190 24080 7196 24132
rect 7248 24120 7254 24132
rect 7650 24120 7656 24132
rect 7248 24092 7656 24120
rect 7248 24080 7254 24092
rect 7650 24080 7656 24092
rect 7708 24080 7714 24132
rect 7834 24080 7840 24132
rect 7892 24080 7898 24132
rect 2774 24012 2780 24064
rect 2832 24012 2838 24064
rect 4246 24012 4252 24064
rect 4304 24052 4310 24064
rect 5445 24055 5503 24061
rect 5445 24052 5457 24055
rect 4304 24024 5457 24052
rect 4304 24012 4310 24024
rect 5445 24021 5457 24024
rect 5491 24052 5503 24055
rect 5736 24052 5764 24080
rect 5491 24024 5764 24052
rect 5491 24021 5503 24024
rect 5445 24015 5503 24021
rect 5810 24012 5816 24064
rect 5868 24052 5874 24064
rect 6932 24052 6960 24080
rect 5868 24024 6960 24052
rect 8036 24052 8064 24160
rect 8110 24148 8116 24200
rect 8168 24188 8174 24200
rect 8496 24197 8524 24228
rect 8481 24191 8539 24197
rect 8481 24188 8493 24191
rect 8168 24160 8493 24188
rect 8168 24148 8174 24160
rect 8481 24157 8493 24160
rect 8527 24157 8539 24191
rect 8481 24151 8539 24157
rect 8573 24191 8631 24197
rect 8573 24157 8585 24191
rect 8619 24157 8631 24191
rect 8573 24151 8631 24157
rect 8294 24080 8300 24132
rect 8352 24080 8358 24132
rect 8588 24120 8616 24151
rect 8662 24148 8668 24200
rect 8720 24188 8726 24200
rect 8941 24191 8999 24197
rect 8941 24188 8953 24191
rect 8720 24160 8953 24188
rect 8720 24148 8726 24160
rect 8941 24157 8953 24160
rect 8987 24157 8999 24191
rect 8941 24151 8999 24157
rect 9030 24148 9036 24200
rect 9088 24188 9094 24200
rect 9232 24197 9260 24228
rect 9950 24216 9956 24268
rect 10008 24256 10014 24268
rect 11790 24256 11796 24268
rect 10008 24228 11796 24256
rect 10008 24216 10014 24228
rect 11790 24216 11796 24228
rect 11848 24216 11854 24268
rect 11992 24200 12020 24296
rect 12526 24284 12532 24296
rect 12584 24284 12590 24336
rect 12894 24284 12900 24336
rect 12952 24324 12958 24336
rect 13170 24324 13176 24336
rect 12952 24296 13176 24324
rect 12952 24284 12958 24296
rect 13170 24284 13176 24296
rect 13228 24284 13234 24336
rect 13630 24324 13636 24336
rect 13285 24296 13636 24324
rect 12802 24216 12808 24268
rect 12860 24216 12866 24268
rect 9125 24191 9183 24197
rect 9125 24188 9137 24191
rect 9088 24160 9137 24188
rect 9088 24148 9094 24160
rect 9125 24157 9137 24160
rect 9171 24157 9183 24191
rect 9125 24151 9183 24157
rect 9217 24191 9275 24197
rect 9217 24157 9229 24191
rect 9263 24157 9275 24191
rect 9217 24151 9275 24157
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24188 9367 24191
rect 9582 24188 9588 24200
rect 9355 24160 9588 24188
rect 9355 24157 9367 24160
rect 9309 24151 9367 24157
rect 9582 24148 9588 24160
rect 9640 24148 9646 24200
rect 10226 24148 10232 24200
rect 10284 24188 10290 24200
rect 11517 24191 11575 24197
rect 11517 24188 11529 24191
rect 10284 24160 11529 24188
rect 10284 24148 10290 24160
rect 11517 24157 11529 24160
rect 11563 24157 11575 24191
rect 11517 24151 11575 24157
rect 11974 24148 11980 24200
rect 12032 24148 12038 24200
rect 12342 24148 12348 24200
rect 12400 24188 12406 24200
rect 13081 24191 13139 24197
rect 13081 24188 13093 24191
rect 12400 24160 13093 24188
rect 12400 24148 12406 24160
rect 13081 24157 13093 24160
rect 13127 24188 13139 24191
rect 13285 24188 13313 24296
rect 13630 24284 13636 24296
rect 13688 24324 13694 24336
rect 15194 24324 15200 24336
rect 13688 24296 15200 24324
rect 13688 24284 13694 24296
rect 15194 24284 15200 24296
rect 15252 24324 15258 24336
rect 15252 24296 15700 24324
rect 15252 24284 15258 24296
rect 13127 24160 13313 24188
rect 13127 24157 13139 24160
rect 13081 24151 13139 24157
rect 13354 24148 13360 24200
rect 13412 24197 13418 24200
rect 13412 24191 13461 24197
rect 13412 24157 13415 24191
rect 13449 24157 13461 24191
rect 13412 24151 13461 24157
rect 13541 24191 13599 24197
rect 13541 24157 13553 24191
rect 13587 24157 13599 24191
rect 13541 24151 13599 24157
rect 13412 24148 13418 24151
rect 8754 24120 8760 24132
rect 8588 24092 8760 24120
rect 8588 24052 8616 24092
rect 8754 24080 8760 24092
rect 8812 24120 8818 24132
rect 13556 24120 13584 24151
rect 14366 24148 14372 24200
rect 14424 24188 14430 24200
rect 15672 24197 15700 24296
rect 17037 24259 17095 24265
rect 17037 24225 17049 24259
rect 17083 24256 17095 24259
rect 17328 24256 17356 24352
rect 17788 24256 17816 24352
rect 20898 24284 20904 24336
rect 20956 24324 20962 24336
rect 21358 24324 21364 24336
rect 20956 24296 21364 24324
rect 20956 24284 20962 24296
rect 21358 24284 21364 24296
rect 21416 24284 21422 24336
rect 23308 24324 23336 24352
rect 22940 24296 23336 24324
rect 24029 24327 24087 24333
rect 18233 24259 18291 24265
rect 18233 24256 18245 24259
rect 17083 24228 17356 24256
rect 17696 24228 18245 24256
rect 17083 24225 17095 24228
rect 17037 24219 17095 24225
rect 15473 24191 15531 24197
rect 15473 24188 15485 24191
rect 14424 24160 15485 24188
rect 14424 24148 14430 24160
rect 15473 24157 15485 24160
rect 15519 24157 15531 24191
rect 15473 24151 15531 24157
rect 15657 24191 15715 24197
rect 15657 24157 15669 24191
rect 15703 24157 15715 24191
rect 15657 24151 15715 24157
rect 15933 24191 15991 24197
rect 15933 24157 15945 24191
rect 15979 24188 15991 24191
rect 16206 24188 16212 24200
rect 15979 24160 16212 24188
rect 15979 24157 15991 24160
rect 15933 24151 15991 24157
rect 16206 24148 16212 24160
rect 16264 24188 16270 24200
rect 16482 24188 16488 24200
rect 16264 24160 16488 24188
rect 16264 24148 16270 24160
rect 16482 24148 16488 24160
rect 16540 24148 16546 24200
rect 17221 24191 17279 24197
rect 17221 24157 17233 24191
rect 17267 24188 17279 24191
rect 17696 24188 17724 24228
rect 18233 24225 18245 24228
rect 18279 24225 18291 24259
rect 18233 24219 18291 24225
rect 19889 24259 19947 24265
rect 19889 24225 19901 24259
rect 19935 24256 19947 24259
rect 20622 24256 20628 24268
rect 19935 24228 20628 24256
rect 19935 24225 19947 24228
rect 19889 24219 19947 24225
rect 20622 24216 20628 24228
rect 20680 24216 20686 24268
rect 21726 24216 21732 24268
rect 21784 24256 21790 24268
rect 21784 24228 22692 24256
rect 21784 24216 21790 24228
rect 22480 24200 22508 24228
rect 17267 24160 17724 24188
rect 17773 24191 17831 24197
rect 17267 24157 17279 24160
rect 17221 24151 17279 24157
rect 17773 24157 17785 24191
rect 17819 24188 17831 24191
rect 18138 24188 18144 24200
rect 17819 24160 18144 24188
rect 17819 24157 17831 24160
rect 17773 24151 17831 24157
rect 18138 24148 18144 24160
rect 18196 24148 18202 24200
rect 18322 24148 18328 24200
rect 18380 24148 18386 24200
rect 18693 24191 18751 24197
rect 18693 24157 18705 24191
rect 18739 24157 18751 24191
rect 18693 24151 18751 24157
rect 13998 24120 14004 24132
rect 8812 24092 14004 24120
rect 8812 24080 8818 24092
rect 13998 24080 14004 24092
rect 14056 24080 14062 24132
rect 14461 24123 14519 24129
rect 14461 24089 14473 24123
rect 14507 24120 14519 24123
rect 14642 24120 14648 24132
rect 14507 24092 14648 24120
rect 14507 24089 14519 24092
rect 14461 24083 14519 24089
rect 14642 24080 14648 24092
rect 14700 24080 14706 24132
rect 17405 24123 17463 24129
rect 15764 24092 16620 24120
rect 8036 24024 8616 24052
rect 5868 24012 5874 24024
rect 12986 24012 12992 24064
rect 13044 24052 13050 24064
rect 13725 24055 13783 24061
rect 13725 24052 13737 24055
rect 13044 24024 13737 24052
rect 13044 24012 13050 24024
rect 13725 24021 13737 24024
rect 13771 24021 13783 24055
rect 13725 24015 13783 24021
rect 15378 24012 15384 24064
rect 15436 24052 15442 24064
rect 15764 24052 15792 24092
rect 15436 24024 15792 24052
rect 15436 24012 15442 24024
rect 15838 24012 15844 24064
rect 15896 24012 15902 24064
rect 16592 24052 16620 24092
rect 17405 24089 17417 24123
rect 17451 24120 17463 24123
rect 18046 24120 18052 24132
rect 17451 24092 18052 24120
rect 17451 24089 17463 24092
rect 17405 24083 17463 24089
rect 18046 24080 18052 24092
rect 18104 24080 18110 24132
rect 18156 24120 18184 24148
rect 18708 24120 18736 24151
rect 19978 24148 19984 24200
rect 20036 24188 20042 24200
rect 20073 24191 20131 24197
rect 20073 24188 20085 24191
rect 20036 24160 20085 24188
rect 20036 24148 20042 24160
rect 20073 24157 20085 24160
rect 20119 24157 20131 24191
rect 20073 24151 20131 24157
rect 22462 24148 22468 24200
rect 22520 24148 22526 24200
rect 22664 24197 22692 24228
rect 22557 24191 22615 24197
rect 22557 24157 22569 24191
rect 22603 24157 22615 24191
rect 22557 24151 22615 24157
rect 22649 24191 22707 24197
rect 22649 24157 22661 24191
rect 22695 24157 22707 24191
rect 22649 24151 22707 24157
rect 18156 24092 18736 24120
rect 19794 24080 19800 24132
rect 19852 24120 19858 24132
rect 22572 24120 22600 24151
rect 22738 24148 22744 24200
rect 22796 24188 22802 24200
rect 22940 24197 22968 24296
rect 24029 24293 24041 24327
rect 24075 24293 24087 24327
rect 24029 24287 24087 24293
rect 23290 24216 23296 24268
rect 23348 24216 23354 24268
rect 22833 24191 22891 24197
rect 22833 24188 22845 24191
rect 22796 24160 22845 24188
rect 22796 24148 22802 24160
rect 22833 24157 22845 24160
rect 22879 24157 22891 24191
rect 22833 24151 22891 24157
rect 22925 24191 22983 24197
rect 22925 24157 22937 24191
rect 22971 24188 22983 24191
rect 23014 24188 23020 24200
rect 22971 24160 23020 24188
rect 22971 24157 22983 24160
rect 22925 24151 22983 24157
rect 23014 24148 23020 24160
rect 23072 24148 23078 24200
rect 23109 24191 23167 24197
rect 23109 24157 23121 24191
rect 23155 24188 23167 24191
rect 24044 24188 24072 24287
rect 23155 24160 24072 24188
rect 24320 24188 24348 24364
rect 24394 24352 24400 24404
rect 24452 24352 24458 24404
rect 24946 24352 24952 24404
rect 25004 24352 25010 24404
rect 25130 24352 25136 24404
rect 25188 24392 25194 24404
rect 25406 24392 25412 24404
rect 25188 24364 25412 24392
rect 25188 24352 25194 24364
rect 25406 24352 25412 24364
rect 25464 24392 25470 24404
rect 25685 24395 25743 24401
rect 25685 24392 25697 24395
rect 25464 24364 25697 24392
rect 25464 24352 25470 24364
rect 25685 24361 25697 24364
rect 25731 24361 25743 24395
rect 25685 24355 25743 24361
rect 27430 24352 27436 24404
rect 27488 24392 27494 24404
rect 27893 24395 27951 24401
rect 27893 24392 27905 24395
rect 27488 24364 27905 24392
rect 27488 24352 27494 24364
rect 27893 24361 27905 24364
rect 27939 24361 27951 24395
rect 27893 24355 27951 24361
rect 28534 24352 28540 24404
rect 28592 24392 28598 24404
rect 28721 24395 28779 24401
rect 28721 24392 28733 24395
rect 28592 24364 28733 24392
rect 28592 24352 28598 24364
rect 28721 24361 28733 24364
rect 28767 24361 28779 24395
rect 28721 24355 28779 24361
rect 28810 24352 28816 24404
rect 28868 24392 28874 24404
rect 29638 24392 29644 24404
rect 28868 24364 29644 24392
rect 28868 24352 28874 24364
rect 29638 24352 29644 24364
rect 29696 24352 29702 24404
rect 29917 24395 29975 24401
rect 29917 24361 29929 24395
rect 29963 24392 29975 24395
rect 30006 24392 30012 24404
rect 29963 24364 30012 24392
rect 29963 24361 29975 24364
rect 29917 24355 29975 24361
rect 30006 24352 30012 24364
rect 30064 24352 30070 24404
rect 31478 24352 31484 24404
rect 31536 24352 31542 24404
rect 31757 24395 31815 24401
rect 31757 24361 31769 24395
rect 31803 24392 31815 24395
rect 31846 24392 31852 24404
rect 31803 24364 31852 24392
rect 31803 24361 31815 24364
rect 31757 24355 31815 24361
rect 31846 24352 31852 24364
rect 31904 24352 31910 24404
rect 32490 24352 32496 24404
rect 32548 24392 32554 24404
rect 33594 24392 33600 24404
rect 32548 24364 33600 24392
rect 32548 24352 32554 24364
rect 33594 24352 33600 24364
rect 33652 24352 33658 24404
rect 35342 24392 35348 24404
rect 34164 24364 35348 24392
rect 34164 24336 34192 24364
rect 35342 24352 35348 24364
rect 35400 24392 35406 24404
rect 35526 24392 35532 24404
rect 35400 24364 35532 24392
rect 35400 24352 35406 24364
rect 35526 24352 35532 24364
rect 35584 24352 35590 24404
rect 38286 24352 38292 24404
rect 38344 24352 38350 24404
rect 39574 24352 39580 24404
rect 39632 24392 39638 24404
rect 40129 24395 40187 24401
rect 40129 24392 40141 24395
rect 39632 24364 40141 24392
rect 39632 24352 39638 24364
rect 40129 24361 40141 24364
rect 40175 24361 40187 24395
rect 40129 24355 40187 24361
rect 25869 24327 25927 24333
rect 25869 24324 25881 24327
rect 24596 24296 25881 24324
rect 24596 24268 24624 24296
rect 25869 24293 25881 24296
rect 25915 24293 25927 24327
rect 25869 24287 25927 24293
rect 27341 24327 27399 24333
rect 27341 24293 27353 24327
rect 27387 24324 27399 24327
rect 27614 24324 27620 24336
rect 27387 24296 27620 24324
rect 27387 24293 27399 24296
rect 27341 24287 27399 24293
rect 27614 24284 27620 24296
rect 27672 24284 27678 24336
rect 28169 24327 28227 24333
rect 28169 24293 28181 24327
rect 28215 24324 28227 24327
rect 28258 24324 28264 24336
rect 28215 24296 28264 24324
rect 28215 24293 28227 24296
rect 28169 24287 28227 24293
rect 28258 24284 28264 24296
rect 28316 24324 28322 24336
rect 30285 24327 30343 24333
rect 30285 24324 30297 24327
rect 28316 24296 30297 24324
rect 28316 24284 28322 24296
rect 30285 24293 30297 24296
rect 30331 24293 30343 24327
rect 30285 24287 30343 24293
rect 30834 24284 30840 24336
rect 30892 24284 30898 24336
rect 30929 24327 30987 24333
rect 30929 24293 30941 24327
rect 30975 24324 30987 24327
rect 32214 24324 32220 24336
rect 30975 24296 32220 24324
rect 30975 24293 30987 24296
rect 30929 24287 30987 24293
rect 32214 24284 32220 24296
rect 32272 24284 32278 24336
rect 33502 24284 33508 24336
rect 33560 24284 33566 24336
rect 33870 24284 33876 24336
rect 33928 24324 33934 24336
rect 34057 24327 34115 24333
rect 34057 24324 34069 24327
rect 33928 24296 34069 24324
rect 33928 24284 33934 24296
rect 34057 24293 34069 24296
rect 34103 24293 34115 24327
rect 34057 24287 34115 24293
rect 34146 24284 34152 24336
rect 34204 24284 34210 24336
rect 38304 24324 38332 24352
rect 35084 24296 38332 24324
rect 24578 24216 24584 24268
rect 24636 24216 24642 24268
rect 25317 24259 25375 24265
rect 25317 24256 25329 24259
rect 24964 24228 25329 24256
rect 24964 24200 24992 24228
rect 25317 24225 25329 24228
rect 25363 24225 25375 24259
rect 25317 24219 25375 24225
rect 25409 24259 25467 24265
rect 25409 24225 25421 24259
rect 25455 24256 25467 24259
rect 25958 24256 25964 24268
rect 25455 24228 25964 24256
rect 25455 24225 25467 24228
rect 25409 24219 25467 24225
rect 25958 24216 25964 24228
rect 26016 24216 26022 24268
rect 27249 24259 27307 24265
rect 27249 24225 27261 24259
rect 27295 24256 27307 24259
rect 28718 24256 28724 24268
rect 27295 24228 28724 24256
rect 27295 24225 27307 24228
rect 27249 24219 27307 24225
rect 28718 24216 28724 24228
rect 28776 24216 28782 24268
rect 29089 24259 29147 24265
rect 29089 24225 29101 24259
rect 29135 24256 29147 24259
rect 30852 24256 30880 24284
rect 29135 24228 29776 24256
rect 30852 24228 31616 24256
rect 29135 24225 29147 24228
rect 29089 24219 29147 24225
rect 29748 24200 29776 24228
rect 24320 24160 24624 24188
rect 23155 24157 23167 24160
rect 23109 24151 23167 24157
rect 23290 24120 23296 24132
rect 19852 24092 20392 24120
rect 22572 24092 23296 24120
rect 19852 24080 19858 24092
rect 17494 24052 17500 24064
rect 16592 24024 17500 24052
rect 17494 24012 17500 24024
rect 17552 24052 17558 24064
rect 17589 24055 17647 24061
rect 17589 24052 17601 24055
rect 17552 24024 17601 24052
rect 17552 24012 17558 24024
rect 17589 24021 17601 24024
rect 17635 24021 17647 24055
rect 17589 24015 17647 24021
rect 17678 24012 17684 24064
rect 17736 24052 17742 24064
rect 18877 24055 18935 24061
rect 18877 24052 18889 24055
rect 17736 24024 18889 24052
rect 17736 24012 17742 24024
rect 18877 24021 18889 24024
rect 18923 24021 18935 24055
rect 18877 24015 18935 24021
rect 20254 24012 20260 24064
rect 20312 24012 20318 24064
rect 20364 24052 20392 24092
rect 23290 24080 23296 24092
rect 23348 24080 23354 24132
rect 23658 24080 23664 24132
rect 23716 24080 23722 24132
rect 23768 24092 24164 24120
rect 23768 24052 23796 24092
rect 20364 24024 23796 24052
rect 23842 24012 23848 24064
rect 23900 24061 23906 24064
rect 23900 24055 23919 24061
rect 23907 24021 23919 24055
rect 24136 24052 24164 24092
rect 24394 24080 24400 24132
rect 24452 24080 24458 24132
rect 24596 24120 24624 24160
rect 24670 24148 24676 24200
rect 24728 24148 24734 24200
rect 24946 24148 24952 24200
rect 25004 24148 25010 24200
rect 25133 24191 25191 24197
rect 25133 24157 25145 24191
rect 25179 24188 25191 24191
rect 25179 24160 26372 24188
rect 25179 24157 25191 24160
rect 25133 24151 25191 24157
rect 25332 24132 25360 24160
rect 25222 24120 25228 24132
rect 24596 24092 25228 24120
rect 25222 24080 25228 24092
rect 25280 24080 25286 24132
rect 25314 24080 25320 24132
rect 25372 24080 25378 24132
rect 25498 24080 25504 24132
rect 25556 24080 25562 24132
rect 25682 24080 25688 24132
rect 25740 24129 25746 24132
rect 25740 24123 25759 24129
rect 25747 24089 25759 24123
rect 25740 24083 25759 24089
rect 25740 24080 25746 24083
rect 26050 24080 26056 24132
rect 26108 24080 26114 24132
rect 26344 24120 26372 24160
rect 26970 24148 26976 24200
rect 27028 24188 27034 24200
rect 27157 24191 27215 24197
rect 27157 24188 27169 24191
rect 27028 24160 27169 24188
rect 27028 24148 27034 24160
rect 27157 24157 27169 24160
rect 27203 24157 27215 24191
rect 27157 24151 27215 24157
rect 27422 24191 27480 24197
rect 27422 24157 27434 24191
rect 27468 24188 27480 24191
rect 27522 24188 27528 24200
rect 27468 24160 27528 24188
rect 27468 24157 27480 24160
rect 27422 24151 27480 24157
rect 27522 24148 27528 24160
rect 27580 24148 27586 24200
rect 27614 24148 27620 24200
rect 27672 24148 27678 24200
rect 27890 24148 27896 24200
rect 27948 24148 27954 24200
rect 28077 24191 28135 24197
rect 28077 24157 28089 24191
rect 28123 24188 28135 24191
rect 28166 24188 28172 24200
rect 28123 24160 28172 24188
rect 28123 24157 28135 24160
rect 28077 24151 28135 24157
rect 28166 24148 28172 24160
rect 28224 24148 28230 24200
rect 28258 24148 28264 24200
rect 28316 24148 28322 24200
rect 28353 24191 28411 24197
rect 28353 24157 28365 24191
rect 28399 24157 28411 24191
rect 28353 24151 28411 24157
rect 27908 24120 27936 24148
rect 28368 24120 28396 24151
rect 28442 24148 28448 24200
rect 28500 24148 28506 24200
rect 28905 24191 28963 24197
rect 28905 24157 28917 24191
rect 28951 24157 28963 24191
rect 28905 24151 28963 24157
rect 29181 24191 29239 24197
rect 29181 24157 29193 24191
rect 29227 24188 29239 24191
rect 29454 24188 29460 24200
rect 29227 24160 29460 24188
rect 29227 24157 29239 24160
rect 29181 24151 29239 24157
rect 26344 24092 28396 24120
rect 28460 24120 28488 24148
rect 28920 24120 28948 24151
rect 29454 24148 29460 24160
rect 29512 24148 29518 24200
rect 29730 24148 29736 24200
rect 29788 24148 29794 24200
rect 30009 24191 30067 24197
rect 30009 24157 30021 24191
rect 30055 24157 30067 24191
rect 30009 24151 30067 24157
rect 28460 24092 28948 24120
rect 29086 24080 29092 24132
rect 29144 24080 29150 24132
rect 29825 24123 29883 24129
rect 29825 24089 29837 24123
rect 29871 24089 29883 24123
rect 30024 24120 30052 24151
rect 30098 24148 30104 24200
rect 30156 24148 30162 24200
rect 30282 24148 30288 24200
rect 30340 24148 30346 24200
rect 30374 24148 30380 24200
rect 30432 24148 30438 24200
rect 30745 24191 30803 24197
rect 30745 24157 30757 24191
rect 30791 24188 30803 24191
rect 30834 24188 30840 24200
rect 30791 24160 30840 24188
rect 30791 24157 30803 24160
rect 30745 24151 30803 24157
rect 30834 24148 30840 24160
rect 30892 24148 30898 24200
rect 31021 24191 31079 24197
rect 31021 24157 31033 24191
rect 31067 24188 31079 24191
rect 31067 24160 31432 24188
rect 31067 24157 31079 24160
rect 31021 24151 31079 24157
rect 30300 24120 30328 24148
rect 30024 24092 30328 24120
rect 30392 24120 30420 24148
rect 31036 24120 31064 24151
rect 30392 24092 31064 24120
rect 29825 24083 29883 24089
rect 24857 24055 24915 24061
rect 24857 24052 24869 24055
rect 24136 24024 24869 24052
rect 23900 24015 23919 24021
rect 24857 24021 24869 24024
rect 24903 24021 24915 24055
rect 25516 24052 25544 24080
rect 26068 24052 26096 24080
rect 25516 24024 26096 24052
rect 24857 24015 24915 24021
rect 23900 24012 23906 24015
rect 26142 24012 26148 24064
rect 26200 24052 26206 24064
rect 26694 24052 26700 24064
rect 26200 24024 26700 24052
rect 26200 24012 26206 24024
rect 26694 24012 26700 24024
rect 26752 24012 26758 24064
rect 26973 24055 27031 24061
rect 26973 24021 26985 24055
rect 27019 24052 27031 24055
rect 27246 24052 27252 24064
rect 27019 24024 27252 24052
rect 27019 24021 27031 24024
rect 26973 24015 27031 24021
rect 27246 24012 27252 24024
rect 27304 24012 27310 24064
rect 27338 24012 27344 24064
rect 27396 24052 27402 24064
rect 27709 24055 27767 24061
rect 27709 24052 27721 24055
rect 27396 24024 27721 24052
rect 27396 24012 27402 24024
rect 27709 24021 27721 24024
rect 27755 24021 27767 24055
rect 27709 24015 27767 24021
rect 28350 24012 28356 24064
rect 28408 24052 28414 24064
rect 29104 24052 29132 24080
rect 28408 24024 29132 24052
rect 29840 24052 29868 24083
rect 31294 24080 31300 24132
rect 31352 24080 31358 24132
rect 31404 24120 31432 24160
rect 31478 24148 31484 24200
rect 31536 24148 31542 24200
rect 31588 24197 31616 24228
rect 33318 24216 33324 24268
rect 33376 24256 33382 24268
rect 34241 24259 34299 24265
rect 34241 24256 34253 24259
rect 33376 24228 34253 24256
rect 33376 24216 33382 24228
rect 34241 24225 34253 24228
rect 34287 24225 34299 24259
rect 35084 24256 35112 24296
rect 34241 24219 34299 24225
rect 34808 24228 35112 24256
rect 31573 24191 31631 24197
rect 31573 24157 31585 24191
rect 31619 24157 31631 24191
rect 31573 24151 31631 24157
rect 32858 24148 32864 24200
rect 32916 24148 32922 24200
rect 33505 24191 33563 24197
rect 33505 24157 33517 24191
rect 33551 24157 33563 24191
rect 33505 24151 33563 24157
rect 32876 24120 32904 24148
rect 31404 24092 32904 24120
rect 29914 24052 29920 24064
rect 29840 24024 29920 24052
rect 28408 24012 28414 24024
rect 29914 24012 29920 24024
rect 29972 24052 29978 24064
rect 30098 24052 30104 24064
rect 29972 24024 30104 24052
rect 29972 24012 29978 24024
rect 30098 24012 30104 24024
rect 30156 24012 30162 24064
rect 30374 24012 30380 24064
rect 30432 24052 30438 24064
rect 30561 24055 30619 24061
rect 30561 24052 30573 24055
rect 30432 24024 30573 24052
rect 30432 24012 30438 24024
rect 30561 24021 30573 24024
rect 30607 24021 30619 24055
rect 30561 24015 30619 24021
rect 32490 24012 32496 24064
rect 32548 24052 32554 24064
rect 33226 24052 33232 24064
rect 32548 24024 33232 24052
rect 32548 24012 32554 24024
rect 33226 24012 33232 24024
rect 33284 24012 33290 24064
rect 33520 24052 33548 24151
rect 33962 24148 33968 24200
rect 34020 24188 34026 24200
rect 34808 24188 34836 24228
rect 35084 24197 35112 24228
rect 37550 24216 37556 24268
rect 37608 24216 37614 24268
rect 38304 24256 38332 24296
rect 38304 24228 38516 24256
rect 34020 24160 34836 24188
rect 34885 24191 34943 24197
rect 34020 24148 34026 24160
rect 34885 24157 34897 24191
rect 34931 24157 34943 24191
rect 34885 24151 34943 24157
rect 35069 24191 35127 24197
rect 35069 24157 35081 24191
rect 35115 24157 35127 24191
rect 35069 24151 35127 24157
rect 33873 24123 33931 24129
rect 33873 24089 33885 24123
rect 33919 24120 33931 24123
rect 34241 24123 34299 24129
rect 34241 24120 34253 24123
rect 33919 24092 34253 24120
rect 33919 24089 33931 24092
rect 33873 24083 33931 24089
rect 34241 24089 34253 24092
rect 34287 24089 34299 24123
rect 34241 24083 34299 24089
rect 34422 24080 34428 24132
rect 34480 24120 34486 24132
rect 34900 24120 34928 24151
rect 37274 24148 37280 24200
rect 37332 24188 37338 24200
rect 37645 24191 37703 24197
rect 37645 24188 37657 24191
rect 37332 24160 37657 24188
rect 37332 24148 37338 24160
rect 37645 24157 37657 24160
rect 37691 24188 37703 24191
rect 37734 24188 37740 24200
rect 37691 24160 37740 24188
rect 37691 24157 37703 24160
rect 37645 24151 37703 24157
rect 37734 24148 37740 24160
rect 37792 24148 37798 24200
rect 37826 24148 37832 24200
rect 37884 24188 37890 24200
rect 38289 24191 38347 24197
rect 38289 24188 38301 24191
rect 37884 24160 38301 24188
rect 37884 24148 37890 24160
rect 38289 24157 38301 24160
rect 38335 24188 38347 24191
rect 38378 24188 38384 24200
rect 38335 24160 38384 24188
rect 38335 24157 38347 24160
rect 38289 24151 38347 24157
rect 38378 24148 38384 24160
rect 38436 24148 38442 24200
rect 38488 24197 38516 24228
rect 38473 24191 38531 24197
rect 38473 24157 38485 24191
rect 38519 24157 38531 24191
rect 38473 24151 38531 24157
rect 40310 24148 40316 24200
rect 40368 24148 40374 24200
rect 35158 24120 35164 24132
rect 34480 24092 35164 24120
rect 34480 24080 34486 24092
rect 35158 24080 35164 24092
rect 35216 24080 35222 24132
rect 36722 24080 36728 24132
rect 36780 24120 36786 24132
rect 37921 24123 37979 24129
rect 37921 24120 37933 24123
rect 36780 24092 37933 24120
rect 36780 24080 36786 24092
rect 37921 24089 37933 24092
rect 37967 24089 37979 24123
rect 37921 24083 37979 24089
rect 38013 24123 38071 24129
rect 38013 24089 38025 24123
rect 38059 24120 38071 24123
rect 38654 24120 38660 24132
rect 38059 24092 38660 24120
rect 38059 24089 38071 24092
rect 38013 24083 38071 24089
rect 38654 24080 38660 24092
rect 38712 24080 38718 24132
rect 34977 24055 35035 24061
rect 34977 24052 34989 24055
rect 33520 24024 34989 24052
rect 34977 24021 34989 24024
rect 35023 24052 35035 24055
rect 35986 24052 35992 24064
rect 35023 24024 35992 24052
rect 35023 24021 35035 24024
rect 34977 24015 35035 24021
rect 35986 24012 35992 24024
rect 36044 24012 36050 24064
rect 37366 24012 37372 24064
rect 37424 24012 37430 24064
rect 38381 24055 38439 24061
rect 38381 24021 38393 24055
rect 38427 24052 38439 24055
rect 38470 24052 38476 24064
rect 38427 24024 38476 24052
rect 38427 24021 38439 24024
rect 38381 24015 38439 24021
rect 38470 24012 38476 24024
rect 38528 24012 38534 24064
rect 1104 23962 41400 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 41400 23962
rect 1104 23888 41400 23910
rect 2774 23848 2780 23860
rect 2700 23820 2780 23848
rect 2700 23789 2728 23820
rect 2774 23808 2780 23820
rect 2832 23808 2838 23860
rect 3050 23808 3056 23860
rect 3108 23808 3114 23860
rect 4062 23808 4068 23860
rect 4120 23848 4126 23860
rect 5810 23848 5816 23860
rect 4120 23820 5816 23848
rect 4120 23808 4126 23820
rect 5810 23808 5816 23820
rect 5868 23808 5874 23860
rect 7190 23808 7196 23860
rect 7248 23808 7254 23860
rect 8846 23848 8852 23860
rect 7576 23820 8852 23848
rect 2685 23783 2743 23789
rect 2685 23749 2697 23783
rect 2731 23749 2743 23783
rect 3068 23780 3096 23808
rect 3068 23752 3174 23780
rect 2685 23743 2743 23749
rect 4246 23740 4252 23792
rect 4304 23740 4310 23792
rect 5258 23740 5264 23792
rect 5316 23780 5322 23792
rect 5534 23780 5540 23792
rect 5316 23752 5540 23780
rect 5316 23740 5322 23752
rect 5534 23740 5540 23752
rect 5592 23740 5598 23792
rect 2406 23604 2412 23656
rect 2464 23604 2470 23656
rect 4157 23647 4215 23653
rect 4157 23613 4169 23647
rect 4203 23644 4215 23647
rect 4264 23644 4292 23740
rect 7374 23672 7380 23724
rect 7432 23672 7438 23724
rect 7576 23721 7604 23820
rect 8846 23808 8852 23820
rect 8904 23808 8910 23860
rect 9141 23820 9352 23848
rect 9141 23780 9169 23820
rect 7668 23752 9169 23780
rect 9324 23780 9352 23820
rect 9490 23808 9496 23860
rect 9548 23848 9554 23860
rect 9950 23848 9956 23860
rect 9548 23820 9956 23848
rect 9548 23808 9554 23820
rect 9950 23808 9956 23820
rect 10008 23808 10014 23860
rect 10045 23851 10103 23857
rect 10045 23817 10057 23851
rect 10091 23848 10103 23851
rect 11054 23848 11060 23860
rect 10091 23820 11060 23848
rect 10091 23817 10103 23820
rect 10045 23811 10103 23817
rect 11054 23808 11060 23820
rect 11112 23808 11118 23860
rect 12621 23851 12679 23857
rect 12621 23817 12633 23851
rect 12667 23848 12679 23851
rect 13078 23848 13084 23860
rect 12667 23820 13084 23848
rect 12667 23817 12679 23820
rect 12621 23811 12679 23817
rect 13078 23808 13084 23820
rect 13136 23808 13142 23860
rect 13630 23808 13636 23860
rect 13688 23848 13694 23860
rect 13688 23820 14688 23848
rect 13688 23808 13694 23820
rect 9324 23752 14412 23780
rect 7668 23721 7696 23752
rect 7561 23715 7619 23721
rect 7561 23681 7573 23715
rect 7607 23681 7619 23715
rect 7561 23675 7619 23681
rect 7653 23715 7711 23721
rect 7653 23681 7665 23715
rect 7699 23681 7711 23715
rect 7653 23675 7711 23681
rect 8478 23672 8484 23724
rect 8536 23672 8542 23724
rect 9030 23672 9036 23724
rect 9088 23672 9094 23724
rect 9126 23715 9184 23721
rect 9126 23681 9138 23715
rect 9172 23681 9184 23715
rect 9126 23675 9184 23681
rect 9309 23715 9367 23721
rect 9309 23681 9321 23715
rect 9355 23681 9367 23715
rect 9309 23675 9367 23681
rect 4203 23616 4292 23644
rect 8496 23644 8524 23672
rect 9141 23644 9169 23675
rect 8496 23616 9169 23644
rect 9324 23644 9352 23675
rect 9398 23672 9404 23724
rect 9456 23672 9462 23724
rect 9582 23721 9588 23724
rect 9539 23715 9588 23721
rect 9539 23681 9551 23715
rect 9585 23681 9588 23715
rect 9539 23675 9588 23681
rect 9582 23672 9588 23675
rect 9640 23672 9646 23724
rect 9674 23672 9680 23724
rect 9732 23712 9738 23724
rect 10229 23715 10287 23721
rect 10229 23712 10241 23715
rect 9732 23684 10241 23712
rect 9732 23672 9738 23684
rect 10229 23681 10241 23684
rect 10275 23681 10287 23715
rect 10229 23675 10287 23681
rect 10413 23715 10471 23721
rect 10413 23681 10425 23715
rect 10459 23712 10471 23715
rect 10502 23712 10508 23724
rect 10459 23684 10508 23712
rect 10459 23681 10471 23684
rect 10413 23675 10471 23681
rect 10502 23672 10508 23684
rect 10560 23672 10566 23724
rect 12820 23721 12848 23752
rect 14384 23724 14412 23752
rect 14550 23740 14556 23792
rect 14608 23740 14614 23792
rect 10781 23715 10839 23721
rect 10781 23681 10793 23715
rect 10827 23712 10839 23715
rect 10965 23715 11023 23721
rect 10827 23684 10916 23712
rect 10827 23681 10839 23684
rect 10781 23675 10839 23681
rect 9953 23647 10011 23653
rect 9953 23644 9965 23647
rect 9324 23616 9536 23644
rect 4203 23613 4215 23616
rect 4157 23607 4215 23613
rect 9508 23588 9536 23616
rect 9692 23616 9965 23644
rect 7466 23536 7472 23588
rect 7524 23536 7530 23588
rect 9490 23536 9496 23588
rect 9548 23536 9554 23588
rect 9692 23585 9720 23616
rect 9953 23613 9965 23616
rect 9999 23613 10011 23647
rect 9953 23607 10011 23613
rect 9677 23579 9735 23585
rect 9677 23545 9689 23579
rect 9723 23545 9735 23579
rect 9677 23539 9735 23545
rect 7098 23468 7104 23520
rect 7156 23508 7162 23520
rect 10888 23508 10916 23684
rect 10965 23681 10977 23715
rect 11011 23712 11023 23715
rect 12805 23715 12863 23721
rect 11011 23684 11284 23712
rect 11011 23681 11023 23684
rect 10965 23675 11023 23681
rect 11256 23656 11284 23684
rect 12805 23681 12817 23715
rect 12851 23681 12863 23715
rect 12805 23675 12863 23681
rect 12986 23672 12992 23724
rect 13044 23672 13050 23724
rect 13078 23672 13084 23724
rect 13136 23721 13142 23724
rect 13136 23715 13151 23721
rect 13139 23681 13151 23715
rect 13136 23675 13151 23681
rect 13136 23672 13142 23675
rect 14366 23672 14372 23724
rect 14424 23672 14430 23724
rect 14458 23672 14464 23724
rect 14516 23672 14522 23724
rect 14660 23721 14688 23820
rect 15010 23808 15016 23860
rect 15068 23848 15074 23860
rect 15068 23820 17080 23848
rect 15068 23808 15074 23820
rect 15378 23780 15384 23792
rect 14752 23752 15384 23780
rect 14645 23715 14703 23721
rect 14645 23681 14657 23715
rect 14691 23681 14703 23715
rect 14645 23675 14703 23681
rect 11238 23604 11244 23656
rect 11296 23604 11302 23656
rect 12158 23536 12164 23588
rect 12216 23576 12222 23588
rect 13814 23576 13820 23588
rect 12216 23548 13820 23576
rect 12216 23536 12222 23548
rect 13814 23536 13820 23548
rect 13872 23576 13878 23588
rect 14752 23576 14780 23752
rect 15378 23740 15384 23752
rect 15436 23740 15442 23792
rect 15654 23740 15660 23792
rect 15712 23780 15718 23792
rect 16945 23783 17003 23789
rect 16945 23780 16957 23783
rect 15712 23752 16957 23780
rect 15712 23740 15718 23752
rect 16945 23749 16957 23752
rect 16991 23749 17003 23783
rect 16945 23743 17003 23749
rect 15102 23672 15108 23724
rect 15160 23672 15166 23724
rect 15470 23672 15476 23724
rect 15528 23672 15534 23724
rect 15838 23672 15844 23724
rect 15896 23672 15902 23724
rect 16574 23672 16580 23724
rect 16632 23712 16638 23724
rect 17052 23721 17080 23820
rect 17310 23808 17316 23860
rect 17368 23848 17374 23860
rect 18322 23848 18328 23860
rect 17368 23820 17540 23848
rect 17368 23808 17374 23820
rect 17512 23789 17540 23820
rect 18064 23820 18328 23848
rect 17497 23783 17555 23789
rect 17497 23749 17509 23783
rect 17543 23749 17555 23783
rect 17497 23743 17555 23749
rect 16669 23715 16727 23721
rect 16669 23712 16681 23715
rect 16632 23684 16681 23712
rect 16632 23672 16638 23684
rect 16669 23681 16681 23684
rect 16715 23681 16727 23715
rect 16669 23675 16727 23681
rect 16853 23715 16911 23721
rect 16853 23681 16865 23715
rect 16899 23681 16911 23715
rect 16853 23675 16911 23681
rect 17037 23715 17095 23721
rect 17037 23681 17049 23715
rect 17083 23712 17095 23715
rect 17678 23712 17684 23724
rect 17083 23684 17684 23712
rect 17083 23681 17095 23684
rect 17037 23675 17095 23681
rect 13872 23548 14780 23576
rect 16868 23644 16896 23675
rect 17678 23672 17684 23684
rect 17736 23672 17742 23724
rect 18064 23644 18092 23820
rect 18322 23808 18328 23820
rect 18380 23808 18386 23860
rect 18598 23808 18604 23860
rect 18656 23808 18662 23860
rect 20162 23808 20168 23860
rect 20220 23808 20226 23860
rect 20438 23808 20444 23860
rect 20496 23848 20502 23860
rect 20625 23851 20683 23857
rect 20625 23848 20637 23851
rect 20496 23820 20637 23848
rect 20496 23808 20502 23820
rect 20625 23817 20637 23820
rect 20671 23817 20683 23851
rect 20625 23811 20683 23817
rect 20714 23808 20720 23860
rect 20772 23808 20778 23860
rect 21266 23848 21272 23860
rect 21100 23820 21272 23848
rect 18233 23783 18291 23789
rect 18233 23749 18245 23783
rect 18279 23780 18291 23783
rect 18616 23780 18644 23808
rect 18279 23752 18644 23780
rect 20180 23780 20208 23808
rect 20901 23783 20959 23789
rect 20901 23780 20913 23783
rect 20180 23752 20913 23780
rect 18279 23749 18291 23752
rect 18233 23743 18291 23749
rect 20901 23749 20913 23752
rect 20947 23749 20959 23783
rect 20901 23743 20959 23749
rect 21100 23721 21128 23820
rect 21266 23808 21272 23820
rect 21324 23808 21330 23860
rect 21450 23808 21456 23860
rect 21508 23808 21514 23860
rect 21726 23808 21732 23860
rect 21784 23848 21790 23860
rect 22922 23848 22928 23860
rect 21784 23820 22928 23848
rect 21784 23808 21790 23820
rect 22922 23808 22928 23820
rect 22980 23848 22986 23860
rect 22980 23820 24992 23848
rect 22980 23808 22986 23820
rect 21468 23780 21496 23808
rect 21192 23752 21496 23780
rect 21192 23724 21220 23752
rect 21818 23740 21824 23792
rect 21876 23780 21882 23792
rect 23474 23780 23480 23792
rect 21876 23752 23480 23780
rect 21876 23740 21882 23752
rect 20257 23715 20315 23721
rect 20257 23681 20269 23715
rect 20303 23712 20315 23715
rect 21085 23715 21143 23721
rect 20303 23684 20392 23712
rect 20303 23681 20315 23684
rect 20257 23675 20315 23681
rect 16868 23616 18092 23644
rect 13872 23536 13878 23548
rect 7156 23480 10916 23508
rect 7156 23468 7162 23480
rect 12710 23468 12716 23520
rect 12768 23508 12774 23520
rect 16868 23508 16896 23616
rect 17494 23536 17500 23588
rect 17552 23536 17558 23588
rect 17770 23536 17776 23588
rect 17828 23536 17834 23588
rect 17954 23536 17960 23588
rect 18012 23536 18018 23588
rect 20162 23536 20168 23588
rect 20220 23576 20226 23588
rect 20364 23576 20392 23684
rect 21085 23681 21097 23715
rect 21131 23681 21143 23715
rect 21085 23675 21143 23681
rect 21174 23672 21180 23724
rect 21232 23672 21238 23724
rect 21358 23672 21364 23724
rect 21416 23672 21422 23724
rect 22204 23721 22232 23752
rect 23474 23740 23480 23752
rect 23532 23780 23538 23792
rect 24964 23780 24992 23820
rect 25222 23808 25228 23860
rect 25280 23848 25286 23860
rect 26513 23851 26571 23857
rect 26513 23848 26525 23851
rect 25280 23820 26525 23848
rect 25280 23808 25286 23820
rect 26513 23817 26525 23820
rect 26559 23817 26571 23851
rect 26513 23811 26571 23817
rect 26602 23808 26608 23860
rect 26660 23848 26666 23860
rect 28166 23848 28172 23860
rect 26660 23820 27384 23848
rect 26660 23808 26666 23820
rect 23532 23752 23888 23780
rect 23532 23740 23538 23752
rect 23860 23724 23888 23752
rect 24504 23752 24716 23780
rect 24504 23724 24532 23752
rect 21453 23715 21511 23721
rect 21453 23681 21465 23715
rect 21499 23712 21511 23715
rect 22005 23715 22063 23721
rect 22005 23712 22017 23715
rect 21499 23684 22017 23712
rect 21499 23681 21511 23684
rect 21453 23675 21511 23681
rect 22005 23681 22017 23684
rect 22051 23681 22063 23715
rect 22005 23675 22063 23681
rect 22189 23715 22247 23721
rect 22189 23681 22201 23715
rect 22235 23681 22247 23715
rect 22189 23675 22247 23681
rect 22296 23684 23796 23712
rect 20516 23647 20574 23653
rect 20516 23613 20528 23647
rect 20562 23644 20574 23647
rect 20714 23644 20720 23656
rect 20562 23616 20720 23644
rect 20562 23613 20574 23616
rect 20516 23607 20574 23613
rect 20714 23604 20720 23616
rect 20772 23604 20778 23656
rect 20809 23647 20867 23653
rect 20809 23613 20821 23647
rect 20855 23644 20867 23647
rect 22296 23644 22324 23684
rect 20855 23616 22324 23644
rect 20855 23613 20867 23616
rect 20809 23607 20867 23613
rect 22462 23604 22468 23656
rect 22520 23604 22526 23656
rect 23768 23644 23796 23684
rect 23842 23672 23848 23724
rect 23900 23672 23906 23724
rect 24486 23672 24492 23724
rect 24544 23672 24550 23724
rect 24578 23672 24584 23724
rect 24636 23672 24642 23724
rect 24688 23721 24716 23752
rect 24964 23752 25452 23780
rect 24674 23715 24732 23721
rect 24674 23681 24686 23715
rect 24720 23681 24732 23715
rect 24674 23675 24732 23681
rect 24854 23672 24860 23724
rect 24912 23672 24918 23724
rect 24964 23721 24992 23752
rect 25424 23724 25452 23752
rect 26234 23740 26240 23792
rect 26292 23740 26298 23792
rect 26694 23780 26700 23792
rect 26344 23752 26700 23780
rect 24949 23715 25007 23721
rect 24949 23681 24961 23715
rect 24995 23681 25007 23715
rect 24949 23675 25007 23681
rect 25038 23672 25044 23724
rect 25096 23721 25102 23724
rect 25096 23712 25104 23721
rect 25096 23684 25141 23712
rect 25096 23675 25104 23684
rect 25096 23672 25102 23675
rect 25406 23672 25412 23724
rect 25464 23672 25470 23724
rect 26344 23721 26372 23752
rect 26694 23740 26700 23752
rect 26752 23740 26758 23792
rect 26053 23715 26111 23721
rect 26053 23681 26065 23715
rect 26099 23681 26111 23715
rect 26053 23675 26111 23681
rect 26329 23715 26387 23721
rect 26329 23681 26341 23715
rect 26375 23681 26387 23715
rect 26329 23675 26387 23681
rect 26421 23715 26479 23721
rect 26421 23681 26433 23715
rect 26467 23681 26479 23715
rect 26421 23675 26479 23681
rect 25314 23644 25320 23656
rect 23768 23616 25320 23644
rect 25314 23604 25320 23616
rect 25372 23604 25378 23656
rect 25958 23604 25964 23656
rect 26016 23644 26022 23656
rect 26068 23644 26096 23675
rect 26436 23644 26464 23675
rect 26602 23672 26608 23724
rect 26660 23672 26666 23724
rect 26016 23616 26096 23644
rect 26344 23616 26464 23644
rect 26016 23604 26022 23616
rect 26344 23588 26372 23616
rect 20220 23548 20392 23576
rect 20220 23536 20226 23548
rect 12768 23480 16896 23508
rect 12768 23468 12774 23480
rect 17218 23468 17224 23520
rect 17276 23468 17282 23520
rect 17512 23508 17540 23536
rect 18138 23508 18144 23520
rect 17512 23480 18144 23508
rect 18138 23468 18144 23480
rect 18196 23468 18202 23520
rect 20254 23468 20260 23520
rect 20312 23468 20318 23520
rect 20364 23508 20392 23548
rect 20990 23536 20996 23588
rect 21048 23576 21054 23588
rect 21048 23548 22508 23576
rect 21048 23536 21054 23548
rect 21542 23508 21548 23520
rect 20364 23480 21548 23508
rect 21542 23468 21548 23480
rect 21600 23468 21606 23520
rect 22370 23468 22376 23520
rect 22428 23468 22434 23520
rect 22480 23508 22508 23548
rect 23474 23536 23480 23588
rect 23532 23576 23538 23588
rect 26053 23579 26111 23585
rect 23532 23548 26013 23576
rect 23532 23536 23538 23548
rect 23750 23508 23756 23520
rect 22480 23480 23756 23508
rect 23750 23468 23756 23480
rect 23808 23468 23814 23520
rect 25225 23511 25283 23517
rect 25225 23477 25237 23511
rect 25271 23508 25283 23511
rect 25774 23508 25780 23520
rect 25271 23480 25780 23508
rect 25271 23477 25283 23480
rect 25225 23471 25283 23477
rect 25774 23468 25780 23480
rect 25832 23468 25838 23520
rect 25985 23508 26013 23548
rect 26053 23545 26065 23579
rect 26099 23576 26111 23579
rect 26326 23576 26332 23588
rect 26099 23548 26332 23576
rect 26099 23545 26111 23548
rect 26053 23539 26111 23545
rect 26326 23536 26332 23548
rect 26384 23536 26390 23588
rect 26878 23508 26884 23520
rect 25985 23480 26884 23508
rect 26878 23468 26884 23480
rect 26936 23468 26942 23520
rect 27356 23508 27384 23820
rect 27632 23820 28172 23848
rect 27632 23576 27660 23820
rect 28166 23808 28172 23820
rect 28224 23808 28230 23860
rect 28258 23808 28264 23860
rect 28316 23848 28322 23860
rect 30009 23851 30067 23857
rect 30009 23848 30021 23851
rect 28316 23820 30021 23848
rect 28316 23808 28322 23820
rect 30009 23817 30021 23820
rect 30055 23817 30067 23851
rect 30009 23811 30067 23817
rect 31294 23808 31300 23860
rect 31352 23848 31358 23860
rect 31481 23851 31539 23857
rect 31481 23848 31493 23851
rect 31352 23820 31493 23848
rect 31352 23808 31358 23820
rect 31481 23817 31493 23820
rect 31527 23817 31539 23851
rect 31481 23811 31539 23817
rect 31662 23808 31668 23860
rect 31720 23848 31726 23860
rect 32582 23848 32588 23860
rect 31720 23820 32588 23848
rect 31720 23808 31726 23820
rect 32582 23808 32588 23820
rect 32640 23808 32646 23860
rect 32674 23808 32680 23860
rect 32732 23848 32738 23860
rect 34054 23848 34060 23860
rect 32732 23820 34060 23848
rect 32732 23808 32738 23820
rect 34054 23808 34060 23820
rect 34112 23808 34118 23860
rect 37826 23848 37832 23860
rect 34164 23820 37832 23848
rect 28074 23740 28080 23792
rect 28132 23780 28138 23792
rect 28442 23780 28448 23792
rect 28132 23752 28448 23780
rect 28132 23740 28138 23752
rect 28442 23740 28448 23752
rect 28500 23740 28506 23792
rect 28810 23740 28816 23792
rect 28868 23780 28874 23792
rect 28868 23752 29684 23780
rect 28868 23740 28874 23752
rect 29656 23724 29684 23752
rect 27706 23672 27712 23724
rect 27764 23672 27770 23724
rect 28166 23672 28172 23724
rect 28224 23712 28230 23724
rect 28721 23715 28779 23721
rect 28721 23712 28733 23715
rect 28224 23684 28733 23712
rect 28224 23672 28230 23684
rect 28721 23681 28733 23684
rect 28767 23712 28779 23715
rect 28902 23712 28908 23724
rect 28767 23684 28908 23712
rect 28767 23681 28779 23684
rect 28721 23675 28779 23681
rect 28902 23672 28908 23684
rect 28960 23672 28966 23724
rect 28994 23672 29000 23724
rect 29052 23712 29058 23724
rect 29362 23712 29368 23724
rect 29052 23684 29368 23712
rect 29052 23672 29058 23684
rect 29362 23672 29368 23684
rect 29420 23672 29426 23724
rect 29454 23672 29460 23724
rect 29512 23712 29518 23724
rect 29549 23715 29607 23721
rect 29549 23712 29561 23715
rect 29512 23684 29561 23712
rect 29512 23672 29518 23684
rect 29549 23681 29561 23684
rect 29595 23681 29607 23715
rect 29549 23675 29607 23681
rect 29638 23672 29644 23724
rect 29696 23712 29702 23724
rect 29733 23715 29791 23721
rect 29733 23712 29745 23715
rect 29696 23684 29745 23712
rect 29696 23672 29702 23684
rect 29733 23681 29745 23684
rect 29779 23681 29791 23715
rect 29733 23675 29791 23681
rect 29825 23715 29883 23721
rect 29825 23681 29837 23715
rect 29871 23712 29883 23715
rect 30098 23712 30104 23724
rect 29871 23684 30104 23712
rect 29871 23681 29883 23684
rect 29825 23675 29883 23681
rect 30098 23672 30104 23684
rect 30156 23672 30162 23724
rect 30190 23672 30196 23724
rect 30248 23712 30254 23724
rect 31021 23715 31079 23721
rect 31021 23712 31033 23715
rect 30248 23684 31033 23712
rect 30248 23672 30254 23684
rect 31021 23681 31033 23684
rect 31067 23681 31079 23715
rect 31021 23675 31079 23681
rect 27724 23644 27752 23672
rect 28258 23644 28264 23656
rect 27724 23616 28264 23644
rect 28258 23604 28264 23616
rect 28316 23644 28322 23656
rect 28813 23647 28871 23653
rect 28316 23616 28764 23644
rect 28316 23604 28322 23616
rect 27706 23576 27712 23588
rect 27632 23548 27712 23576
rect 27706 23536 27712 23548
rect 27764 23536 27770 23588
rect 28736 23576 28764 23616
rect 28813 23613 28825 23647
rect 28859 23644 28871 23647
rect 31036 23644 31064 23675
rect 31202 23672 31208 23724
rect 31260 23672 31266 23724
rect 31294 23672 31300 23724
rect 31352 23712 31358 23724
rect 31352 23684 32536 23712
rect 31352 23672 31358 23684
rect 32398 23644 32404 23656
rect 28859 23616 30972 23644
rect 31036 23616 32404 23644
rect 28859 23613 28871 23616
rect 28813 23607 28871 23613
rect 28905 23579 28963 23585
rect 28905 23576 28917 23579
rect 28000 23548 28672 23576
rect 28736 23548 28917 23576
rect 28000 23520 28028 23548
rect 27430 23508 27436 23520
rect 27356 23480 27436 23508
rect 27430 23468 27436 23480
rect 27488 23468 27494 23520
rect 27982 23468 27988 23520
rect 28040 23468 28046 23520
rect 28350 23468 28356 23520
rect 28408 23508 28414 23520
rect 28537 23511 28595 23517
rect 28537 23508 28549 23511
rect 28408 23480 28549 23508
rect 28408 23468 28414 23480
rect 28537 23477 28549 23480
rect 28583 23477 28595 23511
rect 28644 23508 28672 23548
rect 28905 23545 28917 23548
rect 28951 23545 28963 23579
rect 30944 23576 30972 23616
rect 32398 23604 32404 23616
rect 32456 23604 32462 23656
rect 31202 23576 31208 23588
rect 28905 23539 28963 23545
rect 29656 23548 29868 23576
rect 30944 23548 31208 23576
rect 29656 23508 29684 23548
rect 28644 23480 29684 23508
rect 28537 23471 28595 23477
rect 29730 23468 29736 23520
rect 29788 23468 29794 23520
rect 29840 23508 29868 23548
rect 31202 23536 31208 23548
rect 31260 23536 31266 23588
rect 32508 23576 32536 23684
rect 32582 23672 32588 23724
rect 32640 23672 32646 23724
rect 32950 23672 32956 23724
rect 33008 23672 33014 23724
rect 33505 23715 33563 23721
rect 33505 23681 33517 23715
rect 33551 23681 33563 23715
rect 33505 23675 33563 23681
rect 32600 23644 32628 23672
rect 33520 23644 33548 23675
rect 33686 23672 33692 23724
rect 33744 23672 33750 23724
rect 33870 23672 33876 23724
rect 33928 23712 33934 23724
rect 33965 23715 34023 23721
rect 33965 23712 33977 23715
rect 33928 23684 33977 23712
rect 33928 23672 33934 23684
rect 33965 23681 33977 23684
rect 34011 23712 34023 23715
rect 34164 23712 34192 23820
rect 34514 23740 34520 23792
rect 34572 23780 34578 23792
rect 35713 23783 35771 23789
rect 35713 23780 35725 23783
rect 34572 23752 35725 23780
rect 34572 23740 34578 23752
rect 35713 23749 35725 23752
rect 35759 23749 35771 23783
rect 35713 23743 35771 23749
rect 34011 23684 34192 23712
rect 35069 23715 35127 23721
rect 34011 23681 34023 23684
rect 33965 23675 34023 23681
rect 35069 23681 35081 23715
rect 35115 23681 35127 23715
rect 35069 23675 35127 23681
rect 32600 23616 33548 23644
rect 32582 23576 32588 23588
rect 32508 23548 32588 23576
rect 32582 23536 32588 23548
rect 32640 23536 32646 23588
rect 32674 23536 32680 23588
rect 32732 23576 32738 23588
rect 33045 23579 33103 23585
rect 33045 23576 33057 23579
rect 32732 23548 33057 23576
rect 32732 23536 32738 23548
rect 33045 23545 33057 23548
rect 33091 23545 33103 23579
rect 33045 23539 33103 23545
rect 31297 23511 31355 23517
rect 31297 23508 31309 23511
rect 29840 23480 31309 23508
rect 31297 23477 31309 23480
rect 31343 23508 31355 23511
rect 33704 23508 33732 23672
rect 35084 23644 35112 23675
rect 35158 23672 35164 23724
rect 35216 23672 35222 23724
rect 36924 23721 36952 23820
rect 37826 23808 37832 23820
rect 37884 23808 37890 23860
rect 38010 23808 38016 23860
rect 38068 23808 38074 23860
rect 38580 23820 39068 23848
rect 38028 23780 38056 23808
rect 37108 23752 37412 23780
rect 37108 23721 37136 23752
rect 36909 23715 36967 23721
rect 35268 23684 36584 23712
rect 35268 23644 35296 23684
rect 35084 23616 35296 23644
rect 35345 23647 35403 23653
rect 35345 23613 35357 23647
rect 35391 23644 35403 23647
rect 35526 23644 35532 23656
rect 35391 23616 35532 23644
rect 35391 23613 35403 23616
rect 35345 23607 35403 23613
rect 35526 23604 35532 23616
rect 35584 23604 35590 23656
rect 36446 23604 36452 23656
rect 36504 23604 36510 23656
rect 36556 23644 36584 23684
rect 36909 23681 36921 23715
rect 36955 23681 36967 23715
rect 36909 23675 36967 23681
rect 37093 23715 37151 23721
rect 37093 23681 37105 23715
rect 37139 23681 37151 23715
rect 37093 23675 37151 23681
rect 37277 23715 37335 23721
rect 37277 23681 37289 23715
rect 37323 23681 37335 23715
rect 37384 23712 37412 23752
rect 37660 23752 38056 23780
rect 37458 23712 37464 23724
rect 37384 23684 37464 23712
rect 37277 23675 37335 23681
rect 37108 23644 37136 23675
rect 37292 23644 37320 23675
rect 37458 23672 37464 23684
rect 37516 23712 37522 23724
rect 37553 23715 37611 23721
rect 37553 23712 37565 23715
rect 37516 23684 37565 23712
rect 37516 23672 37522 23684
rect 37553 23681 37565 23684
rect 37599 23681 37611 23715
rect 37553 23675 37611 23681
rect 37660 23644 37688 23752
rect 37737 23715 37795 23721
rect 37737 23681 37749 23715
rect 37783 23681 37795 23715
rect 37737 23675 37795 23681
rect 37921 23715 37979 23721
rect 37921 23681 37933 23715
rect 37967 23712 37979 23715
rect 38286 23712 38292 23724
rect 37967 23684 38292 23712
rect 37967 23681 37979 23684
rect 37921 23675 37979 23681
rect 36556 23616 37136 23644
rect 37246 23616 37688 23644
rect 37246 23576 37274 23616
rect 35452 23548 37274 23576
rect 31343 23480 33732 23508
rect 31343 23477 31355 23480
rect 31297 23471 31355 23477
rect 34054 23468 34060 23520
rect 34112 23508 34118 23520
rect 34422 23508 34428 23520
rect 34112 23480 34428 23508
rect 34112 23468 34118 23480
rect 34422 23468 34428 23480
rect 34480 23508 34486 23520
rect 35452 23508 35480 23548
rect 37550 23536 37556 23588
rect 37608 23536 37614 23588
rect 37752 23576 37780 23675
rect 38286 23672 38292 23684
rect 38344 23672 38350 23724
rect 38378 23672 38384 23724
rect 38436 23712 38442 23724
rect 38580 23721 38608 23820
rect 38746 23740 38752 23792
rect 38804 23740 38810 23792
rect 39040 23780 39068 23820
rect 39114 23808 39120 23860
rect 39172 23848 39178 23860
rect 39172 23820 39528 23848
rect 39172 23808 39178 23820
rect 39500 23789 39528 23820
rect 39485 23783 39543 23789
rect 39040 23752 39252 23780
rect 38565 23715 38623 23721
rect 38565 23712 38577 23715
rect 38436 23684 38577 23712
rect 38436 23672 38442 23684
rect 38565 23681 38577 23684
rect 38611 23681 38623 23715
rect 38565 23675 38623 23681
rect 38841 23715 38899 23721
rect 38841 23681 38853 23715
rect 38887 23681 38899 23715
rect 38841 23675 38899 23681
rect 38470 23604 38476 23656
rect 38528 23604 38534 23656
rect 37660 23548 37780 23576
rect 38488 23576 38516 23604
rect 38856 23576 38884 23675
rect 38930 23672 38936 23724
rect 38988 23672 38994 23724
rect 39224 23721 39252 23752
rect 39485 23749 39497 23783
rect 39531 23749 39543 23783
rect 39485 23743 39543 23749
rect 39209 23715 39267 23721
rect 39209 23681 39221 23715
rect 39255 23681 39267 23715
rect 39209 23675 39267 23681
rect 39393 23715 39451 23721
rect 39393 23681 39405 23715
rect 39439 23681 39451 23715
rect 39393 23675 39451 23681
rect 38488 23548 38884 23576
rect 34480 23480 35480 23508
rect 34480 23468 34486 23480
rect 36538 23468 36544 23520
rect 36596 23508 36602 23520
rect 36909 23511 36967 23517
rect 36909 23508 36921 23511
rect 36596 23480 36921 23508
rect 36596 23468 36602 23480
rect 36909 23477 36921 23480
rect 36955 23477 36967 23511
rect 36909 23471 36967 23477
rect 36998 23468 37004 23520
rect 37056 23508 37062 23520
rect 37660 23508 37688 23548
rect 39114 23536 39120 23588
rect 39172 23536 39178 23588
rect 37056 23480 37688 23508
rect 37056 23468 37062 23480
rect 37734 23468 37740 23520
rect 37792 23468 37798 23520
rect 38746 23468 38752 23520
rect 38804 23508 38810 23520
rect 39408 23508 39436 23675
rect 39574 23672 39580 23724
rect 39632 23672 39638 23724
rect 38804 23480 39436 23508
rect 38804 23468 38810 23480
rect 39758 23468 39764 23520
rect 39816 23468 39822 23520
rect 1104 23418 41400 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 41400 23418
rect 1104 23344 41400 23366
rect 5074 23264 5080 23316
rect 5132 23304 5138 23316
rect 7098 23304 7104 23316
rect 5132 23276 7104 23304
rect 5132 23264 5138 23276
rect 7098 23264 7104 23276
rect 7156 23264 7162 23316
rect 7466 23264 7472 23316
rect 7524 23304 7530 23316
rect 7745 23307 7803 23313
rect 7745 23304 7757 23307
rect 7524 23276 7757 23304
rect 7524 23264 7530 23276
rect 7745 23273 7757 23276
rect 7791 23273 7803 23307
rect 7745 23267 7803 23273
rect 8110 23264 8116 23316
rect 8168 23304 8174 23316
rect 8168 23276 11284 23304
rect 8168 23264 8174 23276
rect 3142 23196 3148 23248
rect 3200 23236 3206 23248
rect 9398 23236 9404 23248
rect 3200 23208 9404 23236
rect 3200 23196 3206 23208
rect 1397 23171 1455 23177
rect 1397 23137 1409 23171
rect 1443 23168 1455 23171
rect 2406 23168 2412 23180
rect 1443 23140 2412 23168
rect 1443 23137 1455 23140
rect 1397 23131 1455 23137
rect 2406 23128 2412 23140
rect 2464 23128 2470 23180
rect 3050 23100 3056 23112
rect 2806 23072 3056 23100
rect 3050 23060 3056 23072
rect 3108 23060 3114 23112
rect 5074 23060 5080 23112
rect 5132 23060 5138 23112
rect 1670 22992 1676 23044
rect 1728 22992 1734 23044
rect 5184 23032 5212 23208
rect 9398 23196 9404 23208
rect 9456 23196 9462 23248
rect 9585 23239 9643 23245
rect 9585 23205 9597 23239
rect 9631 23205 9643 23239
rect 9585 23199 9643 23205
rect 10229 23239 10287 23245
rect 10229 23205 10241 23239
rect 10275 23236 10287 23239
rect 10275 23208 11009 23236
rect 10275 23205 10287 23208
rect 10229 23199 10287 23205
rect 5276 23140 7420 23168
rect 5276 23112 5304 23140
rect 5258 23060 5264 23112
rect 5316 23060 5322 23112
rect 5353 23103 5411 23109
rect 5353 23069 5365 23103
rect 5399 23069 5411 23103
rect 5353 23063 5411 23069
rect 5445 23103 5503 23109
rect 5445 23069 5457 23103
rect 5491 23100 5503 23103
rect 5994 23100 6000 23112
rect 5491 23072 6000 23100
rect 5491 23069 5503 23072
rect 5445 23063 5503 23069
rect 5368 23032 5396 23063
rect 5994 23060 6000 23072
rect 6052 23060 6058 23112
rect 7098 23060 7104 23112
rect 7156 23100 7162 23112
rect 7392 23109 7420 23140
rect 7484 23140 9352 23168
rect 7484 23112 7512 23140
rect 7193 23103 7251 23109
rect 7193 23100 7205 23103
rect 7156 23072 7205 23100
rect 7156 23060 7162 23072
rect 7193 23069 7205 23072
rect 7239 23069 7251 23103
rect 7193 23063 7251 23069
rect 7377 23103 7435 23109
rect 7377 23069 7389 23103
rect 7423 23069 7435 23103
rect 7377 23063 7435 23069
rect 5184 23004 5396 23032
rect 7208 23032 7236 23063
rect 7466 23060 7472 23112
rect 7524 23060 7530 23112
rect 7561 23103 7619 23109
rect 7561 23069 7573 23103
rect 7607 23100 7619 23103
rect 7926 23100 7932 23112
rect 7607 23072 7932 23100
rect 7607 23069 7619 23072
rect 7561 23063 7619 23069
rect 7926 23060 7932 23072
rect 7984 23060 7990 23112
rect 8570 23060 8576 23112
rect 8628 23060 8634 23112
rect 8846 23060 8852 23112
rect 8904 23100 8910 23112
rect 9324 23109 9352 23140
rect 8941 23103 8999 23109
rect 8941 23100 8953 23103
rect 8904 23072 8953 23100
rect 8904 23060 8910 23072
rect 8941 23069 8953 23072
rect 8987 23069 8999 23103
rect 8941 23063 8999 23069
rect 9034 23103 9092 23109
rect 9034 23069 9046 23103
rect 9080 23069 9092 23103
rect 9034 23063 9092 23069
rect 9309 23103 9367 23109
rect 9309 23069 9321 23103
rect 9355 23069 9367 23103
rect 9309 23063 9367 23069
rect 9406 23103 9464 23109
rect 9406 23069 9418 23103
rect 9452 23100 9464 23103
rect 9600 23100 9628 23199
rect 10594 23128 10600 23180
rect 10652 23168 10658 23180
rect 10689 23171 10747 23177
rect 10689 23168 10701 23171
rect 10652 23140 10701 23168
rect 10652 23128 10658 23140
rect 10689 23137 10701 23140
rect 10735 23137 10747 23171
rect 10689 23131 10747 23137
rect 9953 23103 10011 23109
rect 9953 23100 9965 23103
rect 9452 23072 9536 23100
rect 9600 23072 9965 23100
rect 9452 23069 9464 23072
rect 9406 23063 9464 23069
rect 8110 23032 8116 23044
rect 7208 23004 8116 23032
rect 8110 22992 8116 23004
rect 8168 22992 8174 23044
rect 8588 23032 8616 23060
rect 9048 23032 9076 23063
rect 8588 23004 9076 23032
rect 9217 23035 9275 23041
rect 9217 23001 9229 23035
rect 9263 23001 9275 23035
rect 9508 23032 9536 23072
rect 9953 23069 9965 23072
rect 9999 23069 10011 23103
rect 9953 23063 10011 23069
rect 10502 23060 10508 23112
rect 10560 23100 10566 23112
rect 10873 23103 10931 23109
rect 10873 23100 10885 23103
rect 10560 23072 10885 23100
rect 10560 23060 10566 23072
rect 10873 23069 10885 23072
rect 10919 23069 10931 23103
rect 10873 23063 10931 23069
rect 9508 23004 9628 23032
rect 9217 22995 9275 23001
rect 4798 22924 4804 22976
rect 4856 22964 4862 22976
rect 5629 22967 5687 22973
rect 5629 22964 5641 22967
rect 4856 22936 5641 22964
rect 4856 22924 4862 22936
rect 5629 22933 5641 22936
rect 5675 22933 5687 22967
rect 9232 22964 9260 22995
rect 9600 22976 9628 23004
rect 9490 22964 9496 22976
rect 9232 22936 9496 22964
rect 5629 22927 5687 22933
rect 9490 22924 9496 22936
rect 9548 22924 9554 22976
rect 9582 22924 9588 22976
rect 9640 22924 9646 22976
rect 10888 22964 10916 23063
rect 10981 23032 11009 23208
rect 11256 23109 11284 23276
rect 11974 23264 11980 23316
rect 12032 23264 12038 23316
rect 14458 23264 14464 23316
rect 14516 23304 14522 23316
rect 14829 23307 14887 23313
rect 14829 23304 14841 23307
rect 14516 23276 14841 23304
rect 14516 23264 14522 23276
rect 14829 23273 14841 23276
rect 14875 23273 14887 23307
rect 14829 23267 14887 23273
rect 15838 23264 15844 23316
rect 15896 23264 15902 23316
rect 17678 23264 17684 23316
rect 17736 23304 17742 23316
rect 22186 23304 22192 23316
rect 17736 23276 22192 23304
rect 17736 23264 17742 23276
rect 22186 23264 22192 23276
rect 22244 23264 22250 23316
rect 22738 23264 22744 23316
rect 22796 23304 22802 23316
rect 23569 23307 23627 23313
rect 23569 23304 23581 23307
rect 22796 23276 23581 23304
rect 22796 23264 22802 23276
rect 23569 23273 23581 23276
rect 23615 23273 23627 23307
rect 23569 23267 23627 23273
rect 23934 23264 23940 23316
rect 23992 23304 23998 23316
rect 26418 23304 26424 23316
rect 23992 23276 26424 23304
rect 23992 23264 23998 23276
rect 26418 23264 26424 23276
rect 26476 23264 26482 23316
rect 26878 23264 26884 23316
rect 26936 23304 26942 23316
rect 27338 23304 27344 23316
rect 26936 23276 27344 23304
rect 26936 23264 26942 23276
rect 27338 23264 27344 23276
rect 27396 23264 27402 23316
rect 27614 23264 27620 23316
rect 27672 23304 27678 23316
rect 28261 23307 28319 23313
rect 28261 23304 28273 23307
rect 27672 23276 28273 23304
rect 27672 23264 27678 23276
rect 28261 23273 28273 23276
rect 28307 23273 28319 23307
rect 28261 23267 28319 23273
rect 30006 23264 30012 23316
rect 30064 23304 30070 23316
rect 30064 23276 32720 23304
rect 30064 23264 30070 23276
rect 15856 23236 15884 23264
rect 32692 23248 32720 23276
rect 39850 23264 39856 23316
rect 39908 23304 39914 23316
rect 40218 23304 40224 23316
rect 39908 23276 40224 23304
rect 39908 23264 39914 23276
rect 40218 23264 40224 23276
rect 40276 23264 40282 23316
rect 40310 23264 40316 23316
rect 40368 23264 40374 23316
rect 14476 23208 15884 23236
rect 13998 23128 14004 23180
rect 14056 23168 14062 23180
rect 14476 23177 14504 23208
rect 17494 23196 17500 23248
rect 17552 23236 17558 23248
rect 24670 23236 24676 23248
rect 17552 23208 24676 23236
rect 17552 23196 17558 23208
rect 14461 23171 14519 23177
rect 14056 23140 14412 23168
rect 14056 23128 14062 23140
rect 11241 23103 11299 23109
rect 11241 23069 11253 23103
rect 11287 23069 11299 23103
rect 11241 23063 11299 23069
rect 11793 23103 11851 23109
rect 11793 23069 11805 23103
rect 11839 23069 11851 23103
rect 11793 23063 11851 23069
rect 11885 23103 11943 23109
rect 11885 23069 11897 23103
rect 11931 23069 11943 23103
rect 11885 23063 11943 23069
rect 11606 23032 11612 23044
rect 10981 23004 11612 23032
rect 11606 22992 11612 23004
rect 11664 22992 11670 23044
rect 11146 22964 11152 22976
rect 10888 22936 11152 22964
rect 11146 22924 11152 22936
rect 11204 22924 11210 22976
rect 11238 22924 11244 22976
rect 11296 22964 11302 22976
rect 11808 22964 11836 23063
rect 11900 23032 11928 23063
rect 11974 23060 11980 23112
rect 12032 23100 12038 23112
rect 14384 23109 14412 23140
rect 14461 23137 14473 23171
rect 14507 23137 14519 23171
rect 15565 23171 15623 23177
rect 15565 23168 15577 23171
rect 14461 23131 14519 23137
rect 14936 23140 15577 23168
rect 12069 23103 12127 23109
rect 12069 23100 12081 23103
rect 12032 23072 12081 23100
rect 12032 23060 12038 23072
rect 12069 23069 12081 23072
rect 12115 23069 12127 23103
rect 12069 23063 12127 23069
rect 14369 23103 14427 23109
rect 14369 23069 14381 23103
rect 14415 23069 14427 23103
rect 14369 23063 14427 23069
rect 14553 23103 14611 23109
rect 14553 23069 14565 23103
rect 14599 23069 14611 23103
rect 14553 23063 14611 23069
rect 12342 23032 12348 23044
rect 11900 23004 12348 23032
rect 12342 22992 12348 23004
rect 12400 22992 12406 23044
rect 13354 22964 13360 22976
rect 11296 22936 13360 22964
rect 11296 22924 11302 22936
rect 13354 22924 13360 22936
rect 13412 22924 13418 22976
rect 14384 22964 14412 23063
rect 14568 23032 14596 23063
rect 14642 23060 14648 23112
rect 14700 23100 14706 23112
rect 14936 23100 14964 23140
rect 15565 23137 15577 23140
rect 15611 23137 15623 23171
rect 15565 23131 15623 23137
rect 15841 23171 15899 23177
rect 15841 23137 15853 23171
rect 15887 23168 15899 23171
rect 16114 23168 16120 23180
rect 15887 23140 16120 23168
rect 15887 23137 15899 23140
rect 15841 23131 15899 23137
rect 16114 23128 16120 23140
rect 16172 23128 16178 23180
rect 16298 23128 16304 23180
rect 16356 23168 16362 23180
rect 19334 23168 19340 23180
rect 16356 23140 19340 23168
rect 16356 23128 16362 23140
rect 19334 23128 19340 23140
rect 19392 23128 19398 23180
rect 21085 23171 21143 23177
rect 21085 23168 21097 23171
rect 20640 23140 21097 23168
rect 14700 23072 14964 23100
rect 15013 23103 15071 23109
rect 14700 23060 14706 23072
rect 15013 23069 15025 23103
rect 15059 23100 15071 23103
rect 15059 23072 15700 23100
rect 15059 23069 15071 23072
rect 15013 23063 15071 23069
rect 14826 23032 14832 23044
rect 14568 23004 14832 23032
rect 14826 22992 14832 23004
rect 14884 22992 14890 23044
rect 15194 22992 15200 23044
rect 15252 23032 15258 23044
rect 15289 23035 15347 23041
rect 15289 23032 15301 23035
rect 15252 23004 15301 23032
rect 15252 22992 15258 23004
rect 15289 23001 15301 23004
rect 15335 23001 15347 23035
rect 15672 23032 15700 23072
rect 15746 23060 15752 23112
rect 15804 23060 15810 23112
rect 15930 23060 15936 23112
rect 15988 23060 15994 23112
rect 16025 23103 16083 23109
rect 16025 23069 16037 23103
rect 16071 23100 16083 23103
rect 17310 23100 17316 23112
rect 16071 23072 17316 23100
rect 16071 23069 16083 23072
rect 16025 23063 16083 23069
rect 17310 23060 17316 23072
rect 17368 23060 17374 23112
rect 17402 23060 17408 23112
rect 17460 23060 17466 23112
rect 18046 23060 18052 23112
rect 18104 23060 18110 23112
rect 18322 23060 18328 23112
rect 18380 23100 18386 23112
rect 20530 23100 20536 23112
rect 18380 23072 20536 23100
rect 18380 23060 18386 23072
rect 20530 23060 20536 23072
rect 20588 23060 20594 23112
rect 16482 23032 16488 23044
rect 15672 23004 16488 23032
rect 15289 22995 15347 23001
rect 16482 22992 16488 23004
rect 16540 22992 16546 23044
rect 16666 22992 16672 23044
rect 16724 23032 16730 23044
rect 17218 23032 17224 23044
rect 16724 23004 17224 23032
rect 16724 22992 16730 23004
rect 17218 22992 17224 23004
rect 17276 22992 17282 23044
rect 17957 23035 18015 23041
rect 17957 23001 17969 23035
rect 18003 23032 18015 23035
rect 18064 23032 18092 23060
rect 18003 23004 18092 23032
rect 18003 23001 18015 23004
rect 17957 22995 18015 23001
rect 18690 22992 18696 23044
rect 18748 23032 18754 23044
rect 20640 23032 20668 23140
rect 21085 23137 21097 23140
rect 21131 23137 21143 23171
rect 21085 23131 21143 23137
rect 20901 23103 20959 23109
rect 20901 23069 20913 23103
rect 20947 23100 20959 23103
rect 21100 23100 21128 23131
rect 21174 23128 21180 23180
rect 21232 23128 21238 23180
rect 22848 23177 22876 23208
rect 24670 23196 24676 23208
rect 24728 23196 24734 23248
rect 29454 23236 29460 23248
rect 24780 23208 29460 23236
rect 22833 23171 22891 23177
rect 22833 23137 22845 23171
rect 22879 23137 22891 23171
rect 22833 23131 22891 23137
rect 22922 23128 22928 23180
rect 22980 23168 22986 23180
rect 24780 23168 24808 23208
rect 29454 23196 29460 23208
rect 29512 23236 29518 23248
rect 29822 23236 29828 23248
rect 29512 23208 29828 23236
rect 29512 23196 29518 23208
rect 29822 23196 29828 23208
rect 29880 23236 29886 23248
rect 30190 23236 30196 23248
rect 29880 23208 30196 23236
rect 29880 23196 29886 23208
rect 30190 23196 30196 23208
rect 30248 23196 30254 23248
rect 32674 23196 32680 23248
rect 32732 23196 32738 23248
rect 39022 23236 39028 23248
rect 32876 23208 38700 23236
rect 32876 23180 32904 23208
rect 22980 23140 24808 23168
rect 22980 23128 22986 23140
rect 25038 23128 25044 23180
rect 25096 23168 25102 23180
rect 25685 23171 25743 23177
rect 25685 23168 25697 23171
rect 25096 23140 25697 23168
rect 25096 23128 25102 23140
rect 25685 23137 25697 23140
rect 25731 23137 25743 23171
rect 26510 23168 26516 23180
rect 25685 23131 25743 23137
rect 25884 23140 26516 23168
rect 21450 23100 21456 23112
rect 20947 23072 21036 23100
rect 21100 23072 21456 23100
rect 20947 23069 20959 23072
rect 20901 23063 20959 23069
rect 18748 23004 20668 23032
rect 18748 22992 18754 23004
rect 14550 22964 14556 22976
rect 14384 22936 14556 22964
rect 14550 22924 14556 22936
rect 14608 22924 14614 22976
rect 16117 22967 16175 22973
rect 16117 22933 16129 22967
rect 16163 22964 16175 22967
rect 16206 22964 16212 22976
rect 16163 22936 16212 22964
rect 16163 22933 16175 22936
rect 16117 22927 16175 22933
rect 16206 22924 16212 22936
rect 16264 22924 16270 22976
rect 17402 22924 17408 22976
rect 17460 22964 17466 22976
rect 17497 22967 17555 22973
rect 17497 22964 17509 22967
rect 17460 22936 17509 22964
rect 17460 22924 17466 22936
rect 17497 22933 17509 22936
rect 17543 22933 17555 22967
rect 17497 22927 17555 22933
rect 18046 22924 18052 22976
rect 18104 22924 18110 22976
rect 20714 22924 20720 22976
rect 20772 22924 20778 22976
rect 21008 22964 21036 23072
rect 21450 23060 21456 23072
rect 21508 23060 21514 23112
rect 21542 23060 21548 23112
rect 21600 23100 21606 23112
rect 23201 23103 23259 23109
rect 23201 23100 23213 23103
rect 21600 23072 23213 23100
rect 21600 23060 21606 23072
rect 23201 23069 23213 23072
rect 23247 23069 23259 23103
rect 23201 23063 23259 23069
rect 21266 22992 21272 23044
rect 21324 22992 21330 23044
rect 23216 23032 23244 23063
rect 23382 23060 23388 23112
rect 23440 23060 23446 23112
rect 25884 23109 25912 23140
rect 26510 23128 26516 23140
rect 26568 23128 26574 23180
rect 26712 23140 30420 23168
rect 25869 23103 25927 23109
rect 25869 23069 25881 23103
rect 25915 23069 25927 23103
rect 25869 23063 25927 23069
rect 26050 23060 26056 23112
rect 26108 23060 26114 23112
rect 26712 23109 26740 23140
rect 30392 23112 30420 23140
rect 31496 23140 31984 23168
rect 26697 23103 26755 23109
rect 26697 23069 26709 23103
rect 26743 23069 26755 23103
rect 26697 23063 26755 23069
rect 26878 23060 26884 23112
rect 26936 23060 26942 23112
rect 27246 23060 27252 23112
rect 27304 23060 27310 23112
rect 27614 23060 27620 23112
rect 27672 23100 27678 23112
rect 27890 23100 27896 23112
rect 27672 23072 27896 23100
rect 27672 23060 27678 23072
rect 27890 23060 27896 23072
rect 27948 23060 27954 23112
rect 28261 23103 28319 23109
rect 28261 23069 28273 23103
rect 28307 23100 28319 23103
rect 28350 23100 28356 23112
rect 28307 23072 28356 23100
rect 28307 23069 28319 23072
rect 28261 23063 28319 23069
rect 28350 23060 28356 23072
rect 28408 23060 28414 23112
rect 28445 23103 28503 23109
rect 28445 23069 28457 23103
rect 28491 23100 28503 23103
rect 28534 23100 28540 23112
rect 28491 23072 28540 23100
rect 28491 23069 28503 23072
rect 28445 23063 28503 23069
rect 25498 23032 25504 23044
rect 23216 23004 25504 23032
rect 25498 22992 25504 23004
rect 25556 22992 25562 23044
rect 28460 23032 28488 23063
rect 28534 23060 28540 23072
rect 28592 23060 28598 23112
rect 30374 23060 30380 23112
rect 30432 23060 30438 23112
rect 31496 23109 31524 23140
rect 31481 23103 31539 23109
rect 31481 23069 31493 23103
rect 31527 23069 31539 23103
rect 31481 23063 31539 23069
rect 31662 23060 31668 23112
rect 31720 23060 31726 23112
rect 31754 23060 31760 23112
rect 31812 23060 31818 23112
rect 31956 23109 31984 23140
rect 32582 23128 32588 23180
rect 32640 23168 32646 23180
rect 32769 23171 32827 23177
rect 32769 23168 32781 23171
rect 32640 23140 32781 23168
rect 32640 23128 32646 23140
rect 32769 23137 32781 23140
rect 32815 23137 32827 23171
rect 32769 23131 32827 23137
rect 32858 23128 32864 23180
rect 32916 23128 32922 23180
rect 36170 23128 36176 23180
rect 36228 23128 36234 23180
rect 31941 23103 31999 23109
rect 31941 23069 31953 23103
rect 31987 23100 31999 23103
rect 32030 23100 32036 23112
rect 31987 23072 32036 23100
rect 31987 23069 31999 23072
rect 31941 23063 31999 23069
rect 32030 23060 32036 23072
rect 32088 23060 32094 23112
rect 32493 23103 32551 23109
rect 32493 23069 32505 23103
rect 32539 23069 32551 23103
rect 32493 23063 32551 23069
rect 32677 23103 32735 23109
rect 32677 23069 32689 23103
rect 32723 23100 32735 23103
rect 33226 23100 33232 23112
rect 32723 23072 33232 23100
rect 32723 23069 32735 23072
rect 32677 23063 32735 23069
rect 26988 23004 28488 23032
rect 22830 22964 22836 22976
rect 21008 22936 22836 22964
rect 22830 22924 22836 22936
rect 22888 22924 22894 22976
rect 23566 22924 23572 22976
rect 23624 22964 23630 22976
rect 24854 22964 24860 22976
rect 23624 22936 24860 22964
rect 23624 22924 23630 22936
rect 24854 22924 24860 22936
rect 24912 22924 24918 22976
rect 26878 22924 26884 22976
rect 26936 22964 26942 22976
rect 26988 22964 27016 23004
rect 26936 22936 27016 22964
rect 26936 22924 26942 22936
rect 28074 22924 28080 22976
rect 28132 22924 28138 22976
rect 30558 22924 30564 22976
rect 30616 22964 30622 22976
rect 31573 22967 31631 22973
rect 31573 22964 31585 22967
rect 30616 22936 31585 22964
rect 30616 22924 30622 22936
rect 31573 22933 31585 22936
rect 31619 22933 31631 22967
rect 31573 22927 31631 22933
rect 31846 22924 31852 22976
rect 31904 22924 31910 22976
rect 32048 22964 32076 23060
rect 32214 22992 32220 23044
rect 32272 23032 32278 23044
rect 32508 23032 32536 23063
rect 33226 23060 33232 23072
rect 33284 23060 33290 23112
rect 34241 23103 34299 23109
rect 34241 23100 34253 23103
rect 33428 23072 34253 23100
rect 32950 23032 32956 23044
rect 32272 23004 32956 23032
rect 32272 22992 32278 23004
rect 32950 22992 32956 23004
rect 33008 22992 33014 23044
rect 32674 22964 32680 22976
rect 32048 22936 32680 22964
rect 32674 22924 32680 22936
rect 32732 22964 32738 22976
rect 33428 22964 33456 23072
rect 34241 23069 34253 23072
rect 34287 23069 34299 23103
rect 34241 23063 34299 23069
rect 34256 23032 34284 23063
rect 34422 23060 34428 23112
rect 34480 23060 34486 23112
rect 36262 23060 36268 23112
rect 36320 23100 36326 23112
rect 37182 23100 37188 23112
rect 36320 23072 37188 23100
rect 36320 23060 36326 23072
rect 37182 23060 37188 23072
rect 37240 23060 37246 23112
rect 38562 23060 38568 23112
rect 38620 23100 38626 23112
rect 38672 23109 38700 23208
rect 38948 23208 39028 23236
rect 38948 23109 38976 23208
rect 39022 23196 39028 23208
rect 39080 23196 39086 23248
rect 38657 23103 38715 23109
rect 38657 23100 38669 23103
rect 38620 23072 38669 23100
rect 38620 23060 38626 23072
rect 38657 23069 38669 23072
rect 38703 23069 38715 23103
rect 38657 23063 38715 23069
rect 38933 23103 38991 23109
rect 38933 23069 38945 23103
rect 38979 23069 38991 23103
rect 38933 23063 38991 23069
rect 39025 23103 39083 23109
rect 39025 23069 39037 23103
rect 39071 23100 39083 23103
rect 39574 23100 39580 23112
rect 39071 23072 39580 23100
rect 39071 23069 39083 23072
rect 39025 23063 39083 23069
rect 34514 23032 34520 23044
rect 34256 23004 34520 23032
rect 34514 22992 34520 23004
rect 34572 22992 34578 23044
rect 35802 22992 35808 23044
rect 35860 23032 35866 23044
rect 36541 23035 36599 23041
rect 36541 23032 36553 23035
rect 35860 23004 36553 23032
rect 35860 22992 35866 23004
rect 36541 23001 36553 23004
rect 36587 23001 36599 23035
rect 36541 22995 36599 23001
rect 36630 22992 36636 23044
rect 36688 22992 36694 23044
rect 38746 22992 38752 23044
rect 38804 23032 38810 23044
rect 38841 23035 38899 23041
rect 38841 23032 38853 23035
rect 38804 23004 38853 23032
rect 38804 22992 38810 23004
rect 38841 23001 38853 23004
rect 38887 23001 38899 23035
rect 38841 22995 38899 23001
rect 32732 22936 33456 22964
rect 32732 22924 32738 22936
rect 33502 22924 33508 22976
rect 33560 22964 33566 22976
rect 34333 22967 34391 22973
rect 34333 22964 34345 22967
rect 33560 22936 34345 22964
rect 33560 22924 33566 22936
rect 34333 22933 34345 22936
rect 34379 22933 34391 22967
rect 34333 22927 34391 22933
rect 35989 22967 36047 22973
rect 35989 22933 36001 22967
rect 36035 22964 36047 22967
rect 37274 22964 37280 22976
rect 36035 22936 37280 22964
rect 36035 22933 36047 22936
rect 35989 22927 36047 22933
rect 37274 22924 37280 22936
rect 37332 22924 37338 22976
rect 37458 22924 37464 22976
rect 37516 22964 37522 22976
rect 39040 22964 39068 23063
rect 39574 23060 39580 23072
rect 39632 23060 39638 23112
rect 39942 22992 39948 23044
rect 40000 22992 40006 23044
rect 40129 23035 40187 23041
rect 40129 23001 40141 23035
rect 40175 23032 40187 23035
rect 40586 23032 40592 23044
rect 40175 23004 40592 23032
rect 40175 23001 40187 23004
rect 40129 22995 40187 23001
rect 40586 22992 40592 23004
rect 40644 22992 40650 23044
rect 37516 22936 39068 22964
rect 37516 22924 37522 22936
rect 39206 22924 39212 22976
rect 39264 22924 39270 22976
rect 1104 22874 41400 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 41400 22874
rect 1104 22800 41400 22822
rect 1670 22720 1676 22772
rect 1728 22760 1734 22772
rect 1857 22763 1915 22769
rect 1857 22760 1869 22763
rect 1728 22732 1869 22760
rect 1728 22720 1734 22732
rect 1857 22729 1869 22732
rect 1903 22729 1915 22763
rect 1857 22723 1915 22729
rect 2866 22720 2872 22772
rect 2924 22720 2930 22772
rect 2961 22763 3019 22769
rect 2961 22729 2973 22763
rect 3007 22760 3019 22763
rect 3142 22760 3148 22772
rect 3007 22732 3148 22760
rect 3007 22729 3019 22732
rect 2961 22723 3019 22729
rect 3142 22720 3148 22732
rect 3200 22720 3206 22772
rect 5902 22720 5908 22772
rect 5960 22760 5966 22772
rect 7466 22760 7472 22772
rect 5960 22732 7472 22760
rect 5960 22720 5966 22732
rect 7466 22720 7472 22732
rect 7524 22720 7530 22772
rect 8297 22763 8355 22769
rect 8297 22729 8309 22763
rect 8343 22760 8355 22763
rect 8849 22763 8907 22769
rect 8849 22760 8861 22763
rect 8343 22732 8861 22760
rect 8343 22729 8355 22732
rect 8297 22723 8355 22729
rect 8849 22729 8861 22732
rect 8895 22760 8907 22763
rect 11882 22760 11888 22772
rect 8895 22732 11888 22760
rect 8895 22729 8907 22732
rect 8849 22723 8907 22729
rect 11882 22720 11888 22732
rect 11940 22760 11946 22772
rect 11940 22732 12434 22760
rect 11940 22720 11946 22732
rect 5810 22692 5816 22704
rect 5658 22664 5816 22692
rect 5810 22652 5816 22664
rect 5868 22652 5874 22704
rect 7282 22652 7288 22704
rect 7340 22652 7346 22704
rect 8757 22695 8815 22701
rect 8757 22661 8769 22695
rect 8803 22692 8815 22695
rect 9122 22692 9128 22704
rect 8803 22664 9128 22692
rect 8803 22661 8815 22664
rect 8757 22655 8815 22661
rect 9122 22652 9128 22664
rect 9180 22652 9186 22704
rect 10229 22695 10287 22701
rect 10229 22692 10241 22695
rect 9232 22664 10241 22692
rect 2041 22627 2099 22633
rect 2041 22593 2053 22627
rect 2087 22624 2099 22627
rect 2087 22596 2544 22624
rect 2087 22593 2099 22596
rect 2041 22587 2099 22593
rect 2516 22497 2544 22596
rect 6362 22584 6368 22636
rect 6420 22624 6426 22636
rect 6549 22627 6607 22633
rect 6549 22624 6561 22627
rect 6420 22596 6561 22624
rect 6420 22584 6426 22596
rect 6549 22593 6561 22596
rect 6595 22593 6607 22627
rect 6549 22587 6607 22593
rect 8202 22584 8208 22636
rect 8260 22624 8266 22636
rect 9232 22624 9260 22664
rect 10229 22661 10241 22664
rect 10275 22661 10287 22695
rect 12406 22692 12434 22732
rect 15304 22732 16436 22760
rect 12805 22695 12863 22701
rect 12805 22692 12817 22695
rect 12406 22664 12817 22692
rect 10229 22655 10287 22661
rect 12805 22661 12817 22664
rect 12851 22661 12863 22695
rect 12805 22655 12863 22661
rect 12912 22664 15056 22692
rect 9766 22624 9772 22636
rect 8260 22596 9260 22624
rect 9646 22596 9772 22624
rect 8260 22584 8266 22596
rect 3145 22559 3203 22565
rect 3145 22525 3157 22559
rect 3191 22525 3203 22559
rect 3145 22519 3203 22525
rect 2501 22491 2559 22497
rect 2501 22457 2513 22491
rect 2547 22457 2559 22491
rect 2501 22451 2559 22457
rect 3160 22432 3188 22519
rect 4154 22516 4160 22568
rect 4212 22516 4218 22568
rect 4433 22559 4491 22565
rect 4433 22525 4445 22559
rect 4479 22556 4491 22559
rect 4522 22556 4528 22568
rect 4479 22528 4528 22556
rect 4479 22525 4491 22528
rect 4433 22519 4491 22525
rect 4522 22516 4528 22528
rect 4580 22516 4586 22568
rect 6825 22559 6883 22565
rect 6825 22525 6837 22559
rect 6871 22556 6883 22559
rect 7190 22556 7196 22568
rect 6871 22528 7196 22556
rect 6871 22525 6883 22528
rect 6825 22519 6883 22525
rect 7190 22516 7196 22528
rect 7248 22516 7254 22568
rect 9033 22559 9091 22565
rect 9033 22525 9045 22559
rect 9079 22556 9091 22559
rect 9398 22556 9404 22568
rect 9079 22528 9404 22556
rect 9079 22525 9091 22528
rect 9033 22519 9091 22525
rect 9398 22516 9404 22528
rect 9456 22516 9462 22568
rect 9490 22516 9496 22568
rect 9548 22556 9554 22568
rect 9646 22556 9674 22596
rect 9766 22584 9772 22596
rect 9824 22584 9830 22636
rect 9953 22627 10011 22633
rect 9953 22593 9965 22627
rect 9999 22624 10011 22627
rect 10042 22624 10048 22636
rect 9999 22596 10048 22624
rect 9999 22593 10011 22596
rect 9953 22587 10011 22593
rect 10042 22584 10048 22596
rect 10100 22584 10106 22636
rect 10137 22627 10195 22633
rect 10137 22593 10149 22627
rect 10183 22593 10195 22627
rect 10137 22587 10195 22593
rect 10321 22627 10379 22633
rect 10321 22593 10333 22627
rect 10367 22593 10379 22627
rect 10321 22587 10379 22593
rect 11517 22627 11575 22633
rect 11517 22593 11529 22627
rect 11563 22624 11575 22627
rect 12066 22624 12072 22636
rect 11563 22596 12072 22624
rect 11563 22593 11575 22596
rect 11517 22587 11575 22593
rect 10152 22556 10180 22587
rect 9548 22528 10180 22556
rect 10336 22556 10364 22587
rect 12066 22584 12072 22596
rect 12124 22584 12130 22636
rect 12158 22584 12164 22636
rect 12216 22584 12222 22636
rect 12526 22584 12532 22636
rect 12584 22584 12590 22636
rect 12710 22584 12716 22636
rect 12768 22584 12774 22636
rect 12912 22633 12940 22664
rect 15028 22636 15056 22664
rect 12897 22627 12955 22633
rect 12897 22593 12909 22627
rect 12943 22593 12955 22627
rect 12897 22587 12955 22593
rect 12434 22556 12440 22568
rect 10336 22528 12440 22556
rect 9548 22516 9554 22528
rect 9582 22448 9588 22500
rect 9640 22488 9646 22500
rect 10336 22488 10364 22528
rect 12434 22516 12440 22528
rect 12492 22556 12498 22568
rect 12912 22556 12940 22587
rect 13722 22584 13728 22636
rect 13780 22624 13786 22636
rect 14090 22624 14096 22636
rect 13780 22596 14096 22624
rect 13780 22584 13786 22596
rect 14090 22584 14096 22596
rect 14148 22584 14154 22636
rect 14645 22627 14703 22633
rect 14645 22593 14657 22627
rect 14691 22593 14703 22627
rect 14645 22587 14703 22593
rect 12492 22528 12940 22556
rect 14660 22556 14688 22587
rect 14734 22584 14740 22636
rect 14792 22584 14798 22636
rect 15010 22584 15016 22636
rect 15068 22584 15074 22636
rect 15304 22633 15332 22732
rect 15470 22652 15476 22704
rect 15528 22692 15534 22704
rect 15565 22695 15623 22701
rect 15565 22692 15577 22695
rect 15528 22664 15577 22692
rect 15528 22652 15534 22664
rect 15565 22661 15577 22664
rect 15611 22661 15623 22695
rect 15565 22655 15623 22661
rect 16022 22652 16028 22704
rect 16080 22692 16086 22704
rect 16408 22692 16436 22732
rect 16482 22720 16488 22772
rect 16540 22720 16546 22772
rect 17034 22760 17040 22772
rect 16961 22732 17040 22760
rect 16758 22692 16764 22704
rect 16080 22664 16252 22692
rect 16408 22664 16764 22692
rect 16080 22652 16086 22664
rect 15289 22627 15347 22633
rect 15289 22593 15301 22627
rect 15335 22593 15347 22627
rect 15289 22587 15347 22593
rect 15381 22627 15439 22633
rect 15381 22593 15393 22627
rect 15427 22593 15439 22627
rect 15381 22587 15439 22593
rect 15396 22556 15424 22587
rect 15654 22584 15660 22636
rect 15712 22584 15718 22636
rect 15838 22584 15844 22636
rect 15896 22584 15902 22636
rect 15930 22584 15936 22636
rect 15988 22584 15994 22636
rect 16117 22627 16175 22633
rect 16117 22624 16129 22627
rect 16040 22596 16129 22624
rect 15856 22556 15884 22584
rect 14660 22528 14780 22556
rect 15396 22528 15884 22556
rect 12492 22516 12498 22528
rect 9640 22460 10364 22488
rect 9640 22448 9646 22460
rect 11698 22448 11704 22500
rect 11756 22488 11762 22500
rect 11793 22491 11851 22497
rect 11793 22488 11805 22491
rect 11756 22460 11805 22488
rect 11756 22448 11762 22460
rect 11793 22457 11805 22460
rect 11839 22457 11851 22491
rect 13906 22488 13912 22500
rect 11793 22451 11851 22457
rect 13096 22460 13912 22488
rect 3142 22380 3148 22432
rect 3200 22380 3206 22432
rect 8386 22380 8392 22432
rect 8444 22380 8450 22432
rect 10505 22423 10563 22429
rect 10505 22389 10517 22423
rect 10551 22420 10563 22423
rect 10778 22420 10784 22432
rect 10551 22392 10784 22420
rect 10551 22389 10563 22392
rect 10505 22383 10563 22389
rect 10778 22380 10784 22392
rect 10836 22380 10842 22432
rect 13096 22429 13124 22460
rect 13906 22448 13912 22460
rect 13964 22448 13970 22500
rect 13081 22423 13139 22429
rect 13081 22389 13093 22423
rect 13127 22389 13139 22423
rect 13081 22383 13139 22389
rect 14001 22423 14059 22429
rect 14001 22389 14013 22423
rect 14047 22420 14059 22423
rect 14182 22420 14188 22432
rect 14047 22392 14188 22420
rect 14047 22389 14059 22392
rect 14001 22383 14059 22389
rect 14182 22380 14188 22392
rect 14240 22380 14246 22432
rect 14752 22420 14780 22528
rect 14829 22491 14887 22497
rect 14829 22457 14841 22491
rect 14875 22488 14887 22491
rect 14918 22488 14924 22500
rect 14875 22460 14924 22488
rect 14875 22457 14887 22460
rect 14829 22451 14887 22457
rect 14918 22448 14924 22460
rect 14976 22448 14982 22500
rect 15746 22448 15752 22500
rect 15804 22488 15810 22500
rect 16040 22488 16068 22596
rect 16117 22593 16129 22596
rect 16163 22593 16175 22627
rect 16117 22587 16175 22593
rect 16224 22565 16252 22664
rect 16758 22652 16764 22664
rect 16816 22652 16822 22704
rect 16666 22584 16672 22636
rect 16724 22624 16730 22636
rect 16961 22633 16989 22732
rect 17034 22720 17040 22732
rect 17092 22720 17098 22772
rect 17310 22720 17316 22772
rect 17368 22760 17374 22772
rect 20162 22760 20168 22772
rect 17368 22732 20168 22760
rect 17368 22720 17374 22732
rect 20162 22720 20168 22732
rect 20220 22720 20226 22772
rect 21450 22720 21456 22772
rect 21508 22760 21514 22772
rect 21508 22732 22324 22760
rect 21508 22720 21514 22732
rect 18046 22652 18052 22704
rect 18104 22652 18110 22704
rect 18138 22652 18144 22704
rect 18196 22692 18202 22704
rect 18626 22695 18684 22701
rect 18626 22692 18638 22695
rect 18196 22664 18638 22692
rect 18196 22652 18202 22664
rect 18626 22661 18638 22664
rect 18672 22661 18684 22695
rect 18626 22655 18684 22661
rect 19886 22652 19892 22704
rect 19944 22692 19950 22704
rect 21542 22692 21548 22704
rect 19944 22664 21548 22692
rect 19944 22652 19950 22664
rect 21542 22652 21548 22664
rect 21600 22652 21606 22704
rect 22094 22652 22100 22704
rect 22152 22652 22158 22704
rect 22296 22692 22324 22732
rect 22922 22720 22928 22772
rect 22980 22760 22986 22772
rect 23658 22760 23664 22772
rect 22980 22732 23664 22760
rect 22980 22720 22986 22732
rect 23658 22720 23664 22732
rect 23716 22720 23722 22772
rect 24670 22760 24676 22772
rect 24320 22732 24676 22760
rect 23014 22692 23020 22704
rect 22296 22664 22416 22692
rect 16853 22627 16911 22633
rect 16853 22624 16865 22627
rect 16724 22596 16865 22624
rect 16724 22584 16730 22596
rect 16853 22593 16865 22596
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 16946 22627 17004 22633
rect 16946 22593 16958 22627
rect 16992 22593 17004 22627
rect 17129 22627 17187 22633
rect 17129 22624 17141 22627
rect 16946 22587 17004 22593
rect 17052 22596 17141 22624
rect 16209 22559 16267 22565
rect 16209 22525 16221 22559
rect 16255 22556 16267 22559
rect 16298 22556 16304 22568
rect 16255 22528 16304 22556
rect 16255 22525 16267 22528
rect 16209 22519 16267 22525
rect 16298 22516 16304 22528
rect 16356 22516 16362 22568
rect 16482 22516 16488 22568
rect 16540 22556 16546 22568
rect 17052 22556 17080 22596
rect 17129 22593 17141 22596
rect 17175 22593 17187 22627
rect 17129 22587 17187 22593
rect 17218 22584 17224 22636
rect 17276 22584 17282 22636
rect 17402 22633 17408 22636
rect 17359 22627 17408 22633
rect 17359 22593 17371 22627
rect 17405 22593 17408 22627
rect 17359 22587 17408 22593
rect 17402 22584 17408 22587
rect 17460 22584 17466 22636
rect 18064 22556 18092 22652
rect 18156 22596 18736 22624
rect 18156 22565 18184 22596
rect 18708 22568 18736 22596
rect 18874 22584 18880 22636
rect 18932 22624 18938 22636
rect 21266 22624 21272 22636
rect 18932 22596 21272 22624
rect 18932 22584 18938 22596
rect 21266 22584 21272 22596
rect 21324 22584 21330 22636
rect 22112 22624 22140 22652
rect 22388 22633 22416 22664
rect 22664 22664 23020 22692
rect 22664 22633 22692 22664
rect 23014 22652 23020 22664
rect 23072 22652 23078 22704
rect 23676 22692 23704 22720
rect 23845 22695 23903 22701
rect 23676 22664 23796 22692
rect 22281 22627 22339 22633
rect 22112 22614 22232 22624
rect 22281 22614 22293 22627
rect 22112 22596 22293 22614
rect 22204 22593 22293 22596
rect 22327 22593 22339 22627
rect 22204 22587 22339 22593
rect 22373 22627 22431 22633
rect 22373 22593 22385 22627
rect 22419 22593 22431 22627
rect 22373 22587 22431 22593
rect 22557 22627 22615 22633
rect 22557 22593 22569 22627
rect 22603 22593 22615 22627
rect 22557 22587 22615 22593
rect 22649 22627 22707 22633
rect 22649 22593 22661 22627
rect 22695 22593 22707 22627
rect 22649 22587 22707 22593
rect 22204 22586 22324 22587
rect 16540 22528 18092 22556
rect 18141 22559 18199 22565
rect 16540 22516 16546 22528
rect 18141 22525 18153 22559
rect 18187 22525 18199 22559
rect 18141 22519 18199 22525
rect 18414 22516 18420 22568
rect 18472 22516 18478 22568
rect 18509 22559 18567 22565
rect 18509 22525 18521 22559
rect 18555 22525 18567 22559
rect 18509 22519 18567 22525
rect 18524 22488 18552 22519
rect 18690 22516 18696 22568
rect 18748 22516 18754 22568
rect 20714 22516 20720 22568
rect 20772 22556 20778 22568
rect 21358 22556 21364 22568
rect 20772 22528 21364 22556
rect 20772 22516 20778 22528
rect 21358 22516 21364 22528
rect 21416 22556 21422 22568
rect 22572 22556 22600 22587
rect 22830 22584 22836 22636
rect 22888 22624 22894 22636
rect 23661 22627 23719 22633
rect 23661 22624 23673 22627
rect 22888 22596 23673 22624
rect 22888 22584 22894 22596
rect 23661 22593 23673 22596
rect 23707 22593 23719 22627
rect 23768 22624 23796 22664
rect 23845 22661 23857 22695
rect 23891 22692 23903 22695
rect 24210 22692 24216 22704
rect 23891 22664 24216 22692
rect 23891 22661 23903 22664
rect 23845 22655 23903 22661
rect 24210 22652 24216 22664
rect 24268 22652 24274 22704
rect 24320 22701 24348 22732
rect 24670 22720 24676 22732
rect 24728 22720 24734 22772
rect 27522 22720 27528 22772
rect 27580 22720 27586 22772
rect 30834 22760 30840 22772
rect 28092 22732 30840 22760
rect 24305 22695 24363 22701
rect 24305 22661 24317 22695
rect 24351 22661 24363 22695
rect 24305 22655 24363 22661
rect 24486 22652 24492 22704
rect 24544 22692 24550 22704
rect 25038 22692 25044 22704
rect 24544 22664 25044 22692
rect 24544 22652 24550 22664
rect 25038 22652 25044 22664
rect 25096 22652 25102 22704
rect 23937 22627 23995 22633
rect 23937 22624 23949 22627
rect 23768 22596 23949 22624
rect 23661 22587 23719 22593
rect 23937 22593 23949 22596
rect 23983 22593 23995 22627
rect 23937 22587 23995 22593
rect 24026 22584 24032 22636
rect 24084 22584 24090 22636
rect 27540 22624 27568 22720
rect 28092 22633 28120 22732
rect 30834 22720 30840 22732
rect 30892 22720 30898 22772
rect 31754 22720 31760 22772
rect 31812 22760 31818 22772
rect 32490 22760 32496 22772
rect 31812 22732 32496 22760
rect 31812 22720 31818 22732
rect 32490 22720 32496 22732
rect 32548 22720 32554 22772
rect 34793 22763 34851 22769
rect 34793 22729 34805 22763
rect 34839 22760 34851 22763
rect 34882 22760 34888 22772
rect 34839 22732 34888 22760
rect 34839 22729 34851 22732
rect 34793 22723 34851 22729
rect 34882 22720 34888 22732
rect 34940 22720 34946 22772
rect 37458 22760 37464 22772
rect 36214 22732 37464 22760
rect 28442 22652 28448 22704
rect 28500 22652 28506 22704
rect 31202 22692 31208 22704
rect 29196 22664 29960 22692
rect 29196 22636 29224 22664
rect 28077 22627 28135 22633
rect 28077 22624 28089 22627
rect 26252 22596 28089 22624
rect 26252 22568 26280 22596
rect 28077 22593 28089 22596
rect 28123 22593 28135 22627
rect 28077 22587 28135 22593
rect 28258 22584 28264 22636
rect 28316 22584 28322 22636
rect 28626 22584 28632 22636
rect 28684 22624 28690 22636
rect 28684 22596 29145 22624
rect 28684 22584 28690 22596
rect 21416 22528 22600 22556
rect 22940 22528 23980 22556
rect 21416 22516 21422 22528
rect 22940 22488 22968 22528
rect 23952 22500 23980 22528
rect 24486 22516 24492 22568
rect 24544 22556 24550 22568
rect 25041 22559 25099 22565
rect 25041 22556 25053 22559
rect 24544 22528 25053 22556
rect 24544 22516 24550 22528
rect 25041 22525 25053 22528
rect 25087 22525 25099 22559
rect 25041 22519 25099 22525
rect 25590 22516 25596 22568
rect 25648 22516 25654 22568
rect 26234 22516 26240 22568
rect 26292 22516 26298 22568
rect 28276 22556 28304 22584
rect 27586 22528 28304 22556
rect 15804 22460 16068 22488
rect 16132 22460 17632 22488
rect 18524 22460 22968 22488
rect 15804 22448 15810 22460
rect 16132 22420 16160 22460
rect 14752 22392 16160 22420
rect 16206 22380 16212 22432
rect 16264 22380 16270 22432
rect 16758 22380 16764 22432
rect 16816 22420 16822 22432
rect 17218 22420 17224 22432
rect 16816 22392 17224 22420
rect 16816 22380 16822 22392
rect 17218 22380 17224 22392
rect 17276 22380 17282 22432
rect 17402 22380 17408 22432
rect 17460 22420 17466 22432
rect 17497 22423 17555 22429
rect 17497 22420 17509 22423
rect 17460 22392 17509 22420
rect 17460 22380 17466 22392
rect 17497 22389 17509 22392
rect 17543 22389 17555 22423
rect 17604 22420 17632 22460
rect 23014 22448 23020 22500
rect 23072 22488 23078 22500
rect 23842 22488 23848 22500
rect 23072 22460 23848 22488
rect 23072 22448 23078 22460
rect 23842 22448 23848 22460
rect 23900 22448 23906 22500
rect 23934 22448 23940 22500
rect 23992 22448 23998 22500
rect 25608 22488 25636 22516
rect 27586 22488 27614 22528
rect 28718 22516 28724 22568
rect 28776 22556 28782 22568
rect 28776 22528 28994 22556
rect 28776 22516 28782 22528
rect 25608 22460 27614 22488
rect 18785 22423 18843 22429
rect 18785 22420 18797 22423
rect 17604 22392 18797 22420
rect 17497 22383 17555 22389
rect 18785 22389 18797 22392
rect 18831 22389 18843 22423
rect 18785 22383 18843 22389
rect 20806 22380 20812 22432
rect 20864 22420 20870 22432
rect 21266 22420 21272 22432
rect 20864 22392 21272 22420
rect 20864 22380 20870 22392
rect 21266 22380 21272 22392
rect 21324 22380 21330 22432
rect 22094 22380 22100 22432
rect 22152 22380 22158 22432
rect 22186 22380 22192 22432
rect 22244 22420 22250 22432
rect 22738 22420 22744 22432
rect 22244 22392 22744 22420
rect 22244 22380 22250 22392
rect 22738 22380 22744 22392
rect 22796 22380 22802 22432
rect 24210 22380 24216 22432
rect 24268 22380 24274 22432
rect 28966 22420 28994 22528
rect 29117 22488 29145 22596
rect 29178 22584 29184 22636
rect 29236 22584 29242 22636
rect 29638 22584 29644 22636
rect 29696 22584 29702 22636
rect 29932 22633 29960 22664
rect 30116 22664 31208 22692
rect 29917 22627 29975 22633
rect 29917 22593 29929 22627
rect 29963 22593 29975 22627
rect 29917 22587 29975 22593
rect 29454 22516 29460 22568
rect 29512 22516 29518 22568
rect 29733 22559 29791 22565
rect 29733 22525 29745 22559
rect 29779 22556 29791 22559
rect 30116 22556 30144 22664
rect 31202 22652 31208 22664
rect 31260 22652 31266 22704
rect 31297 22695 31355 22701
rect 31297 22661 31309 22695
rect 31343 22692 31355 22695
rect 31662 22692 31668 22704
rect 31343 22664 31668 22692
rect 31343 22661 31355 22664
rect 31297 22655 31355 22661
rect 31662 22652 31668 22664
rect 31720 22692 31726 22704
rect 32214 22692 32220 22704
rect 31720 22664 32220 22692
rect 31720 22652 31726 22664
rect 32214 22652 32220 22664
rect 32272 22652 32278 22704
rect 34054 22652 34060 22704
rect 34112 22692 34118 22704
rect 36214 22701 36242 22732
rect 37458 22720 37464 22732
rect 37516 22720 37522 22772
rect 39853 22763 39911 22769
rect 39853 22729 39865 22763
rect 39899 22760 39911 22763
rect 39942 22760 39948 22772
rect 39899 22732 39948 22760
rect 39899 22729 39911 22732
rect 39853 22723 39911 22729
rect 39942 22720 39948 22732
rect 40000 22720 40006 22772
rect 36199 22695 36257 22701
rect 36199 22692 36211 22695
rect 34112 22664 36211 22692
rect 34112 22652 34118 22664
rect 36199 22661 36211 22664
rect 36245 22661 36257 22695
rect 36199 22655 36257 22661
rect 36630 22652 36636 22704
rect 36688 22692 36694 22704
rect 38654 22692 38660 22704
rect 36688 22664 38660 22692
rect 36688 22652 36694 22664
rect 38654 22652 38660 22664
rect 38712 22692 38718 22704
rect 38749 22695 38807 22701
rect 38749 22692 38761 22695
rect 38712 22664 38761 22692
rect 38712 22652 38718 22664
rect 38749 22661 38761 22664
rect 38795 22661 38807 22695
rect 38749 22655 38807 22661
rect 38838 22652 38844 22704
rect 38896 22652 38902 22704
rect 39316 22664 40724 22692
rect 30190 22584 30196 22636
rect 30248 22584 30254 22636
rect 30285 22627 30343 22633
rect 30285 22593 30297 22627
rect 30331 22593 30343 22627
rect 30285 22587 30343 22593
rect 29779 22528 30144 22556
rect 29779 22525 29791 22528
rect 29733 22519 29791 22525
rect 29748 22488 29776 22519
rect 29117 22460 29776 22488
rect 29825 22491 29883 22497
rect 29825 22457 29837 22491
rect 29871 22488 29883 22491
rect 30006 22488 30012 22500
rect 29871 22460 30012 22488
rect 29871 22457 29883 22460
rect 29825 22451 29883 22457
rect 30006 22448 30012 22460
rect 30064 22448 30070 22500
rect 30208 22488 30236 22584
rect 30300 22556 30328 22587
rect 30374 22584 30380 22636
rect 30432 22624 30438 22636
rect 30561 22627 30619 22633
rect 30561 22624 30573 22627
rect 30432 22596 30573 22624
rect 30432 22584 30438 22596
rect 30561 22593 30573 22596
rect 30607 22624 30619 22627
rect 30650 22624 30656 22636
rect 30607 22596 30656 22624
rect 30607 22593 30619 22596
rect 30561 22587 30619 22593
rect 30650 22584 30656 22596
rect 30708 22584 30714 22636
rect 30742 22584 30748 22636
rect 30800 22584 30806 22636
rect 30837 22627 30895 22633
rect 30837 22593 30849 22627
rect 30883 22624 30895 22627
rect 30926 22624 30932 22636
rect 30883 22596 30932 22624
rect 30883 22593 30895 22596
rect 30837 22587 30895 22593
rect 30926 22584 30932 22596
rect 30984 22624 30990 22636
rect 31386 22624 31392 22636
rect 30984 22596 31392 22624
rect 30984 22584 30990 22596
rect 31386 22584 31392 22596
rect 31444 22584 31450 22636
rect 31481 22627 31539 22633
rect 31481 22593 31493 22627
rect 31527 22593 31539 22627
rect 31481 22587 31539 22593
rect 30760 22556 30788 22584
rect 31018 22556 31024 22568
rect 30300 22528 30788 22556
rect 30944 22528 31024 22556
rect 30377 22491 30435 22497
rect 30377 22488 30389 22491
rect 30208 22460 30389 22488
rect 30377 22457 30389 22460
rect 30423 22457 30435 22491
rect 30377 22451 30435 22457
rect 30466 22448 30472 22500
rect 30524 22448 30530 22500
rect 30101 22423 30159 22429
rect 30101 22420 30113 22423
rect 28966 22392 30113 22420
rect 30101 22389 30113 22392
rect 30147 22389 30159 22423
rect 30101 22383 30159 22389
rect 30190 22380 30196 22432
rect 30248 22420 30254 22432
rect 30576 22420 30604 22528
rect 30248 22392 30604 22420
rect 30248 22380 30254 22392
rect 30650 22380 30656 22432
rect 30708 22420 30714 22432
rect 30944 22429 30972 22528
rect 31018 22516 31024 22528
rect 31076 22516 31082 22568
rect 31496 22556 31524 22587
rect 31570 22584 31576 22636
rect 31628 22584 31634 22636
rect 31846 22584 31852 22636
rect 31904 22624 31910 22636
rect 32122 22624 32128 22636
rect 31904 22596 32128 22624
rect 31904 22584 31910 22596
rect 32122 22584 32128 22596
rect 32180 22584 32186 22636
rect 32493 22627 32551 22633
rect 32493 22593 32505 22627
rect 32539 22593 32551 22627
rect 32493 22587 32551 22593
rect 32508 22556 32536 22587
rect 32674 22584 32680 22636
rect 32732 22584 32738 22636
rect 33226 22584 33232 22636
rect 33284 22584 33290 22636
rect 34514 22584 34520 22636
rect 34572 22624 34578 22636
rect 34701 22627 34759 22633
rect 34701 22624 34713 22627
rect 34572 22596 34713 22624
rect 34572 22584 34578 22596
rect 34701 22593 34713 22596
rect 34747 22593 34759 22627
rect 34701 22587 34759 22593
rect 34885 22627 34943 22633
rect 34885 22593 34897 22627
rect 34931 22624 34943 22627
rect 35342 22624 35348 22636
rect 34931 22596 35348 22624
rect 34931 22593 34943 22596
rect 34885 22587 34943 22593
rect 35342 22584 35348 22596
rect 35400 22584 35406 22636
rect 35802 22624 35808 22636
rect 35452 22596 35808 22624
rect 33244 22556 33272 22584
rect 31496 22528 31616 22556
rect 32508 22528 33272 22556
rect 31588 22488 31616 22528
rect 33870 22516 33876 22568
rect 33928 22556 33934 22568
rect 35452 22556 35480 22596
rect 35802 22584 35808 22596
rect 35860 22624 35866 22636
rect 35897 22627 35955 22633
rect 35897 22624 35909 22627
rect 35860 22596 35909 22624
rect 35860 22584 35866 22596
rect 35897 22593 35909 22596
rect 35943 22593 35955 22627
rect 35897 22587 35955 22593
rect 35989 22627 36047 22633
rect 35989 22593 36001 22627
rect 36035 22593 36047 22627
rect 35989 22587 36047 22593
rect 36081 22627 36139 22633
rect 36081 22593 36093 22627
rect 36127 22593 36139 22627
rect 36081 22587 36139 22593
rect 33928 22528 35480 22556
rect 33928 22516 33934 22528
rect 35526 22516 35532 22568
rect 35584 22556 35590 22568
rect 36004 22556 36032 22587
rect 35584 22528 36032 22556
rect 35584 22516 35590 22528
rect 31588 22460 32628 22488
rect 30929 22423 30987 22429
rect 30929 22420 30941 22423
rect 30708 22392 30941 22420
rect 30708 22380 30714 22392
rect 30929 22389 30941 22392
rect 30975 22389 30987 22423
rect 30929 22383 30987 22389
rect 31018 22380 31024 22432
rect 31076 22420 31082 22432
rect 31297 22423 31355 22429
rect 31297 22420 31309 22423
rect 31076 22392 31309 22420
rect 31076 22380 31082 22392
rect 31297 22389 31309 22392
rect 31343 22389 31355 22423
rect 31297 22383 31355 22389
rect 32490 22380 32496 22432
rect 32548 22380 32554 22432
rect 32600 22420 32628 22460
rect 33226 22448 33232 22500
rect 33284 22488 33290 22500
rect 33778 22488 33784 22500
rect 33284 22460 33784 22488
rect 33284 22448 33290 22460
rect 33778 22448 33784 22460
rect 33836 22448 33842 22500
rect 34422 22448 34428 22500
rect 34480 22488 34486 22500
rect 36096 22488 36124 22587
rect 36354 22584 36360 22636
rect 36412 22584 36418 22636
rect 38473 22627 38531 22633
rect 38473 22593 38485 22627
rect 38519 22593 38531 22627
rect 38473 22587 38531 22593
rect 38488 22556 38516 22587
rect 38562 22584 38568 22636
rect 38620 22624 38626 22636
rect 39022 22633 39028 22636
rect 38979 22627 39028 22633
rect 38620 22596 38665 22624
rect 38620 22584 38626 22596
rect 38979 22593 38991 22627
rect 39025 22593 39028 22627
rect 38979 22587 39028 22593
rect 39022 22584 39028 22587
rect 39080 22584 39086 22636
rect 39114 22556 39120 22568
rect 38488 22528 39120 22556
rect 39114 22516 39120 22528
rect 39172 22556 39178 22568
rect 39316 22556 39344 22664
rect 39390 22584 39396 22636
rect 39448 22584 39454 22636
rect 39669 22627 39727 22633
rect 39669 22593 39681 22627
rect 39715 22593 39727 22627
rect 39669 22587 39727 22593
rect 39172 22528 39344 22556
rect 39172 22516 39178 22528
rect 39482 22516 39488 22568
rect 39540 22516 39546 22568
rect 34480 22460 36124 22488
rect 34480 22448 34486 22460
rect 38838 22448 38844 22500
rect 38896 22488 38902 22500
rect 39684 22488 39712 22587
rect 40696 22568 40724 22664
rect 40678 22516 40684 22568
rect 40736 22516 40742 22568
rect 38896 22460 39712 22488
rect 38896 22448 38902 22460
rect 35342 22420 35348 22432
rect 32600 22392 35348 22420
rect 35342 22380 35348 22392
rect 35400 22380 35406 22432
rect 35713 22423 35771 22429
rect 35713 22389 35725 22423
rect 35759 22420 35771 22423
rect 37826 22420 37832 22432
rect 35759 22392 37832 22420
rect 35759 22389 35771 22392
rect 35713 22383 35771 22389
rect 37826 22380 37832 22392
rect 37884 22380 37890 22432
rect 39114 22380 39120 22432
rect 39172 22380 39178 22432
rect 39206 22380 39212 22432
rect 39264 22420 39270 22432
rect 39393 22423 39451 22429
rect 39393 22420 39405 22423
rect 39264 22392 39405 22420
rect 39264 22380 39270 22392
rect 39393 22389 39405 22392
rect 39439 22420 39451 22423
rect 39850 22420 39856 22432
rect 39439 22392 39856 22420
rect 39439 22389 39451 22392
rect 39393 22383 39451 22389
rect 39850 22380 39856 22392
rect 39908 22380 39914 22432
rect 1104 22330 41400 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 41400 22330
rect 1104 22256 41400 22278
rect 4525 22219 4583 22225
rect 4525 22185 4537 22219
rect 4571 22216 4583 22219
rect 4614 22216 4620 22228
rect 4571 22188 4620 22216
rect 4571 22185 4583 22188
rect 4525 22179 4583 22185
rect 4614 22176 4620 22188
rect 4672 22176 4678 22228
rect 5810 22176 5816 22228
rect 5868 22216 5874 22228
rect 6086 22216 6092 22228
rect 5868 22188 6092 22216
rect 5868 22176 5874 22188
rect 6086 22176 6092 22188
rect 6144 22176 6150 22228
rect 7190 22176 7196 22228
rect 7248 22176 7254 22228
rect 9214 22176 9220 22228
rect 9272 22176 9278 22228
rect 11422 22176 11428 22228
rect 11480 22216 11486 22228
rect 12158 22216 12164 22228
rect 11480 22188 12164 22216
rect 11480 22176 11486 22188
rect 12158 22176 12164 22188
rect 12216 22176 12222 22228
rect 12710 22176 12716 22228
rect 12768 22176 12774 22228
rect 13633 22219 13691 22225
rect 13633 22185 13645 22219
rect 13679 22216 13691 22219
rect 13814 22216 13820 22228
rect 13679 22188 13820 22216
rect 13679 22185 13691 22188
rect 13633 22179 13691 22185
rect 13814 22176 13820 22188
rect 13872 22176 13878 22228
rect 14734 22176 14740 22228
rect 14792 22176 14798 22228
rect 21634 22216 21640 22228
rect 14844 22188 21640 22216
rect 3142 22108 3148 22160
rect 3200 22148 3206 22160
rect 3200 22120 5488 22148
rect 3200 22108 3206 22120
rect 3053 22083 3111 22089
rect 3053 22049 3065 22083
rect 3099 22080 3111 22083
rect 3160 22080 3188 22108
rect 5460 22092 5488 22120
rect 5442 22080 5448 22092
rect 3099 22052 3188 22080
rect 5403 22052 5448 22080
rect 3099 22049 3111 22052
rect 3053 22043 3111 22049
rect 5442 22040 5448 22052
rect 5500 22040 5506 22092
rect 5902 22040 5908 22092
rect 5960 22040 5966 22092
rect 7098 22040 7104 22092
rect 7156 22080 7162 22092
rect 7466 22080 7472 22092
rect 7156 22052 7472 22080
rect 7156 22040 7162 22052
rect 7466 22040 7472 22052
rect 7524 22040 7530 22092
rect 4709 22015 4767 22021
rect 4709 21981 4721 22015
rect 4755 21981 4767 22015
rect 4709 21975 4767 21981
rect 5261 22015 5319 22021
rect 5261 21981 5273 22015
rect 5307 22012 5319 22015
rect 5920 22012 5948 22040
rect 5307 21984 5948 22012
rect 7377 22015 7435 22021
rect 5307 21981 5319 21984
rect 5261 21975 5319 21981
rect 7377 21981 7389 22015
rect 7423 22012 7435 22015
rect 8386 22012 8392 22024
rect 7423 21984 8392 22012
rect 7423 21981 7435 21984
rect 7377 21975 7435 21981
rect 4614 21944 4620 21956
rect 2884 21916 4620 21944
rect 2884 21888 2912 21916
rect 4614 21904 4620 21916
rect 4672 21904 4678 21956
rect 2498 21836 2504 21888
rect 2556 21836 2562 21888
rect 2866 21836 2872 21888
rect 2924 21836 2930 21888
rect 2961 21879 3019 21885
rect 2961 21845 2973 21879
rect 3007 21876 3019 21879
rect 3142 21876 3148 21888
rect 3007 21848 3148 21876
rect 3007 21845 3019 21848
rect 2961 21839 3019 21845
rect 3142 21836 3148 21848
rect 3200 21836 3206 21888
rect 4724 21876 4752 21975
rect 8386 21972 8392 21984
rect 8444 21972 8450 22024
rect 8846 21972 8852 22024
rect 8904 22012 8910 22024
rect 9232 22021 9260 22176
rect 9766 22108 9772 22160
rect 9824 22148 9830 22160
rect 12728 22148 12756 22176
rect 9824 22120 12756 22148
rect 9824 22108 9830 22120
rect 9861 22083 9919 22089
rect 9861 22049 9873 22083
rect 9907 22080 9919 22083
rect 10134 22080 10140 22092
rect 9907 22052 10140 22080
rect 9907 22049 9919 22052
rect 9861 22043 9919 22049
rect 10134 22040 10140 22052
rect 10192 22040 10198 22092
rect 10686 22040 10692 22092
rect 10744 22080 10750 22092
rect 10744 22052 11009 22080
rect 10744 22040 10750 22052
rect 9033 22015 9091 22021
rect 9033 22012 9045 22015
rect 8904 21984 9045 22012
rect 8904 21972 8910 21984
rect 9033 21981 9045 21984
rect 9079 21981 9091 22015
rect 9033 21975 9091 21981
rect 9181 22015 9260 22021
rect 9181 21981 9193 22015
rect 9227 21984 9260 22015
rect 9227 21981 9239 21984
rect 9181 21975 9239 21981
rect 9306 21972 9312 22024
rect 9364 21972 9370 22024
rect 9582 22021 9588 22024
rect 9539 22015 9588 22021
rect 9539 21981 9551 22015
rect 9585 21981 9588 22015
rect 9539 21975 9588 21981
rect 9582 21972 9588 21975
rect 9640 21972 9646 22024
rect 9766 21972 9772 22024
rect 9824 21972 9830 22024
rect 10042 21972 10048 22024
rect 10100 21972 10106 22024
rect 10229 22015 10287 22021
rect 10229 21981 10241 22015
rect 10275 21981 10287 22015
rect 10229 21975 10287 21981
rect 5350 21944 5356 21956
rect 5184 21916 5356 21944
rect 4801 21879 4859 21885
rect 4801 21876 4813 21879
rect 4724 21848 4813 21876
rect 4801 21845 4813 21848
rect 4847 21845 4859 21879
rect 4801 21839 4859 21845
rect 4982 21836 4988 21888
rect 5040 21876 5046 21888
rect 5184 21885 5212 21916
rect 5350 21904 5356 21916
rect 5408 21904 5414 21956
rect 5721 21947 5779 21953
rect 5721 21913 5733 21947
rect 5767 21913 5779 21947
rect 5721 21907 5779 21913
rect 5169 21879 5227 21885
rect 5169 21876 5181 21879
rect 5040 21848 5181 21876
rect 5040 21836 5046 21848
rect 5169 21845 5181 21848
rect 5215 21845 5227 21879
rect 5169 21839 5227 21845
rect 5626 21836 5632 21888
rect 5684 21876 5690 21888
rect 5736 21876 5764 21907
rect 5810 21904 5816 21956
rect 5868 21944 5874 21956
rect 9401 21947 9459 21953
rect 9401 21944 9413 21947
rect 5868 21916 9413 21944
rect 5868 21904 5874 21916
rect 9401 21913 9413 21916
rect 9447 21913 9459 21947
rect 9401 21907 9459 21913
rect 7282 21876 7288 21888
rect 5684 21848 7288 21876
rect 5684 21836 5690 21848
rect 7282 21836 7288 21848
rect 7340 21836 7346 21888
rect 9674 21836 9680 21888
rect 9732 21836 9738 21888
rect 10244 21876 10272 21975
rect 10594 21972 10600 22024
rect 10652 21972 10658 22024
rect 10781 22015 10839 22021
rect 10781 21981 10793 22015
rect 10827 21981 10839 22015
rect 10781 21975 10839 21981
rect 10686 21904 10692 21956
rect 10744 21944 10750 21956
rect 10796 21944 10824 21975
rect 10870 21972 10876 22024
rect 10928 21972 10934 22024
rect 10981 22021 11009 22052
rect 11238 22040 11244 22092
rect 11296 22080 11302 22092
rect 11296 22052 11381 22080
rect 11296 22040 11302 22052
rect 11353 22021 11381 22052
rect 10966 22015 11024 22021
rect 10966 21981 10978 22015
rect 11012 21981 11024 22015
rect 11338 22015 11396 22021
rect 11338 22012 11350 22015
rect 10966 21975 11024 21981
rect 11072 21984 11350 22012
rect 11072 21944 11100 21984
rect 11338 21981 11350 21984
rect 11384 21981 11396 22015
rect 11338 21975 11396 21981
rect 11974 21972 11980 22024
rect 12032 21972 12038 22024
rect 12158 22021 12164 22024
rect 12125 22015 12164 22021
rect 12125 21981 12137 22015
rect 12125 21975 12164 21981
rect 12158 21972 12164 21975
rect 12216 21972 12222 22024
rect 12268 22021 12296 22120
rect 12802 22108 12808 22160
rect 12860 22148 12866 22160
rect 13078 22148 13084 22160
rect 12860 22120 13084 22148
rect 12860 22108 12866 22120
rect 13078 22108 13084 22120
rect 13136 22108 13142 22160
rect 13357 22151 13415 22157
rect 13357 22117 13369 22151
rect 13403 22117 13415 22151
rect 13357 22111 13415 22117
rect 12636 22052 13032 22080
rect 12253 22015 12311 22021
rect 12253 21981 12265 22015
rect 12299 21981 12311 22015
rect 12253 21975 12311 21981
rect 12434 21972 12440 22024
rect 12492 22021 12498 22024
rect 12492 22012 12500 22021
rect 12492 21984 12537 22012
rect 12492 21975 12500 21984
rect 12492 21972 12498 21975
rect 10744 21916 11100 21944
rect 10744 21904 10750 21916
rect 11146 21904 11152 21956
rect 11204 21904 11210 21956
rect 11238 21904 11244 21956
rect 11296 21904 11302 21956
rect 11348 21916 11836 21944
rect 10410 21876 10416 21888
rect 10244 21848 10416 21876
rect 10410 21836 10416 21848
rect 10468 21876 10474 21888
rect 11164 21876 11192 21904
rect 11348 21876 11376 21916
rect 10468 21848 11376 21876
rect 10468 21836 10474 21848
rect 11514 21836 11520 21888
rect 11572 21836 11578 21888
rect 11808 21876 11836 21916
rect 11882 21904 11888 21956
rect 11940 21944 11946 21956
rect 12345 21947 12403 21953
rect 12345 21944 12357 21947
rect 11940 21916 12357 21944
rect 11940 21904 11946 21916
rect 12345 21913 12357 21916
rect 12391 21913 12403 21947
rect 12636 21944 12664 22052
rect 12713 22015 12771 22021
rect 12713 21981 12725 22015
rect 12759 21981 12771 22015
rect 12713 21975 12771 21981
rect 12806 22015 12864 22021
rect 12806 21981 12818 22015
rect 12852 21981 12864 22015
rect 12806 21975 12864 21981
rect 12345 21907 12403 21913
rect 12452 21916 12664 21944
rect 12452 21876 12480 21916
rect 11808 21848 12480 21876
rect 12621 21879 12679 21885
rect 12621 21845 12633 21879
rect 12667 21876 12679 21879
rect 12728 21876 12756 21975
rect 12667 21848 12756 21876
rect 12820 21876 12848 21975
rect 13004 21953 13032 22052
rect 13178 22015 13236 22021
rect 13178 21981 13190 22015
rect 13224 21981 13236 22015
rect 13372 22012 13400 22111
rect 13722 22108 13728 22160
rect 13780 22148 13786 22160
rect 14844 22148 14872 22188
rect 21634 22176 21640 22188
rect 21692 22176 21698 22228
rect 22002 22176 22008 22228
rect 22060 22176 22066 22228
rect 22278 22176 22284 22228
rect 22336 22216 22342 22228
rect 26145 22219 26203 22225
rect 26145 22216 26157 22219
rect 22336 22188 26157 22216
rect 22336 22176 22342 22188
rect 26145 22185 26157 22188
rect 26191 22185 26203 22219
rect 26145 22179 26203 22185
rect 29086 22176 29092 22228
rect 29144 22216 29150 22228
rect 29270 22216 29276 22228
rect 29144 22188 29276 22216
rect 29144 22176 29150 22188
rect 29270 22176 29276 22188
rect 29328 22176 29334 22228
rect 29454 22176 29460 22228
rect 29512 22216 29518 22228
rect 29917 22219 29975 22225
rect 29917 22216 29929 22219
rect 29512 22188 29929 22216
rect 29512 22176 29518 22188
rect 29917 22185 29929 22188
rect 29963 22185 29975 22219
rect 29917 22179 29975 22185
rect 30466 22176 30472 22228
rect 30524 22216 30530 22228
rect 30650 22216 30656 22228
rect 30524 22188 30656 22216
rect 30524 22176 30530 22188
rect 30650 22176 30656 22188
rect 30708 22176 30714 22228
rect 30834 22176 30840 22228
rect 30892 22216 30898 22228
rect 31202 22216 31208 22228
rect 30892 22188 31208 22216
rect 30892 22176 30898 22188
rect 31202 22176 31208 22188
rect 31260 22176 31266 22228
rect 31570 22176 31576 22228
rect 31628 22176 31634 22228
rect 35526 22176 35532 22228
rect 35584 22216 35590 22228
rect 35802 22216 35808 22228
rect 35584 22188 35808 22216
rect 35584 22176 35590 22188
rect 35802 22176 35808 22188
rect 35860 22176 35866 22228
rect 39390 22176 39396 22228
rect 39448 22176 39454 22228
rect 13780 22120 14872 22148
rect 13780 22108 13786 22120
rect 19334 22108 19340 22160
rect 19392 22108 19398 22160
rect 22020 22148 22048 22176
rect 20318 22120 22048 22148
rect 13556 22052 14642 22080
rect 13449 22015 13507 22021
rect 13449 22012 13461 22015
rect 13372 21984 13461 22012
rect 13178 21975 13236 21981
rect 13449 21981 13461 21984
rect 13495 21981 13507 22015
rect 13449 21975 13507 21981
rect 12989 21947 13047 21953
rect 12989 21913 13001 21947
rect 13035 21913 13047 21947
rect 12989 21907 13047 21913
rect 12894 21876 12900 21888
rect 12820 21848 12900 21876
rect 12667 21845 12679 21848
rect 12621 21839 12679 21845
rect 12894 21836 12900 21848
rect 12952 21836 12958 21888
rect 13004 21876 13032 21907
rect 13078 21904 13084 21956
rect 13136 21904 13142 21956
rect 13193 21944 13221 21975
rect 13354 21944 13360 21956
rect 13193 21916 13360 21944
rect 13354 21904 13360 21916
rect 13412 21944 13418 21956
rect 13556 21944 13584 22052
rect 14090 21972 14096 22024
rect 14148 21972 14154 22024
rect 14614 22021 14642 22052
rect 17402 22040 17408 22092
rect 17460 22040 17466 22092
rect 19352 22080 19380 22108
rect 19797 22083 19855 22089
rect 19797 22080 19809 22083
rect 18708 22052 19012 22080
rect 19352 22052 19809 22080
rect 18708 22024 18736 22052
rect 14186 22015 14244 22021
rect 14186 21981 14198 22015
rect 14232 21981 14244 22015
rect 14186 21975 14244 21981
rect 14599 22015 14657 22021
rect 14599 21981 14611 22015
rect 14645 22012 14657 22015
rect 17310 22012 17316 22024
rect 14645 21984 17316 22012
rect 14645 21981 14657 21984
rect 14599 21975 14657 21981
rect 14200 21944 14228 21975
rect 17310 21972 17316 21984
rect 17368 21972 17374 22024
rect 17770 21972 17776 22024
rect 17828 21972 17834 22024
rect 17954 21972 17960 22024
rect 18012 21972 18018 22024
rect 18046 21972 18052 22024
rect 18104 21972 18110 22024
rect 18325 22015 18383 22021
rect 18325 21981 18337 22015
rect 18371 22012 18383 22015
rect 18414 22012 18420 22024
rect 18371 21984 18420 22012
rect 18371 21981 18383 21984
rect 18325 21975 18383 21981
rect 18414 21972 18420 21984
rect 18472 21972 18478 22024
rect 18506 21972 18512 22024
rect 18564 21972 18570 22024
rect 18690 21972 18696 22024
rect 18748 21972 18754 22024
rect 18874 21972 18880 22024
rect 18932 21972 18938 22024
rect 18984 22021 19012 22052
rect 19797 22049 19809 22052
rect 19843 22049 19855 22083
rect 19797 22043 19855 22049
rect 19886 22040 19892 22092
rect 19944 22080 19950 22092
rect 19944 22052 20116 22080
rect 19944 22040 19950 22052
rect 18969 22015 19027 22021
rect 18969 21981 18981 22015
rect 19015 21981 19027 22015
rect 18969 21975 19027 21981
rect 14274 21944 14280 21956
rect 13412 21916 13584 21944
rect 13648 21916 14044 21944
rect 14200 21916 14280 21944
rect 13412 21904 13418 21916
rect 13648 21876 13676 21916
rect 13004 21848 13676 21876
rect 13906 21836 13912 21888
rect 13964 21836 13970 21888
rect 14016 21876 14044 21916
rect 14274 21904 14280 21916
rect 14332 21904 14338 21956
rect 14369 21947 14427 21953
rect 14369 21913 14381 21947
rect 14415 21913 14427 21947
rect 14369 21907 14427 21913
rect 14384 21876 14412 21907
rect 14458 21904 14464 21956
rect 14516 21904 14522 21956
rect 16482 21904 16488 21956
rect 16540 21904 16546 21956
rect 17402 21904 17408 21956
rect 17460 21904 17466 21956
rect 17972 21944 18000 21972
rect 18141 21947 18199 21953
rect 18141 21944 18153 21947
rect 17972 21916 18153 21944
rect 18141 21913 18153 21916
rect 18187 21913 18199 21947
rect 18524 21944 18552 21972
rect 19150 21944 19156 21956
rect 18524 21916 19156 21944
rect 18141 21907 18199 21913
rect 19150 21904 19156 21916
rect 19208 21944 19214 21956
rect 19904 21944 19932 22040
rect 20088 22021 20116 22052
rect 20318 22021 20346 22120
rect 20441 22083 20499 22089
rect 20441 22049 20453 22083
rect 20487 22080 20499 22083
rect 20487 22052 20853 22080
rect 20487 22049 20499 22052
rect 20441 22043 20499 22049
rect 19981 22015 20039 22021
rect 19981 21981 19993 22015
rect 20027 21981 20039 22015
rect 19981 21975 20039 21981
rect 20073 22015 20131 22021
rect 20073 21981 20085 22015
rect 20119 21981 20131 22015
rect 20073 21975 20131 21981
rect 20303 22015 20361 22021
rect 20303 21981 20315 22015
rect 20349 21981 20361 22015
rect 20303 21975 20361 21981
rect 19208 21916 19932 21944
rect 19208 21904 19214 21916
rect 16500 21876 16528 21904
rect 14016 21848 16528 21876
rect 17420 21876 17448 21904
rect 19996 21888 20024 21975
rect 20622 21972 20628 22024
rect 20680 22012 20686 22024
rect 20825 22021 20853 22052
rect 20990 22021 20996 22024
rect 20717 22015 20775 22021
rect 20717 22012 20729 22015
rect 20680 21984 20729 22012
rect 20680 21972 20686 21984
rect 20717 21981 20729 21984
rect 20763 21981 20775 22015
rect 20717 21975 20775 21981
rect 20810 22015 20868 22021
rect 20810 21981 20822 22015
rect 20856 21981 20868 22015
rect 20947 22015 20996 22021
rect 20947 22014 20959 22015
rect 20916 21984 20959 22014
rect 20810 21975 20868 21981
rect 20947 21981 20959 21984
rect 20993 21981 20996 22015
rect 20947 21975 20996 21981
rect 20162 21904 20168 21956
rect 20220 21904 20226 21956
rect 17497 21879 17555 21885
rect 17497 21876 17509 21879
rect 17420 21848 17509 21876
rect 17497 21845 17509 21848
rect 17543 21845 17555 21879
rect 17497 21839 17555 21845
rect 19978 21836 19984 21888
rect 20036 21836 20042 21888
rect 20438 21836 20444 21888
rect 20496 21876 20502 21888
rect 20825 21876 20853 21975
rect 20990 21972 20996 21975
rect 21048 21972 21054 22024
rect 21201 22015 21259 22021
rect 21201 21981 21213 22015
rect 21247 22012 21259 22015
rect 21247 22009 21266 22012
rect 21376 22009 21404 22120
rect 22094 22108 22100 22160
rect 22152 22148 22158 22160
rect 22833 22151 22891 22157
rect 22833 22148 22845 22151
rect 22152 22120 22845 22148
rect 22152 22108 22158 22120
rect 22833 22117 22845 22120
rect 22879 22117 22891 22151
rect 22833 22111 22891 22117
rect 22925 22151 22983 22157
rect 22925 22117 22937 22151
rect 22971 22148 22983 22151
rect 23014 22148 23020 22160
rect 22971 22120 23020 22148
rect 22971 22117 22983 22120
rect 22925 22111 22983 22117
rect 23014 22108 23020 22120
rect 23072 22108 23078 22160
rect 23198 22108 23204 22160
rect 23256 22108 23262 22160
rect 24118 22108 24124 22160
rect 24176 22108 24182 22160
rect 24673 22151 24731 22157
rect 24673 22117 24685 22151
rect 24719 22148 24731 22151
rect 24854 22148 24860 22160
rect 24719 22120 24860 22148
rect 24719 22117 24731 22120
rect 24673 22111 24731 22117
rect 24854 22108 24860 22120
rect 24912 22108 24918 22160
rect 25314 22108 25320 22160
rect 25372 22108 25378 22160
rect 25498 22148 25504 22160
rect 25424 22120 25504 22148
rect 22741 22083 22799 22089
rect 22741 22049 22753 22083
rect 22787 22080 22799 22083
rect 23216 22080 23244 22108
rect 22787 22052 23244 22080
rect 24136 22080 24164 22108
rect 24765 22083 24823 22089
rect 24765 22080 24777 22083
rect 24136 22052 24777 22080
rect 22787 22049 22799 22052
rect 22741 22043 22799 22049
rect 24765 22049 24777 22052
rect 24811 22049 24823 22083
rect 24765 22043 24823 22049
rect 21247 21981 21404 22009
rect 21453 22015 21511 22021
rect 21453 21981 21465 22015
rect 21499 22012 21511 22015
rect 21818 22012 21824 22024
rect 21499 21984 21824 22012
rect 21499 21981 21511 21984
rect 21201 21975 21259 21981
rect 21453 21975 21511 21981
rect 21818 21972 21824 21984
rect 21876 22012 21882 22024
rect 22097 22015 22155 22021
rect 22097 22012 22109 22015
rect 21876 21984 22109 22012
rect 21876 21972 21882 21984
rect 22097 21981 22109 21984
rect 22143 21981 22155 22015
rect 22097 21975 22155 21981
rect 22281 22015 22339 22021
rect 22281 21981 22293 22015
rect 22327 21981 22339 22015
rect 22281 21975 22339 21981
rect 22373 22015 22431 22021
rect 22373 21981 22385 22015
rect 22419 22012 22431 22015
rect 22462 22012 22468 22024
rect 22419 21984 22468 22012
rect 22419 21981 22431 21984
rect 22373 21975 22431 21981
rect 21085 21947 21143 21953
rect 21085 21913 21097 21947
rect 21131 21913 21143 21947
rect 22296 21944 22324 21975
rect 22462 21972 22468 21984
rect 22520 21972 22526 22024
rect 22830 21972 22836 22024
rect 22888 22012 22894 22024
rect 23017 22015 23075 22021
rect 23017 22012 23029 22015
rect 22888 21984 23029 22012
rect 22888 21972 22894 21984
rect 23017 21981 23029 21984
rect 23063 21981 23075 22015
rect 23017 21975 23075 21981
rect 23201 22015 23259 22021
rect 23201 21981 23213 22015
rect 23247 22012 23259 22015
rect 23290 22012 23296 22024
rect 23247 21984 23296 22012
rect 23247 21981 23259 21984
rect 23201 21975 23259 21981
rect 23290 21972 23296 21984
rect 23348 21972 23354 22024
rect 23934 21972 23940 22024
rect 23992 21972 23998 22024
rect 24394 21972 24400 22024
rect 24452 22012 24458 22024
rect 24581 22015 24639 22021
rect 24581 22012 24593 22015
rect 24452 21984 24593 22012
rect 24452 21972 24458 21984
rect 24581 21981 24593 21984
rect 24627 21981 24639 22015
rect 24581 21975 24639 21981
rect 24857 22015 24915 22021
rect 24857 21981 24869 22015
rect 24903 22012 24915 22015
rect 25424 22012 25452 22120
rect 25498 22108 25504 22120
rect 25556 22108 25562 22160
rect 25593 22151 25651 22157
rect 25593 22117 25605 22151
rect 25639 22148 25651 22151
rect 26050 22148 26056 22160
rect 25639 22120 26056 22148
rect 25639 22117 25651 22120
rect 25593 22111 25651 22117
rect 26050 22108 26056 22120
rect 26108 22108 26114 22160
rect 27062 22148 27068 22160
rect 26712 22120 27068 22148
rect 26712 22080 26740 22120
rect 27062 22108 27068 22120
rect 27120 22108 27126 22160
rect 29546 22148 29552 22160
rect 29288 22120 29552 22148
rect 25516 22052 26096 22080
rect 25516 22021 25544 22052
rect 24903 21984 25452 22012
rect 25501 22015 25559 22021
rect 24903 21981 24915 21984
rect 24857 21975 24915 21981
rect 25501 21981 25513 22015
rect 25547 21981 25559 22015
rect 25501 21975 25559 21981
rect 25685 22015 25743 22021
rect 25685 21981 25697 22015
rect 25731 21981 25743 22015
rect 25685 21975 25743 21981
rect 23566 21944 23572 21956
rect 21085 21907 21143 21913
rect 21652 21916 22048 21944
rect 22296 21916 23572 21944
rect 20496 21848 20853 21876
rect 20496 21836 20502 21848
rect 20990 21836 20996 21888
rect 21048 21876 21054 21888
rect 21100 21876 21128 21907
rect 21652 21888 21680 21916
rect 22020 21888 22048 21916
rect 23566 21904 23572 21916
rect 23624 21904 23630 21956
rect 23753 21947 23811 21953
rect 23753 21913 23765 21947
rect 23799 21944 23811 21947
rect 23842 21944 23848 21956
rect 23799 21916 23848 21944
rect 23799 21913 23811 21916
rect 23753 21907 23811 21913
rect 23842 21904 23848 21916
rect 23900 21904 23906 21956
rect 25222 21904 25228 21956
rect 25280 21904 25286 21956
rect 21048 21848 21128 21876
rect 21361 21879 21419 21885
rect 21048 21836 21054 21848
rect 21361 21845 21373 21879
rect 21407 21876 21419 21879
rect 21542 21876 21548 21888
rect 21407 21848 21548 21876
rect 21407 21845 21419 21848
rect 21361 21839 21419 21845
rect 21542 21836 21548 21848
rect 21600 21836 21606 21888
rect 21634 21836 21640 21888
rect 21692 21836 21698 21888
rect 21726 21836 21732 21888
rect 21784 21876 21790 21888
rect 21913 21879 21971 21885
rect 21913 21876 21925 21879
rect 21784 21848 21925 21876
rect 21784 21836 21790 21848
rect 21913 21845 21925 21848
rect 21959 21845 21971 21879
rect 21913 21839 21971 21845
rect 22002 21836 22008 21888
rect 22060 21836 22066 21888
rect 22462 21836 22468 21888
rect 22520 21836 22526 21888
rect 23014 21836 23020 21888
rect 23072 21876 23078 21888
rect 24121 21879 24179 21885
rect 24121 21876 24133 21879
rect 23072 21848 24133 21876
rect 23072 21836 23078 21848
rect 24121 21845 24133 21848
rect 24167 21845 24179 21879
rect 24121 21839 24179 21845
rect 24394 21836 24400 21888
rect 24452 21836 24458 21888
rect 25240 21876 25268 21904
rect 25590 21876 25596 21888
rect 25240 21848 25596 21876
rect 25590 21836 25596 21848
rect 25648 21836 25654 21888
rect 25700 21876 25728 21975
rect 25774 21972 25780 22024
rect 25832 21972 25838 22024
rect 25958 21972 25964 22024
rect 26016 21972 26022 22024
rect 26068 21956 26096 22052
rect 26344 22052 26740 22080
rect 26344 22024 26372 22052
rect 26326 21972 26332 22024
rect 26384 21972 26390 22024
rect 26418 21972 26424 22024
rect 26476 21972 26482 22024
rect 26712 22021 26740 22052
rect 26789 22083 26847 22089
rect 26789 22049 26801 22083
rect 26835 22080 26847 22083
rect 27540 22080 27844 22094
rect 29288 22092 29316 22120
rect 29546 22108 29552 22120
rect 29604 22148 29610 22160
rect 30101 22151 30159 22157
rect 30101 22148 30113 22151
rect 29604 22120 30113 22148
rect 29604 22108 29610 22120
rect 30101 22117 30113 22120
rect 30147 22117 30159 22151
rect 30101 22111 30159 22117
rect 28721 22083 28779 22089
rect 28721 22080 28733 22083
rect 26835 22066 28733 22080
rect 26835 22052 27568 22066
rect 27816 22052 28733 22066
rect 26835 22049 26847 22052
rect 26789 22043 26847 22049
rect 28721 22049 28733 22052
rect 28767 22049 28779 22083
rect 28721 22043 28779 22049
rect 29270 22040 29276 22092
rect 29328 22040 29334 22092
rect 30926 22080 30932 22092
rect 29840 22052 30932 22080
rect 26697 22015 26755 22021
rect 26697 21981 26709 22015
rect 26743 21981 26755 22015
rect 26697 21975 26755 21981
rect 27062 21972 27068 22024
rect 27120 21972 27126 22024
rect 27157 22015 27215 22021
rect 27157 21981 27169 22015
rect 27203 21981 27215 22015
rect 27157 21975 27215 21981
rect 26050 21904 26056 21956
rect 26108 21904 26114 21956
rect 26436 21944 26464 21972
rect 27172 21944 27200 21975
rect 27338 21972 27344 22024
rect 27396 22012 27402 22024
rect 27525 22015 27583 22021
rect 27525 22012 27537 22015
rect 27396 21984 27537 22012
rect 27396 21972 27402 21984
rect 27525 21981 27537 21984
rect 27571 21981 27583 22015
rect 27525 21975 27583 21981
rect 27893 22015 27951 22021
rect 27893 21981 27905 22015
rect 27939 21981 27951 22015
rect 27893 21975 27951 21981
rect 26436 21916 27200 21944
rect 27430 21904 27436 21956
rect 27488 21904 27494 21956
rect 27614 21904 27620 21956
rect 27672 21904 27678 21956
rect 27709 21947 27767 21953
rect 27709 21913 27721 21947
rect 27755 21913 27767 21947
rect 27908 21944 27936 21975
rect 27982 21972 27988 22024
rect 28040 22012 28046 22024
rect 28040 21984 28212 22012
rect 28040 21972 28046 21984
rect 28184 21944 28212 21984
rect 28258 21972 28264 22024
rect 28316 21972 28322 22024
rect 28534 21972 28540 22024
rect 28592 21972 28598 22024
rect 28626 21972 28632 22024
rect 28684 21972 28690 22024
rect 29840 22021 29868 22052
rect 30926 22040 30932 22052
rect 30984 22040 30990 22092
rect 31588 22080 31616 22176
rect 32030 22108 32036 22160
rect 32088 22148 32094 22160
rect 33318 22148 33324 22160
rect 32088 22120 33324 22148
rect 32088 22108 32094 22120
rect 33318 22108 33324 22120
rect 33376 22108 33382 22160
rect 39408 22148 39436 22176
rect 35866 22120 39436 22148
rect 33689 22083 33747 22089
rect 31404 22052 31708 22080
rect 28813 22015 28871 22021
rect 28813 21981 28825 22015
rect 28859 22012 28871 22015
rect 29549 22015 29607 22021
rect 29549 22012 29561 22015
rect 28859 21984 29561 22012
rect 28859 21981 28871 21984
rect 28813 21975 28871 21981
rect 29549 21981 29561 21984
rect 29595 21981 29607 22015
rect 29549 21975 29607 21981
rect 29825 22015 29883 22021
rect 29825 21981 29837 22015
rect 29871 21981 29883 22015
rect 29825 21975 29883 21981
rect 30009 22015 30067 22021
rect 30009 21981 30021 22015
rect 30055 21981 30067 22015
rect 30009 21975 30067 21981
rect 28718 21944 28724 21956
rect 27908 21916 28120 21944
rect 28184 21916 28724 21944
rect 27709 21907 27767 21913
rect 27341 21879 27399 21885
rect 27341 21876 27353 21879
rect 25700 21848 27353 21876
rect 27341 21845 27353 21848
rect 27387 21845 27399 21879
rect 27448 21876 27476 21904
rect 27724 21876 27752 21907
rect 28092 21888 28120 21916
rect 28718 21904 28724 21916
rect 28776 21904 28782 21956
rect 29086 21904 29092 21956
rect 29144 21944 29150 21956
rect 30024 21944 30052 21975
rect 30098 21972 30104 22024
rect 30156 22012 30162 22024
rect 30285 22015 30343 22021
rect 30285 22012 30297 22015
rect 30156 21984 30297 22012
rect 30156 21972 30162 21984
rect 30285 21981 30297 21984
rect 30331 21981 30343 22015
rect 30285 21975 30343 21981
rect 30374 21972 30380 22024
rect 30432 21972 30438 22024
rect 31404 22021 31432 22052
rect 31389 22015 31447 22021
rect 31389 21981 31401 22015
rect 31435 21981 31447 22015
rect 31389 21975 31447 21981
rect 31570 21972 31576 22024
rect 31628 21972 31634 22024
rect 31680 22021 31708 22052
rect 33689 22049 33701 22083
rect 33735 22080 33747 22083
rect 35866 22080 35894 22120
rect 33735 22052 35894 22080
rect 33735 22049 33747 22052
rect 33689 22043 33747 22049
rect 31665 22015 31723 22021
rect 31665 21981 31677 22015
rect 31711 21981 31723 22015
rect 31665 21975 31723 21981
rect 31849 22015 31907 22021
rect 31849 21981 31861 22015
rect 31895 22012 31907 22015
rect 32674 22012 32680 22024
rect 31895 21984 32680 22012
rect 31895 21981 31907 21984
rect 31849 21975 31907 21981
rect 32674 21972 32680 21984
rect 32732 21972 32738 22024
rect 33870 21972 33876 22024
rect 33928 21972 33934 22024
rect 34330 21972 34336 22024
rect 34388 21972 34394 22024
rect 29144 21916 30052 21944
rect 29144 21904 29150 21916
rect 27448 21848 27752 21876
rect 27341 21839 27399 21845
rect 28074 21836 28080 21888
rect 28132 21836 28138 21888
rect 28445 21879 28503 21885
rect 28445 21845 28457 21879
rect 28491 21876 28503 21879
rect 29546 21876 29552 21888
rect 28491 21848 29552 21876
rect 28491 21845 28503 21848
rect 28445 21839 28503 21845
rect 29546 21836 29552 21848
rect 29604 21876 29610 21888
rect 30392 21876 30420 21972
rect 30650 21904 30656 21956
rect 30708 21944 30714 21956
rect 31757 21947 31815 21953
rect 31757 21944 31769 21947
rect 30708 21916 31769 21944
rect 30708 21904 30714 21916
rect 31757 21913 31769 21916
rect 31803 21913 31815 21947
rect 31757 21907 31815 21913
rect 33318 21904 33324 21956
rect 33376 21904 33382 21956
rect 33962 21904 33968 21956
rect 34020 21904 34026 21956
rect 34057 21947 34115 21953
rect 34057 21913 34069 21947
rect 34103 21913 34115 21947
rect 34057 21907 34115 21913
rect 34195 21947 34253 21953
rect 34195 21913 34207 21947
rect 34241 21944 34253 21947
rect 34241 21916 36400 21944
rect 34241 21913 34253 21916
rect 34195 21907 34253 21913
rect 29604 21848 30420 21876
rect 29604 21836 29610 21848
rect 31294 21836 31300 21888
rect 31352 21876 31358 21888
rect 31481 21879 31539 21885
rect 31481 21876 31493 21879
rect 31352 21848 31493 21876
rect 31352 21836 31358 21848
rect 31481 21845 31493 21848
rect 31527 21876 31539 21879
rect 31938 21876 31944 21888
rect 31527 21848 31944 21876
rect 31527 21845 31539 21848
rect 31481 21839 31539 21845
rect 31938 21836 31944 21848
rect 31996 21836 32002 21888
rect 33336 21876 33364 21904
rect 34072 21876 34100 21907
rect 36372 21888 36400 21916
rect 34514 21876 34520 21888
rect 33336 21848 34520 21876
rect 34514 21836 34520 21848
rect 34572 21836 34578 21888
rect 36354 21836 36360 21888
rect 36412 21836 36418 21888
rect 1104 21786 41400 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 41400 21786
rect 1104 21712 41400 21734
rect 2498 21632 2504 21684
rect 2556 21632 2562 21684
rect 5626 21672 5632 21684
rect 5092 21644 5632 21672
rect 2041 21539 2099 21545
rect 2041 21505 2053 21539
rect 2087 21536 2099 21539
rect 2516 21536 2544 21632
rect 3234 21604 3240 21616
rect 2608 21576 3240 21604
rect 2608 21545 2636 21576
rect 3234 21564 3240 21576
rect 3292 21564 3298 21616
rect 5092 21604 5120 21644
rect 5626 21632 5632 21644
rect 5684 21632 5690 21684
rect 7193 21675 7251 21681
rect 7193 21641 7205 21675
rect 7239 21672 7251 21675
rect 7650 21672 7656 21684
rect 7239 21644 7656 21672
rect 7239 21641 7251 21644
rect 7193 21635 7251 21641
rect 7650 21632 7656 21644
rect 7708 21672 7714 21684
rect 8202 21672 8208 21684
rect 7708 21644 8208 21672
rect 7708 21632 7714 21644
rect 8202 21632 8208 21644
rect 8260 21632 8266 21684
rect 9214 21672 9220 21684
rect 8312 21644 9220 21672
rect 4186 21576 5120 21604
rect 5166 21564 5172 21616
rect 5224 21604 5230 21616
rect 5442 21604 5448 21616
rect 5224 21576 5448 21604
rect 5224 21564 5230 21576
rect 5442 21564 5448 21576
rect 5500 21604 5506 21616
rect 5500 21576 6868 21604
rect 5500 21564 5506 21576
rect 2087 21508 2544 21536
rect 2593 21539 2651 21545
rect 2087 21505 2099 21508
rect 2041 21499 2099 21505
rect 2593 21505 2605 21539
rect 2639 21505 2651 21539
rect 2593 21499 2651 21505
rect 6549 21539 6607 21545
rect 6549 21505 6561 21539
rect 6595 21536 6607 21539
rect 6595 21508 6776 21536
rect 6595 21505 6607 21508
rect 6549 21499 6607 21505
rect 2682 21428 2688 21480
rect 2740 21428 2746 21480
rect 2961 21471 3019 21477
rect 2961 21468 2973 21471
rect 2792 21440 2973 21468
rect 2409 21403 2467 21409
rect 2409 21369 2421 21403
rect 2455 21400 2467 21403
rect 2792 21400 2820 21440
rect 2961 21437 2973 21440
rect 3007 21437 3019 21471
rect 2961 21431 3019 21437
rect 2455 21372 2820 21400
rect 2455 21369 2467 21372
rect 2409 21363 2467 21369
rect 4062 21360 4068 21412
rect 4120 21400 4126 21412
rect 6748 21409 6776 21508
rect 6840 21468 6868 21576
rect 7101 21539 7159 21545
rect 7101 21505 7113 21539
rect 7147 21536 7159 21539
rect 7558 21536 7564 21548
rect 7147 21508 7564 21536
rect 7147 21505 7159 21508
rect 7101 21499 7159 21505
rect 7558 21496 7564 21508
rect 7616 21496 7622 21548
rect 7377 21471 7435 21477
rect 7377 21468 7389 21471
rect 6840 21440 7389 21468
rect 7377 21437 7389 21440
rect 7423 21468 7435 21471
rect 8312 21468 8340 21644
rect 9214 21632 9220 21644
rect 9272 21632 9278 21684
rect 9306 21632 9312 21684
rect 9364 21632 9370 21684
rect 9493 21675 9551 21681
rect 9493 21641 9505 21675
rect 9539 21672 9551 21675
rect 9766 21672 9772 21684
rect 9539 21644 9772 21672
rect 9539 21641 9551 21644
rect 9493 21635 9551 21641
rect 9766 21632 9772 21644
rect 9824 21632 9830 21684
rect 10781 21675 10839 21681
rect 10781 21641 10793 21675
rect 10827 21672 10839 21675
rect 11422 21672 11428 21684
rect 10827 21644 11428 21672
rect 10827 21641 10839 21644
rect 10781 21635 10839 21641
rect 11422 21632 11428 21644
rect 11480 21632 11486 21684
rect 11514 21632 11520 21684
rect 11572 21672 11578 21684
rect 15381 21675 15439 21681
rect 11572 21644 15148 21672
rect 11572 21632 11578 21644
rect 8478 21564 8484 21616
rect 8536 21604 8542 21616
rect 9125 21607 9183 21613
rect 8536 21576 8985 21604
rect 8536 21564 8542 21576
rect 8846 21496 8852 21548
rect 8904 21496 8910 21548
rect 8957 21545 8985 21576
rect 9125 21573 9137 21607
rect 9171 21604 9183 21607
rect 9324 21604 9352 21632
rect 10870 21604 10876 21616
rect 9171 21576 9352 21604
rect 10336 21576 10876 21604
rect 9171 21573 9183 21576
rect 9125 21567 9183 21573
rect 8942 21539 9000 21545
rect 8942 21505 8954 21539
rect 8988 21505 9000 21539
rect 9217 21539 9275 21545
rect 9217 21536 9229 21539
rect 8942 21499 9000 21505
rect 9048 21508 9229 21536
rect 7423 21440 8340 21468
rect 7423 21437 7435 21440
rect 7377 21431 7435 21437
rect 4433 21403 4491 21409
rect 4433 21400 4445 21403
rect 4120 21372 4445 21400
rect 4120 21360 4126 21372
rect 4433 21369 4445 21372
rect 4479 21400 4491 21403
rect 6733 21403 6791 21409
rect 4479 21372 6500 21400
rect 4479 21369 4491 21372
rect 4433 21363 4491 21369
rect 1854 21292 1860 21344
rect 1912 21292 1918 21344
rect 2682 21292 2688 21344
rect 2740 21332 2746 21344
rect 4154 21332 4160 21344
rect 2740 21304 4160 21332
rect 2740 21292 2746 21304
rect 4154 21292 4160 21304
rect 4212 21332 4218 21344
rect 5902 21332 5908 21344
rect 4212 21304 5908 21332
rect 4212 21292 4218 21304
rect 5902 21292 5908 21304
rect 5960 21292 5966 21344
rect 6270 21292 6276 21344
rect 6328 21332 6334 21344
rect 6365 21335 6423 21341
rect 6365 21332 6377 21335
rect 6328 21304 6377 21332
rect 6328 21292 6334 21304
rect 6365 21301 6377 21304
rect 6411 21301 6423 21335
rect 6472 21332 6500 21372
rect 6733 21369 6745 21403
rect 6779 21369 6791 21403
rect 6733 21363 6791 21369
rect 6914 21360 6920 21412
rect 6972 21400 6978 21412
rect 9048 21400 9076 21508
rect 9217 21505 9229 21508
rect 9263 21505 9275 21539
rect 9217 21499 9275 21505
rect 9355 21539 9413 21545
rect 9355 21505 9367 21539
rect 9401 21536 9413 21539
rect 9582 21536 9588 21548
rect 9401 21508 9588 21536
rect 9401 21505 9413 21508
rect 9355 21499 9413 21505
rect 9582 21496 9588 21508
rect 9640 21496 9646 21548
rect 9674 21496 9680 21548
rect 9732 21536 9738 21548
rect 10336 21545 10364 21576
rect 10870 21564 10876 21576
rect 10928 21564 10934 21616
rect 13906 21604 13912 21616
rect 13464 21576 13912 21604
rect 10137 21539 10195 21545
rect 10137 21536 10149 21539
rect 9732 21508 10149 21536
rect 9732 21496 9738 21508
rect 10137 21505 10149 21508
rect 10183 21505 10195 21539
rect 10137 21499 10195 21505
rect 10285 21539 10364 21545
rect 10285 21505 10297 21539
rect 10331 21508 10364 21539
rect 10331 21505 10343 21508
rect 10285 21499 10343 21505
rect 10410 21496 10416 21548
rect 10468 21496 10474 21548
rect 10502 21496 10508 21548
rect 10560 21496 10566 21548
rect 10686 21545 10692 21548
rect 10643 21539 10692 21545
rect 10643 21505 10655 21539
rect 10689 21505 10692 21539
rect 10643 21499 10692 21505
rect 10686 21496 10692 21499
rect 10744 21496 10750 21548
rect 13464 21545 13492 21576
rect 13906 21564 13912 21576
rect 13964 21564 13970 21616
rect 15013 21607 15071 21613
rect 15013 21573 15025 21607
rect 15059 21573 15071 21607
rect 15013 21567 15071 21573
rect 13449 21539 13507 21545
rect 13449 21505 13461 21539
rect 13495 21505 13507 21539
rect 13449 21499 13507 21505
rect 13998 21496 14004 21548
rect 14056 21536 14062 21548
rect 14274 21536 14280 21548
rect 14056 21508 14280 21536
rect 14056 21496 14062 21508
rect 14274 21496 14280 21508
rect 14332 21496 14338 21548
rect 11606 21428 11612 21480
rect 11664 21468 11670 21480
rect 12066 21468 12072 21480
rect 11664 21440 12072 21468
rect 11664 21428 11670 21440
rect 12066 21428 12072 21440
rect 12124 21428 12130 21480
rect 15028 21468 15056 21567
rect 15120 21536 15148 21644
rect 15381 21641 15393 21675
rect 15427 21672 15439 21675
rect 15746 21672 15752 21684
rect 15427 21644 15752 21672
rect 15427 21641 15439 21644
rect 15381 21635 15439 21641
rect 15746 21632 15752 21644
rect 15804 21632 15810 21684
rect 16390 21632 16396 21684
rect 16448 21672 16454 21684
rect 17405 21675 17463 21681
rect 17405 21672 17417 21675
rect 16448 21644 17417 21672
rect 16448 21632 16454 21644
rect 17405 21641 17417 21644
rect 17451 21641 17463 21675
rect 17405 21635 17463 21641
rect 17770 21632 17776 21684
rect 17828 21672 17834 21684
rect 18877 21675 18935 21681
rect 18877 21672 18889 21675
rect 17828 21644 18889 21672
rect 17828 21632 17834 21644
rect 18877 21641 18889 21644
rect 18923 21641 18935 21675
rect 18877 21635 18935 21641
rect 19058 21632 19064 21684
rect 19116 21672 19122 21684
rect 19518 21672 19524 21684
rect 19116 21644 19524 21672
rect 19116 21632 19122 21644
rect 19518 21632 19524 21644
rect 19576 21632 19582 21684
rect 20990 21632 20996 21684
rect 21048 21672 21054 21684
rect 21174 21672 21180 21684
rect 21048 21644 21180 21672
rect 21048 21632 21054 21644
rect 15229 21607 15287 21613
rect 15229 21573 15241 21607
rect 15275 21604 15287 21607
rect 15654 21604 15660 21616
rect 15275 21576 15660 21604
rect 15275 21573 15287 21576
rect 15229 21567 15287 21573
rect 15654 21564 15660 21576
rect 15712 21604 15718 21616
rect 15841 21607 15899 21613
rect 15841 21604 15853 21607
rect 15712 21576 15853 21604
rect 15712 21564 15718 21576
rect 15841 21573 15853 21576
rect 15887 21573 15899 21607
rect 15841 21567 15899 21573
rect 18417 21607 18475 21613
rect 18417 21573 18429 21607
rect 18463 21604 18475 21607
rect 19334 21604 19340 21616
rect 18463 21576 19340 21604
rect 18463 21573 18475 21576
rect 18417 21567 18475 21573
rect 17313 21539 17371 21545
rect 17313 21536 17325 21539
rect 15120 21508 17325 21536
rect 17313 21505 17325 21508
rect 17359 21505 17371 21539
rect 17313 21499 17371 21505
rect 17681 21539 17739 21545
rect 17681 21505 17693 21539
rect 17727 21536 17739 21539
rect 17954 21536 17960 21548
rect 17727 21508 17960 21536
rect 17727 21505 17739 21508
rect 17681 21499 17739 21505
rect 17954 21496 17960 21508
rect 18012 21496 18018 21548
rect 15378 21468 15384 21480
rect 15028 21440 15384 21468
rect 15378 21428 15384 21440
rect 15436 21428 15442 21480
rect 15470 21428 15476 21480
rect 15528 21428 15534 21480
rect 15746 21428 15752 21480
rect 15804 21428 15810 21480
rect 15958 21471 16016 21477
rect 15958 21468 15970 21471
rect 15948 21437 15970 21468
rect 16004 21437 16016 21471
rect 15948 21431 16016 21437
rect 17865 21471 17923 21477
rect 17865 21437 17877 21471
rect 17911 21468 17923 21471
rect 18432 21468 18460 21567
rect 19334 21564 19340 21576
rect 19392 21564 19398 21616
rect 20162 21564 20168 21616
rect 20220 21604 20226 21616
rect 20533 21607 20591 21613
rect 20220 21576 20484 21604
rect 20220 21564 20226 21576
rect 18966 21496 18972 21548
rect 19024 21496 19030 21548
rect 19153 21539 19211 21545
rect 19153 21505 19165 21539
rect 19199 21536 19211 21539
rect 19426 21536 19432 21548
rect 19199 21508 19432 21536
rect 19199 21505 19211 21508
rect 19153 21499 19211 21505
rect 19426 21496 19432 21508
rect 19484 21496 19490 21548
rect 20257 21539 20315 21545
rect 20257 21505 20269 21539
rect 20303 21505 20315 21539
rect 20257 21499 20315 21505
rect 20349 21539 20407 21545
rect 20349 21505 20361 21539
rect 20395 21505 20407 21539
rect 20456 21536 20484 21576
rect 20533 21573 20545 21607
rect 20579 21604 20591 21607
rect 20714 21604 20720 21616
rect 20579 21576 20720 21604
rect 20579 21573 20591 21576
rect 20533 21567 20591 21573
rect 20714 21564 20720 21576
rect 20772 21564 20778 21616
rect 21100 21545 21128 21644
rect 21174 21632 21180 21644
rect 21232 21632 21238 21684
rect 22465 21675 22523 21681
rect 22465 21672 22477 21675
rect 21284 21644 22477 21672
rect 21284 21604 21312 21644
rect 22465 21641 22477 21644
rect 22511 21641 22523 21675
rect 22465 21635 22523 21641
rect 22922 21632 22928 21684
rect 22980 21632 22986 21684
rect 23842 21632 23848 21684
rect 23900 21632 23906 21684
rect 24394 21632 24400 21684
rect 24452 21632 24458 21684
rect 27154 21632 27160 21684
rect 27212 21672 27218 21684
rect 27430 21672 27436 21684
rect 27212 21644 27436 21672
rect 27212 21632 27218 21644
rect 27430 21632 27436 21644
rect 27488 21632 27494 21684
rect 28353 21675 28411 21681
rect 28353 21641 28365 21675
rect 28399 21672 28411 21675
rect 28626 21672 28632 21684
rect 28399 21644 28632 21672
rect 28399 21641 28411 21644
rect 28353 21635 28411 21641
rect 28626 21632 28632 21644
rect 28684 21632 28690 21684
rect 29178 21632 29184 21684
rect 29236 21632 29242 21684
rect 29730 21632 29736 21684
rect 29788 21672 29794 21684
rect 30834 21672 30840 21684
rect 29788 21644 30840 21672
rect 29788 21632 29794 21644
rect 30834 21632 30840 21644
rect 30892 21632 30898 21684
rect 33965 21675 34023 21681
rect 33965 21641 33977 21675
rect 34011 21672 34023 21675
rect 34054 21672 34060 21684
rect 34011 21644 34060 21672
rect 34011 21641 34023 21644
rect 33965 21635 34023 21641
rect 34054 21632 34060 21644
rect 34112 21632 34118 21684
rect 34716 21644 35480 21672
rect 22097 21607 22155 21613
rect 21192 21576 21312 21604
rect 21744 21576 22048 21604
rect 21192 21545 21220 21576
rect 20901 21539 20959 21545
rect 20456 21508 20852 21536
rect 20349 21499 20407 21505
rect 17911 21440 18460 21468
rect 17911 21437 17923 21440
rect 17865 21431 17923 21437
rect 11974 21400 11980 21412
rect 6972 21372 9076 21400
rect 9646 21372 11980 21400
rect 6972 21360 6978 21372
rect 6932 21332 6960 21360
rect 6472 21304 6960 21332
rect 6365 21295 6423 21301
rect 8846 21292 8852 21344
rect 8904 21332 8910 21344
rect 9646 21332 9674 21372
rect 11974 21360 11980 21372
rect 12032 21360 12038 21412
rect 12986 21360 12992 21412
rect 13044 21400 13050 21412
rect 13630 21400 13636 21412
rect 13044 21372 13636 21400
rect 13044 21360 13050 21372
rect 13630 21360 13636 21372
rect 13688 21360 13694 21412
rect 15396 21400 15424 21428
rect 15948 21400 15976 21431
rect 18506 21428 18512 21480
rect 18564 21468 18570 21480
rect 18564 21440 20208 21468
rect 18564 21428 18570 21440
rect 15396 21372 15976 21400
rect 18785 21403 18843 21409
rect 18785 21369 18797 21403
rect 18831 21400 18843 21403
rect 19058 21400 19064 21412
rect 18831 21372 19064 21400
rect 18831 21369 18843 21372
rect 18785 21363 18843 21369
rect 19058 21360 19064 21372
rect 19116 21360 19122 21412
rect 19168 21372 20116 21400
rect 8904 21304 9674 21332
rect 8904 21292 8910 21304
rect 13814 21292 13820 21344
rect 13872 21332 13878 21344
rect 14458 21332 14464 21344
rect 13872 21304 14464 21332
rect 13872 21292 13878 21304
rect 14458 21292 14464 21304
rect 14516 21292 14522 21344
rect 15197 21335 15255 21341
rect 15197 21301 15209 21335
rect 15243 21332 15255 21335
rect 15746 21332 15752 21344
rect 15243 21304 15752 21332
rect 15243 21301 15255 21304
rect 15197 21295 15255 21301
rect 15746 21292 15752 21304
rect 15804 21292 15810 21344
rect 16114 21292 16120 21344
rect 16172 21292 16178 21344
rect 19168 21341 19196 21372
rect 20088 21344 20116 21372
rect 19153 21335 19211 21341
rect 19153 21301 19165 21335
rect 19199 21301 19211 21335
rect 19153 21295 19211 21301
rect 19242 21292 19248 21344
rect 19300 21332 19306 21344
rect 19337 21335 19395 21341
rect 19337 21332 19349 21335
rect 19300 21304 19349 21332
rect 19300 21292 19306 21304
rect 19337 21301 19349 21304
rect 19383 21301 19395 21335
rect 19337 21295 19395 21301
rect 20070 21292 20076 21344
rect 20128 21292 20134 21344
rect 20180 21332 20208 21440
rect 20272 21400 20300 21499
rect 20364 21468 20392 21499
rect 20714 21468 20720 21480
rect 20364 21440 20720 21468
rect 20714 21428 20720 21440
rect 20772 21428 20778 21480
rect 20824 21468 20852 21508
rect 20901 21505 20913 21539
rect 20947 21536 20959 21539
rect 21066 21539 21128 21545
rect 20947 21508 21036 21536
rect 20947 21505 20959 21508
rect 20901 21499 20959 21505
rect 21008 21468 21036 21508
rect 21066 21505 21078 21539
rect 21112 21508 21128 21539
rect 21177 21539 21235 21545
rect 21112 21505 21124 21508
rect 21066 21499 21124 21505
rect 21177 21505 21189 21539
rect 21223 21505 21235 21539
rect 21177 21499 21235 21505
rect 21266 21496 21272 21548
rect 21324 21496 21330 21548
rect 21744 21468 21772 21576
rect 21818 21496 21824 21548
rect 21876 21496 21882 21548
rect 21914 21539 21972 21545
rect 21914 21505 21926 21539
rect 21960 21505 21972 21539
rect 21914 21499 21972 21505
rect 20824 21440 20908 21468
rect 21008 21440 21772 21468
rect 20438 21400 20444 21412
rect 20272 21372 20444 21400
rect 20438 21360 20444 21372
rect 20496 21400 20502 21412
rect 20880 21400 20908 21440
rect 21929 21400 21957 21499
rect 22020 21468 22048 21576
rect 22097 21573 22109 21607
rect 22143 21604 22155 21607
rect 22940 21604 22968 21632
rect 23566 21604 23572 21616
rect 22143 21576 23572 21604
rect 22143 21573 22155 21576
rect 22097 21567 22155 21573
rect 23566 21564 23572 21576
rect 23624 21564 23630 21616
rect 23860 21604 23888 21632
rect 23860 21576 23980 21604
rect 22186 21496 22192 21548
rect 22244 21496 22250 21548
rect 22327 21539 22385 21545
rect 22327 21505 22339 21539
rect 22373 21536 22385 21539
rect 22738 21536 22744 21548
rect 22373 21508 22744 21536
rect 22373 21505 22385 21508
rect 22327 21499 22385 21505
rect 22738 21496 22744 21508
rect 22796 21536 22802 21548
rect 23842 21536 23848 21548
rect 22796 21508 23848 21536
rect 22796 21496 22802 21508
rect 23842 21496 23848 21508
rect 23900 21496 23906 21548
rect 23952 21468 23980 21576
rect 24029 21539 24087 21545
rect 24029 21505 24041 21539
rect 24075 21536 24087 21539
rect 24412 21536 24440 21632
rect 25869 21607 25927 21613
rect 25869 21604 25881 21607
rect 25424 21576 25881 21604
rect 25424 21548 25452 21576
rect 25869 21573 25881 21576
rect 25915 21573 25927 21607
rect 25869 21567 25927 21573
rect 25958 21564 25964 21616
rect 26016 21564 26022 21616
rect 27062 21604 27068 21616
rect 26068 21576 27068 21604
rect 24075 21508 24440 21536
rect 24075 21505 24087 21508
rect 24029 21499 24087 21505
rect 25406 21496 25412 21548
rect 25464 21496 25470 21548
rect 25685 21539 25743 21545
rect 25685 21536 25697 21539
rect 25608 21508 25697 21536
rect 24121 21471 24179 21477
rect 24121 21468 24133 21471
rect 22020 21440 23904 21468
rect 23952 21440 24133 21468
rect 20496 21372 20852 21400
rect 20880 21372 21957 21400
rect 20496 21360 20502 21372
rect 20717 21335 20775 21341
rect 20717 21332 20729 21335
rect 20180 21304 20729 21332
rect 20717 21301 20729 21304
rect 20763 21301 20775 21335
rect 20824 21332 20852 21372
rect 21634 21332 21640 21344
rect 20824 21304 21640 21332
rect 20717 21295 20775 21301
rect 21634 21292 21640 21304
rect 21692 21292 21698 21344
rect 21929 21332 21957 21372
rect 22738 21360 22744 21412
rect 22796 21400 22802 21412
rect 23014 21400 23020 21412
rect 22796 21372 23020 21400
rect 22796 21360 22802 21372
rect 23014 21360 23020 21372
rect 23072 21360 23078 21412
rect 23876 21400 23904 21440
rect 24121 21437 24133 21440
rect 24167 21468 24179 21471
rect 24394 21468 24400 21480
rect 24167 21440 24400 21468
rect 24167 21437 24179 21440
rect 24121 21431 24179 21437
rect 24394 21428 24400 21440
rect 24452 21428 24458 21480
rect 25498 21468 25504 21480
rect 24780 21440 25504 21468
rect 24780 21400 24808 21440
rect 25498 21428 25504 21440
rect 25556 21428 25562 21480
rect 23876 21372 24808 21400
rect 24854 21360 24860 21412
rect 24912 21400 24918 21412
rect 25608 21400 25636 21508
rect 25685 21505 25697 21508
rect 25731 21505 25743 21539
rect 25976 21535 26004 21564
rect 26068 21545 26096 21576
rect 27062 21564 27068 21576
rect 27120 21564 27126 21616
rect 27798 21604 27804 21616
rect 27356 21576 27804 21604
rect 26053 21539 26111 21545
rect 25685 21499 25743 21505
rect 25957 21529 26015 21535
rect 25957 21495 25969 21529
rect 26003 21495 26015 21529
rect 26053 21505 26065 21539
rect 26099 21505 26111 21539
rect 26053 21499 26111 21505
rect 25957 21489 26015 21495
rect 24912 21372 25636 21400
rect 25685 21403 25743 21409
rect 24912 21360 24918 21372
rect 25685 21369 25697 21403
rect 25731 21400 25743 21403
rect 26068 21400 26096 21499
rect 26326 21428 26332 21480
rect 26384 21468 26390 21480
rect 26694 21468 26700 21480
rect 26384 21440 26700 21468
rect 26384 21428 26390 21440
rect 26694 21428 26700 21440
rect 26752 21428 26758 21480
rect 25731 21372 26096 21400
rect 25731 21369 25743 21372
rect 25685 21363 25743 21369
rect 23934 21332 23940 21344
rect 21929 21304 23940 21332
rect 23934 21292 23940 21304
rect 23992 21292 23998 21344
rect 24210 21292 24216 21344
rect 24268 21292 24274 21344
rect 24394 21292 24400 21344
rect 24452 21292 24458 21344
rect 25038 21292 25044 21344
rect 25096 21332 25102 21344
rect 25774 21332 25780 21344
rect 25096 21304 25780 21332
rect 25096 21292 25102 21304
rect 25774 21292 25780 21304
rect 25832 21332 25838 21344
rect 26145 21335 26203 21341
rect 26145 21332 26157 21335
rect 25832 21304 26157 21332
rect 25832 21292 25838 21304
rect 26145 21301 26157 21304
rect 26191 21301 26203 21335
rect 26145 21295 26203 21301
rect 27062 21292 27068 21344
rect 27120 21332 27126 21344
rect 27356 21332 27384 21576
rect 27798 21564 27804 21576
rect 27856 21564 27862 21616
rect 27893 21607 27951 21613
rect 27893 21573 27905 21607
rect 27939 21604 27951 21607
rect 27982 21604 27988 21616
rect 27939 21576 27988 21604
rect 27939 21573 27951 21576
rect 27893 21567 27951 21573
rect 27982 21564 27988 21576
rect 28040 21564 28046 21616
rect 29196 21604 29224 21632
rect 28736 21576 29224 21604
rect 34072 21604 34100 21632
rect 34716 21616 34744 21644
rect 34330 21604 34336 21616
rect 34072 21576 34336 21604
rect 27433 21539 27491 21545
rect 27433 21505 27445 21539
rect 27479 21536 27491 21539
rect 27706 21536 27712 21548
rect 27479 21508 27712 21536
rect 27479 21505 27491 21508
rect 27433 21499 27491 21505
rect 27706 21496 27712 21508
rect 27764 21496 27770 21548
rect 28074 21496 28080 21548
rect 28132 21496 28138 21548
rect 28169 21539 28227 21545
rect 28169 21505 28181 21539
rect 28215 21536 28227 21539
rect 28445 21539 28503 21545
rect 28445 21536 28457 21539
rect 28215 21508 28457 21536
rect 28215 21505 28227 21508
rect 28169 21499 28227 21505
rect 28445 21505 28457 21508
rect 28491 21505 28503 21539
rect 28445 21499 28503 21505
rect 28534 21496 28540 21548
rect 28592 21536 28598 21548
rect 28736 21545 28764 21576
rect 34330 21564 34336 21576
rect 34388 21564 34394 21616
rect 34698 21564 34704 21616
rect 34756 21564 34762 21616
rect 35342 21564 35348 21616
rect 35400 21564 35406 21616
rect 35452 21604 35480 21644
rect 36354 21632 36360 21684
rect 36412 21672 36418 21684
rect 38010 21672 38016 21684
rect 36412 21644 38016 21672
rect 36412 21632 36418 21644
rect 38010 21632 38016 21644
rect 38068 21672 38074 21684
rect 39022 21672 39028 21684
rect 38068 21644 39028 21672
rect 38068 21632 38074 21644
rect 39022 21632 39028 21644
rect 39080 21672 39086 21684
rect 39942 21672 39948 21684
rect 39080 21644 39948 21672
rect 39080 21632 39086 21644
rect 39942 21632 39948 21644
rect 40000 21632 40006 21684
rect 40862 21632 40868 21684
rect 40920 21632 40926 21684
rect 35555 21607 35613 21613
rect 35555 21604 35567 21607
rect 35452 21576 35567 21604
rect 35555 21573 35567 21576
rect 35601 21573 35613 21607
rect 36630 21604 36636 21616
rect 35555 21567 35613 21573
rect 35728 21576 36636 21604
rect 28721 21539 28779 21545
rect 28721 21536 28733 21539
rect 28592 21508 28733 21536
rect 28592 21496 28598 21508
rect 28721 21505 28733 21508
rect 28767 21505 28779 21539
rect 28721 21499 28779 21505
rect 29181 21539 29239 21545
rect 29181 21505 29193 21539
rect 29227 21536 29239 21539
rect 30098 21536 30104 21548
rect 29227 21508 30104 21536
rect 29227 21505 29239 21508
rect 29181 21499 29239 21505
rect 30098 21496 30104 21508
rect 30156 21536 30162 21548
rect 31386 21536 31392 21548
rect 30156 21508 31392 21536
rect 30156 21496 30162 21508
rect 31386 21496 31392 21508
rect 31444 21496 31450 21548
rect 33134 21496 33140 21548
rect 33192 21536 33198 21548
rect 35728 21545 35756 21576
rect 36630 21564 36636 21576
rect 36688 21564 36694 21616
rect 37274 21564 37280 21616
rect 37332 21604 37338 21616
rect 37332 21576 39068 21604
rect 37332 21564 37338 21576
rect 33689 21539 33747 21545
rect 33689 21536 33701 21539
rect 33192 21508 33701 21536
rect 33192 21496 33198 21508
rect 33689 21505 33701 21508
rect 33735 21536 33747 21539
rect 35253 21539 35311 21545
rect 35253 21536 35265 21539
rect 33735 21508 35265 21536
rect 33735 21505 33747 21508
rect 33689 21499 33747 21505
rect 27724 21468 27752 21496
rect 28258 21468 28264 21480
rect 27724 21440 28264 21468
rect 28258 21428 28264 21440
rect 28316 21428 28322 21480
rect 31754 21428 31760 21480
rect 31812 21428 31818 21480
rect 28442 21360 28448 21412
rect 28500 21400 28506 21412
rect 28813 21403 28871 21409
rect 28813 21400 28825 21403
rect 28500 21372 28825 21400
rect 28500 21360 28506 21372
rect 28813 21369 28825 21372
rect 28859 21369 28871 21403
rect 28813 21363 28871 21369
rect 29454 21360 29460 21412
rect 29512 21400 29518 21412
rect 31110 21400 31116 21412
rect 29512 21372 31116 21400
rect 29512 21360 29518 21372
rect 31110 21360 31116 21372
rect 31168 21360 31174 21412
rect 31294 21360 31300 21412
rect 31352 21360 31358 21412
rect 31386 21360 31392 21412
rect 31444 21400 31450 21412
rect 31772 21400 31800 21428
rect 31444 21372 31800 21400
rect 31444 21360 31450 21372
rect 27525 21335 27583 21341
rect 27525 21332 27537 21335
rect 27120 21304 27537 21332
rect 27120 21292 27126 21304
rect 27525 21301 27537 21304
rect 27571 21301 27583 21335
rect 27525 21295 27583 21301
rect 27798 21292 27804 21344
rect 27856 21332 27862 21344
rect 27893 21335 27951 21341
rect 27893 21332 27905 21335
rect 27856 21304 27905 21332
rect 27856 21292 27862 21304
rect 27893 21301 27905 21304
rect 27939 21301 27951 21335
rect 27893 21295 27951 21301
rect 28902 21292 28908 21344
rect 28960 21292 28966 21344
rect 28997 21335 29055 21341
rect 28997 21301 29009 21335
rect 29043 21332 29055 21335
rect 31312 21332 31340 21360
rect 29043 21304 31340 21332
rect 34992 21332 35020 21508
rect 35253 21505 35265 21508
rect 35299 21505 35311 21539
rect 35437 21539 35495 21545
rect 35437 21536 35449 21539
rect 35253 21499 35311 21505
rect 35360 21508 35449 21536
rect 35360 21480 35388 21508
rect 35437 21505 35449 21508
rect 35483 21505 35495 21539
rect 35437 21499 35495 21505
rect 35713 21539 35771 21545
rect 35713 21505 35725 21539
rect 35759 21505 35771 21539
rect 37458 21536 37464 21548
rect 35713 21499 35771 21505
rect 36648 21508 37464 21536
rect 35342 21428 35348 21480
rect 35400 21468 35406 21480
rect 35618 21468 35624 21480
rect 35400 21440 35624 21468
rect 35400 21428 35406 21440
rect 35618 21428 35624 21440
rect 35676 21428 35682 21480
rect 35069 21403 35127 21409
rect 35069 21369 35081 21403
rect 35115 21400 35127 21403
rect 36648 21400 36676 21508
rect 37458 21496 37464 21508
rect 37516 21536 37522 21548
rect 37553 21539 37611 21545
rect 37553 21536 37565 21539
rect 37516 21508 37565 21536
rect 37516 21496 37522 21508
rect 37553 21505 37565 21508
rect 37599 21505 37611 21539
rect 37553 21499 37611 21505
rect 38838 21496 38844 21548
rect 38896 21536 38902 21548
rect 39040 21545 39068 21576
rect 38933 21539 38991 21545
rect 38933 21536 38945 21539
rect 38896 21508 38945 21536
rect 38896 21496 38902 21508
rect 38933 21505 38945 21508
rect 38979 21505 38991 21539
rect 38933 21499 38991 21505
rect 39025 21539 39083 21545
rect 39025 21505 39037 21539
rect 39071 21505 39083 21539
rect 39025 21499 39083 21505
rect 41049 21539 41107 21545
rect 41049 21505 41061 21539
rect 41095 21536 41107 21539
rect 41414 21536 41420 21548
rect 41095 21508 41420 21536
rect 41095 21505 41107 21508
rect 41049 21499 41107 21505
rect 41414 21496 41420 21508
rect 41472 21496 41478 21548
rect 37366 21428 37372 21480
rect 37424 21468 37430 21480
rect 38654 21468 38660 21480
rect 37424 21440 38660 21468
rect 37424 21428 37430 21440
rect 38654 21428 38660 21440
rect 38712 21428 38718 21480
rect 35115 21372 36676 21400
rect 35115 21369 35127 21372
rect 35069 21363 35127 21369
rect 38470 21360 38476 21412
rect 38528 21400 38534 21412
rect 38528 21372 39252 21400
rect 38528 21360 38534 21372
rect 39224 21344 39252 21372
rect 35434 21332 35440 21344
rect 34992 21304 35440 21332
rect 29043 21301 29055 21304
rect 28997 21295 29055 21301
rect 35434 21292 35440 21304
rect 35492 21292 35498 21344
rect 35526 21292 35532 21344
rect 35584 21332 35590 21344
rect 37277 21335 37335 21341
rect 37277 21332 37289 21335
rect 35584 21304 37289 21332
rect 35584 21292 35590 21304
rect 37277 21301 37289 21304
rect 37323 21301 37335 21335
rect 37277 21295 37335 21301
rect 37642 21292 37648 21344
rect 37700 21332 37706 21344
rect 37737 21335 37795 21341
rect 37737 21332 37749 21335
rect 37700 21304 37749 21332
rect 37700 21292 37706 21304
rect 37737 21301 37749 21304
rect 37783 21301 37795 21335
rect 37737 21295 37795 21301
rect 37826 21292 37832 21344
rect 37884 21332 37890 21344
rect 38562 21332 38568 21344
rect 37884 21304 38568 21332
rect 37884 21292 37890 21304
rect 38562 21292 38568 21304
rect 38620 21332 38626 21344
rect 38933 21335 38991 21341
rect 38933 21332 38945 21335
rect 38620 21304 38945 21332
rect 38620 21292 38626 21304
rect 38933 21301 38945 21304
rect 38979 21301 38991 21335
rect 38933 21295 38991 21301
rect 39206 21292 39212 21344
rect 39264 21292 39270 21344
rect 39298 21292 39304 21344
rect 39356 21292 39362 21344
rect 1104 21242 41400 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 41400 21242
rect 1104 21168 41400 21190
rect 1660 21131 1718 21137
rect 1660 21097 1672 21131
rect 1706 21128 1718 21131
rect 1854 21128 1860 21140
rect 1706 21100 1860 21128
rect 1706 21097 1718 21100
rect 1660 21091 1718 21097
rect 1854 21088 1860 21100
rect 1912 21088 1918 21140
rect 3234 21088 3240 21140
rect 3292 21128 3298 21140
rect 3789 21131 3847 21137
rect 3789 21128 3801 21131
rect 3292 21100 3801 21128
rect 3292 21088 3298 21100
rect 3789 21097 3801 21100
rect 3835 21097 3847 21131
rect 3789 21091 3847 21097
rect 5368 21100 7236 21128
rect 1394 20952 1400 21004
rect 1452 20992 1458 21004
rect 2682 20992 2688 21004
rect 1452 20964 2688 20992
rect 1452 20952 1458 20964
rect 2682 20952 2688 20964
rect 2740 20952 2746 21004
rect 3142 20952 3148 21004
rect 3200 20992 3206 21004
rect 3200 20964 4016 20992
rect 3200 20952 3206 20964
rect 3050 20856 3056 20868
rect 2898 20828 3056 20856
rect 3050 20816 3056 20828
rect 3108 20816 3114 20868
rect 3988 20856 4016 20964
rect 4062 20952 4068 21004
rect 4120 20952 4126 21004
rect 4433 20995 4491 21001
rect 4433 20961 4445 20995
rect 4479 20961 4491 20995
rect 5368 20992 5396 21100
rect 7208 21060 7236 21100
rect 7650 21088 7656 21140
rect 7708 21088 7714 21140
rect 10502 21088 10508 21140
rect 10560 21088 10566 21140
rect 11514 21088 11520 21140
rect 11572 21128 11578 21140
rect 14550 21128 14556 21140
rect 11572 21100 14556 21128
rect 11572 21088 11578 21100
rect 14550 21088 14556 21100
rect 14608 21088 14614 21140
rect 15562 21128 15568 21140
rect 14660 21100 15568 21128
rect 7926 21060 7932 21072
rect 7208 21032 7932 21060
rect 7926 21020 7932 21032
rect 7984 21060 7990 21072
rect 10520 21060 10548 21088
rect 7984 21032 10548 21060
rect 7984 21020 7990 21032
rect 4433 20955 4491 20961
rect 5276 20964 5396 20992
rect 5552 20964 5856 20992
rect 4080 20924 4108 20952
rect 4249 20927 4307 20933
rect 4249 20924 4261 20927
rect 4080 20896 4261 20924
rect 4249 20893 4261 20896
rect 4295 20893 4307 20927
rect 4448 20924 4476 20955
rect 5166 20924 5172 20936
rect 4448 20896 5172 20924
rect 4249 20887 4307 20893
rect 5166 20884 5172 20896
rect 5224 20884 5230 20936
rect 5276 20933 5304 20964
rect 5261 20927 5319 20933
rect 5261 20893 5273 20927
rect 5307 20893 5319 20927
rect 5261 20887 5319 20893
rect 5350 20884 5356 20936
rect 5408 20924 5414 20936
rect 5552 20933 5580 20964
rect 5828 20936 5856 20964
rect 5902 20952 5908 21004
rect 5960 20952 5966 21004
rect 6181 20995 6239 21001
rect 6181 20961 6193 20995
rect 6227 20992 6239 20995
rect 6270 20992 6276 21004
rect 6227 20964 6276 20992
rect 6227 20961 6239 20964
rect 6181 20955 6239 20961
rect 6270 20952 6276 20964
rect 6328 20952 6334 21004
rect 9398 20952 9404 21004
rect 9456 20992 9462 21004
rect 11885 20995 11943 21001
rect 11885 20992 11897 20995
rect 9456 20964 11897 20992
rect 9456 20952 9462 20964
rect 11885 20961 11897 20964
rect 11931 20992 11943 20995
rect 14660 20992 14688 21100
rect 15562 21088 15568 21100
rect 15620 21088 15626 21140
rect 16850 21128 16856 21140
rect 15672 21100 16856 21128
rect 15013 21063 15071 21069
rect 15013 21029 15025 21063
rect 15059 21060 15071 21063
rect 15470 21060 15476 21072
rect 15059 21032 15476 21060
rect 15059 21029 15071 21032
rect 15013 21023 15071 21029
rect 15470 21020 15476 21032
rect 15528 21060 15534 21072
rect 15672 21060 15700 21100
rect 16850 21088 16856 21100
rect 16908 21128 16914 21140
rect 17678 21128 17684 21140
rect 16908 21100 17684 21128
rect 16908 21088 16914 21100
rect 17678 21088 17684 21100
rect 17736 21088 17742 21140
rect 18966 21088 18972 21140
rect 19024 21088 19030 21140
rect 19429 21131 19487 21137
rect 19429 21097 19441 21131
rect 19475 21128 19487 21131
rect 20070 21128 20076 21140
rect 19475 21100 20076 21128
rect 19475 21097 19487 21100
rect 19429 21091 19487 21097
rect 20070 21088 20076 21100
rect 20128 21088 20134 21140
rect 21453 21131 21511 21137
rect 21453 21097 21465 21131
rect 21499 21128 21511 21131
rect 21726 21128 21732 21140
rect 21499 21100 21732 21128
rect 21499 21097 21511 21100
rect 21453 21091 21511 21097
rect 21726 21088 21732 21100
rect 21784 21088 21790 21140
rect 21910 21088 21916 21140
rect 21968 21128 21974 21140
rect 21968 21100 23336 21128
rect 21968 21088 21974 21100
rect 15528 21032 15700 21060
rect 15528 21020 15534 21032
rect 15746 21020 15752 21072
rect 15804 21060 15810 21072
rect 15933 21063 15991 21069
rect 15933 21060 15945 21063
rect 15804 21032 15945 21060
rect 15804 21020 15810 21032
rect 15933 21029 15945 21032
rect 15979 21029 15991 21063
rect 15933 21023 15991 21029
rect 16022 21020 16028 21072
rect 16080 21060 16086 21072
rect 16206 21060 16212 21072
rect 16080 21032 16212 21060
rect 16080 21020 16086 21032
rect 16206 21020 16212 21032
rect 16264 21060 16270 21072
rect 17221 21063 17279 21069
rect 17221 21060 17233 21063
rect 16264 21032 17233 21060
rect 16264 21020 16270 21032
rect 17221 21029 17233 21032
rect 17267 21029 17279 21063
rect 18984 21060 19012 21088
rect 23198 21060 23204 21072
rect 18984 21032 23204 21060
rect 17221 21023 17279 21029
rect 23198 21020 23204 21032
rect 23256 21020 23262 21072
rect 23308 21060 23336 21100
rect 24210 21088 24216 21140
rect 24268 21128 24274 21140
rect 24394 21128 24400 21140
rect 24268 21100 24400 21128
rect 24268 21088 24274 21100
rect 24394 21088 24400 21100
rect 24452 21088 24458 21140
rect 27338 21128 27344 21140
rect 26988 21100 27344 21128
rect 26988 21060 27016 21100
rect 27338 21088 27344 21100
rect 27396 21088 27402 21140
rect 27522 21088 27528 21140
rect 27580 21128 27586 21140
rect 28166 21128 28172 21140
rect 27580 21100 28172 21128
rect 27580 21088 27586 21100
rect 28166 21088 28172 21100
rect 28224 21088 28230 21140
rect 30926 21088 30932 21140
rect 30984 21128 30990 21140
rect 31754 21128 31760 21140
rect 30984 21100 31760 21128
rect 30984 21088 30990 21100
rect 31754 21088 31760 21100
rect 31812 21088 31818 21140
rect 32490 21088 32496 21140
rect 32548 21128 32554 21140
rect 32858 21128 32864 21140
rect 32548 21100 32864 21128
rect 32548 21088 32554 21100
rect 32858 21088 32864 21100
rect 32916 21088 32922 21140
rect 33045 21131 33103 21137
rect 33045 21097 33057 21131
rect 33091 21128 33103 21131
rect 36078 21128 36084 21140
rect 33091 21100 36084 21128
rect 33091 21097 33103 21100
rect 33045 21091 33103 21097
rect 36078 21088 36084 21100
rect 36136 21088 36142 21140
rect 36262 21088 36268 21140
rect 36320 21128 36326 21140
rect 36722 21128 36728 21140
rect 36320 21100 36728 21128
rect 36320 21088 36326 21100
rect 36722 21088 36728 21100
rect 36780 21088 36786 21140
rect 36906 21088 36912 21140
rect 36964 21128 36970 21140
rect 36964 21100 37596 21128
rect 36964 21088 36970 21100
rect 23308 21032 27016 21060
rect 27065 21063 27123 21069
rect 11931 20964 14688 20992
rect 11931 20961 11943 20964
rect 11885 20955 11943 20961
rect 15378 20952 15384 21004
rect 15436 20992 15442 21004
rect 15565 20995 15623 21001
rect 15565 20992 15577 20995
rect 15436 20964 15577 20992
rect 15436 20952 15442 20964
rect 15565 20961 15577 20964
rect 15611 20992 15623 20995
rect 16393 20995 16451 21001
rect 16393 20992 16405 20995
rect 15611 20964 16405 20992
rect 15611 20961 15623 20964
rect 15565 20955 15623 20961
rect 16393 20961 16405 20964
rect 16439 20992 16451 20995
rect 19150 20992 19156 21004
rect 16439 20964 19156 20992
rect 16439 20961 16451 20964
rect 16393 20955 16451 20961
rect 5445 20927 5503 20933
rect 5445 20924 5457 20927
rect 5408 20896 5457 20924
rect 5408 20884 5414 20896
rect 5445 20893 5457 20896
rect 5491 20893 5503 20927
rect 5445 20887 5503 20893
rect 5537 20927 5595 20933
rect 5537 20893 5549 20927
rect 5583 20893 5595 20927
rect 5537 20887 5595 20893
rect 5629 20927 5687 20933
rect 5629 20893 5641 20927
rect 5675 20893 5687 20927
rect 5629 20887 5687 20893
rect 5552 20856 5580 20887
rect 3988 20828 5580 20856
rect 5644 20856 5672 20887
rect 5810 20884 5816 20936
rect 5868 20884 5874 20936
rect 7282 20884 7288 20936
rect 7340 20884 7346 20936
rect 10870 20884 10876 20936
rect 10928 20924 10934 20936
rect 11330 20924 11336 20936
rect 10928 20896 11336 20924
rect 10928 20884 10934 20896
rect 11330 20884 11336 20896
rect 11388 20884 11394 20936
rect 11609 20927 11667 20933
rect 11609 20893 11621 20927
rect 11655 20924 11667 20927
rect 12434 20924 12440 20936
rect 11655 20896 12440 20924
rect 11655 20893 11667 20896
rect 11609 20887 11667 20893
rect 12434 20884 12440 20896
rect 12492 20884 12498 20936
rect 14461 20927 14519 20933
rect 14461 20893 14473 20927
rect 14507 20924 14519 20927
rect 15749 20927 15807 20933
rect 15749 20924 15761 20927
rect 14507 20896 15761 20924
rect 14507 20893 14519 20896
rect 14461 20887 14519 20893
rect 15749 20893 15761 20896
rect 15795 20893 15807 20927
rect 15749 20887 15807 20893
rect 16485 20927 16543 20933
rect 16485 20893 16497 20927
rect 16531 20924 16543 20927
rect 16761 20927 16819 20933
rect 16761 20924 16773 20927
rect 16531 20896 16773 20924
rect 16531 20893 16543 20896
rect 16485 20887 16543 20893
rect 16761 20893 16773 20896
rect 16807 20924 16819 20927
rect 16850 20924 16856 20936
rect 16807 20896 16856 20924
rect 16807 20893 16819 20896
rect 16761 20887 16819 20893
rect 16850 20884 16856 20896
rect 16908 20884 16914 20936
rect 16960 20933 16988 20964
rect 19150 20952 19156 20964
rect 19208 20952 19214 21004
rect 19337 20995 19395 21001
rect 19337 20961 19349 20995
rect 19383 20992 19395 20995
rect 19426 20992 19432 21004
rect 19383 20964 19432 20992
rect 19383 20961 19395 20964
rect 19337 20955 19395 20961
rect 19426 20952 19432 20964
rect 19484 20952 19490 21004
rect 20254 20952 20260 21004
rect 20312 20952 20318 21004
rect 21361 20995 21419 21001
rect 21361 20961 21373 20995
rect 21407 20992 21419 20995
rect 21818 20992 21824 21004
rect 21407 20964 21824 20992
rect 21407 20961 21419 20964
rect 21361 20955 21419 20961
rect 21818 20952 21824 20964
rect 21876 20992 21882 21004
rect 22094 20992 22100 21004
rect 21876 20964 22100 20992
rect 21876 20952 21882 20964
rect 22094 20952 22100 20964
rect 22152 20952 22158 21004
rect 22278 20952 22284 21004
rect 22336 20992 22342 21004
rect 22741 20995 22799 21001
rect 22741 20992 22753 20995
rect 22336 20964 22753 20992
rect 22336 20952 22342 20964
rect 22741 20961 22753 20964
rect 22787 20961 22799 20995
rect 23308 20992 23336 21032
rect 27065 21029 27077 21063
rect 27111 21060 27123 21063
rect 30561 21063 30619 21069
rect 30561 21060 30573 21063
rect 27111 21032 30573 21060
rect 27111 21029 27123 21032
rect 27065 21023 27123 21029
rect 30561 21029 30573 21032
rect 30607 21029 30619 21063
rect 35437 21063 35495 21069
rect 30561 21023 30619 21029
rect 31220 21032 35204 21060
rect 22741 20955 22799 20961
rect 23216 20964 23336 20992
rect 16945 20927 17003 20933
rect 16945 20893 16957 20927
rect 16991 20893 17003 20927
rect 17313 20927 17371 20933
rect 17313 20924 17325 20927
rect 16945 20887 17003 20893
rect 17052 20896 17325 20924
rect 15013 20859 15071 20865
rect 5644 20828 6040 20856
rect 6012 20800 6040 20828
rect 15013 20825 15025 20859
rect 15059 20825 15071 20859
rect 15013 20819 15071 20825
rect 15473 20859 15531 20865
rect 15473 20825 15485 20859
rect 15519 20856 15531 20859
rect 15654 20856 15660 20868
rect 15519 20828 15660 20856
rect 15519 20825 15531 20828
rect 15473 20819 15531 20825
rect 4157 20791 4215 20797
rect 4157 20757 4169 20791
rect 4203 20788 4215 20791
rect 4706 20788 4712 20800
rect 4203 20760 4712 20788
rect 4203 20757 4215 20760
rect 4157 20751 4215 20757
rect 4706 20748 4712 20760
rect 4764 20788 4770 20800
rect 5074 20788 5080 20800
rect 4764 20760 5080 20788
rect 4764 20748 4770 20760
rect 5074 20748 5080 20760
rect 5132 20748 5138 20800
rect 5626 20748 5632 20800
rect 5684 20788 5690 20800
rect 5813 20791 5871 20797
rect 5813 20788 5825 20791
rect 5684 20760 5825 20788
rect 5684 20748 5690 20760
rect 5813 20757 5825 20760
rect 5859 20757 5871 20791
rect 5813 20751 5871 20757
rect 5994 20748 6000 20800
rect 6052 20748 6058 20800
rect 7742 20748 7748 20800
rect 7800 20788 7806 20800
rect 8386 20788 8392 20800
rect 7800 20760 8392 20788
rect 7800 20748 7806 20760
rect 8386 20748 8392 20760
rect 8444 20748 8450 20800
rect 10962 20748 10968 20800
rect 11020 20788 11026 20800
rect 11241 20791 11299 20797
rect 11241 20788 11253 20791
rect 11020 20760 11253 20788
rect 11020 20748 11026 20760
rect 11241 20757 11253 20760
rect 11287 20757 11299 20791
rect 11241 20751 11299 20757
rect 11701 20791 11759 20797
rect 11701 20757 11713 20791
rect 11747 20788 11759 20791
rect 11882 20788 11888 20800
rect 11747 20760 11888 20788
rect 11747 20757 11759 20760
rect 11701 20751 11759 20757
rect 11882 20748 11888 20760
rect 11940 20788 11946 20800
rect 12158 20788 12164 20800
rect 11940 20760 12164 20788
rect 11940 20748 11946 20760
rect 12158 20748 12164 20760
rect 12216 20748 12222 20800
rect 15028 20788 15056 20819
rect 15654 20816 15660 20828
rect 15712 20856 15718 20868
rect 15933 20859 15991 20865
rect 15933 20856 15945 20859
rect 15712 20828 15945 20856
rect 15712 20816 15718 20828
rect 15933 20825 15945 20828
rect 15979 20856 15991 20859
rect 16206 20856 16212 20868
rect 15979 20828 16212 20856
rect 15979 20825 15991 20828
rect 15933 20819 15991 20825
rect 16206 20816 16212 20828
rect 16264 20816 16270 20868
rect 16666 20816 16672 20868
rect 16724 20816 16730 20868
rect 15746 20788 15752 20800
rect 15028 20760 15752 20788
rect 15746 20748 15752 20760
rect 15804 20788 15810 20800
rect 17052 20788 17080 20896
rect 17313 20893 17325 20896
rect 17359 20893 17371 20927
rect 17313 20887 17371 20893
rect 17328 20856 17356 20887
rect 19242 20884 19248 20936
rect 19300 20884 19306 20936
rect 20272 20856 20300 20952
rect 20622 20884 20628 20936
rect 20680 20924 20686 20936
rect 21177 20927 21235 20933
rect 21177 20924 21189 20927
rect 20680 20896 21189 20924
rect 20680 20884 20686 20896
rect 21177 20893 21189 20896
rect 21223 20893 21235 20927
rect 21177 20887 21235 20893
rect 21453 20927 21511 20933
rect 21453 20893 21465 20927
rect 21499 20924 21511 20927
rect 22002 20924 22008 20936
rect 21499 20896 22008 20924
rect 21499 20893 21511 20896
rect 21453 20887 21511 20893
rect 22002 20884 22008 20896
rect 22060 20884 22066 20936
rect 22465 20927 22523 20933
rect 22465 20893 22477 20927
rect 22511 20893 22523 20927
rect 22465 20887 22523 20893
rect 17328 20828 20300 20856
rect 22370 20816 22376 20868
rect 22428 20856 22434 20868
rect 22480 20856 22508 20887
rect 22922 20884 22928 20936
rect 22980 20884 22986 20936
rect 23106 20884 23112 20936
rect 23164 20884 23170 20936
rect 23216 20924 23244 20964
rect 23658 20952 23664 21004
rect 23716 20992 23722 21004
rect 24854 20992 24860 21004
rect 23716 20964 24860 20992
rect 23716 20952 23722 20964
rect 24854 20952 24860 20964
rect 24912 20952 24918 21004
rect 25774 20952 25780 21004
rect 25832 20992 25838 21004
rect 27249 20995 27307 21001
rect 25832 20964 27016 20992
rect 25832 20952 25838 20964
rect 23293 20927 23351 20933
rect 23293 20924 23305 20927
rect 23216 20896 23305 20924
rect 23293 20893 23305 20896
rect 23339 20893 23351 20927
rect 23293 20887 23351 20893
rect 23477 20927 23535 20933
rect 23477 20893 23489 20927
rect 23523 20893 23535 20927
rect 23477 20887 23535 20893
rect 22428 20828 22508 20856
rect 23124 20856 23152 20884
rect 23492 20856 23520 20887
rect 23934 20884 23940 20936
rect 23992 20924 23998 20936
rect 26510 20924 26516 20936
rect 23992 20896 26516 20924
rect 23992 20884 23998 20896
rect 26510 20884 26516 20896
rect 26568 20884 26574 20936
rect 26988 20933 27016 20964
rect 27249 20961 27261 20995
rect 27295 20992 27307 20995
rect 27982 20992 27988 21004
rect 27295 20964 27988 20992
rect 27295 20961 27307 20964
rect 27249 20955 27307 20961
rect 27982 20952 27988 20964
rect 28040 20952 28046 21004
rect 29917 20995 29975 21001
rect 29917 20961 29929 20995
rect 29963 20992 29975 20995
rect 30190 20992 30196 21004
rect 29963 20964 30196 20992
rect 29963 20961 29975 20964
rect 29917 20955 29975 20961
rect 30190 20952 30196 20964
rect 30248 20992 30254 21004
rect 31220 20992 31248 21032
rect 30248 20964 31248 20992
rect 31312 20964 32168 20992
rect 30248 20952 30254 20964
rect 26973 20927 27031 20933
rect 26973 20893 26985 20927
rect 27019 20924 27031 20927
rect 27062 20924 27068 20936
rect 27019 20896 27068 20924
rect 27019 20893 27031 20896
rect 26973 20887 27031 20893
rect 27062 20884 27068 20896
rect 27120 20884 27126 20936
rect 29822 20884 29828 20936
rect 29880 20884 29886 20936
rect 30009 20927 30067 20933
rect 30009 20893 30021 20927
rect 30055 20893 30067 20927
rect 30009 20887 30067 20893
rect 30101 20927 30159 20933
rect 30101 20893 30113 20927
rect 30147 20924 30159 20927
rect 30282 20924 30288 20936
rect 30147 20896 30288 20924
rect 30147 20893 30159 20896
rect 30101 20887 30159 20893
rect 23124 20828 23520 20856
rect 30024 20856 30052 20887
rect 30282 20884 30288 20896
rect 30340 20884 30346 20936
rect 30374 20884 30380 20936
rect 30432 20924 30438 20936
rect 30650 20924 30656 20936
rect 30432 20896 30656 20924
rect 30432 20884 30438 20896
rect 30650 20884 30656 20896
rect 30708 20884 30714 20936
rect 30837 20927 30895 20933
rect 30837 20893 30849 20927
rect 30883 20893 30895 20927
rect 30837 20887 30895 20893
rect 30392 20856 30420 20884
rect 30024 20828 30420 20856
rect 22428 20816 22434 20828
rect 15804 20760 17080 20788
rect 15804 20748 15810 20760
rect 17126 20748 17132 20800
rect 17184 20788 17190 20800
rect 19613 20791 19671 20797
rect 19613 20788 19625 20791
rect 17184 20760 19625 20788
rect 17184 20748 17190 20760
rect 19613 20757 19625 20760
rect 19659 20757 19671 20791
rect 19613 20751 19671 20757
rect 21634 20748 21640 20800
rect 21692 20748 21698 20800
rect 22462 20748 22468 20800
rect 22520 20788 22526 20800
rect 22557 20791 22615 20797
rect 22557 20788 22569 20791
rect 22520 20760 22569 20788
rect 22520 20748 22526 20760
rect 22557 20757 22569 20760
rect 22603 20757 22615 20791
rect 22557 20751 22615 20757
rect 24946 20748 24952 20800
rect 25004 20788 25010 20800
rect 27249 20791 27307 20797
rect 27249 20788 27261 20791
rect 25004 20760 27261 20788
rect 25004 20748 25010 20760
rect 27249 20757 27261 20760
rect 27295 20757 27307 20791
rect 27249 20751 27307 20757
rect 29638 20748 29644 20800
rect 29696 20748 29702 20800
rect 30852 20788 30880 20887
rect 30926 20884 30932 20936
rect 30984 20924 30990 20936
rect 31021 20927 31079 20933
rect 31021 20924 31033 20927
rect 30984 20896 31033 20924
rect 30984 20884 30990 20896
rect 31021 20893 31033 20896
rect 31067 20893 31079 20927
rect 31021 20887 31079 20893
rect 31113 20927 31171 20933
rect 31113 20893 31125 20927
rect 31159 20924 31171 20927
rect 31202 20924 31208 20936
rect 31159 20896 31208 20924
rect 31159 20893 31171 20896
rect 31113 20887 31171 20893
rect 31036 20856 31064 20887
rect 31202 20884 31208 20896
rect 31260 20884 31266 20936
rect 31312 20933 31340 20964
rect 31297 20927 31355 20933
rect 31297 20893 31309 20927
rect 31343 20893 31355 20927
rect 31297 20887 31355 20893
rect 31389 20927 31447 20933
rect 31389 20893 31401 20927
rect 31435 20924 31447 20927
rect 31435 20896 31984 20924
rect 31435 20893 31447 20896
rect 31389 20887 31447 20893
rect 31956 20868 31984 20896
rect 31036 20828 31248 20856
rect 31110 20788 31116 20800
rect 30852 20760 31116 20788
rect 31110 20748 31116 20760
rect 31168 20748 31174 20800
rect 31220 20788 31248 20828
rect 31570 20816 31576 20868
rect 31628 20816 31634 20868
rect 31938 20816 31944 20868
rect 31996 20816 32002 20868
rect 31386 20788 31392 20800
rect 31220 20760 31392 20788
rect 31386 20748 31392 20760
rect 31444 20788 31450 20800
rect 31757 20791 31815 20797
rect 31757 20788 31769 20791
rect 31444 20760 31769 20788
rect 31444 20748 31450 20760
rect 31757 20757 31769 20760
rect 31803 20757 31815 20791
rect 32140 20788 32168 20964
rect 32692 20964 34928 20992
rect 32490 20884 32496 20936
rect 32548 20884 32554 20936
rect 32214 20816 32220 20868
rect 32272 20856 32278 20868
rect 32692 20865 32720 20964
rect 32769 20927 32827 20933
rect 32769 20893 32781 20927
rect 32815 20893 32827 20927
rect 32769 20887 32827 20893
rect 32861 20927 32919 20933
rect 32861 20893 32873 20927
rect 32907 20924 32919 20927
rect 33134 20924 33140 20936
rect 32907 20896 33140 20924
rect 32907 20893 32919 20896
rect 32861 20887 32919 20893
rect 32677 20859 32735 20865
rect 32677 20856 32689 20859
rect 32272 20828 32689 20856
rect 32272 20816 32278 20828
rect 32677 20825 32689 20828
rect 32723 20825 32735 20859
rect 32677 20819 32735 20825
rect 32582 20788 32588 20800
rect 32140 20760 32588 20788
rect 31757 20751 31815 20757
rect 32582 20748 32588 20760
rect 32640 20788 32646 20800
rect 32784 20788 32812 20887
rect 33134 20884 33140 20896
rect 33192 20884 33198 20936
rect 34900 20933 34928 20964
rect 35176 20933 35204 21032
rect 35437 21029 35449 21063
rect 35483 21060 35495 21063
rect 37274 21060 37280 21072
rect 35483 21032 37280 21060
rect 35483 21029 35495 21032
rect 35437 21023 35495 21029
rect 37274 21020 37280 21032
rect 37332 21020 37338 21072
rect 37458 21020 37464 21072
rect 37516 21020 37522 21072
rect 37476 20992 37504 21020
rect 37384 20964 37504 20992
rect 37568 20992 37596 21100
rect 38562 21088 38568 21140
rect 38620 21128 38626 21140
rect 38749 21131 38807 21137
rect 38749 21128 38761 21131
rect 38620 21100 38761 21128
rect 38620 21088 38626 21100
rect 38749 21097 38761 21100
rect 38795 21097 38807 21131
rect 38749 21091 38807 21097
rect 39206 21088 39212 21140
rect 39264 21128 39270 21140
rect 39853 21131 39911 21137
rect 39853 21128 39865 21131
rect 39264 21100 39865 21128
rect 39264 21088 39270 21100
rect 39853 21097 39865 21100
rect 39899 21097 39911 21131
rect 39853 21091 39911 21097
rect 38286 21020 38292 21072
rect 38344 21060 38350 21072
rect 38344 21032 40632 21060
rect 38344 21020 38350 21032
rect 37568 20964 38884 20992
rect 34885 20927 34943 20933
rect 34885 20893 34897 20927
rect 34931 20893 34943 20927
rect 34885 20887 34943 20893
rect 35161 20927 35219 20933
rect 35161 20893 35173 20927
rect 35207 20893 35219 20927
rect 35161 20887 35219 20893
rect 35253 20927 35311 20933
rect 35253 20893 35265 20927
rect 35299 20924 35311 20927
rect 35434 20924 35440 20936
rect 35299 20896 35440 20924
rect 35299 20893 35311 20896
rect 35253 20887 35311 20893
rect 35434 20884 35440 20896
rect 35492 20884 35498 20936
rect 35526 20884 35532 20936
rect 35584 20884 35590 20936
rect 35622 20927 35680 20933
rect 35622 20893 35634 20927
rect 35668 20893 35680 20927
rect 35622 20887 35680 20893
rect 34698 20856 34704 20868
rect 32876 20828 34704 20856
rect 32876 20800 32904 20828
rect 34698 20816 34704 20828
rect 34756 20856 34762 20868
rect 35069 20859 35127 20865
rect 35069 20856 35081 20859
rect 34756 20828 35081 20856
rect 34756 20816 34762 20828
rect 35069 20825 35081 20828
rect 35115 20825 35127 20859
rect 35069 20819 35127 20825
rect 32640 20760 32812 20788
rect 32640 20748 32646 20760
rect 32858 20748 32864 20800
rect 32916 20748 32922 20800
rect 33410 20748 33416 20800
rect 33468 20788 33474 20800
rect 33870 20788 33876 20800
rect 33468 20760 33876 20788
rect 33468 20748 33474 20760
rect 33870 20748 33876 20760
rect 33928 20748 33934 20800
rect 34514 20748 34520 20800
rect 34572 20788 34578 20800
rect 35636 20788 35664 20887
rect 35894 20884 35900 20936
rect 35952 20884 35958 20936
rect 35994 20927 36052 20933
rect 35994 20893 36006 20927
rect 36040 20924 36052 20927
rect 36354 20924 36360 20936
rect 36040 20896 36360 20924
rect 36040 20893 36052 20896
rect 35994 20887 36052 20893
rect 36354 20884 36360 20896
rect 36412 20884 36418 20936
rect 36722 20884 36728 20936
rect 36780 20924 36786 20936
rect 37384 20933 37412 20964
rect 37369 20927 37427 20933
rect 36780 20896 37320 20924
rect 36780 20884 36786 20896
rect 35710 20816 35716 20868
rect 35768 20856 35774 20868
rect 35805 20859 35863 20865
rect 35805 20856 35817 20859
rect 35768 20828 35817 20856
rect 35768 20816 35774 20828
rect 35805 20825 35817 20828
rect 35851 20825 35863 20859
rect 37182 20856 37188 20868
rect 35805 20819 35863 20825
rect 36188 20828 37188 20856
rect 36188 20797 36216 20828
rect 37182 20816 37188 20828
rect 37240 20816 37246 20868
rect 37292 20856 37320 20896
rect 37369 20893 37381 20927
rect 37415 20893 37427 20927
rect 37369 20887 37427 20893
rect 37458 20884 37464 20936
rect 37516 20884 37522 20936
rect 37734 20884 37740 20936
rect 37792 20884 37798 20936
rect 37875 20927 37933 20933
rect 37875 20893 37887 20927
rect 37921 20924 37933 20927
rect 38010 20924 38016 20936
rect 37921 20896 38016 20924
rect 37921 20893 37933 20896
rect 37875 20887 37933 20893
rect 38010 20884 38016 20896
rect 38068 20884 38074 20936
rect 37645 20859 37703 20865
rect 37645 20856 37657 20859
rect 37292 20828 37657 20856
rect 37645 20825 37657 20828
rect 37691 20825 37703 20859
rect 38749 20859 38807 20865
rect 38749 20856 38761 20859
rect 37645 20819 37703 20825
rect 37752 20828 38761 20856
rect 34572 20760 35664 20788
rect 36173 20791 36231 20797
rect 34572 20748 34578 20760
rect 36173 20757 36185 20791
rect 36219 20757 36231 20791
rect 36173 20751 36231 20757
rect 36630 20748 36636 20800
rect 36688 20788 36694 20800
rect 37752 20788 37780 20828
rect 38749 20825 38761 20828
rect 38795 20825 38807 20859
rect 38856 20856 38884 20964
rect 38930 20952 38936 21004
rect 38988 20992 38994 21004
rect 39482 20992 39488 21004
rect 38988 20964 39488 20992
rect 38988 20952 38994 20964
rect 39482 20952 39488 20964
rect 39540 20952 39546 21004
rect 39758 20952 39764 21004
rect 39816 20992 39822 21004
rect 40037 20995 40095 21001
rect 40037 20992 40049 20995
rect 39816 20964 40049 20992
rect 39816 20952 39822 20964
rect 40037 20961 40049 20964
rect 40083 20961 40095 20995
rect 40037 20955 40095 20961
rect 39025 20927 39083 20933
rect 39025 20893 39037 20927
rect 39071 20924 39083 20927
rect 39666 20924 39672 20936
rect 39071 20896 39672 20924
rect 39071 20893 39083 20896
rect 39025 20887 39083 20893
rect 39666 20884 39672 20896
rect 39724 20884 39730 20936
rect 39850 20884 39856 20936
rect 39908 20884 39914 20936
rect 40604 20933 40632 21032
rect 40129 20927 40187 20933
rect 40129 20893 40141 20927
rect 40175 20893 40187 20927
rect 40129 20887 40187 20893
rect 40589 20927 40647 20933
rect 40589 20893 40601 20927
rect 40635 20893 40647 20927
rect 40589 20887 40647 20893
rect 40144 20856 40172 20887
rect 38856 20828 40172 20856
rect 40405 20859 40463 20865
rect 38749 20819 38807 20825
rect 40405 20825 40417 20859
rect 40451 20825 40463 20859
rect 40405 20819 40463 20825
rect 36688 20760 37780 20788
rect 36688 20748 36694 20760
rect 38010 20748 38016 20800
rect 38068 20748 38074 20800
rect 39206 20748 39212 20800
rect 39264 20748 39270 20800
rect 40313 20791 40371 20797
rect 40313 20757 40325 20791
rect 40359 20788 40371 20791
rect 40420 20788 40448 20819
rect 40359 20760 40448 20788
rect 40359 20757 40371 20760
rect 40313 20751 40371 20757
rect 40770 20748 40776 20800
rect 40828 20748 40834 20800
rect 1104 20698 41400 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 41400 20698
rect 1104 20624 41400 20646
rect 5810 20544 5816 20596
rect 5868 20544 5874 20596
rect 7650 20544 7656 20596
rect 7708 20544 7714 20596
rect 8849 20587 8907 20593
rect 8849 20553 8861 20587
rect 8895 20553 8907 20587
rect 8849 20547 8907 20553
rect 2685 20519 2743 20525
rect 2685 20485 2697 20519
rect 2731 20516 2743 20519
rect 2958 20516 2964 20528
rect 2731 20488 2964 20516
rect 2731 20485 2743 20488
rect 2685 20479 2743 20485
rect 2958 20476 2964 20488
rect 3016 20516 3022 20528
rect 5902 20516 5908 20528
rect 3016 20488 5908 20516
rect 3016 20476 3022 20488
rect 5902 20476 5908 20488
rect 5960 20516 5966 20528
rect 6822 20516 6828 20528
rect 5960 20488 6828 20516
rect 5960 20476 5966 20488
rect 6822 20476 6828 20488
rect 6880 20476 6886 20528
rect 7668 20516 7696 20544
rect 7929 20519 7987 20525
rect 7929 20516 7941 20519
rect 7668 20488 7941 20516
rect 7929 20485 7941 20488
rect 7975 20485 7987 20519
rect 7929 20479 7987 20485
rect 2590 20408 2596 20460
rect 2648 20448 2654 20460
rect 4341 20451 4399 20457
rect 4341 20448 4353 20451
rect 2648 20420 4353 20448
rect 2648 20408 2654 20420
rect 4341 20417 4353 20420
rect 4387 20417 4399 20451
rect 4341 20411 4399 20417
rect 4982 20408 4988 20460
rect 5040 20448 5046 20460
rect 5261 20451 5319 20457
rect 5261 20448 5273 20451
rect 5040 20420 5273 20448
rect 5040 20408 5046 20420
rect 5261 20417 5273 20420
rect 5307 20417 5319 20451
rect 5261 20411 5319 20417
rect 2682 20340 2688 20392
rect 2740 20380 2746 20392
rect 3421 20383 3479 20389
rect 3421 20380 3433 20383
rect 2740 20352 3433 20380
rect 2740 20340 2746 20352
rect 3421 20349 3433 20352
rect 3467 20349 3479 20383
rect 3697 20383 3755 20389
rect 3697 20380 3709 20383
rect 3421 20343 3479 20349
rect 3620 20352 3709 20380
rect 3436 20256 3464 20343
rect 3620 20256 3648 20352
rect 3697 20349 3709 20352
rect 3743 20349 3755 20383
rect 3697 20343 3755 20349
rect 3418 20204 3424 20256
rect 3476 20204 3482 20256
rect 3602 20204 3608 20256
rect 3660 20204 3666 20256
rect 5276 20244 5304 20411
rect 5350 20408 5356 20460
rect 5408 20448 5414 20460
rect 5445 20451 5503 20457
rect 5445 20448 5457 20451
rect 5408 20420 5457 20448
rect 5408 20408 5414 20420
rect 5445 20417 5457 20420
rect 5491 20417 5503 20451
rect 5445 20411 5503 20417
rect 5537 20451 5595 20457
rect 5537 20417 5549 20451
rect 5583 20417 5595 20451
rect 5537 20411 5595 20417
rect 5629 20451 5687 20457
rect 5629 20417 5641 20451
rect 5675 20448 5687 20451
rect 5994 20448 6000 20460
rect 5675 20420 6000 20448
rect 5675 20417 5687 20420
rect 5629 20411 5687 20417
rect 5460 20312 5488 20411
rect 5552 20380 5580 20411
rect 5994 20408 6000 20420
rect 6052 20448 6058 20460
rect 6052 20420 7052 20448
rect 6052 20408 6058 20420
rect 6914 20380 6920 20392
rect 5552 20352 6920 20380
rect 6914 20340 6920 20352
rect 6972 20340 6978 20392
rect 7024 20380 7052 20420
rect 7650 20408 7656 20460
rect 7708 20408 7714 20460
rect 7742 20408 7748 20460
rect 7800 20448 7806 20460
rect 7837 20451 7895 20457
rect 7837 20448 7849 20451
rect 7800 20420 7849 20448
rect 7800 20408 7806 20420
rect 7837 20417 7849 20420
rect 7883 20417 7895 20451
rect 7837 20411 7895 20417
rect 8018 20408 8024 20460
rect 8076 20408 8082 20460
rect 8757 20451 8815 20457
rect 8757 20417 8769 20451
rect 8803 20448 8815 20451
rect 8864 20448 8892 20547
rect 9858 20544 9864 20596
rect 9916 20544 9922 20596
rect 10318 20544 10324 20596
rect 10376 20544 10382 20596
rect 10962 20544 10968 20596
rect 11020 20544 11026 20596
rect 11701 20587 11759 20593
rect 11701 20584 11713 20587
rect 11072 20556 11713 20584
rect 9309 20519 9367 20525
rect 9309 20485 9321 20519
rect 9355 20516 9367 20519
rect 9950 20516 9956 20528
rect 9355 20488 9956 20516
rect 9355 20485 9367 20488
rect 9309 20479 9367 20485
rect 9950 20476 9956 20488
rect 10008 20516 10014 20528
rect 10336 20516 10364 20544
rect 10980 20516 11008 20544
rect 10008 20488 10364 20516
rect 10796 20488 11008 20516
rect 10008 20476 10014 20488
rect 8803 20420 8892 20448
rect 8803 20417 8815 20420
rect 8757 20411 8815 20417
rect 9214 20408 9220 20460
rect 9272 20408 9278 20460
rect 9677 20451 9735 20457
rect 9677 20448 9689 20451
rect 9508 20420 9689 20448
rect 8036 20380 8064 20408
rect 9508 20389 9536 20420
rect 9677 20417 9689 20420
rect 9723 20448 9735 20451
rect 10502 20448 10508 20460
rect 9723 20420 10508 20448
rect 9723 20417 9735 20420
rect 9677 20411 9735 20417
rect 10502 20408 10508 20420
rect 10560 20408 10566 20460
rect 10796 20457 10824 20488
rect 10781 20451 10839 20457
rect 10781 20417 10793 20451
rect 10827 20417 10839 20451
rect 10781 20411 10839 20417
rect 10965 20451 11023 20457
rect 10965 20417 10977 20451
rect 11011 20448 11023 20451
rect 11072 20448 11100 20556
rect 11701 20553 11713 20556
rect 11747 20553 11759 20587
rect 12342 20584 12348 20596
rect 11701 20547 11759 20553
rect 11808 20556 12348 20584
rect 11808 20516 11836 20556
rect 12342 20544 12348 20556
rect 12400 20584 12406 20596
rect 12400 20556 14780 20584
rect 12400 20544 12406 20556
rect 13078 20516 13084 20528
rect 11011 20420 11100 20448
rect 11164 20488 11836 20516
rect 11900 20488 13084 20516
rect 11011 20417 11023 20420
rect 10965 20411 11023 20417
rect 9493 20383 9551 20389
rect 7024 20352 8800 20380
rect 7742 20312 7748 20324
rect 5460 20284 7748 20312
rect 7742 20272 7748 20284
rect 7800 20312 7806 20324
rect 8018 20312 8024 20324
rect 7800 20284 8024 20312
rect 7800 20272 7806 20284
rect 8018 20272 8024 20284
rect 8076 20272 8082 20324
rect 8772 20312 8800 20352
rect 9493 20349 9505 20383
rect 9539 20349 9551 20383
rect 9493 20343 9551 20349
rect 9858 20340 9864 20392
rect 9916 20380 9922 20392
rect 10980 20380 11008 20411
rect 9916 20352 11008 20380
rect 9916 20340 9922 20352
rect 11164 20312 11192 20488
rect 11517 20451 11575 20457
rect 11517 20417 11529 20451
rect 11563 20448 11575 20451
rect 11790 20448 11796 20460
rect 11563 20420 11796 20448
rect 11563 20417 11575 20420
rect 11517 20411 11575 20417
rect 11790 20408 11796 20420
rect 11848 20408 11854 20460
rect 11900 20457 11928 20488
rect 13078 20476 13084 20488
rect 13136 20476 13142 20528
rect 13906 20476 13912 20528
rect 13964 20476 13970 20528
rect 14752 20516 14780 20556
rect 14826 20544 14832 20596
rect 14884 20544 14890 20596
rect 15930 20584 15936 20596
rect 14936 20556 15936 20584
rect 14936 20516 14964 20556
rect 15930 20544 15936 20556
rect 15988 20584 15994 20596
rect 16301 20587 16359 20593
rect 16301 20584 16313 20587
rect 15988 20556 16313 20584
rect 15988 20544 15994 20556
rect 16301 20553 16313 20556
rect 16347 20553 16359 20587
rect 16301 20547 16359 20553
rect 19889 20587 19947 20593
rect 19889 20553 19901 20587
rect 19935 20584 19947 20587
rect 19978 20584 19984 20596
rect 19935 20556 19984 20584
rect 19935 20553 19947 20556
rect 19889 20547 19947 20553
rect 19978 20544 19984 20556
rect 20036 20544 20042 20596
rect 22922 20544 22928 20596
rect 22980 20584 22986 20596
rect 23293 20587 23351 20593
rect 23293 20584 23305 20587
rect 22980 20556 23305 20584
rect 22980 20544 22986 20556
rect 23293 20553 23305 20556
rect 23339 20553 23351 20587
rect 23293 20547 23351 20553
rect 25222 20544 25228 20596
rect 25280 20584 25286 20596
rect 25958 20584 25964 20596
rect 25280 20556 25964 20584
rect 25280 20544 25286 20556
rect 25958 20544 25964 20556
rect 26016 20544 26022 20596
rect 26602 20544 26608 20596
rect 26660 20584 26666 20596
rect 28537 20587 28595 20593
rect 28537 20584 28549 20587
rect 26660 20556 28549 20584
rect 26660 20544 26666 20556
rect 28537 20553 28549 20556
rect 28583 20553 28595 20587
rect 28537 20547 28595 20553
rect 28966 20556 33456 20584
rect 15654 20516 15660 20528
rect 14752 20488 14964 20516
rect 15028 20488 15660 20516
rect 11885 20451 11943 20457
rect 11885 20417 11897 20451
rect 11931 20417 11943 20451
rect 11885 20411 11943 20417
rect 12069 20451 12127 20457
rect 12069 20417 12081 20451
rect 12115 20417 12127 20451
rect 12069 20411 12127 20417
rect 11698 20340 11704 20392
rect 11756 20380 11762 20392
rect 11900 20380 11928 20411
rect 11756 20352 11928 20380
rect 12084 20380 12112 20411
rect 12158 20408 12164 20460
rect 12216 20408 12222 20460
rect 12253 20451 12311 20457
rect 12253 20417 12265 20451
rect 12299 20448 12311 20451
rect 12342 20448 12348 20460
rect 12299 20420 12348 20448
rect 12299 20417 12311 20420
rect 12253 20411 12311 20417
rect 12342 20408 12348 20420
rect 12400 20408 12406 20460
rect 12710 20408 12716 20460
rect 12768 20408 12774 20460
rect 15028 20457 15056 20488
rect 15654 20476 15660 20488
rect 15712 20476 15718 20528
rect 15746 20476 15752 20528
rect 15804 20476 15810 20528
rect 16666 20476 16672 20528
rect 16724 20516 16730 20528
rect 16761 20519 16819 20525
rect 16761 20516 16773 20519
rect 16724 20488 16773 20516
rect 16724 20476 16730 20488
rect 16761 20485 16773 20488
rect 16807 20485 16819 20519
rect 16761 20479 16819 20485
rect 19426 20476 19432 20528
rect 19484 20516 19490 20528
rect 20070 20516 20076 20528
rect 19484 20488 20076 20516
rect 19484 20476 19490 20488
rect 20070 20476 20076 20488
rect 20128 20516 20134 20528
rect 20165 20519 20223 20525
rect 20165 20516 20177 20519
rect 20128 20488 20177 20516
rect 20128 20476 20134 20488
rect 20165 20485 20177 20488
rect 20211 20485 20223 20519
rect 20809 20519 20867 20525
rect 20809 20516 20821 20519
rect 20165 20479 20223 20485
rect 20456 20488 20821 20516
rect 15013 20451 15071 20457
rect 15013 20417 15025 20451
rect 15059 20417 15071 20451
rect 15013 20411 15071 20417
rect 15197 20451 15255 20457
rect 15197 20417 15209 20451
rect 15243 20448 15255 20451
rect 15289 20451 15347 20457
rect 15289 20448 15301 20451
rect 15243 20420 15301 20448
rect 15243 20417 15255 20420
rect 15197 20411 15255 20417
rect 15289 20417 15301 20420
rect 15335 20448 15347 20451
rect 15378 20448 15384 20460
rect 15335 20420 15384 20448
rect 15335 20417 15347 20420
rect 15289 20411 15347 20417
rect 15378 20408 15384 20420
rect 15436 20408 15442 20460
rect 15470 20408 15476 20460
rect 15528 20408 15534 20460
rect 15565 20451 15623 20457
rect 15565 20417 15577 20451
rect 15611 20448 15623 20451
rect 15764 20448 15792 20476
rect 20456 20460 20484 20488
rect 20809 20485 20821 20488
rect 20855 20485 20867 20519
rect 20809 20479 20867 20485
rect 21039 20519 21097 20525
rect 21039 20485 21051 20519
rect 21085 20516 21097 20519
rect 21450 20516 21456 20528
rect 21085 20488 21456 20516
rect 21085 20485 21097 20488
rect 21039 20479 21097 20485
rect 21450 20476 21456 20488
rect 21508 20476 21514 20528
rect 22833 20519 22891 20525
rect 22833 20485 22845 20519
rect 22879 20516 22891 20519
rect 25593 20519 25651 20525
rect 22879 20488 23336 20516
rect 22879 20485 22891 20488
rect 22833 20479 22891 20485
rect 23308 20460 23336 20488
rect 25593 20485 25605 20519
rect 25639 20516 25651 20519
rect 26142 20516 26148 20528
rect 25639 20488 26148 20516
rect 25639 20485 25651 20488
rect 25593 20479 25651 20485
rect 26142 20476 26148 20488
rect 26200 20476 26206 20528
rect 26234 20476 26240 20528
rect 26292 20516 26298 20528
rect 26292 20488 28120 20516
rect 26292 20476 26298 20488
rect 15611 20420 15792 20448
rect 15611 20417 15623 20420
rect 15565 20411 15623 20417
rect 16114 20408 16120 20460
rect 16172 20408 16178 20460
rect 17402 20408 17408 20460
rect 17460 20408 17466 20460
rect 19889 20451 19947 20457
rect 19889 20417 19901 20451
rect 19935 20448 19947 20451
rect 20438 20448 20444 20460
rect 19935 20420 20444 20448
rect 19935 20417 19947 20420
rect 19889 20411 19947 20417
rect 20438 20408 20444 20420
rect 20496 20408 20502 20460
rect 20717 20451 20775 20457
rect 20717 20417 20729 20451
rect 20763 20417 20775 20451
rect 20717 20411 20775 20417
rect 20901 20451 20959 20457
rect 20901 20417 20913 20451
rect 20947 20448 20959 20451
rect 23109 20451 23167 20457
rect 20947 20420 21036 20448
rect 20947 20417 20959 20420
rect 20901 20411 20959 20417
rect 12084 20352 13032 20380
rect 11756 20340 11762 20352
rect 12084 20312 12112 20352
rect 12618 20312 12624 20324
rect 8128 20284 8708 20312
rect 8772 20284 11192 20312
rect 11808 20284 12112 20312
rect 12452 20284 12624 20312
rect 8128 20244 8156 20284
rect 5276 20216 8156 20244
rect 8202 20204 8208 20256
rect 8260 20204 8266 20256
rect 8570 20204 8576 20256
rect 8628 20204 8634 20256
rect 8680 20244 8708 20284
rect 11808 20256 11836 20284
rect 10410 20244 10416 20256
rect 8680 20216 10416 20244
rect 10410 20204 10416 20216
rect 10468 20204 10474 20256
rect 10594 20204 10600 20256
rect 10652 20204 10658 20256
rect 11241 20247 11299 20253
rect 11241 20213 11253 20247
rect 11287 20244 11299 20247
rect 11606 20244 11612 20256
rect 11287 20216 11612 20244
rect 11287 20213 11299 20216
rect 11241 20207 11299 20213
rect 11606 20204 11612 20216
rect 11664 20204 11670 20256
rect 11790 20204 11796 20256
rect 11848 20204 11854 20256
rect 12452 20253 12480 20284
rect 12618 20272 12624 20284
rect 12676 20272 12682 20324
rect 12437 20247 12495 20253
rect 12437 20213 12449 20247
rect 12483 20213 12495 20247
rect 12437 20207 12495 20213
rect 12526 20204 12532 20256
rect 12584 20204 12590 20256
rect 13004 20244 13032 20352
rect 13078 20340 13084 20392
rect 13136 20340 13142 20392
rect 13354 20340 13360 20392
rect 13412 20340 13418 20392
rect 15838 20380 15844 20392
rect 14752 20352 15844 20380
rect 14752 20244 14780 20352
rect 15838 20340 15844 20352
rect 15896 20380 15902 20392
rect 16025 20383 16083 20389
rect 16025 20380 16037 20383
rect 15896 20352 16037 20380
rect 15896 20340 15902 20352
rect 16025 20349 16037 20352
rect 16071 20349 16083 20383
rect 16025 20343 16083 20349
rect 19058 20340 19064 20392
rect 19116 20380 19122 20392
rect 20162 20380 20168 20392
rect 19116 20352 20168 20380
rect 19116 20340 19122 20352
rect 20162 20340 20168 20352
rect 20220 20380 20226 20392
rect 20732 20380 20760 20411
rect 21008 20392 21036 20420
rect 23109 20417 23121 20451
rect 23155 20417 23167 20451
rect 23109 20411 23167 20417
rect 20220 20352 20760 20380
rect 20220 20340 20226 20352
rect 20990 20340 20996 20392
rect 21048 20340 21054 20392
rect 21082 20340 21088 20392
rect 21140 20380 21146 20392
rect 21177 20383 21235 20389
rect 21177 20380 21189 20383
rect 21140 20352 21189 20380
rect 21140 20340 21146 20352
rect 21177 20349 21189 20352
rect 21223 20349 21235 20383
rect 21177 20343 21235 20349
rect 23017 20383 23075 20389
rect 23017 20349 23029 20383
rect 23063 20349 23075 20383
rect 23124 20380 23152 20411
rect 23290 20408 23296 20460
rect 23348 20408 23354 20460
rect 23566 20408 23572 20460
rect 23624 20408 23630 20460
rect 24394 20408 24400 20460
rect 24452 20448 24458 20460
rect 25961 20451 26019 20457
rect 25961 20448 25973 20451
rect 24452 20420 25973 20448
rect 24452 20408 24458 20420
rect 25961 20417 25973 20420
rect 26007 20448 26019 20451
rect 27430 20448 27436 20460
rect 26007 20420 27436 20448
rect 26007 20417 26019 20420
rect 25961 20411 26019 20417
rect 27430 20408 27436 20420
rect 27488 20408 27494 20460
rect 27617 20451 27675 20457
rect 27617 20417 27629 20451
rect 27663 20417 27675 20451
rect 28092 20448 28120 20488
rect 28166 20476 28172 20528
rect 28224 20476 28230 20528
rect 28350 20476 28356 20528
rect 28408 20525 28414 20528
rect 28408 20519 28427 20525
rect 28415 20516 28427 20519
rect 28966 20516 28994 20556
rect 33428 20528 33456 20556
rect 35618 20544 35624 20596
rect 35676 20584 35682 20596
rect 37458 20584 37464 20596
rect 35676 20556 37464 20584
rect 35676 20544 35682 20556
rect 37458 20544 37464 20556
rect 37516 20544 37522 20596
rect 37737 20587 37795 20593
rect 37737 20553 37749 20587
rect 37783 20584 37795 20587
rect 38930 20584 38936 20596
rect 37783 20556 38936 20584
rect 37783 20553 37795 20556
rect 37737 20547 37795 20553
rect 38930 20544 38936 20556
rect 38988 20544 38994 20596
rect 39206 20544 39212 20596
rect 39264 20544 39270 20596
rect 40034 20544 40040 20596
rect 40092 20584 40098 20596
rect 40313 20587 40371 20593
rect 40313 20584 40325 20587
rect 40092 20556 40325 20584
rect 40092 20544 40098 20556
rect 40313 20553 40325 20556
rect 40359 20553 40371 20587
rect 40313 20547 40371 20553
rect 28415 20488 28994 20516
rect 28415 20485 28427 20488
rect 28408 20479 28427 20485
rect 28408 20476 28414 20479
rect 30006 20476 30012 20528
rect 30064 20476 30070 20528
rect 32030 20516 32036 20528
rect 31726 20488 32036 20516
rect 30024 20448 30052 20476
rect 28092 20420 30052 20448
rect 27617 20411 27675 20417
rect 23584 20380 23612 20408
rect 26878 20380 26884 20392
rect 23124 20352 26884 20380
rect 23017 20343 23075 20349
rect 15010 20272 15016 20324
rect 15068 20312 15074 20324
rect 16390 20312 16396 20324
rect 15068 20284 16396 20312
rect 15068 20272 15074 20284
rect 16390 20272 16396 20284
rect 16448 20272 16454 20324
rect 19334 20272 19340 20324
rect 19392 20312 19398 20324
rect 19978 20312 19984 20324
rect 19392 20284 19984 20312
rect 19392 20272 19398 20284
rect 19978 20272 19984 20284
rect 20036 20272 20042 20324
rect 23032 20312 23060 20343
rect 26878 20340 26884 20352
rect 26936 20340 26942 20392
rect 23474 20312 23480 20324
rect 23032 20284 23480 20312
rect 23474 20272 23480 20284
rect 23532 20312 23538 20324
rect 26234 20312 26240 20324
rect 23532 20284 26240 20312
rect 23532 20272 23538 20284
rect 26234 20272 26240 20284
rect 26292 20272 26298 20324
rect 13004 20216 14780 20244
rect 15105 20247 15163 20253
rect 15105 20213 15117 20247
rect 15151 20244 15163 20247
rect 15194 20244 15200 20256
rect 15151 20216 15200 20244
rect 15151 20213 15163 20216
rect 15105 20207 15163 20213
rect 15194 20204 15200 20216
rect 15252 20204 15258 20256
rect 16298 20204 16304 20256
rect 16356 20244 16362 20256
rect 16850 20244 16856 20256
rect 16356 20216 16856 20244
rect 16356 20204 16362 20216
rect 16850 20204 16856 20216
rect 16908 20204 16914 20256
rect 17218 20204 17224 20256
rect 17276 20204 17282 20256
rect 20254 20204 20260 20256
rect 20312 20244 20318 20256
rect 20533 20247 20591 20253
rect 20533 20244 20545 20247
rect 20312 20216 20545 20244
rect 20312 20204 20318 20216
rect 20533 20213 20545 20216
rect 20579 20213 20591 20247
rect 20533 20207 20591 20213
rect 20898 20204 20904 20256
rect 20956 20244 20962 20256
rect 22370 20244 22376 20256
rect 20956 20216 22376 20244
rect 20956 20204 20962 20216
rect 22370 20204 22376 20216
rect 22428 20244 22434 20256
rect 22833 20247 22891 20253
rect 22833 20244 22845 20247
rect 22428 20216 22845 20244
rect 22428 20204 22434 20216
rect 22833 20213 22845 20216
rect 22879 20213 22891 20247
rect 22833 20207 22891 20213
rect 23014 20204 23020 20256
rect 23072 20244 23078 20256
rect 26050 20244 26056 20256
rect 23072 20216 26056 20244
rect 23072 20204 23078 20216
rect 26050 20204 26056 20216
rect 26108 20204 26114 20256
rect 26896 20244 26924 20340
rect 27632 20324 27660 20411
rect 31570 20408 31576 20460
rect 31628 20408 31634 20460
rect 31294 20380 31300 20392
rect 27724 20352 31300 20380
rect 27614 20272 27620 20324
rect 27672 20272 27678 20324
rect 27724 20244 27752 20352
rect 31294 20340 31300 20352
rect 31352 20340 31358 20392
rect 31386 20340 31392 20392
rect 31444 20380 31450 20392
rect 31726 20380 31754 20488
rect 32030 20476 32036 20488
rect 32088 20476 32094 20528
rect 33410 20476 33416 20528
rect 33468 20476 33474 20528
rect 39224 20516 39252 20544
rect 34072 20488 37596 20516
rect 39224 20488 39988 20516
rect 34072 20392 34100 20488
rect 37568 20460 37596 20488
rect 37277 20451 37335 20457
rect 37277 20417 37289 20451
rect 37323 20417 37335 20451
rect 37277 20411 37335 20417
rect 31444 20352 31754 20380
rect 31444 20340 31450 20352
rect 34054 20340 34060 20392
rect 34112 20340 34118 20392
rect 37292 20380 37320 20411
rect 37366 20408 37372 20460
rect 37424 20448 37430 20460
rect 37461 20451 37519 20457
rect 37461 20448 37473 20451
rect 37424 20420 37473 20448
rect 37424 20408 37430 20420
rect 37461 20417 37473 20420
rect 37507 20417 37519 20451
rect 37461 20411 37519 20417
rect 37292 20352 37412 20380
rect 27890 20272 27896 20324
rect 27948 20312 27954 20324
rect 28442 20312 28448 20324
rect 27948 20284 28448 20312
rect 27948 20272 27954 20284
rect 28442 20272 28448 20284
rect 28500 20272 28506 20324
rect 34146 20312 34152 20324
rect 29288 20284 34152 20312
rect 29288 20256 29316 20284
rect 34146 20272 34152 20284
rect 34204 20272 34210 20324
rect 37384 20256 37412 20352
rect 26896 20216 27752 20244
rect 27798 20204 27804 20256
rect 27856 20204 27862 20256
rect 28353 20247 28411 20253
rect 28353 20213 28365 20247
rect 28399 20244 28411 20247
rect 28994 20244 29000 20256
rect 28399 20216 29000 20244
rect 28399 20213 28411 20216
rect 28353 20207 28411 20213
rect 28994 20204 29000 20216
rect 29052 20204 29058 20256
rect 29270 20204 29276 20256
rect 29328 20204 29334 20256
rect 29546 20204 29552 20256
rect 29604 20244 29610 20256
rect 29822 20244 29828 20256
rect 29604 20216 29828 20244
rect 29604 20204 29610 20216
rect 29822 20204 29828 20216
rect 29880 20204 29886 20256
rect 30650 20204 30656 20256
rect 30708 20244 30714 20256
rect 31478 20244 31484 20256
rect 30708 20216 31484 20244
rect 30708 20204 30714 20216
rect 31478 20204 31484 20216
rect 31536 20204 31542 20256
rect 31570 20204 31576 20256
rect 31628 20244 31634 20256
rect 31757 20247 31815 20253
rect 31757 20244 31769 20247
rect 31628 20216 31769 20244
rect 31628 20204 31634 20216
rect 31757 20213 31769 20216
rect 31803 20213 31815 20247
rect 31757 20207 31815 20213
rect 33410 20204 33416 20256
rect 33468 20244 33474 20256
rect 33778 20244 33784 20256
rect 33468 20216 33784 20244
rect 33468 20204 33474 20216
rect 33778 20204 33784 20216
rect 33836 20204 33842 20256
rect 36078 20204 36084 20256
rect 36136 20244 36142 20256
rect 36538 20244 36544 20256
rect 36136 20216 36544 20244
rect 36136 20204 36142 20216
rect 36538 20204 36544 20216
rect 36596 20244 36602 20256
rect 37277 20247 37335 20253
rect 37277 20244 37289 20247
rect 36596 20216 37289 20244
rect 36596 20204 36602 20216
rect 37277 20213 37289 20216
rect 37323 20213 37335 20247
rect 37277 20207 37335 20213
rect 37366 20204 37372 20256
rect 37424 20204 37430 20256
rect 37476 20244 37504 20411
rect 37550 20408 37556 20460
rect 37608 20408 37614 20460
rect 39393 20451 39451 20457
rect 39393 20448 39405 20451
rect 38856 20420 39405 20448
rect 38856 20392 38884 20420
rect 39393 20417 39405 20420
rect 39439 20417 39451 20451
rect 39393 20411 39451 20417
rect 39577 20451 39635 20457
rect 39577 20417 39589 20451
rect 39623 20448 39635 20451
rect 39758 20448 39764 20460
rect 39623 20420 39764 20448
rect 39623 20417 39635 20420
rect 39577 20411 39635 20417
rect 39758 20408 39764 20420
rect 39816 20408 39822 20460
rect 39960 20457 39988 20488
rect 39945 20451 40003 20457
rect 39945 20417 39957 20451
rect 39991 20417 40003 20451
rect 39945 20411 40003 20417
rect 40129 20451 40187 20457
rect 40129 20417 40141 20451
rect 40175 20448 40187 20451
rect 41230 20448 41236 20460
rect 40175 20420 41236 20448
rect 40175 20417 40187 20420
rect 40129 20411 40187 20417
rect 41230 20408 41236 20420
rect 41288 20408 41294 20460
rect 38838 20340 38844 20392
rect 38896 20340 38902 20392
rect 40144 20284 40816 20312
rect 39393 20247 39451 20253
rect 39393 20244 39405 20247
rect 37476 20216 39405 20244
rect 39393 20213 39405 20216
rect 39439 20213 39451 20247
rect 39393 20207 39451 20213
rect 39574 20204 39580 20256
rect 39632 20244 39638 20256
rect 40144 20253 40172 20284
rect 40788 20256 40816 20284
rect 39761 20247 39819 20253
rect 39761 20244 39773 20247
rect 39632 20216 39773 20244
rect 39632 20204 39638 20216
rect 39761 20213 39773 20216
rect 39807 20213 39819 20247
rect 39761 20207 39819 20213
rect 40129 20247 40187 20253
rect 40129 20213 40141 20247
rect 40175 20213 40187 20247
rect 40129 20207 40187 20213
rect 40770 20204 40776 20256
rect 40828 20204 40834 20256
rect 1104 20154 41400 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 41400 20154
rect 1104 20080 41400 20102
rect 3145 20043 3203 20049
rect 3145 20009 3157 20043
rect 3191 20040 3203 20043
rect 3602 20040 3608 20052
rect 3191 20012 3608 20040
rect 3191 20009 3203 20012
rect 3145 20003 3203 20009
rect 3602 20000 3608 20012
rect 3660 20000 3666 20052
rect 3970 20000 3976 20052
rect 4028 20040 4034 20052
rect 4893 20043 4951 20049
rect 4028 20012 4844 20040
rect 4028 20000 4034 20012
rect 1394 19864 1400 19916
rect 1452 19864 1458 19916
rect 3620 19904 3648 20000
rect 3786 19932 3792 19984
rect 3844 19972 3850 19984
rect 4816 19972 4844 20012
rect 4893 20009 4905 20043
rect 4939 20040 4951 20043
rect 5718 20040 5724 20052
rect 4939 20012 5724 20040
rect 4939 20009 4951 20012
rect 4893 20003 4951 20009
rect 5718 20000 5724 20012
rect 5776 20000 5782 20052
rect 5810 20000 5816 20052
rect 5868 20000 5874 20052
rect 8202 20040 8208 20052
rect 7852 20012 8208 20040
rect 5629 19975 5687 19981
rect 5629 19972 5641 19975
rect 3844 19944 4660 19972
rect 4816 19944 5641 19972
rect 3844 19932 3850 19944
rect 3620 19876 4384 19904
rect 3970 19796 3976 19848
rect 4028 19796 4034 19848
rect 4246 19796 4252 19848
rect 4304 19796 4310 19848
rect 4356 19845 4384 19876
rect 4632 19845 4660 19944
rect 5629 19941 5641 19944
rect 5675 19941 5687 19975
rect 5629 19935 5687 19941
rect 5828 19904 5856 20000
rect 7852 19904 7880 20012
rect 8202 20000 8208 20012
rect 8260 20000 8266 20052
rect 8294 20000 8300 20052
rect 8352 20040 8358 20052
rect 8389 20043 8447 20049
rect 8389 20040 8401 20043
rect 8352 20012 8401 20040
rect 8352 20000 8358 20012
rect 8389 20009 8401 20012
rect 8435 20009 8447 20043
rect 8389 20003 8447 20009
rect 8478 20000 8484 20052
rect 8536 20040 8542 20052
rect 13078 20040 13084 20052
rect 8536 20012 10640 20040
rect 8536 20000 8542 20012
rect 8018 19932 8024 19984
rect 8076 19972 8082 19984
rect 9953 19975 10011 19981
rect 8076 19944 9352 19972
rect 8076 19932 8082 19944
rect 9324 19904 9352 19944
rect 9953 19941 9965 19975
rect 9999 19972 10011 19975
rect 10226 19972 10232 19984
rect 9999 19944 10232 19972
rect 9999 19941 10011 19944
rect 9953 19935 10011 19941
rect 10226 19932 10232 19944
rect 10284 19932 10290 19984
rect 10612 19972 10640 20012
rect 11624 20012 13084 20040
rect 11054 19972 11060 19984
rect 10612 19944 11060 19972
rect 5000 19876 5856 19904
rect 7760 19876 7880 19904
rect 8225 19876 8800 19904
rect 5000 19845 5028 19876
rect 4342 19839 4400 19845
rect 4342 19805 4354 19839
rect 4388 19805 4400 19839
rect 4342 19799 4400 19805
rect 4617 19839 4675 19845
rect 4617 19805 4629 19839
rect 4663 19805 4675 19839
rect 4617 19799 4675 19805
rect 4755 19839 4813 19845
rect 4755 19805 4767 19839
rect 4801 19805 4813 19839
rect 4755 19799 4813 19805
rect 4985 19839 5043 19845
rect 4985 19805 4997 19839
rect 5031 19805 5043 19839
rect 4985 19799 5043 19805
rect 1670 19728 1676 19780
rect 1728 19728 1734 19780
rect 3050 19768 3056 19780
rect 2898 19740 3056 19768
rect 3050 19728 3056 19740
rect 3108 19768 3114 19780
rect 4430 19768 4436 19780
rect 3108 19740 4436 19768
rect 3108 19728 3114 19740
rect 4430 19728 4436 19740
rect 4488 19728 4494 19780
rect 4525 19771 4583 19777
rect 4525 19737 4537 19771
rect 4571 19737 4583 19771
rect 4770 19768 4798 19799
rect 5074 19796 5080 19848
rect 5132 19796 5138 19848
rect 5491 19839 5549 19845
rect 5491 19836 5503 19839
rect 5184 19808 5503 19836
rect 5184 19768 5212 19808
rect 5491 19805 5503 19808
rect 5537 19836 5549 19839
rect 5718 19836 5724 19848
rect 5537 19808 5724 19836
rect 5537 19805 5549 19808
rect 5491 19799 5549 19805
rect 5718 19796 5724 19808
rect 5776 19796 5782 19848
rect 7760 19845 7788 19876
rect 7745 19839 7803 19845
rect 7745 19805 7757 19839
rect 7791 19805 7803 19839
rect 7745 19799 7803 19805
rect 7834 19796 7840 19848
rect 7892 19796 7898 19848
rect 8225 19845 8253 19876
rect 8772 19848 8800 19876
rect 9324 19876 9904 19904
rect 8210 19839 8268 19845
rect 8210 19836 8222 19839
rect 7944 19808 8222 19836
rect 4770 19740 5212 19768
rect 5261 19771 5319 19777
rect 4525 19731 4583 19737
rect 5261 19737 5273 19771
rect 5307 19737 5319 19771
rect 5261 19731 5319 19737
rect 3602 19660 3608 19712
rect 3660 19700 3666 19712
rect 3789 19703 3847 19709
rect 3789 19700 3801 19703
rect 3660 19672 3801 19700
rect 3660 19660 3666 19672
rect 3789 19669 3801 19672
rect 3835 19669 3847 19703
rect 4540 19700 4568 19731
rect 5166 19700 5172 19712
rect 4540 19672 5172 19700
rect 3789 19663 3847 19669
rect 5166 19660 5172 19672
rect 5224 19700 5230 19712
rect 5276 19700 5304 19731
rect 5350 19728 5356 19780
rect 5408 19728 5414 19780
rect 5810 19768 5816 19780
rect 5460 19740 5816 19768
rect 5460 19700 5488 19740
rect 5810 19728 5816 19740
rect 5868 19728 5874 19780
rect 7006 19728 7012 19780
rect 7064 19768 7070 19780
rect 7944 19768 7972 19808
rect 8210 19805 8222 19808
rect 8256 19805 8268 19839
rect 8210 19799 8268 19805
rect 8478 19796 8484 19848
rect 8536 19796 8542 19848
rect 8754 19796 8760 19848
rect 8812 19796 8818 19848
rect 9030 19796 9036 19848
rect 9088 19796 9094 19848
rect 9217 19839 9275 19845
rect 9217 19805 9229 19839
rect 9263 19836 9275 19839
rect 9324 19836 9352 19876
rect 9263 19808 9352 19836
rect 9263 19805 9275 19808
rect 9217 19799 9275 19805
rect 9398 19796 9404 19848
rect 9456 19796 9462 19848
rect 9582 19796 9588 19848
rect 9640 19796 9646 19848
rect 9677 19839 9735 19845
rect 9677 19805 9689 19839
rect 9723 19805 9735 19839
rect 9677 19799 9735 19805
rect 7064 19740 7972 19768
rect 8021 19771 8079 19777
rect 7064 19728 7070 19740
rect 8021 19737 8033 19771
rect 8067 19737 8079 19771
rect 8021 19731 8079 19737
rect 5224 19672 5488 19700
rect 5224 19660 5230 19672
rect 6822 19660 6828 19712
rect 6880 19700 6886 19712
rect 8036 19700 8064 19731
rect 8110 19728 8116 19780
rect 8168 19728 8174 19780
rect 8496 19700 8524 19796
rect 8573 19771 8631 19777
rect 8573 19737 8585 19771
rect 8619 19768 8631 19771
rect 8938 19768 8944 19780
rect 8619 19740 8944 19768
rect 8619 19737 8631 19740
rect 8573 19731 8631 19737
rect 8938 19728 8944 19740
rect 8996 19728 9002 19780
rect 9309 19771 9367 19777
rect 9309 19737 9321 19771
rect 9355 19768 9367 19771
rect 9600 19768 9628 19796
rect 9355 19740 9628 19768
rect 9355 19737 9367 19740
rect 9309 19731 9367 19737
rect 6880 19672 8524 19700
rect 8665 19703 8723 19709
rect 6880 19660 6886 19672
rect 8665 19669 8677 19703
rect 8711 19700 8723 19703
rect 9490 19700 9496 19712
rect 8711 19672 9496 19700
rect 8711 19669 8723 19672
rect 8665 19663 8723 19669
rect 9490 19660 9496 19672
rect 9548 19660 9554 19712
rect 9585 19703 9643 19709
rect 9585 19669 9597 19703
rect 9631 19700 9643 19703
rect 9692 19700 9720 19799
rect 9631 19672 9720 19700
rect 9876 19700 9904 19876
rect 10410 19864 10416 19916
rect 10468 19864 10474 19916
rect 9950 19796 9956 19848
rect 10008 19796 10014 19848
rect 10612 19845 10640 19944
rect 11054 19932 11060 19944
rect 11112 19932 11118 19984
rect 11624 19913 11652 20012
rect 13078 20000 13084 20012
rect 13136 20000 13142 20052
rect 13354 20000 13360 20052
rect 13412 20040 13418 20052
rect 17218 20049 17224 20052
rect 13541 20043 13599 20049
rect 13541 20040 13553 20043
rect 13412 20012 13553 20040
rect 13412 20000 13418 20012
rect 13541 20009 13553 20012
rect 13587 20009 13599 20043
rect 13541 20003 13599 20009
rect 17208 20043 17224 20049
rect 17208 20009 17220 20043
rect 17208 20003 17224 20009
rect 17218 20000 17224 20003
rect 17276 20000 17282 20052
rect 17310 20000 17316 20052
rect 17368 20040 17374 20052
rect 21450 20040 21456 20052
rect 17368 20012 18276 20040
rect 17368 20000 17374 20012
rect 14093 19975 14151 19981
rect 14093 19941 14105 19975
rect 14139 19941 14151 19975
rect 14093 19935 14151 19941
rect 11609 19907 11667 19913
rect 11609 19904 11621 19907
rect 10796 19876 11621 19904
rect 10796 19848 10824 19876
rect 11609 19873 11621 19876
rect 11655 19873 11667 19907
rect 11609 19867 11667 19873
rect 11885 19907 11943 19913
rect 11885 19873 11897 19907
rect 11931 19904 11943 19907
rect 12526 19904 12532 19916
rect 11931 19876 12532 19904
rect 11931 19873 11943 19876
rect 11885 19867 11943 19873
rect 12526 19864 12532 19876
rect 12584 19864 12590 19916
rect 10597 19839 10655 19845
rect 10597 19805 10609 19839
rect 10643 19805 10655 19839
rect 10597 19799 10655 19805
rect 10778 19796 10784 19848
rect 10836 19796 10842 19848
rect 10965 19839 11023 19845
rect 10965 19805 10977 19839
rect 11011 19805 11023 19839
rect 10965 19799 11023 19805
rect 9968 19768 9996 19796
rect 10980 19768 11008 19799
rect 11514 19796 11520 19848
rect 11572 19796 11578 19848
rect 13725 19839 13783 19845
rect 13725 19805 13737 19839
rect 13771 19836 13783 19839
rect 14108 19836 14136 19935
rect 14734 19864 14740 19916
rect 14792 19864 14798 19916
rect 14826 19864 14832 19916
rect 14884 19864 14890 19916
rect 16945 19907 17003 19913
rect 16945 19873 16957 19907
rect 16991 19904 17003 19907
rect 17862 19904 17868 19916
rect 16991 19876 17868 19904
rect 16991 19873 17003 19876
rect 16945 19867 17003 19873
rect 17862 19864 17868 19876
rect 17920 19864 17926 19916
rect 18248 19904 18276 20012
rect 19812 20012 21456 20040
rect 19058 19932 19064 19984
rect 19116 19972 19122 19984
rect 19702 19972 19708 19984
rect 19116 19944 19708 19972
rect 19116 19932 19122 19944
rect 19702 19932 19708 19944
rect 19760 19932 19766 19984
rect 19812 19981 19840 20012
rect 21450 20000 21456 20012
rect 21508 20000 21514 20052
rect 22186 20000 22192 20052
rect 22244 20040 22250 20052
rect 23753 20043 23811 20049
rect 23753 20040 23765 20043
rect 22244 20012 23765 20040
rect 22244 20000 22250 20012
rect 23753 20009 23765 20012
rect 23799 20009 23811 20043
rect 23753 20003 23811 20009
rect 19797 19975 19855 19981
rect 19797 19941 19809 19975
rect 19843 19941 19855 19975
rect 23768 19972 23796 20003
rect 24670 20000 24676 20052
rect 24728 20040 24734 20052
rect 25593 20043 25651 20049
rect 25593 20040 25605 20043
rect 24728 20012 25605 20040
rect 24728 20000 24734 20012
rect 25593 20009 25605 20012
rect 25639 20009 25651 20043
rect 25593 20003 25651 20009
rect 27709 20043 27767 20049
rect 27709 20009 27721 20043
rect 27755 20009 27767 20043
rect 27709 20003 27767 20009
rect 27614 19972 27620 19984
rect 19797 19935 19855 19941
rect 20180 19944 20760 19972
rect 23768 19944 27620 19972
rect 20180 19916 20208 19944
rect 18969 19907 19027 19913
rect 18969 19904 18981 19907
rect 18248 19876 18981 19904
rect 18969 19873 18981 19876
rect 19015 19873 19027 19907
rect 18969 19867 19027 19873
rect 19334 19864 19340 19916
rect 19392 19904 19398 19916
rect 20073 19907 20131 19913
rect 20073 19904 20085 19907
rect 19392 19876 20085 19904
rect 19392 19864 19398 19876
rect 20073 19873 20085 19876
rect 20119 19873 20131 19907
rect 20073 19867 20131 19873
rect 20162 19864 20168 19916
rect 20220 19864 20226 19916
rect 20257 19907 20315 19913
rect 20257 19873 20269 19907
rect 20303 19904 20315 19907
rect 20622 19904 20628 19916
rect 20303 19876 20628 19904
rect 20303 19873 20315 19876
rect 20257 19867 20315 19873
rect 20622 19864 20628 19876
rect 20680 19864 20686 19916
rect 20732 19913 20760 19944
rect 27614 19932 27620 19944
rect 27672 19972 27678 19984
rect 27724 19972 27752 20003
rect 28166 20000 28172 20052
rect 28224 20040 28230 20052
rect 28902 20040 28908 20052
rect 28224 20012 28908 20040
rect 28224 20000 28230 20012
rect 28902 20000 28908 20012
rect 28960 20000 28966 20052
rect 30101 20043 30159 20049
rect 30101 20009 30113 20043
rect 30147 20040 30159 20043
rect 30650 20040 30656 20052
rect 30147 20012 30656 20040
rect 30147 20009 30159 20012
rect 30101 20003 30159 20009
rect 30650 20000 30656 20012
rect 30708 20000 30714 20052
rect 31018 20000 31024 20052
rect 31076 20000 31082 20052
rect 31297 20043 31355 20049
rect 31297 20009 31309 20043
rect 31343 20040 31355 20043
rect 34054 20040 34060 20052
rect 31343 20012 34060 20040
rect 31343 20009 31355 20012
rect 31297 20003 31355 20009
rect 34054 20000 34060 20012
rect 34112 20000 34118 20052
rect 34330 20000 34336 20052
rect 34388 20000 34394 20052
rect 34606 20000 34612 20052
rect 34664 20000 34670 20052
rect 28994 19972 29000 19984
rect 27672 19944 27752 19972
rect 28920 19944 29000 19972
rect 27672 19932 27678 19944
rect 20717 19907 20775 19913
rect 20717 19873 20729 19907
rect 20763 19873 20775 19907
rect 20717 19867 20775 19873
rect 20806 19864 20812 19916
rect 20864 19904 20870 19916
rect 24762 19904 24768 19916
rect 20864 19876 24768 19904
rect 20864 19864 20870 19876
rect 24762 19864 24768 19876
rect 24820 19864 24826 19916
rect 25774 19904 25780 19916
rect 24964 19876 25780 19904
rect 13771 19808 14136 19836
rect 14553 19839 14611 19845
rect 13771 19805 13783 19808
rect 13725 19799 13783 19805
rect 14553 19805 14565 19839
rect 14599 19836 14611 19839
rect 14844 19836 14872 19864
rect 14599 19808 14872 19836
rect 14599 19805 14611 19808
rect 14553 19799 14611 19805
rect 15194 19796 15200 19848
rect 15252 19796 15258 19848
rect 15289 19839 15347 19845
rect 15289 19805 15301 19839
rect 15335 19836 15347 19839
rect 16022 19836 16028 19848
rect 15335 19808 16028 19836
rect 15335 19805 15347 19808
rect 15289 19799 15347 19805
rect 16022 19796 16028 19808
rect 16080 19796 16086 19848
rect 19610 19796 19616 19848
rect 19668 19796 19674 19848
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19805 19947 19839
rect 19889 19799 19947 19805
rect 20349 19839 20407 19845
rect 20349 19805 20361 19839
rect 20395 19836 20407 19839
rect 20990 19836 20996 19848
rect 20395 19808 20996 19836
rect 20395 19805 20407 19808
rect 20349 19799 20407 19805
rect 13906 19768 13912 19780
rect 9968 19740 11008 19768
rect 13110 19740 13912 19768
rect 13906 19728 13912 19740
rect 13964 19728 13970 19780
rect 15212 19768 15240 19796
rect 15212 19740 15792 19768
rect 15764 19712 15792 19740
rect 16942 19728 16948 19780
rect 17000 19768 17006 19780
rect 19904 19768 19932 19799
rect 20990 19796 20996 19808
rect 21048 19796 21054 19848
rect 22278 19796 22284 19848
rect 22336 19836 22342 19848
rect 23569 19839 23627 19845
rect 23569 19836 23581 19839
rect 22336 19808 23581 19836
rect 22336 19796 22342 19808
rect 23569 19805 23581 19808
rect 23615 19805 23627 19839
rect 23569 19799 23627 19805
rect 17000 19740 17710 19768
rect 19306 19740 19932 19768
rect 23584 19768 23612 19799
rect 23842 19796 23848 19848
rect 23900 19796 23906 19848
rect 24026 19796 24032 19848
rect 24084 19796 24090 19848
rect 24964 19845 24992 19876
rect 25774 19864 25780 19876
rect 25832 19864 25838 19916
rect 27356 19876 28396 19904
rect 25130 19845 25136 19848
rect 24949 19839 25007 19845
rect 24949 19805 24961 19839
rect 24995 19805 25007 19839
rect 24949 19799 25007 19805
rect 25097 19839 25136 19845
rect 25097 19805 25109 19839
rect 25097 19799 25136 19805
rect 25130 19796 25136 19799
rect 25188 19796 25194 19848
rect 25455 19839 25513 19845
rect 25455 19805 25467 19839
rect 25501 19836 25513 19839
rect 25590 19836 25596 19848
rect 25501 19808 25596 19836
rect 25501 19805 25513 19808
rect 25455 19799 25513 19805
rect 25590 19796 25596 19808
rect 25648 19836 25654 19848
rect 25866 19836 25872 19848
rect 25648 19808 25872 19836
rect 25648 19796 25654 19808
rect 25866 19796 25872 19808
rect 25924 19796 25930 19848
rect 23934 19768 23940 19780
rect 23584 19740 23940 19768
rect 17000 19728 17006 19740
rect 11790 19700 11796 19712
rect 9876 19672 11796 19700
rect 9631 19669 9643 19672
rect 9585 19663 9643 19669
rect 11790 19660 11796 19672
rect 11848 19660 11854 19712
rect 13354 19660 13360 19712
rect 13412 19660 13418 19712
rect 14366 19660 14372 19712
rect 14424 19700 14430 19712
rect 14461 19703 14519 19709
rect 14461 19700 14473 19703
rect 14424 19672 14473 19700
rect 14424 19660 14430 19672
rect 14461 19669 14473 19672
rect 14507 19669 14519 19703
rect 14461 19663 14519 19669
rect 14550 19660 14556 19712
rect 14608 19700 14614 19712
rect 15473 19703 15531 19709
rect 15473 19700 15485 19703
rect 14608 19672 15485 19700
rect 14608 19660 14614 19672
rect 15473 19669 15485 19672
rect 15519 19669 15531 19703
rect 15473 19663 15531 19669
rect 15746 19660 15752 19712
rect 15804 19660 15810 19712
rect 17604 19700 17632 19740
rect 17954 19700 17960 19712
rect 17604 19672 17960 19700
rect 17954 19660 17960 19672
rect 18012 19660 18018 19712
rect 18138 19660 18144 19712
rect 18196 19700 18202 19712
rect 19306 19700 19334 19740
rect 23934 19728 23940 19740
rect 23992 19728 23998 19780
rect 24044 19768 24072 19796
rect 25225 19771 25283 19777
rect 25225 19768 25237 19771
rect 24044 19740 25237 19768
rect 25225 19737 25237 19740
rect 25271 19737 25283 19771
rect 25225 19731 25283 19737
rect 25317 19771 25375 19777
rect 25317 19737 25329 19771
rect 25363 19737 25375 19771
rect 27356 19768 27384 19876
rect 28368 19845 28396 19876
rect 27433 19839 27491 19845
rect 27433 19805 27445 19839
rect 27479 19836 27491 19839
rect 28353 19839 28411 19845
rect 27479 19808 27568 19836
rect 27479 19805 27491 19808
rect 27433 19799 27491 19805
rect 27540 19780 27568 19808
rect 28353 19805 28365 19839
rect 28399 19805 28411 19839
rect 28353 19799 28411 19805
rect 27356 19740 27476 19768
rect 25317 19731 25375 19737
rect 18196 19672 19334 19700
rect 18196 19660 18202 19672
rect 19426 19660 19432 19712
rect 19484 19660 19490 19712
rect 20438 19660 20444 19712
rect 20496 19660 20502 19712
rect 20530 19660 20536 19712
rect 20588 19700 20594 19712
rect 20625 19703 20683 19709
rect 20625 19700 20637 19703
rect 20588 19672 20637 19700
rect 20588 19660 20594 19672
rect 20625 19669 20637 19672
rect 20671 19669 20683 19703
rect 20625 19663 20683 19669
rect 20714 19660 20720 19712
rect 20772 19700 20778 19712
rect 23014 19700 23020 19712
rect 20772 19672 23020 19700
rect 20772 19660 20778 19672
rect 23014 19660 23020 19672
rect 23072 19660 23078 19712
rect 23382 19660 23388 19712
rect 23440 19660 23446 19712
rect 25332 19700 25360 19731
rect 27448 19712 27476 19740
rect 27522 19728 27528 19780
rect 27580 19728 27586 19780
rect 27617 19771 27675 19777
rect 27617 19737 27629 19771
rect 27663 19737 27675 19771
rect 28368 19768 28396 19799
rect 28442 19796 28448 19848
rect 28500 19836 28506 19848
rect 28537 19839 28595 19845
rect 28537 19836 28549 19839
rect 28500 19808 28549 19836
rect 28500 19796 28506 19808
rect 28537 19805 28549 19808
rect 28583 19805 28595 19839
rect 28537 19799 28595 19805
rect 28629 19839 28687 19845
rect 28629 19805 28641 19839
rect 28675 19836 28687 19839
rect 28810 19836 28816 19848
rect 28675 19808 28816 19836
rect 28675 19805 28687 19808
rect 28629 19799 28687 19805
rect 28810 19796 28816 19808
rect 28868 19796 28874 19848
rect 28920 19836 28948 19944
rect 28994 19932 29000 19944
rect 29052 19932 29058 19984
rect 29288 19944 29500 19972
rect 29288 19904 29316 19944
rect 29196 19876 29316 19904
rect 29196 19845 29224 19876
rect 28977 19839 29035 19845
rect 28977 19836 28989 19839
rect 28920 19808 28989 19836
rect 28977 19805 28989 19808
rect 29023 19805 29035 19839
rect 28977 19799 29035 19805
rect 29089 19839 29147 19845
rect 29089 19805 29101 19839
rect 29135 19805 29147 19839
rect 29089 19799 29147 19805
rect 29181 19839 29239 19845
rect 29181 19805 29193 19839
rect 29227 19805 29239 19839
rect 29181 19799 29239 19805
rect 29104 19768 29132 19799
rect 29362 19796 29368 19848
rect 29420 19845 29426 19848
rect 29420 19839 29435 19845
rect 29423 19805 29435 19839
rect 29420 19799 29435 19805
rect 29420 19796 29426 19799
rect 29270 19768 29276 19780
rect 28368 19740 28856 19768
rect 29104 19740 29276 19768
rect 27617 19731 27675 19737
rect 25406 19700 25412 19712
rect 25332 19672 25412 19700
rect 25406 19660 25412 19672
rect 25464 19660 25470 19712
rect 27430 19660 27436 19712
rect 27488 19660 27494 19712
rect 27632 19700 27660 19731
rect 27706 19700 27712 19712
rect 27632 19672 27712 19700
rect 27706 19660 27712 19672
rect 27764 19660 27770 19712
rect 28350 19660 28356 19712
rect 28408 19700 28414 19712
rect 28721 19703 28779 19709
rect 28721 19700 28733 19703
rect 28408 19672 28733 19700
rect 28408 19660 28414 19672
rect 28721 19669 28733 19672
rect 28767 19669 28779 19703
rect 28828 19700 28856 19740
rect 29270 19728 29276 19740
rect 29328 19728 29334 19780
rect 29472 19768 29500 19944
rect 29546 19932 29552 19984
rect 29604 19932 29610 19984
rect 30006 19932 30012 19984
rect 30064 19972 30070 19984
rect 31036 19972 31064 20000
rect 33778 19972 33784 19984
rect 30064 19944 31064 19972
rect 31312 19944 33784 19972
rect 30064 19932 30070 19944
rect 31312 19916 31340 19944
rect 33778 19932 33784 19944
rect 33836 19932 33842 19984
rect 34348 19972 34376 20000
rect 34072 19944 34376 19972
rect 34072 19916 34100 19944
rect 30374 19904 30380 19916
rect 30208 19876 30380 19904
rect 29822 19796 29828 19848
rect 29880 19796 29886 19848
rect 29914 19796 29920 19848
rect 29972 19796 29978 19848
rect 30009 19839 30067 19845
rect 30009 19805 30021 19839
rect 30055 19836 30067 19839
rect 30208 19836 30236 19876
rect 30374 19864 30380 19876
rect 30432 19864 30438 19916
rect 31294 19864 31300 19916
rect 31352 19864 31358 19916
rect 31386 19864 31392 19916
rect 31444 19904 31450 19916
rect 31444 19876 32812 19904
rect 31444 19864 31450 19876
rect 30055 19808 30236 19836
rect 30285 19839 30343 19845
rect 30055 19805 30067 19808
rect 30009 19799 30067 19805
rect 30285 19805 30297 19839
rect 30331 19836 30343 19839
rect 30834 19836 30840 19848
rect 30331 19808 30840 19836
rect 30331 19805 30343 19808
rect 30285 19799 30343 19805
rect 30834 19796 30840 19808
rect 30892 19796 30898 19848
rect 31478 19796 31484 19848
rect 31536 19796 31542 19848
rect 31570 19768 31576 19780
rect 29472 19740 31576 19768
rect 31570 19728 31576 19740
rect 31628 19728 31634 19780
rect 31705 19777 31733 19876
rect 32784 19848 32812 19876
rect 33410 19864 33416 19916
rect 33468 19864 33474 19916
rect 34054 19864 34060 19916
rect 34112 19864 34118 19916
rect 34146 19864 34152 19916
rect 34204 19864 34210 19916
rect 34624 19904 34652 20000
rect 34624 19876 35020 19904
rect 31941 19839 31999 19845
rect 31941 19805 31953 19839
rect 31987 19836 31999 19839
rect 32030 19836 32036 19848
rect 31987 19808 32036 19836
rect 31987 19805 31999 19808
rect 31941 19799 31999 19805
rect 32030 19796 32036 19808
rect 32088 19836 32094 19848
rect 32214 19836 32220 19848
rect 32088 19808 32220 19836
rect 32088 19796 32094 19808
rect 32214 19796 32220 19808
rect 32272 19796 32278 19848
rect 32766 19796 32772 19848
rect 32824 19796 32830 19848
rect 33321 19839 33379 19845
rect 33321 19805 33333 19839
rect 33367 19836 33379 19839
rect 33428 19836 33456 19864
rect 33367 19808 33456 19836
rect 33367 19805 33379 19808
rect 33321 19799 33379 19805
rect 31665 19771 31733 19777
rect 31665 19737 31677 19771
rect 31711 19740 31733 19771
rect 31803 19771 31861 19777
rect 31711 19737 31723 19740
rect 31665 19731 31723 19737
rect 31803 19737 31815 19771
rect 31849 19768 31861 19771
rect 33336 19768 33364 19799
rect 33778 19796 33784 19848
rect 33836 19796 33842 19848
rect 33870 19796 33876 19848
rect 33928 19836 33934 19848
rect 34241 19839 34299 19845
rect 34241 19836 34253 19839
rect 33928 19808 34253 19836
rect 33928 19796 33934 19808
rect 34241 19805 34253 19808
rect 34287 19805 34299 19839
rect 34241 19799 34299 19805
rect 34330 19796 34336 19848
rect 34388 19796 34394 19848
rect 34514 19796 34520 19848
rect 34572 19836 34578 19848
rect 34992 19845 35020 19876
rect 34701 19839 34759 19845
rect 34701 19836 34713 19839
rect 34572 19808 34713 19836
rect 34572 19796 34578 19808
rect 34701 19805 34713 19808
rect 34747 19805 34759 19839
rect 34701 19799 34759 19805
rect 34977 19839 35035 19845
rect 34977 19805 34989 19839
rect 35023 19805 35035 19839
rect 34977 19799 35035 19805
rect 35069 19839 35127 19845
rect 35069 19805 35081 19839
rect 35115 19836 35127 19839
rect 35434 19836 35440 19848
rect 35115 19808 35440 19836
rect 35115 19805 35127 19808
rect 35069 19799 35127 19805
rect 35434 19796 35440 19808
rect 35492 19796 35498 19848
rect 35894 19796 35900 19848
rect 35952 19836 35958 19848
rect 40494 19836 40500 19848
rect 35952 19808 40500 19836
rect 35952 19796 35958 19808
rect 40494 19796 40500 19808
rect 40552 19796 40558 19848
rect 31849 19740 33364 19768
rect 31849 19737 31861 19740
rect 31803 19731 31861 19737
rect 32232 19712 32260 19740
rect 33410 19728 33416 19780
rect 33468 19728 33474 19780
rect 33505 19771 33563 19777
rect 33505 19737 33517 19771
rect 33551 19737 33563 19771
rect 33623 19771 33681 19777
rect 33623 19768 33635 19771
rect 33505 19731 33563 19737
rect 33612 19737 33635 19768
rect 33669 19737 33681 19771
rect 34054 19768 34060 19780
rect 33612 19731 33681 19737
rect 33796 19740 34060 19768
rect 29822 19700 29828 19712
rect 28828 19672 29828 19700
rect 28721 19663 28779 19669
rect 29822 19660 29828 19672
rect 29880 19660 29886 19712
rect 30006 19660 30012 19712
rect 30064 19700 30070 19712
rect 30650 19700 30656 19712
rect 30064 19672 30656 19700
rect 30064 19660 30070 19672
rect 30650 19660 30656 19672
rect 30708 19660 30714 19712
rect 32214 19660 32220 19712
rect 32272 19660 32278 19712
rect 33134 19660 33140 19712
rect 33192 19660 33198 19712
rect 33318 19660 33324 19712
rect 33376 19700 33382 19712
rect 33520 19700 33548 19731
rect 33376 19672 33548 19700
rect 33612 19700 33640 19731
rect 33796 19700 33824 19740
rect 34054 19728 34060 19740
rect 34112 19728 34118 19780
rect 34146 19728 34152 19780
rect 34204 19768 34210 19780
rect 34885 19771 34943 19777
rect 34885 19768 34897 19771
rect 34204 19740 34897 19768
rect 34204 19728 34210 19740
rect 34885 19737 34897 19740
rect 34931 19737 34943 19771
rect 38838 19768 38844 19780
rect 34885 19731 34943 19737
rect 35176 19740 38844 19768
rect 33612 19672 33824 19700
rect 33873 19703 33931 19709
rect 33376 19660 33382 19672
rect 33873 19669 33885 19703
rect 33919 19700 33931 19703
rect 35176 19700 35204 19740
rect 38838 19728 38844 19740
rect 38896 19768 38902 19780
rect 39482 19768 39488 19780
rect 38896 19740 39488 19768
rect 38896 19728 38902 19740
rect 39482 19728 39488 19740
rect 39540 19728 39546 19780
rect 33919 19672 35204 19700
rect 35253 19703 35311 19709
rect 33919 19669 33931 19672
rect 33873 19663 33931 19669
rect 35253 19669 35265 19703
rect 35299 19700 35311 19703
rect 37918 19700 37924 19712
rect 35299 19672 37924 19700
rect 35299 19669 35311 19672
rect 35253 19663 35311 19669
rect 37918 19660 37924 19672
rect 37976 19660 37982 19712
rect 1104 19610 41400 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 41400 19610
rect 1104 19536 41400 19558
rect 1670 19456 1676 19508
rect 1728 19496 1734 19508
rect 1857 19499 1915 19505
rect 1857 19496 1869 19499
rect 1728 19468 1869 19496
rect 1728 19456 1734 19468
rect 1857 19465 1869 19468
rect 1903 19465 1915 19499
rect 1857 19459 1915 19465
rect 2225 19499 2283 19505
rect 2225 19465 2237 19499
rect 2271 19465 2283 19499
rect 2225 19459 2283 19465
rect 2041 19363 2099 19369
rect 2041 19329 2053 19363
rect 2087 19360 2099 19363
rect 2240 19360 2268 19459
rect 2590 19456 2596 19508
rect 2648 19456 2654 19508
rect 3418 19496 3424 19508
rect 3068 19468 3424 19496
rect 2087 19332 2268 19360
rect 2685 19363 2743 19369
rect 2087 19329 2099 19332
rect 2041 19323 2099 19329
rect 2685 19329 2697 19363
rect 2731 19360 2743 19363
rect 2774 19360 2780 19372
rect 2731 19332 2780 19360
rect 2731 19329 2743 19332
rect 2685 19323 2743 19329
rect 2774 19320 2780 19332
rect 2832 19320 2838 19372
rect 3068 19369 3096 19468
rect 3418 19456 3424 19468
rect 3476 19496 3482 19508
rect 4614 19496 4620 19508
rect 3476 19468 4620 19496
rect 3476 19456 3482 19468
rect 4614 19456 4620 19468
rect 4672 19456 4678 19508
rect 4801 19499 4859 19505
rect 4801 19465 4813 19499
rect 4847 19496 4859 19499
rect 5074 19496 5080 19508
rect 4847 19468 5080 19496
rect 4847 19465 4859 19468
rect 4801 19459 4859 19465
rect 5074 19456 5080 19468
rect 5132 19456 5138 19508
rect 5534 19456 5540 19508
rect 5592 19456 5598 19508
rect 7006 19456 7012 19508
rect 7064 19456 7070 19508
rect 8570 19456 8576 19508
rect 8628 19456 8634 19508
rect 8754 19456 8760 19508
rect 8812 19496 8818 19508
rect 9398 19496 9404 19508
rect 8812 19468 9404 19496
rect 8812 19456 8818 19468
rect 9398 19456 9404 19468
rect 9456 19496 9462 19508
rect 9861 19499 9919 19505
rect 9456 19468 9812 19496
rect 9456 19456 9462 19468
rect 3329 19431 3387 19437
rect 3329 19397 3341 19431
rect 3375 19428 3387 19431
rect 3602 19428 3608 19440
rect 3375 19400 3608 19428
rect 3375 19397 3387 19400
rect 3329 19391 3387 19397
rect 3602 19388 3608 19400
rect 3660 19388 3666 19440
rect 7024 19428 7052 19456
rect 4908 19400 5672 19428
rect 3053 19363 3111 19369
rect 3053 19329 3065 19363
rect 3099 19329 3111 19363
rect 3053 19323 3111 19329
rect 4430 19320 4436 19372
rect 4488 19360 4494 19372
rect 4706 19360 4712 19372
rect 4488 19332 4712 19360
rect 4488 19320 4494 19332
rect 4706 19320 4712 19332
rect 4764 19320 4770 19372
rect 4908 19369 4936 19400
rect 5644 19372 5672 19400
rect 5736 19400 7052 19428
rect 7285 19431 7343 19437
rect 5736 19372 5764 19400
rect 7285 19397 7297 19431
rect 7331 19428 7343 19431
rect 8294 19428 8300 19440
rect 7331 19400 8300 19428
rect 7331 19397 7343 19400
rect 7285 19391 7343 19397
rect 8294 19388 8300 19400
rect 8352 19388 8358 19440
rect 8389 19431 8447 19437
rect 8389 19397 8401 19431
rect 8435 19428 8447 19431
rect 8588 19428 8616 19456
rect 8435 19400 8616 19428
rect 8435 19397 8447 19400
rect 8389 19391 8447 19397
rect 4893 19363 4951 19369
rect 4893 19329 4905 19363
rect 4939 19329 4951 19363
rect 4893 19323 4951 19329
rect 4986 19363 5044 19369
rect 4986 19329 4998 19363
rect 5032 19329 5044 19363
rect 4986 19323 5044 19329
rect 2869 19295 2927 19301
rect 2869 19261 2881 19295
rect 2915 19261 2927 19295
rect 2869 19255 2927 19261
rect 2884 19168 2912 19255
rect 4062 19252 4068 19304
rect 4120 19292 4126 19304
rect 5000 19292 5028 19323
rect 5166 19320 5172 19372
rect 5224 19320 5230 19372
rect 5261 19363 5319 19369
rect 5261 19329 5273 19363
rect 5307 19329 5319 19363
rect 5261 19323 5319 19329
rect 5399 19363 5457 19369
rect 5399 19329 5411 19363
rect 5445 19360 5457 19363
rect 5445 19332 5580 19360
rect 5445 19329 5457 19332
rect 5399 19323 5457 19329
rect 4120 19264 5028 19292
rect 4120 19252 4126 19264
rect 2866 19116 2872 19168
rect 2924 19116 2930 19168
rect 3878 19116 3884 19168
rect 3936 19156 3942 19168
rect 5276 19156 5304 19323
rect 5552 19292 5580 19332
rect 5626 19320 5632 19372
rect 5684 19320 5690 19372
rect 5718 19320 5724 19372
rect 5776 19320 5782 19372
rect 7377 19363 7435 19369
rect 7377 19329 7389 19363
rect 7423 19360 7435 19363
rect 7558 19360 7564 19372
rect 7423 19332 7564 19360
rect 7423 19329 7435 19332
rect 7377 19323 7435 19329
rect 7558 19320 7564 19332
rect 7616 19320 7622 19372
rect 8113 19363 8171 19369
rect 8113 19329 8125 19363
rect 8159 19329 8171 19363
rect 8113 19323 8171 19329
rect 5736 19292 5764 19320
rect 5552 19264 5764 19292
rect 7469 19295 7527 19301
rect 7469 19261 7481 19295
rect 7515 19261 7527 19295
rect 7469 19255 7527 19261
rect 5626 19184 5632 19236
rect 5684 19224 5690 19236
rect 5810 19224 5816 19236
rect 5684 19196 5816 19224
rect 5684 19184 5690 19196
rect 5810 19184 5816 19196
rect 5868 19224 5874 19236
rect 6822 19224 6828 19236
rect 5868 19196 6828 19224
rect 5868 19184 5874 19196
rect 6822 19184 6828 19196
rect 6880 19184 6886 19236
rect 3936 19128 5304 19156
rect 3936 19116 3942 19128
rect 6914 19116 6920 19168
rect 6972 19116 6978 19168
rect 7484 19156 7512 19255
rect 8018 19184 8024 19236
rect 8076 19224 8082 19236
rect 8128 19224 8156 19323
rect 9490 19320 9496 19372
rect 9548 19320 9554 19372
rect 9784 19360 9812 19468
rect 9861 19465 9873 19499
rect 9907 19496 9919 19499
rect 9950 19496 9956 19508
rect 9907 19468 9956 19496
rect 9907 19465 9919 19468
rect 9861 19459 9919 19465
rect 9950 19456 9956 19468
rect 10008 19456 10014 19508
rect 12161 19499 12219 19505
rect 12161 19465 12173 19499
rect 12207 19496 12219 19499
rect 12710 19496 12716 19508
rect 12207 19468 12716 19496
rect 12207 19465 12219 19468
rect 12161 19459 12219 19465
rect 12710 19456 12716 19468
rect 12768 19456 12774 19508
rect 13722 19456 13728 19508
rect 13780 19496 13786 19508
rect 16850 19496 16856 19508
rect 13780 19468 16856 19496
rect 13780 19456 13786 19468
rect 10045 19431 10103 19437
rect 10045 19397 10057 19431
rect 10091 19428 10103 19431
rect 10134 19428 10140 19440
rect 10091 19400 10140 19428
rect 10091 19397 10103 19400
rect 10045 19391 10103 19397
rect 10134 19388 10140 19400
rect 10192 19388 10198 19440
rect 11054 19388 11060 19440
rect 11112 19428 11118 19440
rect 12342 19428 12348 19440
rect 11112 19400 12348 19428
rect 11112 19388 11118 19400
rect 12342 19388 12348 19400
rect 12400 19428 12406 19440
rect 14550 19428 14556 19440
rect 12400 19400 14556 19428
rect 12400 19388 12406 19400
rect 14550 19388 14556 19400
rect 14608 19388 14614 19440
rect 9784 19332 12434 19360
rect 8938 19252 8944 19304
rect 8996 19292 9002 19304
rect 9858 19292 9864 19304
rect 8996 19264 9864 19292
rect 8996 19252 9002 19264
rect 9858 19252 9864 19264
rect 9916 19252 9922 19304
rect 9950 19252 9956 19304
rect 10008 19292 10014 19304
rect 10778 19292 10784 19304
rect 10008 19264 10784 19292
rect 10008 19252 10014 19264
rect 10778 19252 10784 19264
rect 10836 19252 10842 19304
rect 8076 19196 8156 19224
rect 12406 19224 12434 19332
rect 12526 19320 12532 19372
rect 12584 19320 12590 19372
rect 12621 19363 12679 19369
rect 12621 19329 12633 19363
rect 12667 19360 12679 19363
rect 13354 19360 13360 19372
rect 12667 19332 13360 19360
rect 12667 19329 12679 19332
rect 12621 19323 12679 19329
rect 13354 19320 13360 19332
rect 13412 19320 13418 19372
rect 14734 19360 14740 19372
rect 13832 19332 14740 19360
rect 12710 19252 12716 19304
rect 12768 19292 12774 19304
rect 12805 19295 12863 19301
rect 12805 19292 12817 19295
rect 12768 19264 12817 19292
rect 12768 19252 12774 19264
rect 12805 19261 12817 19264
rect 12851 19292 12863 19295
rect 13832 19292 13860 19332
rect 14734 19320 14740 19332
rect 14792 19320 14798 19372
rect 15028 19360 15056 19468
rect 16850 19456 16856 19468
rect 16908 19456 16914 19508
rect 16945 19499 17003 19505
rect 16945 19465 16957 19499
rect 16991 19496 17003 19499
rect 17402 19496 17408 19508
rect 16991 19468 17408 19496
rect 16991 19465 17003 19468
rect 16945 19459 17003 19465
rect 17402 19456 17408 19468
rect 17460 19456 17466 19508
rect 17862 19456 17868 19508
rect 17920 19496 17926 19508
rect 24578 19496 24584 19508
rect 17920 19468 24584 19496
rect 17920 19456 17926 19468
rect 24578 19456 24584 19468
rect 24636 19456 24642 19508
rect 25130 19456 25136 19508
rect 25188 19496 25194 19508
rect 25409 19499 25467 19505
rect 25409 19496 25421 19499
rect 25188 19468 25421 19496
rect 25188 19456 25194 19468
rect 25409 19465 25421 19468
rect 25455 19465 25467 19499
rect 25409 19459 25467 19465
rect 25590 19456 25596 19508
rect 25648 19496 25654 19508
rect 27706 19496 27712 19508
rect 25648 19468 27712 19496
rect 25648 19456 25654 19468
rect 16022 19388 16028 19440
rect 16080 19388 16086 19440
rect 16390 19388 16396 19440
rect 16448 19428 16454 19440
rect 16448 19400 17448 19428
rect 16448 19388 16454 19400
rect 15105 19363 15163 19369
rect 15105 19360 15117 19363
rect 15028 19332 15117 19360
rect 15105 19329 15117 19332
rect 15151 19329 15163 19363
rect 15289 19363 15347 19369
rect 15289 19360 15301 19363
rect 15105 19323 15163 19329
rect 15212 19332 15301 19360
rect 12851 19264 13860 19292
rect 12851 19261 12863 19264
rect 12805 19255 12863 19261
rect 14458 19252 14464 19304
rect 14516 19292 14522 19304
rect 15212 19292 15240 19332
rect 15289 19329 15301 19332
rect 15335 19329 15347 19363
rect 15289 19323 15347 19329
rect 15746 19320 15752 19372
rect 15804 19320 15810 19372
rect 16040 19360 16068 19388
rect 16209 19363 16267 19369
rect 16209 19360 16221 19363
rect 16040 19332 16221 19360
rect 16209 19329 16221 19332
rect 16255 19329 16267 19363
rect 16209 19323 16267 19329
rect 17310 19320 17316 19372
rect 17368 19320 17374 19372
rect 17420 19369 17448 19400
rect 17586 19388 17592 19440
rect 17644 19428 17650 19440
rect 18138 19428 18144 19440
rect 17644 19400 18144 19428
rect 17644 19388 17650 19400
rect 18138 19388 18144 19400
rect 18196 19388 18202 19440
rect 18230 19388 18236 19440
rect 18288 19388 18294 19440
rect 20162 19388 20168 19440
rect 20220 19428 20226 19440
rect 20530 19428 20536 19440
rect 20220 19400 20536 19428
rect 20220 19388 20226 19400
rect 20530 19388 20536 19400
rect 20588 19388 20594 19440
rect 21726 19388 21732 19440
rect 21784 19428 21790 19440
rect 21784 19400 22324 19428
rect 21784 19388 21790 19400
rect 17405 19363 17463 19369
rect 17405 19329 17417 19363
rect 17451 19329 17463 19363
rect 17405 19323 17463 19329
rect 18877 19363 18935 19369
rect 18877 19329 18889 19363
rect 18923 19360 18935 19363
rect 20714 19360 20720 19372
rect 18923 19332 20720 19360
rect 18923 19329 18935 19332
rect 18877 19323 18935 19329
rect 20714 19320 20720 19332
rect 20772 19320 20778 19372
rect 22005 19363 22063 19369
rect 22005 19329 22017 19363
rect 22051 19360 22063 19363
rect 22186 19360 22192 19372
rect 22051 19332 22192 19360
rect 22051 19329 22063 19332
rect 22005 19323 22063 19329
rect 22186 19320 22192 19332
rect 22244 19320 22250 19372
rect 22296 19369 22324 19400
rect 22370 19388 22376 19440
rect 22428 19388 22434 19440
rect 24026 19428 24032 19440
rect 23400 19400 24032 19428
rect 22281 19363 22339 19369
rect 22281 19329 22293 19363
rect 22327 19329 22339 19363
rect 22388 19360 22416 19388
rect 22649 19363 22707 19369
rect 22388 19332 22600 19360
rect 22281 19323 22339 19329
rect 14516 19264 15240 19292
rect 17589 19295 17647 19301
rect 14516 19252 14522 19264
rect 17589 19261 17601 19295
rect 17635 19261 17647 19295
rect 17589 19255 17647 19261
rect 18969 19295 19027 19301
rect 18969 19261 18981 19295
rect 19015 19292 19027 19295
rect 19058 19292 19064 19304
rect 19015 19264 19064 19292
rect 19015 19261 19027 19264
rect 18969 19255 19027 19261
rect 12894 19224 12900 19236
rect 12406 19196 12900 19224
rect 8076 19184 8082 19196
rect 12894 19184 12900 19196
rect 12952 19224 12958 19236
rect 13722 19224 13728 19236
rect 12952 19196 13728 19224
rect 12952 19184 12958 19196
rect 13722 19184 13728 19196
rect 13780 19184 13786 19236
rect 14553 19227 14611 19233
rect 14553 19193 14565 19227
rect 14599 19224 14611 19227
rect 14642 19224 14648 19236
rect 14599 19196 14648 19224
rect 14599 19193 14611 19196
rect 14553 19187 14611 19193
rect 14642 19184 14648 19196
rect 14700 19184 14706 19236
rect 14921 19227 14979 19233
rect 14921 19193 14933 19227
rect 14967 19224 14979 19227
rect 15102 19224 15108 19236
rect 14967 19196 15108 19224
rect 14967 19193 14979 19196
rect 14921 19187 14979 19193
rect 15102 19184 15108 19196
rect 15160 19184 15166 19236
rect 17604 19224 17632 19255
rect 19058 19252 19064 19264
rect 19116 19252 19122 19304
rect 19150 19252 19156 19304
rect 19208 19252 19214 19304
rect 19426 19252 19432 19304
rect 19484 19252 19490 19304
rect 21542 19252 21548 19304
rect 21600 19292 21606 19304
rect 21821 19295 21879 19301
rect 21821 19292 21833 19295
rect 21600 19264 21833 19292
rect 21600 19252 21606 19264
rect 21821 19261 21833 19264
rect 21867 19261 21879 19295
rect 21821 19255 21879 19261
rect 22370 19252 22376 19304
rect 22428 19252 22434 19304
rect 22572 19301 22600 19332
rect 22649 19329 22661 19363
rect 22695 19360 22707 19363
rect 23198 19360 23204 19372
rect 22695 19332 23204 19360
rect 22695 19329 22707 19332
rect 22649 19323 22707 19329
rect 23198 19320 23204 19332
rect 23256 19320 23262 19372
rect 23400 19369 23428 19400
rect 24026 19388 24032 19400
rect 24084 19388 24090 19440
rect 24302 19388 24308 19440
rect 24360 19428 24366 19440
rect 24670 19428 24676 19440
rect 24360 19400 24676 19428
rect 24360 19388 24366 19400
rect 24670 19388 24676 19400
rect 24728 19388 24734 19440
rect 25222 19388 25228 19440
rect 25280 19388 25286 19440
rect 25682 19388 25688 19440
rect 25740 19428 25746 19440
rect 25777 19431 25835 19437
rect 25777 19428 25789 19431
rect 25740 19400 25789 19428
rect 25740 19388 25746 19400
rect 25777 19397 25789 19400
rect 25823 19428 25835 19431
rect 25958 19428 25964 19440
rect 25823 19400 25964 19428
rect 25823 19397 25835 19400
rect 25777 19391 25835 19397
rect 25958 19388 25964 19400
rect 26016 19388 26022 19440
rect 27448 19437 27476 19468
rect 27706 19456 27712 19468
rect 27764 19456 27770 19508
rect 27890 19456 27896 19508
rect 27948 19496 27954 19508
rect 29546 19496 29552 19508
rect 27948 19468 29552 19496
rect 27948 19456 27954 19468
rect 28000 19437 28028 19468
rect 29546 19456 29552 19468
rect 29604 19456 29610 19508
rect 29914 19496 29920 19508
rect 29656 19468 29920 19496
rect 27341 19431 27399 19437
rect 27341 19397 27353 19431
rect 27387 19397 27399 19431
rect 27341 19391 27399 19397
rect 27433 19431 27491 19437
rect 27433 19397 27445 19431
rect 27479 19397 27491 19431
rect 27433 19391 27491 19397
rect 27985 19431 28043 19437
rect 27985 19397 27997 19431
rect 28031 19397 28043 19431
rect 27985 19391 28043 19397
rect 23385 19363 23443 19369
rect 23385 19329 23397 19363
rect 23431 19329 23443 19363
rect 23385 19323 23443 19329
rect 23477 19363 23535 19369
rect 23477 19329 23489 19363
rect 23523 19360 23535 19363
rect 23566 19360 23572 19372
rect 23523 19332 23572 19360
rect 23523 19329 23535 19332
rect 23477 19323 23535 19329
rect 23566 19320 23572 19332
rect 23624 19320 23630 19372
rect 23658 19320 23664 19372
rect 23716 19320 23722 19372
rect 23753 19363 23811 19369
rect 23753 19329 23765 19363
rect 23799 19360 23811 19363
rect 23842 19360 23848 19372
rect 23799 19332 23848 19360
rect 23799 19329 23811 19332
rect 23753 19323 23811 19329
rect 23842 19320 23848 19332
rect 23900 19320 23906 19372
rect 24394 19320 24400 19372
rect 24452 19320 24458 19372
rect 25041 19363 25099 19369
rect 24688 19332 24992 19360
rect 22557 19295 22615 19301
rect 22557 19261 22569 19295
rect 22603 19261 22615 19295
rect 22557 19255 22615 19261
rect 24213 19295 24271 19301
rect 24213 19261 24225 19295
rect 24259 19292 24271 19295
rect 24688 19292 24716 19332
rect 24259 19264 24716 19292
rect 24765 19295 24823 19301
rect 24259 19261 24271 19264
rect 24213 19255 24271 19261
rect 24765 19261 24777 19295
rect 24811 19261 24823 19295
rect 24765 19255 24823 19261
rect 19444 19224 19472 19252
rect 17604 19196 19472 19224
rect 20622 19184 20628 19236
rect 20680 19224 20686 19236
rect 20680 19196 24256 19224
rect 20680 19184 20686 19196
rect 9398 19156 9404 19168
rect 7484 19128 9404 19156
rect 9398 19116 9404 19128
rect 9456 19116 9462 19168
rect 12066 19116 12072 19168
rect 12124 19156 12130 19168
rect 15562 19156 15568 19168
rect 12124 19128 15568 19156
rect 12124 19116 12130 19128
rect 15562 19116 15568 19128
rect 15620 19116 15626 19168
rect 16574 19116 16580 19168
rect 16632 19156 16638 19168
rect 17218 19156 17224 19168
rect 16632 19128 17224 19156
rect 16632 19116 16638 19128
rect 17218 19116 17224 19128
rect 17276 19116 17282 19168
rect 18138 19116 18144 19168
rect 18196 19156 18202 19168
rect 18325 19159 18383 19165
rect 18325 19156 18337 19159
rect 18196 19128 18337 19156
rect 18196 19116 18202 19128
rect 18325 19125 18337 19128
rect 18371 19125 18383 19159
rect 18325 19119 18383 19125
rect 19058 19116 19064 19168
rect 19116 19116 19122 19168
rect 21174 19116 21180 19168
rect 21232 19156 21238 19168
rect 22554 19156 22560 19168
rect 21232 19128 22560 19156
rect 21232 19116 21238 19128
rect 22554 19116 22560 19128
rect 22612 19116 22618 19168
rect 23198 19116 23204 19168
rect 23256 19116 23262 19168
rect 24228 19156 24256 19196
rect 24578 19184 24584 19236
rect 24636 19224 24642 19236
rect 24780 19224 24808 19255
rect 24854 19252 24860 19304
rect 24912 19252 24918 19304
rect 24964 19292 24992 19332
rect 25041 19329 25053 19363
rect 25087 19360 25099 19363
rect 25130 19360 25136 19372
rect 25087 19332 25136 19360
rect 25087 19329 25099 19332
rect 25041 19323 25099 19329
rect 25130 19320 25136 19332
rect 25188 19320 25194 19372
rect 25317 19363 25375 19369
rect 25317 19329 25329 19363
rect 25363 19360 25375 19363
rect 25363 19332 25452 19360
rect 25363 19329 25375 19332
rect 25317 19323 25375 19329
rect 25424 19304 25452 19332
rect 25590 19320 25596 19372
rect 25648 19320 25654 19372
rect 25869 19363 25927 19369
rect 25869 19329 25881 19363
rect 25915 19360 25927 19363
rect 25915 19332 26004 19360
rect 25915 19329 25927 19332
rect 25869 19323 25927 19329
rect 25406 19292 25412 19304
rect 24964 19264 25412 19292
rect 25406 19252 25412 19264
rect 25464 19252 25470 19304
rect 25976 19292 26004 19332
rect 26050 19320 26056 19372
rect 26108 19360 26114 19372
rect 26108 19332 26280 19360
rect 26108 19320 26114 19332
rect 26142 19292 26148 19304
rect 25976 19264 26148 19292
rect 26142 19252 26148 19264
rect 26200 19252 26206 19304
rect 26252 19292 26280 19332
rect 26510 19320 26516 19372
rect 26568 19320 26574 19372
rect 26602 19320 26608 19372
rect 26660 19360 26666 19372
rect 27065 19363 27123 19369
rect 27065 19360 27077 19363
rect 26660 19332 27077 19360
rect 26660 19320 26666 19332
rect 27065 19329 27077 19332
rect 27111 19329 27123 19363
rect 27065 19323 27123 19329
rect 27158 19363 27216 19369
rect 27158 19329 27170 19363
rect 27204 19329 27216 19363
rect 27158 19323 27216 19329
rect 26789 19295 26847 19301
rect 26789 19292 26801 19295
rect 26252 19264 26464 19292
rect 26329 19227 26387 19233
rect 26329 19224 26341 19227
rect 24636 19196 24808 19224
rect 24872 19196 26341 19224
rect 24636 19184 24642 19196
rect 24872 19156 24900 19196
rect 26329 19193 26341 19196
rect 26375 19193 26387 19227
rect 26329 19187 26387 19193
rect 24228 19128 24900 19156
rect 24946 19116 24952 19168
rect 25004 19156 25010 19168
rect 25130 19156 25136 19168
rect 25004 19128 25136 19156
rect 25004 19116 25010 19128
rect 25130 19116 25136 19128
rect 25188 19156 25194 19168
rect 25774 19156 25780 19168
rect 25188 19128 25780 19156
rect 25188 19116 25194 19128
rect 25774 19116 25780 19128
rect 25832 19116 25838 19168
rect 26436 19156 26464 19264
rect 26620 19264 26801 19292
rect 26620 19236 26648 19264
rect 26789 19261 26801 19264
rect 26835 19261 26847 19295
rect 26789 19255 26847 19261
rect 26878 19252 26884 19304
rect 26936 19292 26942 19304
rect 27172 19292 27200 19323
rect 27356 19304 27384 19391
rect 28166 19388 28172 19440
rect 28224 19388 28230 19440
rect 29656 19428 29684 19468
rect 29914 19456 29920 19468
rect 29972 19456 29978 19508
rect 30374 19456 30380 19508
rect 30432 19456 30438 19508
rect 31389 19499 31447 19505
rect 31389 19496 31401 19499
rect 30576 19468 31401 19496
rect 30392 19428 30420 19456
rect 28736 19400 29684 19428
rect 29921 19400 30420 19428
rect 27571 19363 27629 19369
rect 27571 19329 27583 19363
rect 27617 19360 27629 19363
rect 27706 19360 27712 19372
rect 27617 19332 27712 19360
rect 27617 19329 27629 19332
rect 27571 19323 27629 19329
rect 27706 19320 27712 19332
rect 27764 19320 27770 19372
rect 27890 19320 27896 19372
rect 27948 19360 27954 19372
rect 28736 19369 28764 19400
rect 28721 19363 28779 19369
rect 27948 19332 28672 19360
rect 27948 19320 27954 19332
rect 26936 19264 27200 19292
rect 26936 19252 26942 19264
rect 27338 19252 27344 19304
rect 27396 19252 27402 19304
rect 28074 19252 28080 19304
rect 28132 19292 28138 19304
rect 28537 19295 28595 19301
rect 28537 19292 28549 19295
rect 28132 19264 28549 19292
rect 28132 19252 28138 19264
rect 28537 19261 28549 19264
rect 28583 19261 28595 19295
rect 28644 19292 28672 19332
rect 28721 19329 28733 19363
rect 28767 19329 28779 19363
rect 28905 19363 28963 19369
rect 28905 19360 28917 19363
rect 28721 19323 28779 19329
rect 28828 19332 28917 19360
rect 28828 19292 28856 19332
rect 28905 19329 28917 19332
rect 28951 19329 28963 19363
rect 28905 19323 28963 19329
rect 29086 19320 29092 19372
rect 29144 19360 29150 19372
rect 29921 19360 29949 19400
rect 30466 19388 30472 19440
rect 30524 19388 30530 19440
rect 30576 19437 30604 19468
rect 31389 19465 31401 19468
rect 31435 19465 31447 19499
rect 31389 19459 31447 19465
rect 33134 19456 33140 19508
rect 33192 19496 33198 19508
rect 39666 19496 39672 19508
rect 33192 19468 39672 19496
rect 33192 19456 33198 19468
rect 39666 19456 39672 19468
rect 39724 19496 39730 19508
rect 40126 19496 40132 19508
rect 39724 19468 40132 19496
rect 39724 19456 39730 19468
rect 40126 19456 40132 19468
rect 40184 19456 40190 19508
rect 30561 19431 30619 19437
rect 30561 19397 30573 19431
rect 30607 19397 30619 19431
rect 33594 19428 33600 19440
rect 30561 19391 30619 19397
rect 31726 19400 33600 19428
rect 29144 19332 29949 19360
rect 30377 19363 30435 19369
rect 29144 19320 29150 19332
rect 30377 19329 30389 19363
rect 30423 19329 30435 19363
rect 30484 19360 30512 19388
rect 30653 19363 30711 19369
rect 30653 19360 30665 19363
rect 30484 19332 30665 19360
rect 30377 19323 30435 19329
rect 30653 19329 30665 19332
rect 30699 19329 30711 19363
rect 30653 19323 30711 19329
rect 30745 19363 30803 19369
rect 30745 19329 30757 19363
rect 30791 19360 30803 19363
rect 30926 19360 30932 19372
rect 30791 19332 30932 19360
rect 30791 19329 30803 19332
rect 30745 19323 30803 19329
rect 28644 19264 28856 19292
rect 30392 19292 30420 19323
rect 30926 19320 30932 19332
rect 30984 19320 30990 19372
rect 31021 19363 31079 19369
rect 31021 19329 31033 19363
rect 31067 19360 31079 19363
rect 31726 19360 31754 19400
rect 33594 19388 33600 19400
rect 33652 19388 33658 19440
rect 34146 19428 34152 19440
rect 33704 19400 34152 19428
rect 31067 19332 31754 19360
rect 31067 19329 31079 19332
rect 31021 19323 31079 19329
rect 33410 19320 33416 19372
rect 33468 19360 33474 19372
rect 33704 19360 33732 19400
rect 34146 19388 34152 19400
rect 34204 19388 34210 19440
rect 34606 19388 34612 19440
rect 34664 19428 34670 19440
rect 35618 19428 35624 19440
rect 34664 19400 35624 19428
rect 34664 19388 34670 19400
rect 35618 19388 35624 19400
rect 35676 19388 35682 19440
rect 39114 19388 39120 19440
rect 39172 19428 39178 19440
rect 39393 19431 39451 19437
rect 39393 19428 39405 19431
rect 39172 19400 39405 19428
rect 39172 19388 39178 19400
rect 39393 19397 39405 19400
rect 39439 19397 39451 19431
rect 39393 19391 39451 19397
rect 33468 19332 33732 19360
rect 33468 19320 33474 19332
rect 33778 19320 33784 19372
rect 33836 19360 33842 19372
rect 35710 19360 35716 19372
rect 33836 19332 35716 19360
rect 33836 19320 33842 19332
rect 35710 19320 35716 19332
rect 35768 19320 35774 19372
rect 39574 19320 39580 19372
rect 39632 19320 39638 19372
rect 39666 19320 39672 19372
rect 39724 19320 39730 19372
rect 30392 19264 30788 19292
rect 28537 19255 28595 19261
rect 26602 19184 26608 19236
rect 26660 19184 26666 19236
rect 26697 19227 26755 19233
rect 26697 19193 26709 19227
rect 26743 19224 26755 19227
rect 26896 19224 26924 19252
rect 30760 19236 30788 19264
rect 31110 19252 31116 19304
rect 31168 19252 31174 19304
rect 32950 19252 32956 19304
rect 33008 19292 33014 19304
rect 33502 19292 33508 19304
rect 33008 19264 33508 19292
rect 33008 19252 33014 19264
rect 33502 19252 33508 19264
rect 33560 19252 33566 19304
rect 38746 19252 38752 19304
rect 38804 19292 38810 19304
rect 39114 19292 39120 19304
rect 38804 19264 39120 19292
rect 38804 19252 38810 19264
rect 39114 19252 39120 19264
rect 39172 19252 39178 19304
rect 28353 19227 28411 19233
rect 28353 19224 28365 19227
rect 26743 19196 26924 19224
rect 27632 19196 28365 19224
rect 26743 19193 26755 19196
rect 26697 19187 26755 19193
rect 27632 19156 27660 19196
rect 28353 19193 28365 19196
rect 28399 19193 28411 19227
rect 28353 19187 28411 19193
rect 30742 19184 30748 19236
rect 30800 19184 30806 19236
rect 31220 19196 31524 19224
rect 26436 19128 27660 19156
rect 27706 19116 27712 19168
rect 27764 19116 27770 19168
rect 30926 19116 30932 19168
rect 30984 19116 30990 19168
rect 31220 19165 31248 19196
rect 31205 19159 31263 19165
rect 31205 19125 31217 19159
rect 31251 19125 31263 19159
rect 31496 19156 31524 19196
rect 31570 19184 31576 19236
rect 31628 19224 31634 19236
rect 37366 19224 37372 19236
rect 31628 19196 37372 19224
rect 31628 19184 31634 19196
rect 37366 19184 37372 19196
rect 37424 19184 37430 19236
rect 32950 19156 32956 19168
rect 31496 19128 32956 19156
rect 31205 19119 31263 19125
rect 32950 19116 32956 19128
rect 33008 19116 33014 19168
rect 33134 19116 33140 19168
rect 33192 19156 33198 19168
rect 37734 19156 37740 19168
rect 33192 19128 37740 19156
rect 33192 19116 33198 19128
rect 37734 19116 37740 19128
rect 37792 19116 37798 19168
rect 39298 19116 39304 19168
rect 39356 19156 39362 19168
rect 39393 19159 39451 19165
rect 39393 19156 39405 19159
rect 39356 19128 39405 19156
rect 39356 19116 39362 19128
rect 39393 19125 39405 19128
rect 39439 19125 39451 19159
rect 39393 19119 39451 19125
rect 39850 19116 39856 19168
rect 39908 19116 39914 19168
rect 1104 19066 41400 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 41400 19066
rect 1104 18992 41400 19014
rect 3789 18955 3847 18961
rect 3789 18921 3801 18955
rect 3835 18952 3847 18955
rect 3970 18952 3976 18964
rect 3835 18924 3976 18952
rect 3835 18921 3847 18924
rect 3789 18915 3847 18921
rect 3970 18912 3976 18924
rect 4028 18912 4034 18964
rect 5718 18912 5724 18964
rect 5776 18912 5782 18964
rect 5997 18955 6055 18961
rect 5997 18921 6009 18955
rect 6043 18952 6055 18955
rect 7374 18952 7380 18964
rect 6043 18924 7380 18952
rect 6043 18921 6055 18924
rect 5997 18915 6055 18921
rect 7374 18912 7380 18924
rect 7432 18912 7438 18964
rect 7834 18912 7840 18964
rect 7892 18912 7898 18964
rect 8294 18912 8300 18964
rect 8352 18952 8358 18964
rect 8573 18955 8631 18961
rect 8573 18952 8585 18955
rect 8352 18924 8585 18952
rect 8352 18912 8358 18924
rect 8573 18921 8585 18924
rect 8619 18921 8631 18955
rect 8573 18915 8631 18921
rect 8754 18912 8760 18964
rect 8812 18952 8818 18964
rect 11977 18955 12035 18961
rect 8812 18924 11928 18952
rect 8812 18912 8818 18924
rect 2866 18776 2872 18828
rect 2924 18816 2930 18828
rect 4341 18819 4399 18825
rect 4341 18816 4353 18819
rect 2924 18788 4353 18816
rect 2924 18776 2930 18788
rect 4341 18785 4353 18788
rect 4387 18816 4399 18819
rect 4709 18819 4767 18825
rect 4387 18788 4476 18816
rect 4387 18785 4399 18788
rect 4341 18779 4399 18785
rect 4448 18760 4476 18788
rect 4709 18785 4721 18819
rect 4755 18816 4767 18819
rect 5074 18816 5080 18828
rect 4755 18788 5080 18816
rect 4755 18785 4767 18788
rect 4709 18779 4767 18785
rect 5074 18776 5080 18788
rect 5132 18776 5138 18828
rect 4430 18708 4436 18760
rect 4488 18708 4494 18760
rect 5445 18751 5503 18757
rect 5445 18717 5457 18751
rect 5491 18748 5503 18751
rect 5534 18748 5540 18760
rect 5491 18720 5540 18748
rect 5491 18717 5503 18720
rect 5445 18711 5503 18717
rect 5534 18708 5540 18720
rect 5592 18708 5598 18760
rect 5626 18708 5632 18760
rect 5684 18708 5690 18760
rect 5736 18748 5764 18912
rect 7852 18816 7880 18912
rect 11900 18884 11928 18924
rect 11977 18921 11989 18955
rect 12023 18952 12035 18955
rect 12158 18952 12164 18964
rect 12023 18924 12164 18952
rect 12023 18921 12035 18924
rect 11977 18915 12035 18921
rect 12158 18912 12164 18924
rect 12216 18912 12222 18964
rect 12713 18955 12771 18961
rect 12713 18921 12725 18955
rect 12759 18952 12771 18955
rect 12802 18952 12808 18964
rect 12759 18924 12808 18952
rect 12759 18921 12771 18924
rect 12713 18915 12771 18921
rect 12802 18912 12808 18924
rect 12860 18912 12866 18964
rect 15930 18912 15936 18964
rect 15988 18952 15994 18964
rect 17954 18952 17960 18964
rect 15988 18924 17960 18952
rect 15988 18912 15994 18924
rect 17954 18912 17960 18924
rect 18012 18912 18018 18964
rect 18782 18912 18788 18964
rect 18840 18952 18846 18964
rect 18840 18924 21404 18952
rect 18840 18912 18846 18924
rect 14826 18884 14832 18896
rect 11900 18856 14832 18884
rect 14826 18844 14832 18856
rect 14884 18844 14890 18896
rect 19150 18884 19156 18896
rect 16960 18856 19156 18884
rect 7929 18819 7987 18825
rect 7929 18816 7941 18819
rect 7852 18788 7941 18816
rect 7929 18785 7941 18788
rect 7975 18785 7987 18819
rect 7929 18779 7987 18785
rect 10505 18819 10563 18825
rect 10505 18785 10517 18819
rect 10551 18816 10563 18819
rect 10594 18816 10600 18828
rect 10551 18788 10600 18816
rect 10551 18785 10563 18788
rect 10505 18779 10563 18785
rect 10594 18776 10600 18788
rect 10652 18776 10658 18828
rect 12710 18816 12716 18828
rect 12084 18788 12716 18816
rect 5813 18751 5871 18757
rect 5813 18748 5825 18751
rect 5736 18720 5825 18748
rect 5813 18717 5825 18720
rect 5859 18717 5871 18751
rect 5813 18711 5871 18717
rect 5994 18708 6000 18760
rect 6052 18748 6058 18760
rect 6089 18751 6147 18757
rect 6089 18748 6101 18751
rect 6052 18720 6101 18748
rect 6052 18708 6058 18720
rect 6089 18717 6101 18720
rect 6135 18717 6147 18751
rect 6089 18711 6147 18717
rect 9950 18708 9956 18760
rect 10008 18748 10014 18760
rect 10229 18751 10287 18757
rect 10229 18748 10241 18751
rect 10008 18720 10241 18748
rect 10008 18708 10014 18720
rect 10229 18717 10241 18720
rect 10275 18717 10287 18751
rect 10229 18711 10287 18717
rect 11606 18708 11612 18760
rect 11664 18708 11670 18760
rect 12084 18757 12112 18788
rect 12710 18776 12716 18788
rect 12768 18776 12774 18828
rect 16850 18776 16856 18828
rect 16908 18816 16914 18828
rect 16960 18825 16988 18856
rect 19150 18844 19156 18856
rect 19208 18844 19214 18896
rect 19306 18856 21036 18884
rect 16945 18819 17003 18825
rect 16945 18816 16957 18819
rect 16908 18788 16957 18816
rect 16908 18776 16914 18788
rect 16945 18785 16957 18788
rect 16991 18785 17003 18819
rect 19306 18816 19334 18856
rect 21008 18828 21036 18856
rect 16945 18779 17003 18785
rect 17144 18788 19334 18816
rect 12069 18751 12127 18757
rect 12069 18717 12081 18751
rect 12115 18717 12127 18751
rect 12069 18711 12127 18717
rect 12158 18708 12164 18760
rect 12216 18748 12222 18760
rect 12216 18720 12261 18748
rect 12216 18708 12222 18720
rect 12342 18708 12348 18760
rect 12400 18708 12406 18760
rect 12575 18751 12633 18757
rect 12575 18717 12587 18751
rect 12621 18748 12633 18751
rect 12894 18748 12900 18760
rect 12621 18720 12900 18748
rect 12621 18717 12633 18720
rect 12575 18711 12633 18717
rect 12894 18708 12900 18720
rect 12952 18708 12958 18760
rect 17144 18757 17172 18788
rect 20622 18776 20628 18828
rect 20680 18776 20686 18828
rect 20898 18776 20904 18828
rect 20956 18776 20962 18828
rect 20990 18776 20996 18828
rect 21048 18776 21054 18828
rect 21174 18776 21180 18828
rect 21232 18776 21238 18828
rect 17129 18751 17187 18757
rect 17129 18717 17141 18751
rect 17175 18717 17187 18751
rect 17129 18711 17187 18717
rect 17954 18708 17960 18760
rect 18012 18748 18018 18760
rect 18322 18748 18328 18760
rect 18012 18720 18328 18748
rect 18012 18708 18018 18720
rect 18322 18708 18328 18720
rect 18380 18708 18386 18760
rect 20441 18751 20499 18757
rect 20441 18717 20453 18751
rect 20487 18748 20499 18751
rect 20640 18748 20668 18776
rect 20487 18720 20668 18748
rect 20717 18751 20775 18757
rect 20487 18717 20499 18720
rect 20441 18711 20499 18717
rect 20717 18717 20729 18751
rect 20763 18748 20775 18751
rect 20916 18748 20944 18776
rect 20763 18720 20944 18748
rect 20763 18717 20775 18720
rect 20717 18711 20775 18717
rect 21082 18708 21088 18760
rect 21140 18708 21146 18760
rect 21269 18751 21327 18757
rect 21269 18717 21281 18751
rect 21315 18717 21327 18751
rect 21376 18748 21404 18924
rect 21450 18912 21456 18964
rect 21508 18912 21514 18964
rect 22925 18955 22983 18961
rect 22925 18921 22937 18955
rect 22971 18952 22983 18955
rect 23198 18952 23204 18964
rect 22971 18924 23204 18952
rect 22971 18921 22983 18924
rect 22925 18915 22983 18921
rect 23198 18912 23204 18924
rect 23256 18912 23262 18964
rect 23750 18912 23756 18964
rect 23808 18952 23814 18964
rect 24578 18952 24584 18964
rect 23808 18924 24584 18952
rect 23808 18912 23814 18924
rect 24578 18912 24584 18924
rect 24636 18912 24642 18964
rect 25501 18955 25559 18961
rect 25501 18921 25513 18955
rect 25547 18952 25559 18955
rect 25590 18952 25596 18964
rect 25547 18924 25596 18952
rect 25547 18921 25559 18924
rect 25501 18915 25559 18921
rect 25590 18912 25596 18924
rect 25648 18912 25654 18964
rect 25682 18912 25688 18964
rect 25740 18952 25746 18964
rect 26513 18955 26571 18961
rect 26513 18952 26525 18955
rect 25740 18924 26525 18952
rect 25740 18912 25746 18924
rect 26513 18921 26525 18924
rect 26559 18921 26571 18955
rect 26513 18915 26571 18921
rect 26602 18912 26608 18964
rect 26660 18952 26666 18964
rect 30926 18952 30932 18964
rect 26660 18924 30932 18952
rect 26660 18912 26666 18924
rect 30926 18912 30932 18924
rect 30984 18912 30990 18964
rect 31297 18955 31355 18961
rect 31297 18921 31309 18955
rect 31343 18952 31355 18955
rect 31570 18952 31576 18964
rect 31343 18924 31576 18952
rect 31343 18921 31355 18924
rect 31297 18915 31355 18921
rect 31570 18912 31576 18924
rect 31628 18912 31634 18964
rect 31662 18912 31668 18964
rect 31720 18952 31726 18964
rect 32490 18952 32496 18964
rect 31720 18924 32496 18952
rect 31720 18912 31726 18924
rect 32490 18912 32496 18924
rect 32548 18912 32554 18964
rect 34054 18952 34060 18964
rect 32876 18924 34060 18952
rect 23109 18887 23167 18893
rect 23109 18853 23121 18887
rect 23155 18853 23167 18887
rect 23109 18847 23167 18853
rect 22002 18776 22008 18828
rect 22060 18776 22066 18828
rect 22830 18776 22836 18828
rect 22888 18776 22894 18828
rect 23124 18816 23152 18847
rect 23845 18819 23903 18825
rect 23124 18788 23704 18816
rect 21729 18751 21787 18757
rect 21729 18748 21741 18751
rect 21376 18720 21741 18748
rect 21269 18711 21327 18717
rect 21729 18717 21741 18720
rect 21775 18717 21787 18751
rect 21729 18711 21787 18717
rect 21913 18751 21971 18757
rect 21913 18717 21925 18751
rect 21959 18748 21971 18751
rect 22925 18751 22983 18757
rect 21959 18720 22094 18748
rect 21959 18717 21971 18720
rect 21913 18711 21971 18717
rect 4157 18683 4215 18689
rect 4157 18649 4169 18683
rect 4203 18680 4215 18683
rect 5261 18683 5319 18689
rect 5261 18680 5273 18683
rect 4203 18652 5273 18680
rect 4203 18649 4215 18652
rect 4157 18643 4215 18649
rect 5261 18649 5273 18652
rect 5307 18649 5319 18683
rect 5261 18643 5319 18649
rect 5721 18683 5779 18689
rect 5721 18649 5733 18683
rect 5767 18680 5779 18683
rect 6365 18683 6423 18689
rect 5767 18652 6224 18680
rect 5767 18649 5779 18652
rect 5721 18643 5779 18649
rect 6196 18624 6224 18652
rect 6365 18649 6377 18683
rect 6411 18649 6423 18683
rect 7590 18652 9352 18680
rect 6365 18643 6423 18649
rect 4249 18615 4307 18621
rect 4249 18581 4261 18615
rect 4295 18612 4307 18615
rect 4798 18612 4804 18624
rect 4295 18584 4804 18612
rect 4295 18581 4307 18584
rect 4249 18575 4307 18581
rect 4798 18572 4804 18584
rect 4856 18572 4862 18624
rect 6178 18572 6184 18624
rect 6236 18572 6242 18624
rect 6380 18612 6408 18643
rect 7098 18612 7104 18624
rect 6380 18584 7104 18612
rect 7098 18572 7104 18584
rect 7156 18572 7162 18624
rect 7282 18572 7288 18624
rect 7340 18612 7346 18624
rect 7668 18612 7696 18652
rect 9324 18624 9352 18652
rect 7340 18584 7696 18612
rect 7340 18572 7346 18584
rect 9306 18572 9312 18624
rect 9364 18612 9370 18624
rect 11624 18612 11652 18708
rect 12437 18683 12495 18689
rect 12437 18649 12449 18683
rect 12483 18649 12495 18683
rect 12437 18643 12495 18649
rect 16485 18683 16543 18689
rect 16485 18649 16497 18683
rect 16531 18680 16543 18683
rect 17313 18683 17371 18689
rect 17313 18680 17325 18683
rect 16531 18652 17325 18680
rect 16531 18649 16543 18652
rect 16485 18643 16543 18649
rect 17313 18649 17325 18652
rect 17359 18649 17371 18683
rect 17313 18643 17371 18649
rect 9364 18584 11652 18612
rect 9364 18572 9370 18584
rect 12250 18572 12256 18624
rect 12308 18612 12314 18624
rect 12452 18612 12480 18643
rect 18598 18640 18604 18692
rect 18656 18640 18662 18692
rect 20809 18683 20867 18689
rect 20809 18680 20821 18683
rect 20548 18652 20821 18680
rect 20548 18624 20576 18652
rect 20809 18649 20821 18652
rect 20855 18649 20867 18683
rect 20809 18643 20867 18649
rect 12308 18584 12480 18612
rect 12308 18572 12314 18584
rect 14734 18572 14740 18624
rect 14792 18612 14798 18624
rect 16577 18615 16635 18621
rect 16577 18612 16589 18615
rect 14792 18584 16589 18612
rect 14792 18572 14798 18584
rect 16577 18581 16589 18584
rect 16623 18581 16635 18615
rect 16577 18575 16635 18581
rect 18690 18572 18696 18624
rect 18748 18572 18754 18624
rect 20530 18612 20536 18624
rect 20588 18621 20594 18624
rect 20449 18584 20536 18612
rect 20530 18572 20536 18584
rect 20588 18575 20597 18621
rect 20625 18615 20683 18621
rect 20625 18581 20637 18615
rect 20671 18612 20683 18615
rect 21100 18612 21128 18708
rect 21284 18680 21312 18711
rect 21284 18652 21772 18680
rect 21744 18624 21772 18652
rect 20671 18584 21128 18612
rect 20671 18581 20683 18584
rect 20625 18575 20683 18581
rect 20588 18572 20594 18575
rect 21542 18572 21548 18624
rect 21600 18572 21606 18624
rect 21726 18572 21732 18624
rect 21784 18572 21790 18624
rect 22066 18612 22094 18720
rect 22925 18717 22937 18751
rect 22971 18748 22983 18751
rect 23382 18748 23388 18760
rect 22971 18720 23388 18748
rect 22971 18717 22983 18720
rect 22925 18711 22983 18717
rect 23382 18708 23388 18720
rect 23440 18708 23446 18760
rect 23474 18708 23480 18760
rect 23532 18748 23538 18760
rect 23676 18757 23704 18788
rect 23845 18785 23857 18819
rect 23891 18785 23903 18819
rect 25597 18816 25625 18912
rect 26697 18887 26755 18893
rect 26697 18853 26709 18887
rect 26743 18853 26755 18887
rect 32674 18884 32680 18896
rect 26697 18847 26755 18853
rect 31680 18856 32680 18884
rect 26712 18816 26740 18847
rect 25597 18788 25729 18816
rect 23845 18779 23903 18785
rect 23569 18751 23627 18757
rect 23569 18748 23581 18751
rect 23532 18720 23581 18748
rect 23532 18708 23538 18720
rect 23569 18717 23581 18720
rect 23615 18717 23627 18751
rect 23569 18711 23627 18717
rect 23661 18751 23719 18757
rect 23661 18717 23673 18751
rect 23707 18717 23719 18751
rect 23661 18711 23719 18717
rect 22186 18640 22192 18692
rect 22244 18680 22250 18692
rect 22649 18683 22707 18689
rect 22649 18680 22661 18683
rect 22244 18652 22661 18680
rect 22244 18640 22250 18652
rect 22649 18649 22661 18652
rect 22695 18680 22707 18683
rect 23750 18680 23756 18692
rect 22695 18652 23756 18680
rect 22695 18649 22707 18652
rect 22649 18643 22707 18649
rect 23750 18640 23756 18652
rect 23808 18640 23814 18692
rect 23290 18612 23296 18624
rect 22066 18584 23296 18612
rect 23290 18572 23296 18584
rect 23348 18572 23354 18624
rect 23382 18572 23388 18624
rect 23440 18572 23446 18624
rect 23860 18612 23888 18779
rect 23937 18751 23995 18757
rect 23937 18717 23949 18751
rect 23983 18748 23995 18751
rect 24762 18748 24768 18760
rect 23983 18720 24768 18748
rect 23983 18717 23995 18720
rect 23937 18711 23995 18717
rect 24762 18708 24768 18720
rect 24820 18708 24826 18760
rect 25130 18708 25136 18760
rect 25188 18708 25194 18760
rect 25701 18757 25729 18788
rect 25976 18788 26740 18816
rect 25593 18751 25651 18757
rect 25593 18717 25605 18751
rect 25639 18717 25651 18751
rect 25593 18711 25651 18717
rect 25686 18751 25744 18757
rect 25686 18717 25698 18751
rect 25732 18717 25744 18751
rect 25976 18748 26004 18788
rect 25686 18711 25744 18717
rect 25792 18720 26004 18748
rect 25314 18640 25320 18692
rect 25372 18680 25378 18692
rect 25498 18680 25504 18692
rect 25372 18652 25504 18680
rect 25372 18640 25378 18652
rect 25498 18640 25504 18652
rect 25556 18640 25562 18692
rect 25608 18680 25636 18711
rect 25792 18680 25820 18720
rect 26050 18708 26056 18760
rect 26108 18757 26114 18760
rect 31680 18757 31708 18856
rect 32674 18844 32680 18856
rect 32732 18844 32738 18896
rect 32876 18884 32904 18924
rect 34054 18912 34060 18924
rect 34112 18952 34118 18964
rect 35434 18952 35440 18964
rect 34112 18924 35440 18952
rect 34112 18912 34118 18924
rect 35434 18912 35440 18924
rect 35492 18912 35498 18964
rect 35989 18955 36047 18961
rect 35989 18921 36001 18955
rect 36035 18952 36047 18955
rect 36449 18955 36507 18961
rect 36449 18952 36461 18955
rect 36035 18924 36461 18952
rect 36035 18921 36047 18924
rect 35989 18915 36047 18921
rect 36449 18921 36461 18924
rect 36495 18952 36507 18955
rect 36495 18924 36952 18952
rect 36495 18921 36507 18924
rect 36449 18915 36507 18921
rect 32784 18856 32904 18884
rect 33413 18887 33471 18893
rect 31941 18819 31999 18825
rect 31941 18785 31953 18819
rect 31987 18816 31999 18819
rect 32582 18816 32588 18828
rect 31987 18788 32588 18816
rect 31987 18785 31999 18788
rect 31941 18779 31999 18785
rect 32582 18776 32588 18788
rect 32640 18816 32646 18828
rect 32784 18816 32812 18856
rect 33413 18853 33425 18887
rect 33459 18884 33471 18887
rect 33459 18856 36584 18884
rect 33459 18853 33471 18856
rect 33413 18847 33471 18853
rect 34422 18816 34428 18828
rect 32640 18788 32812 18816
rect 33060 18788 33456 18816
rect 32640 18776 32646 18788
rect 26108 18748 26116 18757
rect 31481 18751 31539 18757
rect 26108 18720 26153 18748
rect 26108 18711 26116 18720
rect 31481 18717 31493 18751
rect 31527 18717 31539 18751
rect 31481 18711 31539 18717
rect 31665 18751 31723 18757
rect 31665 18717 31677 18751
rect 31711 18717 31723 18751
rect 31665 18711 31723 18717
rect 26108 18708 26114 18711
rect 25608 18652 25820 18680
rect 25866 18640 25872 18692
rect 25924 18640 25930 18692
rect 25961 18683 26019 18689
rect 25961 18649 25973 18683
rect 26007 18680 26019 18683
rect 26142 18680 26148 18692
rect 26007 18652 26148 18680
rect 26007 18649 26019 18652
rect 25961 18643 26019 18649
rect 26142 18640 26148 18652
rect 26200 18640 26206 18692
rect 26326 18640 26332 18692
rect 26384 18640 26390 18692
rect 26237 18615 26295 18621
rect 26237 18612 26249 18615
rect 23860 18584 26249 18612
rect 26237 18581 26249 18584
rect 26283 18581 26295 18615
rect 26237 18575 26295 18581
rect 26510 18572 26516 18624
rect 26568 18621 26574 18624
rect 26568 18615 26587 18621
rect 26575 18581 26587 18615
rect 26568 18575 26587 18581
rect 26568 18572 26574 18575
rect 27338 18572 27344 18624
rect 27396 18612 27402 18624
rect 31386 18612 31392 18624
rect 27396 18584 31392 18612
rect 27396 18572 27402 18584
rect 31386 18572 31392 18584
rect 31444 18572 31450 18624
rect 31496 18612 31524 18711
rect 31754 18708 31760 18760
rect 31812 18757 31818 18760
rect 31812 18751 31841 18757
rect 31829 18717 31841 18751
rect 31812 18711 31841 18717
rect 31812 18708 31818 18711
rect 32766 18708 32772 18760
rect 32824 18742 32830 18760
rect 33060 18757 33088 18788
rect 32861 18751 32919 18757
rect 32861 18742 32873 18751
rect 32824 18717 32873 18742
rect 32907 18717 32919 18751
rect 32824 18714 32919 18717
rect 32824 18708 32830 18714
rect 32861 18711 32919 18714
rect 33045 18751 33103 18757
rect 33045 18717 33057 18751
rect 33091 18717 33103 18751
rect 33045 18711 33103 18717
rect 33134 18708 33140 18760
rect 33192 18708 33198 18760
rect 33229 18751 33287 18757
rect 33229 18717 33241 18751
rect 33275 18717 33287 18751
rect 33229 18711 33287 18717
rect 31573 18683 31631 18689
rect 31573 18649 31585 18683
rect 31619 18680 31631 18683
rect 33244 18680 33272 18711
rect 33428 18692 33456 18788
rect 33796 18788 34428 18816
rect 33796 18757 33824 18788
rect 34422 18776 34428 18788
rect 34480 18776 34486 18828
rect 34882 18776 34888 18828
rect 34940 18816 34946 18828
rect 36265 18819 36323 18825
rect 36265 18816 36277 18819
rect 34940 18788 36277 18816
rect 34940 18776 34946 18788
rect 36265 18785 36277 18788
rect 36311 18785 36323 18819
rect 36265 18779 36323 18785
rect 33505 18751 33563 18757
rect 33505 18717 33517 18751
rect 33551 18717 33563 18751
rect 33505 18711 33563 18717
rect 33781 18751 33839 18757
rect 33781 18717 33793 18751
rect 33827 18717 33839 18751
rect 33781 18711 33839 18717
rect 33873 18751 33931 18757
rect 33873 18717 33885 18751
rect 33919 18748 33931 18751
rect 34054 18748 34060 18760
rect 33919 18720 34060 18748
rect 33919 18717 33931 18720
rect 33873 18711 33931 18717
rect 31619 18652 31892 18680
rect 31619 18649 31631 18652
rect 31573 18643 31631 18649
rect 31662 18612 31668 18624
rect 31496 18584 31668 18612
rect 31662 18572 31668 18584
rect 31720 18572 31726 18624
rect 31864 18612 31892 18652
rect 33152 18652 33272 18680
rect 33152 18624 33180 18652
rect 33410 18640 33416 18692
rect 33468 18640 33474 18692
rect 33520 18624 33548 18711
rect 34054 18708 34060 18720
rect 34112 18708 34118 18760
rect 34698 18708 34704 18760
rect 34756 18748 34762 18760
rect 35437 18751 35495 18757
rect 35437 18748 35449 18751
rect 34756 18720 35449 18748
rect 34756 18708 34762 18720
rect 35437 18717 35449 18720
rect 35483 18717 35495 18751
rect 35437 18711 35495 18717
rect 35710 18708 35716 18760
rect 35768 18708 35774 18760
rect 35802 18708 35808 18760
rect 35860 18708 35866 18760
rect 36449 18751 36507 18757
rect 36449 18717 36461 18751
rect 36495 18717 36507 18751
rect 36556 18748 36584 18856
rect 36630 18844 36636 18896
rect 36688 18844 36694 18896
rect 36924 18757 36952 18924
rect 37274 18912 37280 18964
rect 37332 18912 37338 18964
rect 37826 18912 37832 18964
rect 37884 18912 37890 18964
rect 38010 18912 38016 18964
rect 38068 18952 38074 18964
rect 38473 18955 38531 18961
rect 38473 18952 38485 18955
rect 38068 18924 38485 18952
rect 38068 18912 38074 18924
rect 38473 18921 38485 18924
rect 38519 18921 38531 18955
rect 38473 18915 38531 18921
rect 39850 18912 39856 18964
rect 39908 18912 39914 18964
rect 40037 18955 40095 18961
rect 40037 18921 40049 18955
rect 40083 18921 40095 18955
rect 40037 18915 40095 18921
rect 37292 18884 37320 18912
rect 38286 18884 38292 18896
rect 37292 18856 38292 18884
rect 38286 18844 38292 18856
rect 38344 18884 38350 18896
rect 38344 18856 38516 18884
rect 38344 18844 38350 18856
rect 37093 18819 37151 18825
rect 37093 18785 37105 18819
rect 37139 18816 37151 18819
rect 37550 18816 37556 18828
rect 37139 18788 37556 18816
rect 37139 18785 37151 18788
rect 37093 18779 37151 18785
rect 37550 18776 37556 18788
rect 37608 18816 37614 18828
rect 37608 18788 38240 18816
rect 37608 18776 37614 18788
rect 36725 18751 36783 18757
rect 36725 18748 36737 18751
rect 36556 18720 36737 18748
rect 36449 18711 36507 18717
rect 36725 18717 36737 18720
rect 36771 18717 36783 18751
rect 36725 18711 36783 18717
rect 36909 18751 36967 18757
rect 36909 18717 36921 18751
rect 36955 18717 36967 18751
rect 36909 18711 36967 18717
rect 33686 18640 33692 18692
rect 33744 18640 33750 18692
rect 34716 18680 34744 18708
rect 33796 18652 34744 18680
rect 32490 18612 32496 18624
rect 31864 18584 32496 18612
rect 32490 18572 32496 18584
rect 32548 18572 32554 18624
rect 33134 18572 33140 18624
rect 33192 18572 33198 18624
rect 33502 18572 33508 18624
rect 33560 18612 33566 18624
rect 33796 18612 33824 18652
rect 35158 18640 35164 18692
rect 35216 18680 35222 18692
rect 35621 18683 35679 18689
rect 35621 18680 35633 18683
rect 35216 18652 35633 18680
rect 35216 18640 35222 18652
rect 35621 18649 35633 18652
rect 35667 18649 35679 18683
rect 35621 18643 35679 18649
rect 36173 18683 36231 18689
rect 36173 18649 36185 18683
rect 36219 18680 36231 18683
rect 36354 18680 36360 18692
rect 36219 18652 36360 18680
rect 36219 18649 36231 18652
rect 36173 18643 36231 18649
rect 36354 18640 36360 18652
rect 36412 18640 36418 18692
rect 36464 18624 36492 18711
rect 36740 18680 36768 18711
rect 37366 18708 37372 18760
rect 37424 18748 37430 18760
rect 37829 18751 37887 18757
rect 37829 18748 37841 18751
rect 37424 18720 37841 18748
rect 37424 18708 37430 18720
rect 37829 18717 37841 18720
rect 37875 18717 37887 18751
rect 37829 18711 37887 18717
rect 37918 18708 37924 18760
rect 37976 18748 37982 18760
rect 38013 18751 38071 18757
rect 38013 18748 38025 18751
rect 37976 18720 38025 18748
rect 37976 18708 37982 18720
rect 38013 18717 38025 18720
rect 38059 18717 38071 18751
rect 38013 18711 38071 18717
rect 37274 18680 37280 18692
rect 36740 18652 37280 18680
rect 37274 18640 37280 18652
rect 37332 18640 37338 18692
rect 37553 18683 37611 18689
rect 37553 18649 37565 18683
rect 37599 18680 37611 18683
rect 38102 18680 38108 18692
rect 37599 18652 38108 18680
rect 37599 18649 37611 18652
rect 37553 18643 37611 18649
rect 38102 18640 38108 18652
rect 38160 18640 38166 18692
rect 38212 18680 38240 18788
rect 38488 18757 38516 18856
rect 38473 18751 38531 18757
rect 38473 18717 38485 18751
rect 38519 18717 38531 18751
rect 38473 18711 38531 18717
rect 38657 18751 38715 18757
rect 38657 18717 38669 18751
rect 38703 18717 38715 18751
rect 38657 18711 38715 18717
rect 38672 18680 38700 18711
rect 38746 18708 38752 18760
rect 38804 18708 38810 18760
rect 39868 18757 39896 18912
rect 39858 18751 39916 18757
rect 39858 18717 39870 18751
rect 39904 18717 39916 18751
rect 39858 18711 39916 18717
rect 39945 18751 40003 18757
rect 39945 18717 39957 18751
rect 39991 18717 40003 18751
rect 39945 18711 40003 18717
rect 38212 18652 38700 18680
rect 39022 18640 39028 18692
rect 39080 18680 39086 18692
rect 39960 18680 39988 18711
rect 39080 18652 39988 18680
rect 39080 18640 39086 18652
rect 40052 18624 40080 18915
rect 40218 18912 40224 18964
rect 40276 18912 40282 18964
rect 33560 18584 33824 18612
rect 34057 18615 34115 18621
rect 33560 18572 33566 18584
rect 34057 18581 34069 18615
rect 34103 18612 34115 18615
rect 36446 18612 36452 18624
rect 34103 18584 36452 18612
rect 34103 18581 34115 18584
rect 34057 18575 34115 18581
rect 36446 18572 36452 18584
rect 36504 18572 36510 18624
rect 38194 18572 38200 18624
rect 38252 18572 38258 18624
rect 38933 18615 38991 18621
rect 38933 18581 38945 18615
rect 38979 18612 38991 18615
rect 40034 18612 40040 18624
rect 38979 18584 40040 18612
rect 38979 18581 38991 18584
rect 38933 18575 38991 18581
rect 40034 18572 40040 18584
rect 40092 18572 40098 18624
rect 1104 18522 41400 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 41400 18522
rect 1104 18448 41400 18470
rect 4985 18411 5043 18417
rect 4985 18377 4997 18411
rect 5031 18377 5043 18411
rect 4985 18371 5043 18377
rect 2869 18275 2927 18281
rect 2869 18241 2881 18275
rect 2915 18272 2927 18275
rect 3973 18275 4031 18281
rect 3973 18272 3985 18275
rect 2915 18244 3985 18272
rect 2915 18241 2927 18244
rect 2869 18235 2927 18241
rect 3973 18241 3985 18244
rect 4019 18241 4031 18275
rect 3973 18235 4031 18241
rect 4062 18232 4068 18284
rect 4120 18232 4126 18284
rect 4893 18275 4951 18281
rect 4893 18241 4905 18275
rect 4939 18272 4951 18275
rect 5000 18272 5028 18371
rect 6914 18368 6920 18420
rect 6972 18368 6978 18420
rect 7098 18368 7104 18420
rect 7156 18368 7162 18420
rect 9125 18411 9183 18417
rect 9125 18377 9137 18411
rect 9171 18408 9183 18411
rect 9766 18408 9772 18420
rect 9171 18380 9772 18408
rect 9171 18377 9183 18380
rect 9125 18371 9183 18377
rect 9766 18368 9772 18380
rect 9824 18408 9830 18420
rect 10410 18408 10416 18420
rect 9824 18380 10416 18408
rect 9824 18368 9830 18380
rect 10410 18368 10416 18380
rect 10468 18368 10474 18420
rect 14458 18368 14464 18420
rect 14516 18368 14522 18420
rect 16022 18408 16028 18420
rect 14660 18380 16028 18408
rect 4939 18244 5028 18272
rect 5353 18275 5411 18281
rect 4939 18241 4951 18244
rect 4893 18235 4951 18241
rect 5353 18241 5365 18275
rect 5399 18272 5411 18275
rect 6932 18272 6960 18368
rect 14553 18343 14611 18349
rect 14553 18340 14565 18343
rect 14384 18312 14565 18340
rect 14384 18284 14412 18312
rect 14553 18309 14565 18312
rect 14599 18309 14611 18343
rect 14553 18303 14611 18309
rect 7285 18275 7343 18281
rect 7285 18272 7297 18275
rect 5399 18244 6500 18272
rect 6932 18244 7297 18272
rect 5399 18241 5411 18244
rect 5353 18235 5411 18241
rect 2958 18164 2964 18216
rect 3016 18164 3022 18216
rect 3145 18207 3203 18213
rect 3145 18173 3157 18207
rect 3191 18173 3203 18207
rect 3145 18167 3203 18173
rect 3160 18136 3188 18167
rect 3418 18164 3424 18216
rect 3476 18204 3482 18216
rect 4080 18204 4108 18232
rect 3476 18176 4108 18204
rect 3476 18164 3482 18176
rect 5258 18164 5264 18216
rect 5316 18204 5322 18216
rect 5445 18207 5503 18213
rect 5445 18204 5457 18207
rect 5316 18176 5457 18204
rect 5316 18164 5322 18176
rect 5445 18173 5457 18176
rect 5491 18173 5503 18207
rect 5445 18167 5503 18173
rect 5537 18207 5595 18213
rect 5537 18173 5549 18207
rect 5583 18173 5595 18207
rect 5537 18167 5595 18173
rect 4430 18136 4436 18148
rect 3160 18108 4436 18136
rect 4430 18096 4436 18108
rect 4488 18136 4494 18148
rect 5552 18136 5580 18167
rect 5626 18164 5632 18216
rect 5684 18204 5690 18216
rect 6365 18207 6423 18213
rect 6365 18204 6377 18207
rect 5684 18176 6377 18204
rect 5684 18164 5690 18176
rect 6365 18173 6377 18176
rect 6411 18173 6423 18207
rect 6472 18204 6500 18244
rect 7285 18241 7297 18244
rect 7331 18241 7343 18275
rect 7285 18235 7343 18241
rect 8386 18232 8392 18284
rect 8444 18272 8450 18284
rect 8444 18244 14320 18272
rect 8444 18232 8450 18244
rect 7009 18207 7067 18213
rect 7009 18204 7021 18207
rect 6472 18176 7021 18204
rect 6365 18167 6423 18173
rect 7009 18173 7021 18176
rect 7055 18173 7067 18207
rect 7009 18167 7067 18173
rect 9214 18164 9220 18216
rect 9272 18164 9278 18216
rect 9398 18164 9404 18216
rect 9456 18204 9462 18216
rect 14292 18204 14320 18244
rect 14366 18232 14372 18284
rect 14424 18232 14430 18284
rect 14660 18204 14688 18380
rect 16022 18368 16028 18380
rect 16080 18368 16086 18420
rect 16942 18368 16948 18420
rect 17000 18408 17006 18420
rect 18506 18408 18512 18420
rect 17000 18380 18512 18408
rect 17000 18368 17006 18380
rect 18506 18368 18512 18380
rect 18564 18368 18570 18420
rect 18598 18368 18604 18420
rect 18656 18408 18662 18420
rect 18693 18411 18751 18417
rect 18693 18408 18705 18411
rect 18656 18380 18705 18408
rect 18656 18368 18662 18380
rect 18693 18377 18705 18380
rect 18739 18377 18751 18411
rect 18693 18371 18751 18377
rect 20622 18368 20628 18420
rect 20680 18368 20686 18420
rect 21542 18368 21548 18420
rect 21600 18368 21606 18420
rect 24118 18368 24124 18420
rect 24176 18408 24182 18420
rect 26510 18408 26516 18420
rect 24176 18380 26516 18408
rect 24176 18368 24182 18380
rect 26510 18368 26516 18380
rect 26568 18368 26574 18420
rect 27338 18368 27344 18420
rect 27396 18368 27402 18420
rect 30466 18408 30472 18420
rect 29840 18380 30472 18408
rect 20640 18340 20668 18368
rect 16961 18312 17816 18340
rect 15470 18232 15476 18284
rect 15528 18272 15534 18284
rect 15749 18275 15807 18281
rect 15749 18272 15761 18275
rect 15528 18244 15761 18272
rect 15528 18232 15534 18244
rect 15749 18241 15761 18244
rect 15795 18272 15807 18275
rect 15930 18272 15936 18284
rect 15795 18244 15936 18272
rect 15795 18241 15807 18244
rect 15749 18235 15807 18241
rect 15930 18232 15936 18244
rect 15988 18232 15994 18284
rect 16022 18232 16028 18284
rect 16080 18232 16086 18284
rect 16298 18232 16304 18284
rect 16356 18232 16362 18284
rect 16961 18281 16989 18312
rect 17788 18284 17816 18312
rect 18064 18312 20668 18340
rect 16485 18275 16543 18281
rect 16485 18241 16497 18275
rect 16531 18241 16543 18275
rect 16485 18235 16543 18241
rect 16945 18275 17003 18281
rect 16945 18241 16957 18275
rect 16991 18241 17003 18275
rect 16945 18235 17003 18241
rect 17037 18275 17095 18281
rect 17037 18241 17049 18275
rect 17083 18272 17095 18275
rect 17218 18272 17224 18284
rect 17083 18244 17224 18272
rect 17083 18241 17095 18244
rect 17037 18235 17095 18241
rect 9456 18176 9674 18204
rect 14292 18176 14688 18204
rect 9456 18164 9462 18176
rect 9416 18136 9444 18164
rect 4488 18108 9444 18136
rect 9646 18136 9674 18176
rect 14734 18164 14740 18216
rect 14792 18164 14798 18216
rect 15562 18164 15568 18216
rect 15620 18204 15626 18216
rect 15841 18207 15899 18213
rect 15841 18204 15853 18207
rect 15620 18176 15853 18204
rect 15620 18164 15626 18176
rect 15841 18173 15853 18176
rect 15887 18173 15899 18207
rect 16500 18204 16528 18235
rect 17218 18232 17224 18244
rect 17276 18232 17282 18284
rect 17770 18232 17776 18284
rect 17828 18232 17834 18284
rect 18064 18281 18092 18312
rect 18049 18275 18107 18281
rect 18049 18241 18061 18275
rect 18095 18241 18107 18275
rect 18049 18235 18107 18241
rect 18230 18232 18236 18284
rect 18288 18232 18294 18284
rect 18524 18281 18552 18312
rect 18509 18275 18567 18281
rect 18509 18241 18521 18275
rect 18555 18241 18567 18275
rect 18509 18235 18567 18241
rect 19058 18232 19064 18284
rect 19116 18232 19122 18284
rect 19334 18232 19340 18284
rect 19392 18232 19398 18284
rect 15841 18167 15899 18173
rect 16224 18176 16528 18204
rect 16853 18207 16911 18213
rect 12434 18136 12440 18148
rect 9646 18108 12440 18136
rect 4488 18096 4494 18108
rect 12434 18096 12440 18108
rect 12492 18136 12498 18148
rect 14752 18136 14780 18164
rect 16224 18145 16252 18176
rect 16853 18173 16865 18207
rect 16899 18173 16911 18207
rect 16853 18167 16911 18173
rect 12492 18108 14780 18136
rect 16209 18139 16267 18145
rect 12492 18096 12498 18108
rect 16209 18105 16221 18139
rect 16255 18105 16267 18139
rect 16209 18099 16267 18105
rect 16482 18096 16488 18148
rect 16540 18136 16546 18148
rect 16868 18136 16896 18167
rect 17126 18164 17132 18216
rect 17184 18164 17190 18216
rect 18325 18207 18383 18213
rect 18325 18173 18337 18207
rect 18371 18204 18383 18207
rect 18966 18204 18972 18216
rect 18371 18176 18972 18204
rect 18371 18173 18383 18176
rect 18325 18167 18383 18173
rect 18966 18164 18972 18176
rect 19024 18164 19030 18216
rect 19076 18136 19104 18232
rect 19426 18164 19432 18216
rect 19484 18164 19490 18216
rect 19613 18207 19671 18213
rect 19613 18173 19625 18207
rect 19659 18204 19671 18207
rect 21560 18204 21588 18368
rect 23290 18300 23296 18352
rect 23348 18340 23354 18352
rect 27356 18340 27384 18368
rect 23348 18312 27384 18340
rect 23348 18300 23354 18312
rect 23750 18232 23756 18284
rect 23808 18272 23814 18284
rect 24394 18272 24400 18284
rect 23808 18244 24400 18272
rect 23808 18232 23814 18244
rect 24394 18232 24400 18244
rect 24452 18272 24458 18284
rect 27890 18272 27896 18284
rect 24452 18244 27896 18272
rect 24452 18232 24458 18244
rect 27890 18232 27896 18244
rect 27948 18232 27954 18284
rect 29840 18281 29868 18380
rect 30466 18368 30472 18380
rect 30524 18368 30530 18420
rect 31846 18408 31852 18420
rect 31312 18380 31852 18408
rect 30392 18312 30788 18340
rect 30392 18281 30420 18312
rect 30760 18284 30788 18312
rect 29825 18275 29883 18281
rect 29825 18241 29837 18275
rect 29871 18241 29883 18275
rect 30377 18275 30435 18281
rect 29825 18235 29883 18241
rect 29932 18244 30236 18272
rect 29932 18204 29960 18244
rect 19659 18176 21588 18204
rect 22066 18176 29960 18204
rect 19659 18173 19671 18176
rect 19613 18167 19671 18173
rect 16540 18108 19104 18136
rect 16540 18096 16546 18108
rect 20898 18096 20904 18148
rect 20956 18136 20962 18148
rect 21542 18136 21548 18148
rect 20956 18108 21548 18136
rect 20956 18096 20962 18108
rect 21542 18096 21548 18108
rect 21600 18096 21606 18148
rect 2498 18028 2504 18080
rect 2556 18028 2562 18080
rect 4706 18028 4712 18080
rect 4764 18028 4770 18080
rect 8754 18028 8760 18080
rect 8812 18028 8818 18080
rect 14090 18028 14096 18080
rect 14148 18028 14154 18080
rect 15746 18028 15752 18080
rect 15804 18028 15810 18080
rect 16301 18071 16359 18077
rect 16301 18037 16313 18071
rect 16347 18068 16359 18071
rect 16574 18068 16580 18080
rect 16347 18040 16580 18068
rect 16347 18037 16359 18040
rect 16301 18031 16359 18037
rect 16574 18028 16580 18040
rect 16632 18028 16638 18080
rect 16666 18028 16672 18080
rect 16724 18028 16730 18080
rect 17770 18028 17776 18080
rect 17828 18068 17834 18080
rect 18141 18071 18199 18077
rect 18141 18068 18153 18071
rect 17828 18040 18153 18068
rect 17828 18028 17834 18040
rect 18141 18037 18153 18040
rect 18187 18068 18199 18071
rect 18598 18068 18604 18080
rect 18187 18040 18604 18068
rect 18187 18037 18199 18040
rect 18141 18031 18199 18037
rect 18598 18028 18604 18040
rect 18656 18028 18662 18080
rect 18966 18028 18972 18080
rect 19024 18028 19030 18080
rect 19610 18028 19616 18080
rect 19668 18068 19674 18080
rect 22066 18068 22094 18176
rect 30006 18164 30012 18216
rect 30064 18164 30070 18216
rect 30098 18164 30104 18216
rect 30156 18164 30162 18216
rect 30208 18204 30236 18244
rect 30377 18241 30389 18275
rect 30423 18241 30435 18275
rect 30377 18235 30435 18241
rect 30650 18232 30656 18284
rect 30708 18232 30714 18284
rect 30742 18232 30748 18284
rect 30800 18232 30806 18284
rect 31312 18204 31340 18380
rect 31846 18368 31852 18380
rect 31904 18368 31910 18420
rect 32674 18368 32680 18420
rect 32732 18408 32738 18420
rect 32732 18380 34008 18408
rect 32732 18368 32738 18380
rect 33980 18352 34008 18380
rect 35158 18368 35164 18420
rect 35216 18368 35222 18420
rect 35529 18411 35587 18417
rect 35529 18377 35541 18411
rect 35575 18408 35587 18411
rect 38194 18408 38200 18420
rect 35575 18380 37780 18408
rect 35575 18377 35587 18380
rect 35529 18371 35587 18377
rect 33042 18340 33048 18352
rect 31404 18312 33048 18340
rect 31404 18284 31432 18312
rect 33042 18300 33048 18312
rect 33100 18300 33106 18352
rect 33502 18340 33508 18352
rect 33152 18312 33508 18340
rect 31386 18232 31392 18284
rect 31444 18232 31450 18284
rect 32766 18232 32772 18284
rect 32824 18272 32830 18284
rect 33152 18272 33180 18312
rect 33502 18300 33508 18312
rect 33560 18300 33566 18352
rect 33962 18300 33968 18352
rect 34020 18340 34026 18352
rect 35176 18340 35204 18368
rect 34020 18312 35204 18340
rect 34020 18300 34026 18312
rect 32824 18244 33180 18272
rect 32824 18232 32830 18244
rect 33410 18232 33416 18284
rect 33468 18272 33474 18284
rect 33468 18244 34100 18272
rect 33468 18232 33474 18244
rect 34072 18216 34100 18244
rect 34514 18232 34520 18284
rect 34572 18232 34578 18284
rect 34882 18232 34888 18284
rect 34940 18232 34946 18284
rect 35176 18281 35204 18312
rect 36170 18300 36176 18352
rect 36228 18340 36234 18352
rect 36228 18312 36860 18340
rect 36228 18300 36234 18312
rect 34978 18275 35036 18281
rect 34978 18241 34990 18275
rect 35024 18241 35036 18275
rect 34978 18235 35036 18241
rect 35161 18275 35219 18281
rect 35161 18241 35173 18275
rect 35207 18241 35219 18275
rect 35161 18235 35219 18241
rect 31481 18207 31539 18213
rect 31481 18204 31493 18207
rect 30208 18176 31493 18204
rect 31481 18173 31493 18176
rect 31527 18173 31539 18207
rect 31481 18167 31539 18173
rect 34054 18164 34060 18216
rect 34112 18164 34118 18216
rect 34532 18204 34560 18232
rect 34992 18204 35020 18235
rect 35250 18232 35256 18284
rect 35308 18232 35314 18284
rect 35350 18275 35408 18281
rect 35350 18241 35362 18275
rect 35396 18241 35408 18275
rect 35350 18235 35408 18241
rect 34532 18176 35020 18204
rect 23934 18096 23940 18148
rect 23992 18136 23998 18148
rect 24854 18136 24860 18148
rect 23992 18108 24860 18136
rect 23992 18096 23998 18108
rect 24854 18096 24860 18108
rect 24912 18136 24918 18148
rect 26142 18136 26148 18148
rect 24912 18108 26148 18136
rect 24912 18096 24918 18108
rect 26142 18096 26148 18108
rect 26200 18096 26206 18148
rect 29641 18139 29699 18145
rect 29641 18105 29653 18139
rect 29687 18136 29699 18139
rect 30374 18136 30380 18148
rect 29687 18108 30380 18136
rect 29687 18105 29699 18108
rect 29641 18099 29699 18105
rect 30374 18096 30380 18108
rect 30432 18096 30438 18148
rect 30558 18096 30564 18148
rect 30616 18136 30622 18148
rect 35360 18136 35388 18235
rect 35894 18232 35900 18284
rect 35952 18272 35958 18284
rect 36449 18275 36507 18281
rect 36449 18272 36461 18275
rect 35952 18244 36461 18272
rect 35952 18232 35958 18244
rect 36449 18241 36461 18244
rect 36495 18241 36507 18275
rect 36449 18235 36507 18241
rect 36538 18232 36544 18284
rect 36596 18232 36602 18284
rect 36725 18275 36783 18281
rect 36725 18241 36737 18275
rect 36771 18241 36783 18275
rect 36832 18272 36860 18312
rect 37642 18300 37648 18352
rect 37700 18300 37706 18352
rect 36832 18244 37688 18272
rect 36725 18235 36783 18241
rect 36556 18204 36584 18232
rect 36633 18207 36691 18213
rect 36633 18204 36645 18207
rect 36556 18176 36645 18204
rect 36633 18173 36645 18176
rect 36679 18173 36691 18207
rect 36633 18167 36691 18173
rect 30616 18108 31248 18136
rect 30616 18096 30622 18108
rect 19668 18040 22094 18068
rect 19668 18028 19674 18040
rect 29730 18028 29736 18080
rect 29788 18068 29794 18080
rect 30006 18068 30012 18080
rect 29788 18040 30012 18068
rect 29788 18028 29794 18040
rect 30006 18028 30012 18040
rect 30064 18028 30070 18080
rect 30193 18071 30251 18077
rect 30193 18037 30205 18071
rect 30239 18068 30251 18071
rect 30466 18068 30472 18080
rect 30239 18040 30472 18068
rect 30239 18037 30251 18040
rect 30193 18031 30251 18037
rect 30466 18028 30472 18040
rect 30524 18028 30530 18080
rect 30650 18028 30656 18080
rect 30708 18068 30714 18080
rect 31110 18068 31116 18080
rect 30708 18040 31116 18068
rect 30708 18028 30714 18040
rect 31110 18028 31116 18040
rect 31168 18028 31174 18080
rect 31220 18068 31248 18108
rect 34532 18108 35388 18136
rect 33042 18068 33048 18080
rect 31220 18040 33048 18068
rect 33042 18028 33048 18040
rect 33100 18028 33106 18080
rect 33870 18028 33876 18080
rect 33928 18068 33934 18080
rect 34532 18068 34560 18108
rect 36446 18096 36452 18148
rect 36504 18096 36510 18148
rect 36740 18136 36768 18235
rect 37660 18216 37688 18244
rect 37642 18164 37648 18216
rect 37700 18164 37706 18216
rect 37752 18204 37780 18380
rect 37844 18380 38200 18408
rect 37844 18281 37872 18380
rect 38194 18368 38200 18380
rect 38252 18368 38258 18420
rect 39945 18411 40003 18417
rect 39945 18377 39957 18411
rect 39991 18377 40003 18411
rect 39945 18371 40003 18377
rect 40865 18411 40923 18417
rect 40865 18377 40877 18411
rect 40911 18408 40923 18411
rect 41322 18408 41328 18420
rect 40911 18380 41328 18408
rect 40911 18377 40923 18380
rect 40865 18371 40923 18377
rect 39960 18340 39988 18371
rect 41322 18368 41328 18380
rect 41380 18368 41386 18420
rect 41506 18368 41512 18420
rect 41564 18368 41570 18420
rect 41524 18340 41552 18368
rect 39960 18312 41552 18340
rect 37829 18275 37887 18281
rect 37829 18241 37841 18275
rect 37875 18241 37887 18275
rect 37829 18235 37887 18241
rect 37918 18232 37924 18284
rect 37976 18232 37982 18284
rect 38102 18232 38108 18284
rect 38160 18272 38166 18284
rect 39485 18275 39543 18281
rect 39485 18272 39497 18275
rect 38160 18244 39497 18272
rect 38160 18232 38166 18244
rect 39485 18241 39497 18244
rect 39531 18241 39543 18275
rect 39485 18235 39543 18241
rect 39574 18232 39580 18284
rect 39632 18272 39638 18284
rect 39669 18275 39727 18281
rect 39669 18272 39681 18275
rect 39632 18244 39681 18272
rect 39632 18232 39638 18244
rect 39669 18241 39681 18244
rect 39715 18241 39727 18275
rect 39669 18235 39727 18241
rect 39761 18275 39819 18281
rect 39761 18241 39773 18275
rect 39807 18241 39819 18275
rect 39761 18235 39819 18241
rect 40037 18275 40095 18281
rect 40037 18241 40049 18275
rect 40083 18272 40095 18275
rect 40310 18272 40316 18284
rect 40083 18244 40316 18272
rect 40083 18241 40095 18244
rect 40037 18235 40095 18241
rect 39776 18204 39804 18235
rect 40310 18232 40316 18244
rect 40368 18232 40374 18284
rect 40494 18232 40500 18284
rect 40552 18232 40558 18284
rect 40681 18275 40739 18281
rect 40681 18241 40693 18275
rect 40727 18241 40739 18275
rect 40681 18235 40739 18241
rect 37752 18176 39804 18204
rect 39592 18148 39620 18176
rect 40126 18164 40132 18216
rect 40184 18204 40190 18216
rect 40696 18204 40724 18235
rect 40184 18176 40724 18204
rect 40184 18164 40190 18176
rect 41690 18164 41696 18216
rect 41748 18164 41754 18216
rect 36648 18108 36768 18136
rect 36909 18139 36967 18145
rect 33928 18040 34560 18068
rect 36464 18068 36492 18096
rect 36648 18080 36676 18108
rect 36909 18105 36921 18139
rect 36955 18136 36967 18139
rect 39022 18136 39028 18148
rect 36955 18108 39028 18136
rect 36955 18105 36967 18108
rect 36909 18099 36967 18105
rect 39022 18096 39028 18108
rect 39080 18096 39086 18148
rect 39574 18096 39580 18148
rect 39632 18096 39638 18148
rect 40405 18139 40463 18145
rect 40405 18105 40417 18139
rect 40451 18136 40463 18139
rect 41708 18136 41736 18164
rect 40451 18108 41736 18136
rect 40451 18105 40463 18108
rect 40405 18099 40463 18105
rect 36541 18071 36599 18077
rect 36541 18068 36553 18071
rect 36464 18040 36553 18068
rect 33928 18028 33934 18040
rect 36541 18037 36553 18040
rect 36587 18037 36599 18071
rect 36541 18031 36599 18037
rect 36630 18028 36636 18080
rect 36688 18028 36694 18080
rect 37090 18028 37096 18080
rect 37148 18068 37154 18080
rect 37645 18071 37703 18077
rect 37645 18068 37657 18071
rect 37148 18040 37657 18068
rect 37148 18028 37154 18040
rect 37645 18037 37657 18040
rect 37691 18037 37703 18071
rect 37645 18031 37703 18037
rect 38102 18028 38108 18080
rect 38160 18028 38166 18080
rect 39758 18028 39764 18080
rect 39816 18028 39822 18080
rect 40034 18028 40040 18080
rect 40092 18028 40098 18080
rect 1104 17978 41400 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 41400 17978
rect 1104 17904 41400 17926
rect 5994 17864 6000 17876
rect 1412 17836 6000 17864
rect 1412 17737 1440 17836
rect 5994 17824 6000 17836
rect 6052 17824 6058 17876
rect 6362 17824 6368 17876
rect 6420 17864 6426 17876
rect 6420 17836 11652 17864
rect 6420 17824 6426 17836
rect 3145 17799 3203 17805
rect 3145 17765 3157 17799
rect 3191 17796 3203 17799
rect 3418 17796 3424 17808
rect 3191 17768 3424 17796
rect 3191 17765 3203 17768
rect 3145 17759 3203 17765
rect 3418 17756 3424 17768
rect 3476 17756 3482 17808
rect 5626 17756 5632 17808
rect 5684 17796 5690 17808
rect 5684 17768 6040 17796
rect 5684 17756 5690 17768
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17697 1455 17731
rect 1397 17691 1455 17697
rect 4249 17731 4307 17737
rect 4249 17697 4261 17731
rect 4295 17728 4307 17731
rect 4614 17728 4620 17740
rect 4295 17700 4620 17728
rect 4295 17697 4307 17700
rect 4249 17691 4307 17697
rect 4614 17688 4620 17700
rect 4672 17688 4678 17740
rect 6012 17737 6040 17768
rect 6546 17756 6552 17808
rect 6604 17796 6610 17808
rect 9674 17796 9680 17808
rect 6604 17768 9680 17796
rect 6604 17756 6610 17768
rect 9674 17756 9680 17768
rect 9732 17756 9738 17808
rect 5997 17731 6055 17737
rect 5997 17697 6009 17731
rect 6043 17697 6055 17731
rect 5997 17691 6055 17697
rect 8018 17688 8024 17740
rect 8076 17728 8082 17740
rect 9950 17728 9956 17740
rect 8076 17700 9956 17728
rect 8076 17688 8082 17700
rect 9950 17688 9956 17700
rect 10008 17688 10014 17740
rect 5626 17620 5632 17672
rect 5684 17660 5690 17672
rect 6086 17660 6092 17672
rect 5684 17632 6092 17660
rect 5684 17620 5690 17632
rect 6086 17620 6092 17632
rect 6144 17620 6150 17672
rect 7929 17663 7987 17669
rect 7929 17629 7941 17663
rect 7975 17660 7987 17663
rect 8110 17660 8116 17672
rect 7975 17632 8116 17660
rect 7975 17629 7987 17632
rect 7929 17623 7987 17629
rect 8110 17620 8116 17632
rect 8168 17620 8174 17672
rect 8754 17620 8760 17672
rect 8812 17620 8818 17672
rect 9122 17620 9128 17672
rect 9180 17660 9186 17672
rect 9582 17660 9588 17672
rect 9180 17632 9588 17660
rect 9180 17620 9186 17632
rect 9582 17620 9588 17632
rect 9640 17620 9646 17672
rect 11624 17604 11652 17836
rect 13170 17824 13176 17876
rect 13228 17864 13234 17876
rect 13725 17867 13783 17873
rect 13725 17864 13737 17867
rect 13228 17836 13737 17864
rect 13228 17824 13234 17836
rect 13725 17833 13737 17836
rect 13771 17833 13783 17867
rect 13725 17827 13783 17833
rect 13906 17824 13912 17876
rect 13964 17864 13970 17876
rect 15286 17864 15292 17876
rect 13964 17836 15292 17864
rect 13964 17824 13970 17836
rect 15286 17824 15292 17836
rect 15344 17824 15350 17876
rect 15470 17824 15476 17876
rect 15528 17824 15534 17876
rect 15644 17867 15702 17873
rect 15644 17833 15656 17867
rect 15690 17864 15702 17867
rect 16666 17864 16672 17876
rect 15690 17836 16672 17864
rect 15690 17833 15702 17836
rect 15644 17827 15702 17833
rect 16666 17824 16672 17836
rect 16724 17824 16730 17876
rect 18322 17824 18328 17876
rect 18380 17864 18386 17876
rect 18874 17864 18880 17876
rect 18380 17836 18880 17864
rect 18380 17824 18386 17836
rect 18874 17824 18880 17836
rect 18932 17824 18938 17876
rect 19334 17824 19340 17876
rect 19392 17864 19398 17876
rect 19613 17867 19671 17873
rect 19613 17864 19625 17867
rect 19392 17836 19625 17864
rect 19392 17824 19398 17836
rect 19613 17833 19625 17836
rect 19659 17833 19671 17867
rect 19613 17827 19671 17833
rect 21269 17867 21327 17873
rect 21269 17833 21281 17867
rect 21315 17864 21327 17867
rect 21450 17864 21456 17876
rect 21315 17836 21456 17864
rect 21315 17833 21327 17836
rect 21269 17827 21327 17833
rect 21450 17824 21456 17836
rect 21508 17824 21514 17876
rect 24397 17867 24455 17873
rect 24397 17833 24409 17867
rect 24443 17864 24455 17867
rect 24486 17864 24492 17876
rect 24443 17836 24492 17864
rect 24443 17833 24455 17836
rect 24397 17827 24455 17833
rect 24486 17824 24492 17836
rect 24544 17824 24550 17876
rect 24578 17824 24584 17876
rect 24636 17864 24642 17876
rect 24762 17864 24768 17876
rect 24636 17836 24768 17864
rect 24636 17824 24642 17836
rect 24762 17824 24768 17836
rect 24820 17824 24826 17876
rect 27801 17867 27859 17873
rect 27801 17833 27813 17867
rect 27847 17864 27859 17867
rect 28077 17867 28135 17873
rect 28077 17864 28089 17867
rect 27847 17836 28089 17864
rect 27847 17833 27859 17836
rect 27801 17827 27859 17833
rect 28077 17833 28089 17836
rect 28123 17833 28135 17867
rect 28077 17827 28135 17833
rect 28445 17867 28503 17873
rect 28445 17833 28457 17867
rect 28491 17864 28503 17867
rect 29638 17864 29644 17876
rect 28491 17836 29644 17864
rect 28491 17833 28503 17836
rect 28445 17827 28503 17833
rect 29638 17824 29644 17836
rect 29696 17824 29702 17876
rect 35253 17867 35311 17873
rect 35253 17833 35265 17867
rect 35299 17864 35311 17867
rect 36630 17864 36636 17876
rect 35299 17836 36636 17864
rect 35299 17833 35311 17836
rect 35253 17827 35311 17833
rect 36630 17824 36636 17836
rect 36688 17864 36694 17876
rect 37461 17867 37519 17873
rect 37461 17864 37473 17867
rect 36688 17836 37473 17864
rect 36688 17824 36694 17836
rect 37461 17833 37473 17836
rect 37507 17833 37519 17867
rect 37461 17827 37519 17833
rect 37918 17824 37924 17876
rect 37976 17824 37982 17876
rect 38838 17824 38844 17876
rect 38896 17824 38902 17876
rect 39301 17867 39359 17873
rect 39301 17864 39313 17867
rect 38948 17836 39313 17864
rect 11701 17799 11759 17805
rect 11701 17765 11713 17799
rect 11747 17796 11759 17799
rect 12158 17796 12164 17808
rect 11747 17768 12164 17796
rect 11747 17765 11759 17768
rect 11701 17759 11759 17765
rect 12158 17756 12164 17768
rect 12216 17796 12222 17808
rect 13357 17799 13415 17805
rect 12216 17768 12664 17796
rect 12216 17756 12222 17768
rect 12434 17688 12440 17740
rect 12492 17688 12498 17740
rect 12636 17737 12664 17768
rect 13357 17765 13369 17799
rect 13403 17796 13415 17799
rect 15488 17796 15516 17824
rect 13403 17768 15516 17796
rect 13403 17765 13415 17768
rect 13357 17759 13415 17765
rect 18046 17756 18052 17808
rect 18104 17796 18110 17808
rect 18690 17796 18696 17808
rect 18104 17768 18696 17796
rect 18104 17756 18110 17768
rect 18690 17756 18696 17768
rect 18748 17796 18754 17808
rect 19521 17799 19579 17805
rect 19521 17796 19533 17799
rect 18748 17768 19533 17796
rect 18748 17756 18754 17768
rect 19521 17765 19533 17768
rect 19567 17765 19579 17799
rect 19521 17759 19579 17765
rect 20622 17756 20628 17808
rect 20680 17796 20686 17808
rect 24596 17796 24624 17824
rect 20680 17768 24624 17796
rect 24688 17768 25544 17796
rect 20680 17756 20686 17768
rect 12621 17731 12679 17737
rect 12621 17697 12633 17731
rect 12667 17697 12679 17731
rect 12621 17691 12679 17697
rect 13265 17731 13323 17737
rect 13265 17697 13277 17731
rect 13311 17697 13323 17731
rect 13265 17691 13323 17697
rect 13817 17731 13875 17737
rect 13817 17697 13829 17731
rect 13863 17728 13875 17731
rect 14182 17728 14188 17740
rect 13863 17700 14188 17728
rect 13863 17697 13875 17700
rect 13817 17691 13875 17697
rect 12253 17663 12311 17669
rect 12253 17629 12265 17663
rect 12299 17660 12311 17663
rect 12526 17660 12532 17672
rect 12299 17632 12532 17660
rect 12299 17629 12311 17632
rect 12253 17623 12311 17629
rect 12526 17620 12532 17632
rect 12584 17620 12590 17672
rect 13280 17660 13308 17691
rect 14182 17688 14188 17700
rect 14240 17688 14246 17740
rect 15381 17731 15439 17737
rect 15381 17697 15393 17731
rect 15427 17728 15439 17731
rect 17862 17728 17868 17740
rect 15427 17700 17868 17728
rect 15427 17697 15439 17700
rect 15381 17691 15439 17697
rect 17862 17688 17868 17700
rect 17920 17688 17926 17740
rect 18322 17688 18328 17740
rect 18380 17688 18386 17740
rect 19242 17688 19248 17740
rect 19300 17728 19306 17740
rect 19300 17700 19472 17728
rect 19300 17688 19306 17700
rect 12820 17632 13308 17660
rect 1670 17552 1676 17604
rect 1728 17552 1734 17604
rect 3418 17592 3424 17604
rect 2898 17564 3424 17592
rect 3418 17552 3424 17564
rect 3476 17552 3482 17604
rect 4525 17595 4583 17601
rect 4525 17561 4537 17595
rect 4571 17561 4583 17595
rect 4525 17555 4583 17561
rect 4540 17524 4568 17555
rect 10226 17552 10232 17604
rect 10284 17552 10290 17604
rect 11238 17552 11244 17604
rect 11296 17552 11302 17604
rect 11606 17552 11612 17604
rect 11664 17592 11670 17604
rect 12161 17595 12219 17601
rect 11664 17564 11928 17592
rect 11664 17552 11670 17564
rect 4706 17524 4712 17536
rect 4540 17496 4712 17524
rect 4706 17484 4712 17496
rect 4764 17484 4770 17536
rect 8478 17484 8484 17536
rect 8536 17484 8542 17536
rect 8570 17484 8576 17536
rect 8628 17484 8634 17536
rect 11790 17484 11796 17536
rect 11848 17484 11854 17536
rect 11900 17524 11928 17564
rect 12161 17561 12173 17595
rect 12207 17592 12219 17595
rect 12820 17592 12848 17632
rect 13538 17620 13544 17672
rect 13596 17620 13602 17672
rect 14090 17620 14096 17672
rect 14148 17660 14154 17672
rect 14277 17663 14335 17669
rect 14277 17660 14289 17663
rect 14148 17632 14289 17660
rect 14148 17620 14154 17632
rect 14277 17629 14289 17632
rect 14323 17629 14335 17663
rect 14277 17623 14335 17629
rect 15286 17620 15292 17672
rect 15344 17660 15350 17672
rect 15344 17632 15424 17660
rect 15344 17620 15350 17632
rect 15396 17592 15424 17632
rect 17218 17620 17224 17672
rect 17276 17660 17282 17672
rect 17405 17663 17463 17669
rect 17405 17660 17417 17663
rect 17276 17632 17417 17660
rect 17276 17620 17282 17632
rect 17405 17629 17417 17632
rect 17451 17629 17463 17663
rect 17405 17623 17463 17629
rect 17770 17620 17776 17672
rect 17828 17620 17834 17672
rect 18046 17620 18052 17672
rect 18104 17620 18110 17672
rect 18417 17663 18475 17669
rect 18417 17660 18429 17663
rect 18340 17632 18429 17660
rect 12207 17564 12848 17592
rect 13280 17564 15332 17592
rect 15396 17564 16146 17592
rect 12207 17561 12219 17564
rect 12161 17555 12219 17561
rect 13280 17524 13308 17564
rect 15304 17536 15332 17564
rect 11900 17496 13308 17524
rect 14090 17484 14096 17536
rect 14148 17484 14154 17536
rect 15286 17484 15292 17536
rect 15344 17484 15350 17536
rect 16040 17524 16068 17564
rect 17586 17552 17592 17604
rect 17644 17552 17650 17604
rect 16666 17524 16672 17536
rect 16040 17496 16672 17524
rect 16666 17484 16672 17496
rect 16724 17484 16730 17536
rect 17954 17484 17960 17536
rect 18012 17484 18018 17536
rect 18141 17527 18199 17533
rect 18141 17493 18153 17527
rect 18187 17524 18199 17527
rect 18230 17524 18236 17536
rect 18187 17496 18236 17524
rect 18187 17493 18199 17496
rect 18141 17487 18199 17493
rect 18230 17484 18236 17496
rect 18288 17484 18294 17536
rect 18340 17524 18368 17632
rect 18417 17629 18429 17632
rect 18463 17629 18475 17663
rect 18417 17623 18475 17629
rect 18506 17620 18512 17672
rect 18564 17620 18570 17672
rect 18601 17663 18659 17669
rect 18601 17629 18613 17663
rect 18647 17660 18659 17663
rect 18874 17660 18880 17672
rect 18647 17632 18880 17660
rect 18647 17629 18659 17632
rect 18601 17623 18659 17629
rect 18874 17620 18880 17632
rect 18932 17620 18938 17672
rect 19150 17620 19156 17672
rect 19208 17660 19214 17672
rect 19337 17663 19395 17669
rect 19337 17660 19349 17663
rect 19208 17632 19349 17660
rect 19208 17620 19214 17632
rect 19337 17629 19349 17632
rect 19383 17629 19395 17663
rect 19444 17660 19472 17700
rect 19610 17688 19616 17740
rect 19668 17688 19674 17740
rect 19904 17700 22048 17728
rect 19797 17663 19855 17669
rect 19797 17660 19809 17663
rect 19444 17632 19809 17660
rect 19337 17623 19395 17629
rect 19797 17629 19809 17632
rect 19843 17629 19855 17663
rect 19797 17623 19855 17629
rect 19245 17595 19303 17601
rect 19245 17592 19257 17595
rect 18616 17564 19257 17592
rect 18616 17524 18644 17564
rect 19245 17561 19257 17564
rect 19291 17592 19303 17595
rect 19904 17592 19932 17700
rect 22020 17672 22048 17700
rect 23566 17688 23572 17740
rect 23624 17728 23630 17740
rect 23624 17700 23796 17728
rect 23624 17688 23630 17700
rect 23768 17672 23796 17700
rect 24118 17688 24124 17740
rect 24176 17688 24182 17740
rect 20073 17663 20131 17669
rect 20073 17629 20085 17663
rect 20119 17629 20131 17663
rect 20073 17623 20131 17629
rect 21085 17663 21143 17669
rect 21085 17629 21097 17663
rect 21131 17660 21143 17663
rect 21269 17663 21327 17669
rect 21131 17632 21220 17660
rect 21131 17629 21143 17632
rect 21085 17623 21143 17629
rect 19291 17564 19932 17592
rect 19291 17561 19303 17564
rect 19245 17555 19303 17561
rect 18340 17496 18644 17524
rect 18690 17484 18696 17536
rect 18748 17524 18754 17536
rect 20088 17524 20116 17623
rect 21192 17604 21220 17632
rect 21269 17629 21281 17663
rect 21315 17660 21327 17663
rect 21450 17660 21456 17672
rect 21315 17632 21456 17660
rect 21315 17629 21327 17632
rect 21269 17623 21327 17629
rect 21450 17620 21456 17632
rect 21508 17620 21514 17672
rect 22002 17620 22008 17672
rect 22060 17620 22066 17672
rect 23750 17620 23756 17672
rect 23808 17620 23814 17672
rect 24136 17660 24164 17688
rect 24688 17669 24716 17768
rect 25041 17731 25099 17737
rect 25041 17697 25053 17731
rect 25087 17728 25099 17731
rect 25222 17728 25228 17740
rect 25087 17700 25228 17728
rect 25087 17697 25099 17700
rect 25041 17691 25099 17697
rect 25222 17688 25228 17700
rect 25280 17688 25286 17740
rect 25516 17672 25544 17768
rect 26050 17756 26056 17808
rect 26108 17796 26114 17808
rect 26108 17768 29592 17796
rect 26108 17756 26114 17768
rect 26326 17728 26332 17740
rect 25608 17700 26332 17728
rect 24946 17669 24952 17672
rect 24581 17663 24639 17669
rect 24581 17660 24593 17663
rect 24136 17632 24593 17660
rect 24581 17629 24593 17632
rect 24627 17629 24639 17663
rect 24581 17623 24639 17629
rect 24673 17663 24731 17669
rect 24673 17629 24685 17663
rect 24719 17629 24731 17663
rect 24673 17623 24731 17629
rect 24903 17663 24952 17669
rect 24903 17629 24915 17663
rect 24949 17629 24952 17663
rect 24903 17623 24952 17629
rect 24946 17620 24952 17623
rect 25004 17620 25010 17672
rect 25498 17620 25504 17672
rect 25556 17620 25562 17672
rect 21174 17552 21180 17604
rect 21232 17552 21238 17604
rect 22830 17552 22836 17604
rect 22888 17592 22894 17604
rect 24765 17595 24823 17601
rect 24765 17592 24777 17595
rect 22888 17564 24777 17592
rect 22888 17552 22894 17564
rect 24765 17561 24777 17564
rect 24811 17592 24823 17595
rect 25608 17592 25636 17700
rect 26326 17688 26332 17700
rect 26384 17688 26390 17740
rect 27706 17688 27712 17740
rect 27764 17688 27770 17740
rect 28994 17688 29000 17740
rect 29052 17728 29058 17740
rect 29270 17728 29276 17740
rect 29052 17700 29276 17728
rect 29052 17688 29058 17700
rect 29270 17688 29276 17700
rect 29328 17688 29334 17740
rect 29564 17737 29592 17768
rect 31570 17756 31576 17808
rect 31628 17796 31634 17808
rect 32582 17796 32588 17808
rect 31628 17768 32588 17796
rect 31628 17756 31634 17768
rect 32582 17756 32588 17768
rect 32640 17756 32646 17808
rect 33778 17756 33784 17808
rect 33836 17796 33842 17808
rect 33836 17768 34100 17796
rect 33836 17756 33842 17768
rect 29549 17731 29607 17737
rect 29549 17697 29561 17731
rect 29595 17697 29607 17731
rect 29549 17691 29607 17697
rect 27798 17620 27804 17672
rect 27856 17620 27862 17672
rect 28258 17620 28264 17672
rect 28316 17620 28322 17672
rect 28534 17620 28540 17672
rect 28592 17620 28598 17672
rect 28721 17663 28779 17669
rect 28721 17629 28733 17663
rect 28767 17660 28779 17663
rect 30101 17663 30159 17669
rect 28767 17632 28994 17660
rect 28767 17629 28779 17632
rect 28721 17623 28779 17629
rect 24811 17564 25636 17592
rect 24811 17561 24823 17564
rect 24765 17555 24823 17561
rect 27522 17552 27528 17604
rect 27580 17552 27586 17604
rect 18748 17496 20116 17524
rect 18748 17484 18754 17496
rect 21266 17484 21272 17536
rect 21324 17524 21330 17536
rect 21453 17527 21511 17533
rect 21453 17524 21465 17527
rect 21324 17496 21465 17524
rect 21324 17484 21330 17496
rect 21453 17493 21465 17496
rect 21499 17493 21511 17527
rect 21453 17487 21511 17493
rect 23474 17484 23480 17536
rect 23532 17524 23538 17536
rect 24118 17524 24124 17536
rect 23532 17496 24124 17524
rect 23532 17484 23538 17496
rect 24118 17484 24124 17496
rect 24176 17484 24182 17536
rect 26142 17484 26148 17536
rect 26200 17524 26206 17536
rect 27985 17527 28043 17533
rect 27985 17524 27997 17527
rect 26200 17496 27997 17524
rect 26200 17484 26206 17496
rect 27985 17493 27997 17496
rect 28031 17493 28043 17527
rect 28966 17524 28994 17632
rect 30101 17629 30113 17663
rect 30147 17629 30159 17663
rect 30101 17623 30159 17629
rect 29089 17595 29147 17601
rect 29089 17561 29101 17595
rect 29135 17592 29147 17595
rect 29546 17592 29552 17604
rect 29135 17564 29552 17592
rect 29135 17561 29147 17564
rect 29089 17555 29147 17561
rect 29546 17552 29552 17564
rect 29604 17552 29610 17604
rect 29638 17552 29644 17604
rect 29696 17592 29702 17604
rect 30116 17592 30144 17623
rect 30374 17620 30380 17672
rect 30432 17620 30438 17672
rect 30466 17620 30472 17672
rect 30524 17660 30530 17672
rect 30561 17663 30619 17669
rect 30561 17660 30573 17663
rect 30524 17632 30573 17660
rect 30524 17620 30530 17632
rect 30561 17629 30573 17632
rect 30607 17629 30619 17663
rect 30561 17623 30619 17629
rect 31018 17620 31024 17672
rect 31076 17660 31082 17672
rect 31389 17663 31447 17669
rect 31389 17660 31401 17663
rect 31076 17632 31401 17660
rect 31076 17620 31082 17632
rect 31389 17629 31401 17632
rect 31435 17660 31447 17663
rect 31754 17660 31760 17672
rect 31435 17632 31760 17660
rect 31435 17629 31447 17632
rect 31389 17623 31447 17629
rect 31754 17620 31760 17632
rect 31812 17620 31818 17672
rect 33686 17620 33692 17672
rect 33744 17620 33750 17672
rect 33778 17620 33784 17672
rect 33836 17660 33842 17672
rect 34072 17669 34100 17768
rect 34238 17756 34244 17808
rect 34296 17756 34302 17808
rect 34333 17799 34391 17805
rect 34333 17765 34345 17799
rect 34379 17796 34391 17799
rect 36354 17796 36360 17808
rect 34379 17768 36360 17796
rect 34379 17765 34391 17768
rect 34333 17759 34391 17765
rect 36354 17756 36360 17768
rect 36412 17796 36418 17808
rect 38948 17796 38976 17836
rect 39301 17833 39313 17836
rect 39347 17833 39359 17867
rect 39301 17827 39359 17833
rect 39666 17824 39672 17876
rect 39724 17824 39730 17876
rect 36412 17768 38976 17796
rect 39117 17799 39175 17805
rect 36412 17756 36418 17768
rect 39117 17765 39129 17799
rect 39163 17796 39175 17799
rect 40126 17796 40132 17808
rect 39163 17768 40132 17796
rect 39163 17765 39175 17768
rect 39117 17759 39175 17765
rect 40126 17756 40132 17768
rect 40184 17756 40190 17808
rect 34256 17728 34284 17756
rect 34256 17700 35572 17728
rect 34054 17663 34112 17669
rect 33836 17632 33881 17660
rect 33836 17620 33842 17632
rect 34054 17629 34066 17663
rect 34100 17629 34112 17663
rect 34054 17623 34112 17629
rect 34154 17663 34212 17669
rect 34154 17629 34166 17663
rect 34200 17660 34212 17663
rect 34200 17629 34216 17660
rect 34154 17623 34216 17629
rect 29696 17564 30144 17592
rect 29696 17552 29702 17564
rect 33594 17552 33600 17604
rect 33652 17592 33658 17604
rect 33965 17595 34023 17601
rect 33965 17592 33977 17595
rect 33652 17564 33977 17592
rect 33652 17552 33658 17564
rect 33965 17561 33977 17564
rect 34011 17561 34023 17595
rect 33965 17555 34023 17561
rect 33502 17524 33508 17536
rect 28966 17496 33508 17524
rect 27985 17487 28043 17493
rect 33502 17484 33508 17496
rect 33560 17484 33566 17536
rect 33870 17484 33876 17536
rect 33928 17524 33934 17536
rect 34188 17524 34216 17623
rect 34330 17620 34336 17672
rect 34388 17620 34394 17672
rect 35434 17620 35440 17672
rect 35492 17620 35498 17672
rect 35544 17669 35572 17700
rect 35820 17700 36952 17728
rect 35820 17669 35848 17700
rect 36924 17672 36952 17700
rect 37550 17688 37556 17740
rect 37608 17688 37614 17740
rect 38010 17688 38016 17740
rect 38068 17728 38074 17740
rect 38749 17731 38807 17737
rect 38749 17728 38761 17731
rect 38068 17700 38761 17728
rect 38068 17688 38074 17700
rect 38749 17697 38761 17700
rect 38795 17697 38807 17731
rect 40402 17728 40408 17740
rect 38749 17691 38807 17697
rect 39132 17700 40408 17728
rect 35529 17663 35587 17669
rect 35529 17629 35541 17663
rect 35575 17629 35587 17663
rect 35529 17623 35587 17629
rect 35805 17663 35863 17669
rect 35805 17629 35817 17663
rect 35851 17629 35863 17663
rect 35805 17623 35863 17629
rect 35897 17663 35955 17669
rect 35897 17629 35909 17663
rect 35943 17629 35955 17663
rect 35897 17623 35955 17629
rect 34348 17592 34376 17620
rect 35342 17592 35348 17604
rect 34348 17564 35348 17592
rect 35342 17552 35348 17564
rect 35400 17592 35406 17604
rect 35621 17595 35679 17601
rect 35621 17592 35633 17595
rect 35400 17564 35633 17592
rect 35400 17552 35406 17564
rect 35621 17561 35633 17564
rect 35667 17561 35679 17595
rect 35820 17592 35848 17623
rect 35621 17555 35679 17561
rect 35728 17564 35848 17592
rect 35728 17536 35756 17564
rect 33928 17496 34216 17524
rect 33928 17484 33934 17496
rect 35710 17484 35716 17536
rect 35768 17484 35774 17536
rect 35802 17484 35808 17536
rect 35860 17524 35866 17536
rect 35912 17524 35940 17623
rect 36906 17620 36912 17672
rect 36964 17620 36970 17672
rect 37734 17620 37740 17672
rect 37792 17660 37798 17672
rect 38933 17663 38991 17669
rect 38933 17660 38945 17663
rect 37792 17632 38945 17660
rect 37792 17620 37798 17632
rect 38933 17629 38945 17632
rect 38979 17629 38991 17663
rect 38933 17623 38991 17629
rect 39022 17620 39028 17672
rect 39080 17620 39086 17672
rect 37461 17595 37519 17601
rect 37461 17561 37473 17595
rect 37507 17592 37519 17595
rect 38194 17592 38200 17604
rect 37507 17564 38200 17592
rect 37507 17561 37519 17564
rect 37461 17555 37519 17561
rect 38194 17552 38200 17564
rect 38252 17552 38258 17604
rect 38657 17595 38715 17601
rect 38657 17561 38669 17595
rect 38703 17592 38715 17595
rect 39040 17592 39068 17620
rect 38703 17564 39068 17592
rect 38703 17561 38715 17564
rect 38657 17555 38715 17561
rect 35860 17496 35940 17524
rect 35860 17484 35866 17496
rect 36538 17484 36544 17536
rect 36596 17524 36602 17536
rect 39132 17524 39160 17700
rect 40402 17688 40408 17700
rect 40460 17688 40466 17740
rect 39301 17663 39359 17669
rect 39301 17629 39313 17663
rect 39347 17660 39359 17663
rect 39485 17663 39543 17669
rect 39347 17632 39436 17660
rect 39347 17629 39359 17632
rect 39301 17623 39359 17629
rect 39408 17536 39436 17632
rect 39485 17629 39497 17663
rect 39531 17660 39543 17663
rect 39574 17660 39580 17672
rect 39531 17632 39580 17660
rect 39531 17629 39543 17632
rect 39485 17623 39543 17629
rect 39574 17620 39580 17632
rect 39632 17620 39638 17672
rect 36596 17496 39160 17524
rect 36596 17484 36602 17496
rect 39390 17484 39396 17536
rect 39448 17484 39454 17536
rect 40034 17484 40040 17536
rect 40092 17524 40098 17536
rect 41598 17524 41604 17536
rect 40092 17496 41604 17524
rect 40092 17484 40098 17496
rect 41598 17484 41604 17496
rect 41656 17484 41662 17536
rect 1104 17434 41400 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 41400 17434
rect 1104 17360 41400 17382
rect 1670 17280 1676 17332
rect 1728 17320 1734 17332
rect 1857 17323 1915 17329
rect 1857 17320 1869 17323
rect 1728 17292 1869 17320
rect 1728 17280 1734 17292
rect 1857 17289 1869 17292
rect 1903 17289 1915 17323
rect 1857 17283 1915 17289
rect 2498 17280 2504 17332
rect 2556 17280 2562 17332
rect 7469 17323 7527 17329
rect 7469 17289 7481 17323
rect 7515 17320 7527 17323
rect 8478 17320 8484 17332
rect 7515 17292 8484 17320
rect 7515 17289 7527 17292
rect 7469 17283 7527 17289
rect 8478 17280 8484 17292
rect 8536 17280 8542 17332
rect 8570 17280 8576 17332
rect 8628 17280 8634 17332
rect 9766 17280 9772 17332
rect 9824 17280 9830 17332
rect 10226 17280 10232 17332
rect 10284 17320 10290 17332
rect 10505 17323 10563 17329
rect 10505 17320 10517 17323
rect 10284 17292 10517 17320
rect 10284 17280 10290 17292
rect 10505 17289 10517 17292
rect 10551 17289 10563 17323
rect 10505 17283 10563 17289
rect 11517 17323 11575 17329
rect 11517 17289 11529 17323
rect 11563 17289 11575 17323
rect 11517 17283 11575 17289
rect 2516 17252 2544 17280
rect 2056 17224 2544 17252
rect 2056 17193 2084 17224
rect 2958 17212 2964 17264
rect 3016 17252 3022 17264
rect 3237 17255 3295 17261
rect 3237 17252 3249 17255
rect 3016 17224 3249 17252
rect 3016 17212 3022 17224
rect 3237 17221 3249 17224
rect 3283 17252 3295 17255
rect 3970 17252 3976 17264
rect 3283 17224 3976 17252
rect 3283 17221 3295 17224
rect 3237 17215 3295 17221
rect 3970 17212 3976 17224
rect 4028 17212 4034 17264
rect 8297 17255 8355 17261
rect 6012 17224 7236 17252
rect 6012 17196 6040 17224
rect 2041 17187 2099 17193
rect 2041 17153 2053 17187
rect 2087 17153 2099 17187
rect 2041 17147 2099 17153
rect 2409 17187 2467 17193
rect 2409 17153 2421 17187
rect 2455 17184 2467 17187
rect 3145 17187 3203 17193
rect 2455 17156 2820 17184
rect 2455 17153 2467 17156
rect 2409 17147 2467 17153
rect 2792 17057 2820 17156
rect 3145 17153 3157 17187
rect 3191 17184 3203 17187
rect 4249 17187 4307 17193
rect 4249 17184 4261 17187
rect 3191 17156 4261 17184
rect 3191 17153 3203 17156
rect 3145 17147 3203 17153
rect 4249 17153 4261 17156
rect 4295 17153 4307 17187
rect 4249 17147 4307 17153
rect 5994 17144 6000 17196
rect 6052 17144 6058 17196
rect 6917 17187 6975 17193
rect 6917 17153 6929 17187
rect 6963 17184 6975 17187
rect 7208 17184 7236 17224
rect 8297 17221 8309 17255
rect 8343 17252 8355 17255
rect 8588 17252 8616 17280
rect 8343 17224 8616 17252
rect 8343 17221 8355 17224
rect 8297 17215 8355 17221
rect 9306 17212 9312 17264
rect 9364 17212 9370 17264
rect 8018 17184 8024 17196
rect 6963 17156 7144 17184
rect 7208 17156 8024 17184
rect 6963 17153 6975 17156
rect 6917 17147 6975 17153
rect 3329 17119 3387 17125
rect 3329 17085 3341 17119
rect 3375 17085 3387 17119
rect 3329 17079 3387 17085
rect 3697 17119 3755 17125
rect 3697 17085 3709 17119
rect 3743 17116 3755 17119
rect 3878 17116 3884 17128
rect 3743 17088 3884 17116
rect 3743 17085 3755 17088
rect 3697 17079 3755 17085
rect 2777 17051 2835 17057
rect 2777 17017 2789 17051
rect 2823 17017 2835 17051
rect 2777 17011 2835 17017
rect 3344 16992 3372 17079
rect 3878 17076 3884 17088
rect 3936 17076 3942 17128
rect 7116 17057 7144 17156
rect 8018 17144 8024 17156
rect 8076 17144 8082 17196
rect 9674 17144 9680 17196
rect 9732 17184 9738 17196
rect 10689 17187 10747 17193
rect 9732 17156 9904 17184
rect 9732 17144 9738 17156
rect 7558 17076 7564 17128
rect 7616 17076 7622 17128
rect 7745 17119 7803 17125
rect 7745 17085 7757 17119
rect 7791 17116 7803 17119
rect 7791 17088 9720 17116
rect 7791 17085 7803 17088
rect 7745 17079 7803 17085
rect 7101 17051 7159 17057
rect 7101 17017 7113 17051
rect 7147 17017 7159 17051
rect 7101 17011 7159 17017
rect 2130 16940 2136 16992
rect 2188 16980 2194 16992
rect 2225 16983 2283 16989
rect 2225 16980 2237 16983
rect 2188 16952 2237 16980
rect 2188 16940 2194 16952
rect 2225 16949 2237 16952
rect 2271 16949 2283 16983
rect 2225 16943 2283 16949
rect 3326 16940 3332 16992
rect 3384 16980 3390 16992
rect 4062 16980 4068 16992
rect 3384 16952 4068 16980
rect 3384 16940 3390 16952
rect 4062 16940 4068 16952
rect 4120 16940 4126 16992
rect 6638 16940 6644 16992
rect 6696 16980 6702 16992
rect 6733 16983 6791 16989
rect 6733 16980 6745 16983
rect 6696 16952 6745 16980
rect 6696 16940 6702 16952
rect 6733 16949 6745 16952
rect 6779 16949 6791 16983
rect 6733 16943 6791 16949
rect 6822 16940 6828 16992
rect 6880 16980 6886 16992
rect 7760 16980 7788 17079
rect 9692 16992 9720 17088
rect 9876 17048 9904 17156
rect 10689 17153 10701 17187
rect 10735 17153 10747 17187
rect 10689 17147 10747 17153
rect 11149 17187 11207 17193
rect 11149 17153 11161 17187
rect 11195 17184 11207 17187
rect 11532 17184 11560 17283
rect 11790 17280 11796 17332
rect 11848 17280 11854 17332
rect 11977 17323 12035 17329
rect 11977 17289 11989 17323
rect 12023 17320 12035 17323
rect 12526 17320 12532 17332
rect 12023 17292 12532 17320
rect 12023 17289 12035 17292
rect 11977 17283 12035 17289
rect 12526 17280 12532 17292
rect 12584 17280 12590 17332
rect 14090 17320 14096 17332
rect 13464 17292 14096 17320
rect 11195 17156 11560 17184
rect 11195 17153 11207 17156
rect 11149 17147 11207 17153
rect 10704 17116 10732 17147
rect 11808 17116 11836 17280
rect 13464 17261 13492 17292
rect 14090 17280 14096 17292
rect 14148 17280 14154 17332
rect 14458 17280 14464 17332
rect 14516 17320 14522 17332
rect 14921 17323 14979 17329
rect 14921 17320 14933 17323
rect 14516 17292 14933 17320
rect 14516 17280 14522 17292
rect 14921 17289 14933 17292
rect 14967 17289 14979 17323
rect 14921 17283 14979 17289
rect 16298 17280 16304 17332
rect 16356 17280 16362 17332
rect 16574 17280 16580 17332
rect 16632 17320 16638 17332
rect 17037 17323 17095 17329
rect 17037 17320 17049 17323
rect 16632 17292 17049 17320
rect 16632 17280 16638 17292
rect 17037 17289 17049 17292
rect 17083 17289 17095 17323
rect 18690 17320 18696 17332
rect 17037 17283 17095 17289
rect 17512 17292 18000 17320
rect 13449 17255 13507 17261
rect 13449 17221 13461 17255
rect 13495 17221 13507 17255
rect 13449 17215 13507 17221
rect 13722 17212 13728 17264
rect 13780 17252 13786 17264
rect 13906 17252 13912 17264
rect 13780 17224 13912 17252
rect 13780 17212 13786 17224
rect 13906 17212 13912 17224
rect 13964 17212 13970 17264
rect 15841 17255 15899 17261
rect 15841 17221 15853 17255
rect 15887 17252 15899 17255
rect 16482 17252 16488 17264
rect 15887 17224 16488 17252
rect 15887 17221 15899 17224
rect 15841 17215 15899 17221
rect 16482 17212 16488 17224
rect 16540 17212 16546 17264
rect 16666 17212 16672 17264
rect 16724 17252 16730 17264
rect 17512 17252 17540 17292
rect 17862 17252 17868 17264
rect 16724 17224 17540 17252
rect 17604 17224 17868 17252
rect 16724 17212 16730 17224
rect 11885 17187 11943 17193
rect 11885 17153 11897 17187
rect 11931 17184 11943 17187
rect 12989 17187 13047 17193
rect 12989 17184 13001 17187
rect 11931 17156 13001 17184
rect 11931 17153 11943 17156
rect 11885 17147 11943 17153
rect 12989 17153 13001 17156
rect 13035 17153 13047 17187
rect 12989 17147 13047 17153
rect 15286 17144 15292 17196
rect 15344 17184 15350 17196
rect 16117 17187 16175 17193
rect 16117 17184 16129 17187
rect 15344 17156 16129 17184
rect 15344 17144 15350 17156
rect 16117 17153 16129 17156
rect 16163 17184 16175 17187
rect 16390 17184 16396 17196
rect 16163 17156 16396 17184
rect 16163 17153 16175 17156
rect 16117 17147 16175 17153
rect 16390 17144 16396 17156
rect 16448 17144 16454 17196
rect 17604 17193 17632 17224
rect 17862 17212 17868 17224
rect 17920 17212 17926 17264
rect 17972 17252 18000 17292
rect 18248 17292 18696 17320
rect 18248 17252 18276 17292
rect 18690 17280 18696 17292
rect 18748 17280 18754 17332
rect 21637 17323 21695 17329
rect 20364 17292 21404 17320
rect 17972 17224 18354 17252
rect 19334 17212 19340 17264
rect 19392 17252 19398 17264
rect 19613 17255 19671 17261
rect 19613 17252 19625 17255
rect 19392 17224 19625 17252
rect 19392 17212 19398 17224
rect 19613 17221 19625 17224
rect 19659 17221 19671 17255
rect 20364 17252 20392 17292
rect 19613 17215 19671 17221
rect 19720 17224 20392 17252
rect 17589 17187 17647 17193
rect 17589 17153 17601 17187
rect 17635 17153 17647 17187
rect 17589 17147 17647 17153
rect 10704 17088 11836 17116
rect 12066 17076 12072 17128
rect 12124 17076 12130 17128
rect 12250 17076 12256 17128
rect 12308 17116 12314 17128
rect 12345 17119 12403 17125
rect 12345 17116 12357 17119
rect 12308 17088 12357 17116
rect 12308 17076 12314 17088
rect 12345 17085 12357 17088
rect 12391 17085 12403 17119
rect 12345 17079 12403 17085
rect 13170 17076 13176 17128
rect 13228 17076 13234 17128
rect 15933 17119 15991 17125
rect 15933 17116 15945 17119
rect 13280 17088 15945 17116
rect 10686 17048 10692 17060
rect 9876 17020 10692 17048
rect 10686 17008 10692 17020
rect 10744 17048 10750 17060
rect 13280 17048 13308 17088
rect 15933 17085 15945 17088
rect 15979 17085 15991 17119
rect 15933 17079 15991 17085
rect 17129 17119 17187 17125
rect 17129 17085 17141 17119
rect 17175 17085 17187 17119
rect 17129 17079 17187 17085
rect 10744 17020 13308 17048
rect 17144 17048 17172 17079
rect 17218 17076 17224 17128
rect 17276 17076 17282 17128
rect 17865 17119 17923 17125
rect 17865 17085 17877 17119
rect 17911 17116 17923 17119
rect 18230 17116 18236 17128
rect 17911 17088 18236 17116
rect 17911 17085 17923 17088
rect 17865 17079 17923 17085
rect 18230 17076 18236 17088
rect 18288 17076 18294 17128
rect 18506 17076 18512 17128
rect 18564 17116 18570 17128
rect 19720 17116 19748 17224
rect 20073 17187 20131 17193
rect 20073 17153 20085 17187
rect 20119 17153 20131 17187
rect 20073 17147 20131 17153
rect 20257 17187 20315 17193
rect 20257 17153 20269 17187
rect 20303 17184 20315 17187
rect 20364 17184 20392 17224
rect 20622 17212 20628 17264
rect 20680 17212 20686 17264
rect 21376 17252 21404 17292
rect 21637 17289 21649 17323
rect 21683 17320 21695 17323
rect 23661 17323 23719 17329
rect 23661 17320 23673 17323
rect 21683 17292 23673 17320
rect 21683 17289 21695 17292
rect 21637 17283 21695 17289
rect 23661 17289 23673 17292
rect 23707 17289 23719 17323
rect 23661 17283 23719 17289
rect 23750 17280 23756 17332
rect 23808 17320 23814 17332
rect 24578 17320 24584 17332
rect 23808 17292 24584 17320
rect 23808 17280 23814 17292
rect 24578 17280 24584 17292
rect 24636 17280 24642 17332
rect 26142 17280 26148 17332
rect 26200 17280 26206 17332
rect 26694 17280 26700 17332
rect 26752 17280 26758 17332
rect 27157 17323 27215 17329
rect 27157 17289 27169 17323
rect 27203 17320 27215 17323
rect 27203 17292 27292 17320
rect 27203 17289 27215 17292
rect 27157 17283 27215 17289
rect 23109 17255 23167 17261
rect 21376 17224 22784 17252
rect 22756 17196 22784 17224
rect 23109 17221 23121 17255
rect 23155 17252 23167 17255
rect 23198 17252 23204 17264
rect 23155 17224 23204 17252
rect 23155 17221 23167 17224
rect 23109 17215 23167 17221
rect 23198 17212 23204 17224
rect 23256 17212 23262 17264
rect 23566 17212 23572 17264
rect 23624 17252 23630 17264
rect 24029 17255 24087 17261
rect 24029 17252 24041 17255
rect 23624 17224 24041 17252
rect 23624 17212 23630 17224
rect 24029 17221 24041 17224
rect 24075 17221 24087 17255
rect 26160 17252 26188 17280
rect 24029 17215 24087 17221
rect 24412 17224 26188 17252
rect 20303 17156 20392 17184
rect 20303 17153 20315 17156
rect 20257 17147 20315 17153
rect 18564 17088 19748 17116
rect 20088 17116 20116 17147
rect 20806 17144 20812 17196
rect 20864 17144 20870 17196
rect 21266 17144 21272 17196
rect 21324 17144 21330 17196
rect 21634 17144 21640 17196
rect 21692 17144 21698 17196
rect 21821 17187 21879 17193
rect 21821 17153 21833 17187
rect 21867 17184 21879 17187
rect 22097 17187 22155 17193
rect 21867 17156 22048 17184
rect 21867 17153 21879 17156
rect 21821 17147 21879 17153
rect 20824 17116 20852 17144
rect 20088 17088 20852 17116
rect 18564 17076 18570 17088
rect 21358 17076 21364 17128
rect 21416 17076 21422 17128
rect 21450 17076 21456 17128
rect 21508 17076 21514 17128
rect 21652 17116 21680 17144
rect 21913 17119 21971 17125
rect 21913 17116 21925 17119
rect 21652 17088 21925 17116
rect 21913 17085 21925 17088
rect 21959 17085 21971 17119
rect 22020 17116 22048 17156
rect 22097 17153 22109 17187
rect 22143 17184 22155 17187
rect 22646 17184 22652 17196
rect 22143 17156 22652 17184
rect 22143 17153 22155 17156
rect 22097 17147 22155 17153
rect 22646 17144 22652 17156
rect 22704 17144 22710 17196
rect 22738 17144 22744 17196
rect 22796 17144 22802 17196
rect 23014 17144 23020 17196
rect 23072 17144 23078 17196
rect 23293 17187 23351 17193
rect 23293 17153 23305 17187
rect 23339 17184 23351 17187
rect 23382 17184 23388 17196
rect 23339 17156 23388 17184
rect 23339 17153 23351 17156
rect 23293 17147 23351 17153
rect 23382 17144 23388 17156
rect 23440 17144 23446 17196
rect 23778 17187 23836 17193
rect 23778 17153 23790 17187
rect 23824 17184 23836 17187
rect 23824 17156 24072 17184
rect 23824 17153 23836 17156
rect 23778 17147 23836 17153
rect 23569 17119 23627 17125
rect 22020 17088 22876 17116
rect 21913 17079 21971 17085
rect 20441 17051 20499 17057
rect 17144 17020 17264 17048
rect 10744 17008 10750 17020
rect 6880 16952 7788 16980
rect 6880 16940 6886 16952
rect 9674 16940 9680 16992
rect 9732 16940 9738 16992
rect 10778 16940 10784 16992
rect 10836 16980 10842 16992
rect 10965 16983 11023 16989
rect 10965 16980 10977 16983
rect 10836 16952 10977 16980
rect 10836 16940 10842 16952
rect 10965 16949 10977 16952
rect 11011 16949 11023 16983
rect 10965 16943 11023 16949
rect 11146 16940 11152 16992
rect 11204 16980 11210 16992
rect 15838 16980 15844 16992
rect 11204 16952 15844 16980
rect 11204 16940 11210 16952
rect 15838 16940 15844 16952
rect 15896 16940 15902 16992
rect 16669 16983 16727 16989
rect 16669 16949 16681 16983
rect 16715 16980 16727 16983
rect 17126 16980 17132 16992
rect 16715 16952 17132 16980
rect 16715 16949 16727 16952
rect 16669 16943 16727 16949
rect 17126 16940 17132 16952
rect 17184 16940 17190 16992
rect 17236 16980 17264 17020
rect 20441 17017 20453 17051
rect 20487 17048 20499 17051
rect 21468 17048 21496 17076
rect 22281 17051 22339 17057
rect 22281 17048 22293 17051
rect 20487 17020 21496 17048
rect 21560 17020 22293 17048
rect 20487 17017 20499 17020
rect 20441 17011 20499 17017
rect 17862 16980 17868 16992
rect 17236 16952 17868 16980
rect 17862 16940 17868 16952
rect 17920 16940 17926 16992
rect 19334 16940 19340 16992
rect 19392 16980 19398 16992
rect 20073 16983 20131 16989
rect 20073 16980 20085 16983
rect 19392 16952 20085 16980
rect 19392 16940 19398 16952
rect 20073 16949 20085 16952
rect 20119 16949 20131 16983
rect 20073 16943 20131 16949
rect 20162 16940 20168 16992
rect 20220 16980 20226 16992
rect 20622 16980 20628 16992
rect 20220 16952 20628 16980
rect 20220 16940 20226 16952
rect 20622 16940 20628 16952
rect 20680 16980 20686 16992
rect 20717 16983 20775 16989
rect 20717 16980 20729 16983
rect 20680 16952 20729 16980
rect 20680 16940 20686 16952
rect 20717 16949 20729 16952
rect 20763 16949 20775 16983
rect 20717 16943 20775 16949
rect 21453 16983 21511 16989
rect 21453 16949 21465 16983
rect 21499 16980 21511 16983
rect 21560 16980 21588 17020
rect 22281 17017 22293 17020
rect 22327 17017 22339 17051
rect 22281 17011 22339 17017
rect 21499 16952 21588 16980
rect 22005 16983 22063 16989
rect 21499 16949 21511 16952
rect 21453 16943 21511 16949
rect 22005 16949 22017 16983
rect 22051 16980 22063 16983
rect 22186 16980 22192 16992
rect 22051 16952 22192 16980
rect 22051 16949 22063 16952
rect 22005 16943 22063 16949
rect 22186 16940 22192 16952
rect 22244 16940 22250 16992
rect 22554 16940 22560 16992
rect 22612 16940 22618 16992
rect 22848 16989 22876 17088
rect 23569 17085 23581 17119
rect 23615 17116 23627 17119
rect 24044 17116 24072 17156
rect 24118 17144 24124 17196
rect 24176 17184 24182 17196
rect 24412 17193 24440 17224
rect 24305 17187 24363 17193
rect 24305 17184 24317 17187
rect 24176 17156 24317 17184
rect 24176 17144 24182 17156
rect 24305 17153 24317 17156
rect 24351 17153 24363 17187
rect 24305 17147 24363 17153
rect 24397 17187 24455 17193
rect 24397 17153 24409 17187
rect 24443 17153 24455 17187
rect 24397 17147 24455 17153
rect 24486 17144 24492 17196
rect 24544 17144 24550 17196
rect 24578 17144 24584 17196
rect 24636 17184 24642 17196
rect 24673 17187 24731 17193
rect 24673 17184 24685 17187
rect 24636 17156 24685 17184
rect 24636 17144 24642 17156
rect 24673 17153 24685 17156
rect 24719 17153 24731 17187
rect 24673 17147 24731 17153
rect 26421 17187 26479 17193
rect 26421 17153 26433 17187
rect 26467 17153 26479 17187
rect 26421 17147 26479 17153
rect 25774 17116 25780 17128
rect 23615 17088 23796 17116
rect 24044 17088 25780 17116
rect 23615 17085 23627 17088
rect 23569 17079 23627 17085
rect 23768 17060 23796 17088
rect 25774 17076 25780 17088
rect 25832 17076 25838 17128
rect 26326 17076 26332 17128
rect 26384 17116 26390 17128
rect 26436 17116 26464 17147
rect 26510 17144 26516 17196
rect 26568 17144 26574 17196
rect 26973 17187 27031 17193
rect 26973 17153 26985 17187
rect 27019 17184 27031 17187
rect 27154 17184 27160 17196
rect 27019 17156 27160 17184
rect 27019 17153 27031 17156
rect 26973 17147 27031 17153
rect 27154 17144 27160 17156
rect 27212 17144 27218 17196
rect 27264 17128 27292 17292
rect 27522 17280 27528 17332
rect 27580 17320 27586 17332
rect 27985 17323 28043 17329
rect 27985 17320 27997 17323
rect 27580 17292 27997 17320
rect 27580 17280 27586 17292
rect 27985 17289 27997 17292
rect 28031 17289 28043 17323
rect 28810 17320 28816 17332
rect 27985 17283 28043 17289
rect 28276 17292 28816 17320
rect 27890 17252 27896 17264
rect 27632 17224 27896 17252
rect 27338 17144 27344 17196
rect 27396 17144 27402 17196
rect 27632 17193 27660 17224
rect 27890 17212 27896 17224
rect 27948 17212 27954 17264
rect 27617 17187 27675 17193
rect 27617 17153 27629 17187
rect 27663 17153 27675 17187
rect 27617 17147 27675 17153
rect 28074 17144 28080 17196
rect 28132 17184 28138 17196
rect 28276 17193 28304 17292
rect 28810 17280 28816 17292
rect 28868 17280 28874 17332
rect 29638 17280 29644 17332
rect 29696 17320 29702 17332
rect 30006 17320 30012 17332
rect 29696 17292 30012 17320
rect 29696 17280 29702 17292
rect 30006 17280 30012 17292
rect 30064 17280 30070 17332
rect 32950 17280 32956 17332
rect 33008 17320 33014 17332
rect 33008 17292 35940 17320
rect 33008 17280 33014 17292
rect 35912 17264 35940 17292
rect 36078 17280 36084 17332
rect 36136 17320 36142 17332
rect 39942 17320 39948 17332
rect 36136 17292 39948 17320
rect 36136 17280 36142 17292
rect 39942 17280 39948 17292
rect 40000 17280 40006 17332
rect 40037 17323 40095 17329
rect 40037 17289 40049 17323
rect 40083 17320 40095 17323
rect 40494 17320 40500 17332
rect 40083 17292 40500 17320
rect 40083 17289 40095 17292
rect 40037 17283 40095 17289
rect 40494 17280 40500 17292
rect 40552 17280 40558 17332
rect 29178 17212 29184 17264
rect 29236 17252 29242 17264
rect 34241 17255 34299 17261
rect 34241 17252 34253 17255
rect 29236 17224 34253 17252
rect 29236 17212 29242 17224
rect 34241 17221 34253 17224
rect 34287 17221 34299 17255
rect 34241 17215 34299 17221
rect 35894 17212 35900 17264
rect 35952 17212 35958 17264
rect 39577 17255 39635 17261
rect 39577 17221 39589 17255
rect 39623 17252 39635 17255
rect 39758 17252 39764 17264
rect 39623 17224 39764 17252
rect 39623 17221 39635 17224
rect 39577 17215 39635 17221
rect 39758 17212 39764 17224
rect 39816 17252 39822 17264
rect 39816 17224 40540 17252
rect 39816 17212 39822 17224
rect 28261 17187 28319 17193
rect 28261 17184 28273 17187
rect 28132 17156 28273 17184
rect 28132 17144 28138 17156
rect 28261 17153 28273 17156
rect 28307 17153 28319 17187
rect 28261 17147 28319 17153
rect 28626 17144 28632 17196
rect 28684 17144 28690 17196
rect 28813 17187 28871 17193
rect 28813 17153 28825 17187
rect 28859 17182 28871 17187
rect 28859 17154 28948 17182
rect 28859 17153 28871 17154
rect 28813 17147 28871 17153
rect 26384 17088 26464 17116
rect 26384 17076 26390 17088
rect 27246 17076 27252 17128
rect 27304 17076 27310 17128
rect 27709 17119 27767 17125
rect 27709 17085 27721 17119
rect 27755 17116 27767 17119
rect 28166 17116 28172 17128
rect 27755 17088 28172 17116
rect 27755 17085 27767 17088
rect 27709 17079 27767 17085
rect 28166 17076 28172 17088
rect 28224 17076 28230 17128
rect 28537 17119 28595 17125
rect 28537 17116 28549 17119
rect 28368 17088 28549 17116
rect 22925 17051 22983 17057
rect 22925 17017 22937 17051
rect 22971 17048 22983 17051
rect 23658 17048 23664 17060
rect 22971 17020 23664 17048
rect 22971 17017 22983 17020
rect 22925 17011 22983 17017
rect 23658 17008 23664 17020
rect 23716 17008 23722 17060
rect 23750 17008 23756 17060
rect 23808 17008 23814 17060
rect 28077 17051 28135 17057
rect 28077 17048 28089 17051
rect 23860 17020 28089 17048
rect 22833 16983 22891 16989
rect 22833 16949 22845 16983
rect 22879 16980 22891 16983
rect 23860 16980 23888 17020
rect 28077 17017 28089 17020
rect 28123 17017 28135 17051
rect 28077 17011 28135 17017
rect 22879 16952 23888 16980
rect 22879 16949 22891 16952
rect 22833 16943 22891 16949
rect 23934 16940 23940 16992
rect 23992 16940 23998 16992
rect 26234 16940 26240 16992
rect 26292 16980 26298 16992
rect 26510 16980 26516 16992
rect 26292 16952 26516 16980
rect 26292 16940 26298 16952
rect 26510 16940 26516 16952
rect 26568 16940 26574 16992
rect 27522 16940 27528 16992
rect 27580 16940 27586 16992
rect 27614 16940 27620 16992
rect 27672 16940 27678 16992
rect 28368 16980 28396 17088
rect 28537 17085 28549 17088
rect 28583 17085 28595 17119
rect 28920 17116 28948 17154
rect 28994 17144 29000 17196
rect 29052 17184 29058 17196
rect 29089 17187 29147 17193
rect 29089 17184 29101 17187
rect 29052 17156 29101 17184
rect 29052 17144 29058 17156
rect 29089 17153 29101 17156
rect 29135 17184 29147 17187
rect 29365 17187 29423 17193
rect 29365 17184 29377 17187
rect 29135 17156 29377 17184
rect 29135 17153 29147 17156
rect 29089 17147 29147 17153
rect 29365 17153 29377 17156
rect 29411 17153 29423 17187
rect 29365 17147 29423 17153
rect 29917 17187 29975 17193
rect 29917 17153 29929 17187
rect 29963 17184 29975 17187
rect 30190 17184 30196 17196
rect 29963 17156 30196 17184
rect 29963 17153 29975 17156
rect 29917 17147 29975 17153
rect 29822 17116 29828 17128
rect 28920 17088 29828 17116
rect 28537 17079 28595 17085
rect 29822 17076 29828 17088
rect 29880 17076 29886 17128
rect 28445 17051 28503 17057
rect 28445 17017 28457 17051
rect 28491 17048 28503 17051
rect 28491 17020 28856 17048
rect 28491 17017 28503 17020
rect 28445 17011 28503 17017
rect 28626 16980 28632 16992
rect 28368 16952 28632 16980
rect 28626 16940 28632 16952
rect 28684 16940 28690 16992
rect 28828 16980 28856 17020
rect 28902 17008 28908 17060
rect 28960 17008 28966 17060
rect 28997 17051 29055 17057
rect 28997 17017 29009 17051
rect 29043 17048 29055 17051
rect 29270 17048 29276 17060
rect 29043 17020 29276 17048
rect 29043 17017 29055 17020
rect 28997 17011 29055 17017
rect 29270 17008 29276 17020
rect 29328 17008 29334 17060
rect 29086 16980 29092 16992
rect 28828 16952 29092 16980
rect 29086 16940 29092 16952
rect 29144 16940 29150 16992
rect 29454 16940 29460 16992
rect 29512 16980 29518 16992
rect 29932 16980 29960 17147
rect 30190 17144 30196 17156
rect 30248 17144 30254 17196
rect 33505 17187 33563 17193
rect 33505 17153 33517 17187
rect 33551 17153 33563 17187
rect 33965 17187 34023 17193
rect 33965 17184 33977 17187
rect 33505 17147 33563 17153
rect 33796 17156 33977 17184
rect 33410 17076 33416 17128
rect 33468 17076 33474 17128
rect 32582 17008 32588 17060
rect 32640 17048 32646 17060
rect 33521 17048 33549 17147
rect 33796 17128 33824 17156
rect 33965 17153 33977 17156
rect 34011 17153 34023 17187
rect 33965 17147 34023 17153
rect 34054 17144 34060 17196
rect 34112 17184 34118 17196
rect 34149 17187 34207 17193
rect 34149 17184 34161 17187
rect 34112 17156 34161 17184
rect 34112 17144 34118 17156
rect 34149 17153 34161 17156
rect 34195 17153 34207 17187
rect 34149 17147 34207 17153
rect 34333 17187 34391 17193
rect 34333 17153 34345 17187
rect 34379 17184 34391 17187
rect 35618 17184 35624 17196
rect 34379 17156 35624 17184
rect 34379 17153 34391 17156
rect 34333 17147 34391 17153
rect 35618 17144 35624 17156
rect 35676 17184 35682 17196
rect 39853 17187 39911 17193
rect 35676 17156 35940 17184
rect 35676 17144 35682 17156
rect 33778 17076 33784 17128
rect 33836 17076 33842 17128
rect 33873 17119 33931 17125
rect 33873 17085 33885 17119
rect 33919 17116 33931 17119
rect 33919 17088 34008 17116
rect 33919 17085 33931 17088
rect 33873 17079 33931 17085
rect 32640 17020 33549 17048
rect 32640 17008 32646 17020
rect 33980 16992 34008 17088
rect 35912 17060 35940 17156
rect 39853 17153 39865 17187
rect 39899 17184 39911 17187
rect 40034 17184 40040 17196
rect 39899 17156 40040 17184
rect 39899 17153 39911 17156
rect 39853 17147 39911 17153
rect 40034 17144 40040 17156
rect 40092 17144 40098 17196
rect 40129 17187 40187 17193
rect 40129 17153 40141 17187
rect 40175 17153 40187 17187
rect 40129 17147 40187 17153
rect 39761 17119 39819 17125
rect 39761 17085 39773 17119
rect 39807 17116 39819 17119
rect 39942 17116 39948 17128
rect 39807 17088 39948 17116
rect 39807 17085 39819 17088
rect 39761 17079 39819 17085
rect 39942 17076 39948 17088
rect 40000 17076 40006 17128
rect 35894 17008 35900 17060
rect 35952 17008 35958 17060
rect 40144 17048 40172 17147
rect 40218 17144 40224 17196
rect 40276 17184 40282 17196
rect 40512 17193 40540 17224
rect 40313 17187 40371 17193
rect 40313 17184 40325 17187
rect 40276 17156 40325 17184
rect 40276 17144 40282 17156
rect 40313 17153 40325 17156
rect 40359 17153 40371 17187
rect 40313 17147 40371 17153
rect 40497 17187 40555 17193
rect 40497 17153 40509 17187
rect 40543 17153 40555 17187
rect 40497 17147 40555 17153
rect 39592 17020 40172 17048
rect 39592 16992 39620 17020
rect 29512 16952 29960 16980
rect 29512 16940 29518 16952
rect 31754 16940 31760 16992
rect 31812 16980 31818 16992
rect 32214 16980 32220 16992
rect 31812 16952 32220 16980
rect 31812 16940 31818 16952
rect 32214 16940 32220 16952
rect 32272 16940 32278 16992
rect 33229 16983 33287 16989
rect 33229 16949 33241 16983
rect 33275 16980 33287 16983
rect 33502 16980 33508 16992
rect 33275 16952 33508 16980
rect 33275 16949 33287 16952
rect 33229 16943 33287 16949
rect 33502 16940 33508 16952
rect 33560 16940 33566 16992
rect 33962 16940 33968 16992
rect 34020 16940 34026 16992
rect 34517 16983 34575 16989
rect 34517 16949 34529 16983
rect 34563 16980 34575 16983
rect 37366 16980 37372 16992
rect 34563 16952 37372 16980
rect 34563 16949 34575 16952
rect 34517 16943 34575 16949
rect 37366 16940 37372 16952
rect 37424 16940 37430 16992
rect 39574 16940 39580 16992
rect 39632 16940 39638 16992
rect 39666 16940 39672 16992
rect 39724 16940 39730 16992
rect 1104 16890 41400 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 41400 16890
rect 1104 16816 41400 16838
rect 3510 16776 3516 16788
rect 1780 16748 3516 16776
rect 1780 16649 1808 16748
rect 3510 16736 3516 16748
rect 3568 16736 3574 16788
rect 3878 16736 3884 16788
rect 3936 16736 3942 16788
rect 4062 16736 4068 16788
rect 4120 16776 4126 16788
rect 6730 16776 6736 16788
rect 4120 16748 6736 16776
rect 4120 16736 4126 16748
rect 1765 16643 1823 16649
rect 1765 16609 1777 16643
rect 1811 16609 1823 16643
rect 1765 16603 1823 16609
rect 2041 16643 2099 16649
rect 2041 16609 2053 16643
rect 2087 16640 2099 16643
rect 2130 16640 2136 16652
rect 2087 16612 2136 16640
rect 2087 16609 2099 16612
rect 2041 16603 2099 16609
rect 2130 16600 2136 16612
rect 2188 16600 2194 16652
rect 3513 16643 3571 16649
rect 3513 16609 3525 16643
rect 3559 16640 3571 16643
rect 3896 16640 3924 16736
rect 3559 16612 3924 16640
rect 3559 16609 3571 16612
rect 3513 16603 3571 16609
rect 4798 16600 4804 16652
rect 4856 16600 4862 16652
rect 4908 16649 4936 16748
rect 6730 16736 6736 16748
rect 6788 16736 6794 16788
rect 8021 16779 8079 16785
rect 8021 16745 8033 16779
rect 8067 16776 8079 16779
rect 8110 16776 8116 16788
rect 8067 16748 8116 16776
rect 8067 16745 8079 16748
rect 8021 16739 8079 16745
rect 8110 16736 8116 16748
rect 8168 16736 8174 16788
rect 9674 16736 9680 16788
rect 9732 16776 9738 16788
rect 12161 16779 12219 16785
rect 9732 16748 12112 16776
rect 9732 16736 9738 16748
rect 4893 16643 4951 16649
rect 4893 16609 4905 16643
rect 4939 16609 4951 16643
rect 4893 16603 4951 16609
rect 5261 16643 5319 16649
rect 5261 16609 5273 16643
rect 5307 16640 5319 16643
rect 5350 16640 5356 16652
rect 5307 16612 5356 16640
rect 5307 16609 5319 16612
rect 5261 16603 5319 16609
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 6270 16600 6276 16652
rect 6328 16600 6334 16652
rect 6549 16643 6607 16649
rect 6549 16609 6561 16643
rect 6595 16640 6607 16643
rect 6638 16640 6644 16652
rect 6595 16612 6644 16640
rect 6595 16609 6607 16612
rect 6549 16603 6607 16609
rect 6638 16600 6644 16612
rect 6696 16600 6702 16652
rect 9585 16643 9643 16649
rect 9585 16609 9597 16643
rect 9631 16640 9643 16643
rect 9692 16640 9720 16736
rect 12084 16720 12112 16748
rect 12161 16745 12173 16779
rect 12207 16776 12219 16779
rect 12250 16776 12256 16788
rect 12207 16748 12256 16776
rect 12207 16745 12219 16748
rect 12161 16739 12219 16745
rect 12250 16736 12256 16748
rect 12308 16736 12314 16788
rect 14734 16776 14740 16788
rect 12406 16748 14740 16776
rect 12066 16668 12072 16720
rect 12124 16708 12130 16720
rect 12406 16708 12434 16748
rect 14734 16736 14740 16748
rect 14792 16776 14798 16788
rect 20714 16776 20720 16788
rect 14792 16748 20720 16776
rect 14792 16736 14798 16748
rect 20714 16736 20720 16748
rect 20772 16736 20778 16788
rect 21818 16776 21824 16788
rect 20824 16748 21824 16776
rect 20824 16720 20852 16748
rect 21818 16736 21824 16748
rect 21876 16736 21882 16788
rect 22005 16779 22063 16785
rect 22005 16745 22017 16779
rect 22051 16776 22063 16779
rect 22646 16776 22652 16788
rect 22051 16748 22652 16776
rect 22051 16745 22063 16748
rect 22005 16739 22063 16745
rect 22646 16736 22652 16748
rect 22704 16736 22710 16788
rect 23658 16736 23664 16788
rect 23716 16736 23722 16788
rect 24486 16736 24492 16788
rect 24544 16776 24550 16788
rect 25685 16779 25743 16785
rect 25685 16776 25697 16779
rect 24544 16748 25697 16776
rect 24544 16736 24550 16748
rect 25685 16745 25697 16748
rect 25731 16745 25743 16779
rect 25685 16739 25743 16745
rect 25774 16736 25780 16788
rect 25832 16776 25838 16788
rect 26421 16779 26479 16785
rect 26421 16776 26433 16779
rect 25832 16748 26433 16776
rect 25832 16736 25838 16748
rect 26421 16745 26433 16748
rect 26467 16745 26479 16779
rect 26421 16739 26479 16745
rect 28718 16736 28724 16788
rect 28776 16736 28782 16788
rect 32033 16779 32091 16785
rect 32033 16745 32045 16779
rect 32079 16776 32091 16779
rect 32214 16776 32220 16788
rect 32079 16748 32220 16776
rect 32079 16745 32091 16748
rect 32033 16739 32091 16745
rect 32214 16736 32220 16748
rect 32272 16736 32278 16788
rect 32324 16748 33272 16776
rect 12124 16680 12434 16708
rect 12124 16668 12130 16680
rect 13170 16668 13176 16720
rect 13228 16708 13234 16720
rect 13228 16680 14136 16708
rect 13228 16668 13234 16680
rect 9631 16612 9720 16640
rect 9631 16609 9643 16612
rect 9585 16603 9643 16609
rect 9950 16600 9956 16652
rect 10008 16640 10014 16652
rect 10413 16643 10471 16649
rect 10413 16640 10425 16643
rect 10008 16612 10425 16640
rect 10008 16600 10014 16612
rect 10413 16609 10425 16612
rect 10459 16609 10471 16643
rect 10413 16603 10471 16609
rect 10689 16643 10747 16649
rect 10689 16609 10701 16643
rect 10735 16640 10747 16643
rect 10778 16640 10784 16652
rect 10735 16612 10784 16640
rect 10735 16609 10747 16612
rect 10689 16603 10747 16609
rect 10778 16600 10784 16612
rect 10836 16600 10842 16652
rect 14108 16649 14136 16680
rect 19886 16668 19892 16720
rect 19944 16668 19950 16720
rect 20806 16668 20812 16720
rect 20864 16668 20870 16720
rect 21177 16711 21235 16717
rect 21177 16677 21189 16711
rect 21223 16708 21235 16711
rect 22278 16708 22284 16720
rect 21223 16680 22284 16708
rect 21223 16677 21235 16680
rect 21177 16671 21235 16677
rect 22278 16668 22284 16680
rect 22336 16668 22342 16720
rect 27614 16708 27620 16720
rect 25424 16680 27620 16708
rect 14093 16643 14151 16649
rect 14093 16609 14105 16643
rect 14139 16640 14151 16643
rect 16574 16640 16580 16652
rect 14139 16612 16580 16640
rect 14139 16609 14151 16612
rect 14093 16603 14151 16609
rect 16574 16600 16580 16612
rect 16632 16600 16638 16652
rect 4816 16572 4844 16600
rect 4816 16544 6040 16572
rect 3418 16504 3424 16516
rect 3266 16476 3424 16504
rect 3418 16464 3424 16476
rect 3476 16504 3482 16516
rect 4709 16507 4767 16513
rect 3476 16476 4476 16504
rect 3476 16464 3482 16476
rect 4062 16396 4068 16448
rect 4120 16436 4126 16448
rect 4341 16439 4399 16445
rect 4341 16436 4353 16439
rect 4120 16408 4353 16436
rect 4120 16396 4126 16408
rect 4341 16405 4353 16408
rect 4387 16405 4399 16439
rect 4448 16436 4476 16476
rect 4709 16473 4721 16507
rect 4755 16504 4767 16507
rect 5813 16507 5871 16513
rect 5813 16504 5825 16507
rect 4755 16476 5825 16504
rect 4755 16473 4767 16476
rect 4709 16467 4767 16473
rect 5813 16473 5825 16476
rect 5859 16473 5871 16507
rect 5813 16467 5871 16473
rect 5074 16436 5080 16448
rect 4448 16408 5080 16436
rect 4341 16399 4399 16405
rect 5074 16396 5080 16408
rect 5132 16396 5138 16448
rect 5442 16396 5448 16448
rect 5500 16436 5506 16448
rect 5905 16439 5963 16445
rect 5905 16436 5917 16439
rect 5500 16408 5917 16436
rect 5500 16396 5506 16408
rect 5905 16405 5917 16408
rect 5951 16405 5963 16439
rect 6012 16436 6040 16544
rect 6086 16532 6092 16584
rect 6144 16532 6150 16584
rect 9030 16532 9036 16584
rect 9088 16572 9094 16584
rect 9490 16572 9496 16584
rect 9088 16544 9496 16572
rect 9088 16532 9094 16544
rect 9490 16532 9496 16544
rect 9548 16532 9554 16584
rect 13906 16532 13912 16584
rect 13964 16532 13970 16584
rect 18138 16572 18144 16584
rect 15502 16544 18144 16572
rect 18138 16532 18144 16544
rect 18196 16572 18202 16584
rect 19242 16572 19248 16584
rect 18196 16544 19248 16572
rect 18196 16532 18202 16544
rect 19242 16532 19248 16544
rect 19300 16532 19306 16584
rect 19904 16581 19932 16668
rect 20070 16600 20076 16652
rect 20128 16640 20134 16652
rect 20165 16643 20223 16649
rect 20165 16640 20177 16643
rect 20128 16612 20177 16640
rect 20128 16600 20134 16612
rect 20165 16609 20177 16612
rect 20211 16609 20223 16643
rect 20165 16603 20223 16609
rect 21634 16600 21640 16652
rect 21692 16600 21698 16652
rect 21910 16600 21916 16652
rect 21968 16640 21974 16652
rect 25424 16640 25452 16680
rect 27614 16668 27620 16680
rect 27672 16708 27678 16720
rect 32324 16708 32352 16748
rect 27672 16680 28396 16708
rect 27672 16668 27678 16680
rect 28368 16649 28396 16680
rect 31312 16680 32352 16708
rect 33244 16708 33272 16748
rect 34330 16736 34336 16788
rect 34388 16736 34394 16788
rect 34514 16736 34520 16788
rect 34572 16736 34578 16788
rect 34790 16736 34796 16788
rect 34848 16776 34854 16788
rect 34885 16779 34943 16785
rect 34885 16776 34897 16779
rect 34848 16748 34897 16776
rect 34848 16736 34854 16748
rect 34885 16745 34897 16748
rect 34931 16745 34943 16779
rect 34885 16739 34943 16745
rect 35434 16736 35440 16788
rect 35492 16776 35498 16788
rect 35618 16776 35624 16788
rect 35492 16748 35624 16776
rect 35492 16736 35498 16748
rect 35618 16736 35624 16748
rect 35676 16736 35682 16788
rect 37366 16736 37372 16788
rect 37424 16776 37430 16788
rect 37461 16779 37519 16785
rect 37461 16776 37473 16779
rect 37424 16748 37473 16776
rect 37424 16736 37430 16748
rect 37461 16745 37473 16748
rect 37507 16745 37519 16779
rect 37461 16739 37519 16745
rect 37645 16779 37703 16785
rect 37645 16745 37657 16779
rect 37691 16776 37703 16779
rect 37734 16776 37740 16788
rect 37691 16748 37740 16776
rect 37691 16745 37703 16748
rect 37645 16739 37703 16745
rect 37476 16708 37504 16739
rect 37734 16736 37740 16748
rect 37792 16736 37798 16788
rect 38654 16736 38660 16788
rect 38712 16776 38718 16788
rect 39853 16779 39911 16785
rect 39853 16776 39865 16779
rect 38712 16748 39865 16776
rect 38712 16736 38718 16748
rect 39853 16745 39865 16748
rect 39899 16745 39911 16779
rect 39853 16739 39911 16745
rect 39942 16736 39948 16788
rect 40000 16776 40006 16788
rect 40313 16779 40371 16785
rect 40313 16776 40325 16779
rect 40000 16748 40325 16776
rect 40000 16736 40006 16748
rect 40313 16745 40325 16748
rect 40359 16745 40371 16779
rect 40313 16739 40371 16745
rect 40126 16708 40132 16720
rect 33244 16680 34928 16708
rect 28353 16643 28411 16649
rect 21968 16612 25452 16640
rect 25516 16612 26188 16640
rect 21968 16600 21974 16612
rect 25516 16584 25544 16612
rect 19889 16575 19947 16581
rect 19889 16541 19901 16575
rect 19935 16541 19947 16575
rect 19889 16535 19947 16541
rect 19981 16575 20039 16581
rect 19981 16541 19993 16575
rect 20027 16572 20039 16575
rect 20622 16572 20628 16584
rect 20027 16544 20628 16572
rect 20027 16541 20039 16544
rect 19981 16535 20039 16541
rect 20622 16532 20628 16544
rect 20680 16532 20686 16584
rect 21361 16575 21419 16581
rect 21361 16541 21373 16575
rect 21407 16541 21419 16575
rect 21361 16535 21419 16541
rect 9048 16504 9076 16532
rect 9401 16507 9459 16513
rect 9401 16504 9413 16507
rect 7774 16476 9076 16504
rect 9232 16476 9413 16504
rect 9232 16448 9260 16476
rect 9401 16473 9413 16476
rect 9447 16473 9459 16507
rect 9401 16467 9459 16473
rect 11238 16464 11244 16516
rect 11296 16464 11302 16516
rect 14369 16507 14427 16513
rect 14369 16473 14381 16507
rect 14415 16473 14427 16507
rect 14369 16467 14427 16473
rect 8110 16436 8116 16448
rect 6012 16408 8116 16436
rect 5905 16399 5963 16405
rect 8110 16396 8116 16408
rect 8168 16396 8174 16448
rect 8938 16396 8944 16448
rect 8996 16396 9002 16448
rect 9214 16396 9220 16448
rect 9272 16396 9278 16448
rect 9306 16396 9312 16448
rect 9364 16396 9370 16448
rect 13725 16439 13783 16445
rect 13725 16405 13737 16439
rect 13771 16436 13783 16439
rect 14384 16436 14412 16467
rect 14642 16464 14648 16516
rect 14700 16464 14706 16516
rect 18414 16464 18420 16516
rect 18472 16504 18478 16516
rect 18966 16504 18972 16516
rect 18472 16476 18972 16504
rect 18472 16464 18478 16476
rect 18966 16464 18972 16476
rect 19024 16464 19030 16516
rect 13771 16408 14412 16436
rect 14660 16436 14688 16464
rect 15841 16439 15899 16445
rect 15841 16436 15853 16439
rect 14660 16408 15853 16436
rect 13771 16405 13783 16408
rect 13725 16399 13783 16405
rect 15841 16405 15853 16408
rect 15887 16405 15899 16439
rect 15841 16399 15899 16405
rect 17678 16396 17684 16448
rect 17736 16436 17742 16448
rect 20714 16436 20720 16448
rect 17736 16408 20720 16436
rect 17736 16396 17742 16408
rect 20714 16396 20720 16408
rect 20772 16396 20778 16448
rect 21376 16436 21404 16535
rect 21542 16532 21548 16584
rect 21600 16532 21606 16584
rect 22005 16575 22063 16581
rect 22005 16572 22017 16575
rect 21652 16544 22017 16572
rect 21450 16464 21456 16516
rect 21508 16504 21514 16516
rect 21652 16504 21680 16544
rect 22005 16541 22017 16544
rect 22051 16541 22063 16575
rect 22005 16535 22063 16541
rect 22922 16532 22928 16584
rect 22980 16572 22986 16584
rect 23293 16575 23351 16581
rect 23293 16572 23305 16575
rect 22980 16544 23305 16572
rect 22980 16532 22986 16544
rect 23293 16541 23305 16544
rect 23339 16541 23351 16575
rect 23293 16535 23351 16541
rect 23474 16532 23480 16584
rect 23532 16532 23538 16584
rect 25038 16532 25044 16584
rect 25096 16532 25102 16584
rect 25222 16581 25228 16584
rect 25189 16575 25228 16581
rect 25189 16541 25201 16575
rect 25189 16535 25228 16541
rect 25222 16532 25228 16535
rect 25280 16532 25286 16584
rect 25498 16532 25504 16584
rect 25556 16581 25562 16584
rect 25556 16572 25564 16581
rect 25556 16544 25649 16572
rect 25556 16535 25564 16544
rect 25556 16532 25562 16535
rect 25682 16532 25688 16584
rect 25740 16574 25746 16584
rect 25777 16575 25835 16581
rect 25777 16574 25789 16575
rect 25740 16546 25789 16574
rect 25740 16532 25746 16546
rect 25777 16541 25789 16546
rect 25823 16541 25835 16575
rect 25777 16535 25835 16541
rect 25866 16532 25872 16584
rect 25924 16572 25930 16584
rect 26160 16581 26188 16612
rect 28353 16609 28365 16643
rect 28399 16609 28411 16643
rect 28353 16603 28411 16609
rect 28626 16600 28632 16652
rect 28684 16640 28690 16652
rect 28813 16643 28871 16649
rect 28813 16640 28825 16643
rect 28684 16612 28825 16640
rect 28684 16600 28690 16612
rect 28813 16609 28825 16612
rect 28859 16640 28871 16643
rect 30653 16643 30711 16649
rect 30653 16640 30665 16643
rect 28859 16612 30665 16640
rect 28859 16609 28871 16612
rect 28813 16603 28871 16609
rect 30653 16609 30665 16612
rect 30699 16609 30711 16643
rect 30653 16603 30711 16609
rect 31312 16581 31340 16680
rect 32677 16643 32735 16649
rect 31956 16612 32444 16640
rect 26145 16575 26203 16581
rect 25924 16544 25969 16572
rect 25924 16532 25930 16544
rect 26145 16541 26157 16575
rect 26191 16541 26203 16575
rect 26145 16535 26203 16541
rect 26242 16575 26300 16581
rect 26242 16541 26254 16575
rect 26288 16541 26300 16575
rect 26242 16535 26300 16541
rect 28537 16575 28595 16581
rect 28537 16541 28549 16575
rect 28583 16541 28595 16575
rect 28537 16535 28595 16541
rect 30285 16575 30343 16581
rect 30285 16541 30297 16575
rect 30331 16572 30343 16575
rect 31297 16575 31355 16581
rect 30331 16544 31248 16572
rect 30331 16541 30343 16544
rect 30285 16535 30343 16541
rect 21508 16476 21680 16504
rect 21729 16507 21787 16513
rect 21508 16464 21514 16476
rect 21729 16473 21741 16507
rect 21775 16504 21787 16507
rect 23566 16504 23572 16516
rect 21775 16476 23572 16504
rect 21775 16473 21787 16476
rect 21729 16467 21787 16473
rect 23566 16464 23572 16476
rect 23624 16464 23630 16516
rect 23750 16464 23756 16516
rect 23808 16504 23814 16516
rect 25317 16507 25375 16513
rect 25317 16504 25329 16507
rect 23808 16476 25329 16504
rect 23808 16464 23814 16476
rect 25317 16473 25329 16476
rect 25363 16473 25375 16507
rect 25317 16467 25375 16473
rect 25409 16507 25467 16513
rect 25409 16473 25421 16507
rect 25455 16473 25467 16507
rect 25409 16467 25467 16473
rect 22002 16436 22008 16448
rect 21376 16408 22008 16436
rect 22002 16396 22008 16408
rect 22060 16396 22066 16448
rect 22094 16396 22100 16448
rect 22152 16436 22158 16448
rect 22189 16439 22247 16445
rect 22189 16436 22201 16439
rect 22152 16408 22201 16436
rect 22152 16396 22158 16408
rect 22189 16405 22201 16408
rect 22235 16405 22247 16439
rect 22189 16399 22247 16405
rect 24854 16396 24860 16448
rect 24912 16436 24918 16448
rect 25424 16436 25452 16467
rect 26050 16464 26056 16516
rect 26108 16464 26114 16516
rect 25774 16436 25780 16448
rect 24912 16408 25780 16436
rect 24912 16396 24918 16408
rect 25774 16396 25780 16408
rect 25832 16396 25838 16448
rect 25866 16396 25872 16448
rect 25924 16436 25930 16448
rect 26257 16436 26285 16535
rect 26326 16464 26332 16516
rect 26384 16504 26390 16516
rect 28552 16504 28580 16535
rect 31220 16516 31248 16544
rect 31297 16541 31309 16575
rect 31343 16541 31355 16575
rect 31297 16535 31355 16541
rect 31570 16532 31576 16584
rect 31628 16581 31634 16584
rect 31628 16575 31657 16581
rect 31645 16541 31657 16575
rect 31628 16535 31657 16541
rect 31757 16575 31815 16581
rect 31757 16541 31769 16575
rect 31803 16572 31815 16575
rect 31846 16572 31852 16584
rect 31803 16544 31852 16572
rect 31803 16541 31815 16544
rect 31757 16535 31815 16541
rect 31628 16532 31634 16535
rect 31846 16532 31852 16544
rect 31904 16532 31910 16584
rect 31956 16516 31984 16612
rect 32416 16581 32444 16612
rect 32677 16609 32689 16643
rect 32723 16640 32735 16643
rect 33042 16640 33048 16652
rect 32723 16612 33048 16640
rect 32723 16609 32735 16612
rect 32677 16603 32735 16609
rect 33042 16600 33048 16612
rect 33100 16600 33106 16652
rect 33410 16600 33416 16652
rect 33468 16600 33474 16652
rect 33502 16600 33508 16652
rect 33560 16640 33566 16652
rect 33778 16640 33784 16652
rect 33560 16612 33784 16640
rect 33560 16600 33566 16612
rect 33778 16600 33784 16612
rect 33836 16600 33842 16652
rect 34146 16640 34152 16652
rect 33888 16612 34152 16640
rect 33888 16581 33916 16612
rect 34146 16600 34152 16612
rect 34204 16600 34210 16652
rect 32217 16575 32275 16581
rect 32217 16572 32229 16575
rect 32146 16544 32229 16572
rect 29454 16504 29460 16516
rect 26384 16476 29460 16504
rect 26384 16464 26390 16476
rect 29454 16464 29460 16476
rect 29512 16464 29518 16516
rect 30469 16507 30527 16513
rect 30469 16504 30481 16507
rect 30392 16476 30481 16504
rect 30392 16448 30420 16476
rect 30469 16473 30481 16476
rect 30515 16473 30527 16507
rect 30469 16467 30527 16473
rect 31202 16464 31208 16516
rect 31260 16464 31266 16516
rect 31389 16507 31447 16513
rect 31389 16473 31401 16507
rect 31435 16473 31447 16507
rect 31389 16467 31447 16473
rect 31481 16507 31539 16513
rect 31481 16473 31493 16507
rect 31527 16504 31539 16507
rect 31938 16504 31944 16516
rect 31527 16476 31944 16504
rect 31527 16473 31539 16476
rect 31481 16467 31539 16473
rect 25924 16408 26285 16436
rect 25924 16396 25930 16408
rect 27338 16396 27344 16448
rect 27396 16436 27402 16448
rect 27798 16436 27804 16448
rect 27396 16408 27804 16436
rect 27396 16396 27402 16408
rect 27798 16396 27804 16408
rect 27856 16396 27862 16448
rect 30374 16396 30380 16448
rect 30432 16396 30438 16448
rect 31110 16396 31116 16448
rect 31168 16396 31174 16448
rect 31404 16436 31432 16467
rect 31938 16464 31944 16476
rect 31996 16464 32002 16516
rect 32146 16436 32174 16544
rect 32217 16541 32229 16544
rect 32263 16541 32275 16575
rect 32217 16535 32275 16541
rect 32401 16575 32459 16581
rect 32401 16541 32413 16575
rect 32447 16541 32459 16575
rect 32401 16535 32459 16541
rect 33597 16575 33655 16581
rect 33597 16541 33609 16575
rect 33643 16541 33655 16575
rect 33597 16535 33655 16541
rect 33873 16575 33931 16581
rect 33873 16541 33885 16575
rect 33919 16541 33931 16575
rect 34532 16572 34744 16582
rect 34900 16572 34928 16680
rect 35268 16680 36400 16708
rect 37476 16680 40132 16708
rect 35069 16575 35127 16581
rect 35069 16572 35081 16575
rect 33873 16535 33931 16541
rect 33980 16554 34836 16572
rect 33980 16544 34560 16554
rect 34716 16544 34836 16554
rect 34900 16544 35081 16572
rect 32309 16507 32367 16513
rect 32309 16473 32321 16507
rect 32355 16473 32367 16507
rect 32309 16467 32367 16473
rect 32539 16507 32597 16513
rect 32539 16473 32551 16507
rect 32585 16504 32597 16507
rect 32674 16504 32680 16516
rect 32585 16476 32680 16504
rect 32585 16473 32597 16476
rect 32539 16467 32597 16473
rect 32214 16436 32220 16448
rect 31404 16408 32220 16436
rect 32214 16396 32220 16408
rect 32272 16396 32278 16448
rect 32324 16436 32352 16467
rect 32674 16464 32680 16476
rect 32732 16464 32738 16516
rect 33410 16464 33416 16516
rect 33468 16464 33474 16516
rect 33612 16504 33640 16535
rect 33980 16504 34008 16544
rect 34422 16513 34428 16516
rect 33612 16476 34008 16504
rect 34149 16507 34207 16513
rect 34149 16473 34161 16507
rect 34195 16504 34207 16507
rect 34365 16507 34428 16513
rect 34195 16476 34284 16504
rect 34195 16473 34207 16476
rect 34149 16467 34207 16473
rect 33428 16436 33456 16464
rect 32324 16408 33456 16436
rect 33781 16439 33839 16445
rect 33781 16405 33793 16439
rect 33827 16436 33839 16439
rect 34054 16436 34060 16448
rect 33827 16408 34060 16436
rect 33827 16405 33839 16408
rect 33781 16399 33839 16405
rect 34054 16396 34060 16408
rect 34112 16396 34118 16448
rect 34256 16436 34284 16476
rect 34365 16473 34377 16507
rect 34411 16473 34428 16507
rect 34365 16467 34428 16473
rect 34422 16464 34428 16467
rect 34480 16464 34486 16516
rect 34514 16464 34520 16516
rect 34572 16464 34578 16516
rect 34532 16436 34560 16464
rect 34256 16408 34560 16436
rect 34808 16436 34836 16544
rect 35069 16541 35081 16544
rect 35115 16572 35127 16575
rect 35268 16572 35296 16680
rect 35529 16643 35587 16649
rect 35529 16609 35541 16643
rect 35575 16640 35587 16643
rect 36078 16640 36084 16652
rect 35575 16612 36084 16640
rect 35575 16609 35587 16612
rect 35529 16603 35587 16609
rect 35115 16544 35296 16572
rect 35115 16541 35127 16544
rect 35069 16535 35127 16541
rect 35158 16464 35164 16516
rect 35216 16464 35222 16516
rect 35250 16464 35256 16516
rect 35308 16464 35314 16516
rect 35342 16464 35348 16516
rect 35400 16513 35406 16516
rect 35400 16507 35429 16513
rect 35417 16473 35429 16507
rect 35400 16467 35429 16473
rect 35400 16464 35406 16467
rect 35636 16436 35664 16612
rect 36078 16600 36084 16612
rect 36136 16600 36142 16652
rect 36372 16448 36400 16680
rect 40126 16668 40132 16680
rect 40184 16668 40190 16720
rect 40037 16643 40095 16649
rect 40037 16640 40049 16643
rect 39224 16612 40049 16640
rect 39224 16584 39252 16612
rect 40037 16609 40049 16612
rect 40083 16609 40095 16643
rect 40037 16603 40095 16609
rect 37277 16575 37335 16581
rect 37277 16541 37289 16575
rect 37323 16572 37335 16575
rect 37366 16572 37372 16584
rect 37323 16544 37372 16572
rect 37323 16541 37335 16544
rect 37277 16535 37335 16541
rect 37366 16532 37372 16544
rect 37424 16532 37430 16584
rect 37458 16532 37464 16584
rect 37516 16532 37522 16584
rect 39206 16532 39212 16584
rect 39264 16532 39270 16584
rect 40129 16575 40187 16581
rect 40129 16541 40141 16575
rect 40175 16572 40187 16575
rect 40678 16572 40684 16584
rect 40175 16544 40684 16572
rect 40175 16541 40187 16544
rect 40129 16535 40187 16541
rect 40678 16532 40684 16544
rect 40736 16532 40742 16584
rect 39298 16464 39304 16516
rect 39356 16504 39362 16516
rect 39853 16507 39911 16513
rect 39853 16504 39865 16507
rect 39356 16476 39865 16504
rect 39356 16464 39362 16476
rect 39853 16473 39865 16476
rect 39899 16473 39911 16507
rect 39853 16467 39911 16473
rect 34808 16408 35664 16436
rect 36354 16396 36360 16448
rect 36412 16436 36418 16448
rect 38378 16436 38384 16448
rect 36412 16408 38384 16436
rect 36412 16396 36418 16408
rect 38378 16396 38384 16408
rect 38436 16396 38442 16448
rect 1104 16346 41400 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 41400 16346
rect 1104 16272 41400 16294
rect 5261 16235 5319 16241
rect 5261 16201 5273 16235
rect 5307 16232 5319 16235
rect 5350 16232 5356 16244
rect 5307 16204 5356 16232
rect 5307 16201 5319 16204
rect 5261 16195 5319 16201
rect 5350 16192 5356 16204
rect 5408 16192 5414 16244
rect 5445 16235 5503 16241
rect 5445 16201 5457 16235
rect 5491 16232 5503 16235
rect 6086 16232 6092 16244
rect 5491 16204 6092 16232
rect 5491 16201 5503 16204
rect 5445 16195 5503 16201
rect 6086 16192 6092 16204
rect 6144 16192 6150 16244
rect 9582 16192 9588 16244
rect 9640 16192 9646 16244
rect 9674 16192 9680 16244
rect 9732 16232 9738 16244
rect 10505 16235 10563 16241
rect 10505 16232 10517 16235
rect 9732 16204 10517 16232
rect 9732 16192 9738 16204
rect 10505 16201 10517 16204
rect 10551 16201 10563 16235
rect 10505 16195 10563 16201
rect 12406 16204 13860 16232
rect 5074 16164 5080 16176
rect 5014 16136 5080 16164
rect 5074 16124 5080 16136
rect 5132 16164 5138 16176
rect 5626 16164 5632 16176
rect 5132 16136 5632 16164
rect 5132 16124 5138 16136
rect 5626 16124 5632 16136
rect 5684 16124 5690 16176
rect 9030 16124 9036 16176
rect 9088 16124 9094 16176
rect 9600 16164 9628 16192
rect 11238 16164 11244 16176
rect 9600 16136 11244 16164
rect 11238 16124 11244 16136
rect 11296 16124 11302 16176
rect 3510 16056 3516 16108
rect 3568 16056 3574 16108
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 7009 16099 7067 16105
rect 7009 16096 7021 16099
rect 5859 16068 7021 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 7009 16065 7021 16068
rect 7055 16065 7067 16099
rect 7009 16059 7067 16065
rect 8018 16056 8024 16108
rect 8076 16056 8082 16108
rect 9953 16099 10011 16105
rect 9953 16096 9965 16099
rect 9646 16068 9965 16096
rect 3786 15988 3792 16040
rect 3844 15988 3850 16040
rect 5258 15988 5264 16040
rect 5316 16028 5322 16040
rect 5905 16031 5963 16037
rect 5905 16028 5917 16031
rect 5316 16000 5917 16028
rect 5316 15988 5322 16000
rect 5905 15997 5917 16000
rect 5951 16028 5963 16031
rect 6089 16031 6147 16037
rect 5951 16000 6040 16028
rect 5951 15997 5963 16000
rect 5905 15991 5963 15997
rect 6012 15892 6040 16000
rect 6089 15997 6101 16031
rect 6135 15997 6147 16031
rect 6089 15991 6147 15997
rect 6104 15960 6132 15991
rect 6178 15988 6184 16040
rect 6236 16028 6242 16040
rect 6365 16031 6423 16037
rect 6365 16028 6377 16031
rect 6236 16000 6377 16028
rect 6236 15988 6242 16000
rect 6365 15997 6377 16000
rect 6411 15997 6423 16031
rect 6365 15991 6423 15997
rect 6822 15988 6828 16040
rect 6880 15988 6886 16040
rect 8294 15988 8300 16040
rect 8352 15988 8358 16040
rect 9030 15988 9036 16040
rect 9088 16028 9094 16040
rect 9646 16028 9674 16068
rect 9088 16000 9674 16028
rect 9088 15988 9094 16000
rect 6840 15960 6868 15988
rect 9784 15969 9812 16068
rect 9953 16065 9965 16068
rect 9999 16065 10011 16099
rect 9953 16059 10011 16065
rect 10042 16056 10048 16108
rect 10100 16096 10106 16108
rect 12406 16096 12434 16204
rect 13078 16164 13084 16176
rect 12636 16136 13084 16164
rect 12636 16105 12664 16136
rect 13078 16124 13084 16136
rect 13136 16164 13142 16176
rect 13832 16164 13860 16204
rect 13906 16192 13912 16244
rect 13964 16232 13970 16244
rect 14093 16235 14151 16241
rect 14093 16232 14105 16235
rect 13964 16204 14105 16232
rect 13964 16192 13970 16204
rect 14093 16201 14105 16204
rect 14139 16201 14151 16235
rect 14093 16195 14151 16201
rect 14461 16235 14519 16241
rect 14461 16201 14473 16235
rect 14507 16232 14519 16235
rect 14642 16232 14648 16244
rect 14507 16204 14648 16232
rect 14507 16201 14519 16204
rect 14461 16195 14519 16201
rect 14642 16192 14648 16204
rect 14700 16192 14706 16244
rect 17954 16192 17960 16244
rect 18012 16232 18018 16244
rect 18055 16235 18113 16241
rect 18055 16232 18067 16235
rect 18012 16204 18067 16232
rect 18012 16192 18018 16204
rect 18055 16201 18067 16204
rect 18101 16201 18113 16235
rect 18055 16195 18113 16201
rect 18141 16235 18199 16241
rect 18141 16201 18153 16235
rect 18187 16232 18199 16235
rect 18782 16232 18788 16244
rect 18187 16204 18788 16232
rect 18187 16201 18199 16204
rect 18141 16195 18199 16201
rect 18782 16192 18788 16204
rect 18840 16192 18846 16244
rect 21910 16232 21916 16244
rect 19306 16204 21916 16232
rect 18414 16164 18420 16176
rect 13136 16136 13308 16164
rect 13832 16136 18092 16164
rect 13136 16124 13142 16136
rect 13280 16105 13308 16136
rect 18064 16108 18092 16136
rect 18156 16136 18420 16164
rect 10100 16068 12434 16096
rect 12529 16099 12587 16105
rect 10100 16056 10106 16068
rect 12529 16065 12541 16099
rect 12575 16065 12587 16099
rect 12529 16059 12587 16065
rect 12621 16099 12679 16105
rect 12621 16065 12633 16099
rect 12667 16065 12679 16099
rect 13173 16099 13231 16105
rect 12621 16059 12679 16065
rect 12728 16094 13124 16096
rect 13173 16094 13185 16099
rect 12728 16068 13185 16094
rect 12544 16028 12572 16059
rect 12728 16028 12756 16068
rect 13096 16066 13185 16068
rect 13173 16065 13185 16066
rect 13219 16065 13231 16099
rect 13173 16059 13231 16065
rect 13265 16099 13323 16105
rect 13265 16065 13277 16099
rect 13311 16065 13323 16099
rect 13265 16059 13323 16065
rect 13354 16056 13360 16108
rect 13412 16056 13418 16108
rect 13538 16056 13544 16108
rect 13596 16056 13602 16108
rect 14182 16056 14188 16108
rect 14240 16056 14246 16108
rect 16025 16099 16083 16105
rect 16025 16065 16037 16099
rect 16071 16065 16083 16099
rect 16025 16059 16083 16065
rect 12544 16000 12756 16028
rect 12805 16031 12863 16037
rect 6104 15932 6868 15960
rect 9769 15963 9827 15969
rect 9769 15929 9781 15963
rect 9815 15929 9827 15963
rect 12544 15960 12572 16000
rect 12805 15997 12817 16031
rect 12851 16028 12863 16031
rect 13556 16028 13584 16056
rect 12851 16020 13124 16028
rect 13280 16020 13584 16028
rect 12851 16000 13584 16020
rect 12851 15997 12863 16000
rect 12805 15991 12863 15997
rect 13096 15992 13308 16000
rect 14200 15960 14228 16056
rect 14550 15988 14556 16040
rect 14608 15988 14614 16040
rect 14734 15988 14740 16040
rect 14792 15988 14798 16040
rect 12544 15932 14228 15960
rect 16040 15960 16068 16059
rect 16942 16056 16948 16108
rect 17000 16096 17006 16108
rect 17037 16099 17095 16105
rect 17037 16096 17049 16099
rect 17000 16068 17049 16096
rect 17000 16056 17006 16068
rect 17037 16065 17049 16068
rect 17083 16065 17095 16099
rect 17037 16059 17095 16065
rect 17862 16056 17868 16108
rect 17920 16096 17926 16108
rect 17957 16099 18015 16105
rect 17957 16096 17969 16099
rect 17920 16068 17969 16096
rect 17920 16056 17926 16068
rect 17957 16065 17969 16068
rect 18003 16065 18015 16099
rect 17957 16059 18015 16065
rect 18046 16056 18052 16108
rect 18104 16056 18110 16108
rect 16114 15988 16120 16040
rect 16172 16028 16178 16040
rect 16853 16031 16911 16037
rect 16853 16028 16865 16031
rect 16172 16000 16865 16028
rect 16172 15988 16178 16000
rect 16853 15997 16865 16000
rect 16899 16028 16911 16031
rect 18156 16028 18184 16136
rect 18414 16124 18420 16136
rect 18472 16124 18478 16176
rect 19306 16164 19334 16204
rect 21910 16192 21916 16204
rect 21968 16192 21974 16244
rect 23750 16232 23756 16244
rect 22066 16204 23756 16232
rect 18892 16136 19334 16164
rect 18230 16056 18236 16108
rect 18288 16096 18294 16108
rect 18892 16105 18920 16136
rect 21450 16124 21456 16176
rect 21508 16164 21514 16176
rect 22066 16164 22094 16204
rect 23750 16192 23756 16204
rect 23808 16192 23814 16244
rect 25222 16192 25228 16244
rect 25280 16232 25286 16244
rect 25501 16235 25559 16241
rect 25501 16232 25513 16235
rect 25280 16204 25513 16232
rect 25280 16192 25286 16204
rect 25501 16201 25513 16204
rect 25547 16201 25559 16235
rect 28534 16232 28540 16244
rect 25501 16195 25559 16201
rect 25597 16204 28540 16232
rect 21508 16136 22094 16164
rect 23569 16167 23627 16173
rect 21508 16124 21514 16136
rect 23569 16133 23581 16167
rect 23615 16164 23627 16167
rect 24670 16164 24676 16176
rect 23615 16136 24676 16164
rect 23615 16133 23627 16136
rect 23569 16127 23627 16133
rect 24670 16124 24676 16136
rect 24728 16124 24734 16176
rect 25597 16164 25625 16204
rect 28534 16192 28540 16204
rect 28592 16192 28598 16244
rect 33410 16192 33416 16244
rect 33468 16232 33474 16244
rect 34606 16232 34612 16244
rect 33468 16204 34612 16232
rect 33468 16192 33474 16204
rect 34606 16192 34612 16204
rect 34664 16192 34670 16244
rect 34974 16192 34980 16244
rect 35032 16192 35038 16244
rect 35161 16235 35219 16241
rect 35161 16201 35173 16235
rect 35207 16232 35219 16235
rect 35434 16232 35440 16244
rect 35207 16204 35440 16232
rect 35207 16201 35219 16204
rect 35161 16195 35219 16201
rect 35434 16192 35440 16204
rect 35492 16192 35498 16244
rect 37274 16192 37280 16244
rect 37332 16232 37338 16244
rect 37550 16232 37556 16244
rect 37332 16204 37556 16232
rect 37332 16192 37338 16204
rect 37550 16192 37556 16204
rect 37608 16192 37614 16244
rect 39482 16232 39488 16244
rect 39224 16204 39488 16232
rect 26145 16167 26203 16173
rect 26145 16164 26157 16167
rect 24780 16136 25625 16164
rect 25700 16136 26157 16164
rect 18877 16099 18935 16105
rect 18288 16068 18828 16096
rect 18288 16056 18294 16068
rect 16899 16000 18184 16028
rect 16899 15997 16911 16000
rect 16853 15991 16911 15997
rect 18506 15988 18512 16040
rect 18564 15988 18570 16040
rect 18800 16028 18828 16068
rect 18877 16065 18889 16099
rect 18923 16065 18935 16099
rect 18877 16059 18935 16065
rect 18966 16056 18972 16108
rect 19024 16096 19030 16108
rect 19153 16099 19211 16105
rect 19153 16096 19165 16099
rect 19024 16068 19165 16096
rect 19024 16056 19030 16068
rect 19153 16065 19165 16068
rect 19199 16065 19211 16099
rect 19153 16059 19211 16065
rect 19242 16056 19248 16108
rect 19300 16056 19306 16108
rect 20622 16056 20628 16108
rect 20680 16096 20686 16108
rect 24780 16096 24808 16136
rect 20680 16068 24808 16096
rect 20680 16056 20686 16068
rect 25038 16056 25044 16108
rect 25096 16096 25102 16108
rect 25498 16096 25504 16108
rect 25096 16068 25504 16096
rect 25096 16056 25102 16068
rect 25498 16056 25504 16068
rect 25556 16056 25562 16108
rect 25700 16096 25728 16136
rect 26145 16133 26157 16136
rect 26191 16133 26203 16167
rect 26145 16127 26203 16133
rect 26694 16124 26700 16176
rect 26752 16164 26758 16176
rect 28350 16164 28356 16176
rect 26752 16136 28356 16164
rect 26752 16124 26758 16136
rect 28350 16124 28356 16136
rect 28408 16124 28414 16176
rect 31110 16124 31116 16176
rect 31168 16164 31174 16176
rect 31205 16167 31263 16173
rect 31205 16164 31217 16167
rect 31168 16136 31217 16164
rect 31168 16124 31174 16136
rect 31205 16133 31217 16136
rect 31251 16133 31263 16167
rect 31205 16127 31263 16133
rect 31478 16124 31484 16176
rect 31536 16164 31542 16176
rect 32858 16164 32864 16176
rect 31536 16136 32864 16164
rect 31536 16124 31542 16136
rect 32858 16124 32864 16136
rect 32916 16124 32922 16176
rect 34514 16124 34520 16176
rect 34572 16164 34578 16176
rect 34992 16164 35020 16192
rect 35250 16164 35256 16176
rect 34572 16136 35020 16164
rect 35048 16136 35256 16164
rect 34572 16124 34578 16136
rect 25608 16068 25728 16096
rect 25777 16099 25835 16105
rect 19260 16028 19288 16056
rect 18800 16000 19288 16028
rect 23937 16031 23995 16037
rect 23937 15997 23949 16031
rect 23983 15997 23995 16031
rect 23937 15991 23995 15997
rect 24029 16031 24087 16037
rect 24029 15997 24041 16031
rect 24075 16028 24087 16031
rect 25314 16028 25320 16040
rect 24075 16000 25320 16028
rect 24075 15997 24087 16000
rect 24029 15991 24087 15997
rect 16040 15932 19104 15960
rect 9769 15923 9827 15929
rect 7834 15892 7840 15904
rect 6012 15864 7840 15892
rect 7834 15852 7840 15864
rect 7892 15852 7898 15904
rect 12710 15852 12716 15904
rect 12768 15852 12774 15904
rect 12894 15852 12900 15904
rect 12952 15852 12958 15904
rect 16206 15852 16212 15904
rect 16264 15852 16270 15904
rect 17221 15895 17279 15901
rect 17221 15861 17233 15895
rect 17267 15892 17279 15895
rect 17402 15892 17408 15904
rect 17267 15864 17408 15892
rect 17267 15861 17279 15864
rect 17221 15855 17279 15861
rect 17402 15852 17408 15864
rect 17460 15852 17466 15904
rect 17494 15852 17500 15904
rect 17552 15892 17558 15904
rect 18506 15892 18512 15904
rect 17552 15864 18512 15892
rect 17552 15852 17558 15864
rect 18506 15852 18512 15864
rect 18564 15852 18570 15904
rect 19076 15892 19104 15932
rect 19150 15920 19156 15972
rect 19208 15920 19214 15972
rect 22002 15920 22008 15972
rect 22060 15960 22066 15972
rect 22554 15960 22560 15972
rect 22060 15932 22560 15960
rect 22060 15920 22066 15932
rect 22554 15920 22560 15932
rect 22612 15920 22618 15972
rect 23952 15960 23980 15991
rect 25314 15988 25320 16000
rect 25372 15988 25378 16040
rect 25406 15988 25412 16040
rect 25464 16028 25470 16040
rect 25608 16028 25636 16068
rect 25777 16065 25789 16099
rect 25823 16096 25835 16099
rect 25823 16068 26280 16096
rect 25823 16065 25835 16068
rect 25777 16059 25835 16065
rect 25464 16000 25636 16028
rect 25464 15988 25470 16000
rect 25682 15988 25688 16040
rect 25740 15988 25746 16040
rect 26053 16031 26111 16037
rect 26053 15997 26065 16031
rect 26099 15997 26111 16031
rect 26053 15991 26111 15997
rect 25038 15960 25044 15972
rect 23952 15932 25044 15960
rect 25038 15920 25044 15932
rect 25096 15920 25102 15972
rect 25332 15960 25360 15988
rect 25866 15960 25872 15972
rect 25332 15932 25872 15960
rect 25866 15920 25872 15932
rect 25924 15960 25930 15972
rect 26068 15960 26096 15991
rect 26252 15972 26280 16068
rect 26602 16056 26608 16108
rect 26660 16096 26666 16108
rect 28626 16096 28632 16108
rect 26660 16068 28632 16096
rect 26660 16056 26666 16068
rect 28626 16056 28632 16068
rect 28684 16056 28690 16108
rect 30374 16056 30380 16108
rect 30432 16096 30438 16108
rect 30926 16096 30932 16108
rect 30432 16068 30932 16096
rect 30432 16056 30438 16068
rect 30926 16056 30932 16068
rect 30984 16056 30990 16108
rect 31386 16056 31392 16108
rect 31444 16056 31450 16108
rect 34422 16056 34428 16108
rect 34480 16096 34486 16108
rect 35048 16096 35076 16136
rect 35250 16124 35256 16136
rect 35308 16164 35314 16176
rect 35529 16167 35587 16173
rect 35529 16164 35541 16167
rect 35308 16136 35541 16164
rect 35308 16124 35314 16136
rect 35529 16133 35541 16136
rect 35575 16133 35587 16167
rect 35529 16127 35587 16133
rect 35618 16124 35624 16176
rect 35676 16173 35682 16176
rect 39224 16173 39252 16204
rect 39482 16192 39488 16204
rect 39540 16192 39546 16244
rect 35676 16167 35705 16173
rect 35693 16133 35705 16167
rect 35676 16127 35705 16133
rect 39209 16167 39267 16173
rect 39209 16133 39221 16167
rect 39255 16133 39267 16167
rect 39209 16127 39267 16133
rect 35676 16124 35682 16127
rect 34480 16068 35076 16096
rect 34480 16056 34486 16068
rect 35158 16056 35164 16108
rect 35216 16096 35222 16108
rect 35345 16099 35403 16105
rect 35345 16096 35357 16099
rect 35216 16068 35357 16096
rect 35216 16056 35222 16068
rect 35345 16065 35357 16068
rect 35391 16065 35403 16099
rect 35345 16059 35403 16065
rect 26326 15988 26332 16040
rect 26384 16028 26390 16040
rect 28718 16028 28724 16040
rect 26384 16000 28724 16028
rect 26384 15988 26390 16000
rect 28718 15988 28724 16000
rect 28776 15988 28782 16040
rect 31573 16031 31631 16037
rect 31573 15997 31585 16031
rect 31619 16028 31631 16031
rect 35360 16028 35388 16059
rect 35434 16056 35440 16108
rect 35492 16056 35498 16108
rect 36078 16096 36084 16108
rect 35820 16068 36084 16096
rect 35618 16028 35624 16040
rect 31619 16000 35296 16028
rect 35360 16000 35624 16028
rect 31619 15997 31631 16000
rect 31573 15991 31631 15997
rect 25924 15932 26096 15960
rect 25924 15920 25930 15932
rect 26234 15920 26240 15972
rect 26292 15920 26298 15972
rect 26786 15920 26792 15972
rect 26844 15920 26850 15972
rect 35268 15960 35296 16000
rect 35618 15988 35624 16000
rect 35676 15988 35682 16040
rect 35820 16037 35848 16068
rect 36078 16056 36084 16068
rect 36136 16056 36142 16108
rect 36262 16056 36268 16108
rect 36320 16056 36326 16108
rect 36538 16056 36544 16108
rect 36596 16096 36602 16108
rect 37277 16099 37335 16105
rect 37277 16096 37289 16099
rect 36596 16068 37289 16096
rect 36596 16056 36602 16068
rect 37277 16065 37289 16068
rect 37323 16065 37335 16099
rect 37277 16059 37335 16065
rect 37458 16056 37464 16108
rect 37516 16096 37522 16108
rect 37553 16099 37611 16105
rect 37553 16096 37565 16099
rect 37516 16068 37565 16096
rect 37516 16056 37522 16068
rect 37553 16065 37565 16068
rect 37599 16065 37611 16099
rect 37553 16059 37611 16065
rect 39022 16056 39028 16108
rect 39080 16096 39086 16108
rect 39390 16096 39396 16108
rect 39080 16068 39396 16096
rect 39080 16056 39086 16068
rect 39390 16056 39396 16068
rect 39448 16096 39454 16108
rect 39485 16099 39543 16105
rect 39485 16096 39497 16099
rect 39448 16068 39497 16096
rect 39448 16056 39454 16068
rect 39485 16065 39497 16068
rect 39531 16065 39543 16099
rect 39485 16059 39543 16065
rect 35805 16031 35863 16037
rect 35805 15997 35817 16031
rect 35851 15997 35863 16031
rect 36280 16028 36308 16056
rect 37369 16031 37427 16037
rect 37369 16028 37381 16031
rect 36280 16000 37381 16028
rect 35805 15991 35863 15997
rect 37369 15997 37381 16000
rect 37415 15997 37427 16031
rect 39301 16031 39359 16037
rect 39301 16028 39313 16031
rect 37369 15991 37427 15997
rect 37476 16000 39313 16028
rect 37476 15960 37504 16000
rect 39301 15997 39313 16000
rect 39347 16028 39359 16031
rect 39574 16028 39580 16040
rect 39347 16000 39580 16028
rect 39347 15997 39359 16000
rect 39301 15991 39359 15997
rect 39574 15988 39580 16000
rect 39632 15988 39638 16040
rect 35268 15932 37504 15960
rect 37737 15963 37795 15969
rect 37737 15929 37749 15963
rect 37783 15960 37795 15963
rect 39850 15960 39856 15972
rect 37783 15932 39856 15960
rect 37783 15929 37795 15932
rect 37737 15923 37795 15929
rect 39850 15920 39856 15932
rect 39908 15920 39914 15972
rect 23934 15892 23940 15904
rect 19076 15864 23940 15892
rect 23934 15852 23940 15864
rect 23992 15852 23998 15904
rect 24210 15852 24216 15904
rect 24268 15852 24274 15904
rect 24302 15852 24308 15904
rect 24360 15892 24366 15904
rect 26804 15892 26832 15920
rect 24360 15864 26832 15892
rect 24360 15852 24366 15864
rect 30282 15852 30288 15904
rect 30340 15892 30346 15904
rect 37366 15892 37372 15904
rect 30340 15864 37372 15892
rect 30340 15852 30346 15864
rect 37366 15852 37372 15864
rect 37424 15852 37430 15904
rect 37550 15852 37556 15904
rect 37608 15852 37614 15904
rect 38654 15852 38660 15904
rect 38712 15892 38718 15904
rect 39206 15892 39212 15904
rect 38712 15864 39212 15892
rect 38712 15852 38718 15864
rect 39206 15852 39212 15864
rect 39264 15852 39270 15904
rect 39666 15852 39672 15904
rect 39724 15852 39730 15904
rect 1104 15802 41400 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 41400 15802
rect 1104 15728 41400 15750
rect 3786 15648 3792 15700
rect 3844 15688 3850 15700
rect 3973 15691 4031 15697
rect 3973 15688 3985 15691
rect 3844 15660 3985 15688
rect 3844 15648 3850 15660
rect 3973 15657 3985 15660
rect 4019 15657 4031 15691
rect 3973 15651 4031 15657
rect 4880 15691 4938 15697
rect 4880 15657 4892 15691
rect 4926 15688 4938 15691
rect 5442 15688 5448 15700
rect 4926 15660 5448 15688
rect 4926 15657 4938 15660
rect 4880 15651 4938 15657
rect 5442 15648 5448 15660
rect 5500 15648 5506 15700
rect 6178 15648 6184 15700
rect 6236 15688 6242 15700
rect 6365 15691 6423 15697
rect 6365 15688 6377 15691
rect 6236 15660 6377 15688
rect 6236 15648 6242 15660
rect 6365 15657 6377 15660
rect 6411 15657 6423 15691
rect 6365 15651 6423 15657
rect 8294 15648 8300 15700
rect 8352 15688 8358 15700
rect 8481 15691 8539 15697
rect 8481 15688 8493 15691
rect 8352 15660 8493 15688
rect 8352 15648 8358 15660
rect 8481 15657 8493 15660
rect 8527 15657 8539 15691
rect 8481 15651 8539 15657
rect 8938 15648 8944 15700
rect 8996 15648 9002 15700
rect 12710 15648 12716 15700
rect 12768 15648 12774 15700
rect 12894 15648 12900 15700
rect 12952 15648 12958 15700
rect 17218 15688 17224 15700
rect 13740 15660 17224 15688
rect 2685 15623 2743 15629
rect 2685 15589 2697 15623
rect 2731 15589 2743 15623
rect 2685 15583 2743 15589
rect 2225 15487 2283 15493
rect 2225 15453 2237 15487
rect 2271 15484 2283 15487
rect 2700 15484 2728 15583
rect 3326 15512 3332 15564
rect 3384 15512 3390 15564
rect 3510 15512 3516 15564
rect 3568 15552 3574 15564
rect 4617 15555 4675 15561
rect 4617 15552 4629 15555
rect 3568 15524 4629 15552
rect 3568 15512 3574 15524
rect 4617 15521 4629 15524
rect 4663 15552 4675 15555
rect 4663 15524 6316 15552
rect 4663 15521 4675 15524
rect 4617 15515 4675 15521
rect 6288 15496 6316 15524
rect 8036 15524 8340 15552
rect 2271 15456 2728 15484
rect 3053 15487 3111 15493
rect 2271 15453 2283 15456
rect 2225 15447 2283 15453
rect 3053 15453 3065 15487
rect 3099 15484 3111 15487
rect 3694 15484 3700 15496
rect 3099 15456 3700 15484
rect 3099 15453 3111 15456
rect 3053 15447 3111 15453
rect 3694 15444 3700 15456
rect 3752 15444 3758 15496
rect 4154 15444 4160 15496
rect 4212 15444 4218 15496
rect 6270 15444 6276 15496
rect 6328 15444 6334 15496
rect 7834 15444 7840 15496
rect 7892 15444 7898 15496
rect 8036 15493 8064 15524
rect 8021 15487 8079 15493
rect 8021 15453 8033 15487
rect 8067 15453 8079 15487
rect 8021 15447 8079 15453
rect 8110 15444 8116 15496
rect 8168 15444 8174 15496
rect 8312 15493 8340 15524
rect 8297 15487 8355 15493
rect 8297 15453 8309 15487
rect 8343 15484 8355 15487
rect 8386 15484 8392 15496
rect 8343 15456 8392 15484
rect 8343 15453 8355 15456
rect 8297 15447 8355 15453
rect 8386 15444 8392 15456
rect 8444 15444 8450 15496
rect 8665 15487 8723 15493
rect 8665 15453 8677 15487
rect 8711 15484 8723 15487
rect 8956 15484 8984 15648
rect 11425 15555 11483 15561
rect 11425 15521 11437 15555
rect 11471 15552 11483 15555
rect 11606 15552 11612 15564
rect 11471 15524 11612 15552
rect 11471 15521 11483 15524
rect 11425 15515 11483 15521
rect 11606 15512 11612 15524
rect 11664 15512 11670 15564
rect 8711 15456 8984 15484
rect 12728 15484 12756 15648
rect 12912 15552 12940 15648
rect 13740 15632 13768 15660
rect 17218 15648 17224 15660
rect 17276 15648 17282 15700
rect 17954 15648 17960 15700
rect 18012 15648 18018 15700
rect 18046 15648 18052 15700
rect 18104 15688 18110 15700
rect 18104 15660 18920 15688
rect 18104 15648 18110 15660
rect 13262 15580 13268 15632
rect 13320 15620 13326 15632
rect 13722 15620 13728 15632
rect 13320 15592 13728 15620
rect 13320 15580 13326 15592
rect 13722 15580 13728 15592
rect 13780 15580 13786 15632
rect 15194 15580 15200 15632
rect 15252 15620 15258 15632
rect 17681 15623 17739 15629
rect 17681 15620 17693 15623
rect 15252 15592 17693 15620
rect 15252 15580 15258 15592
rect 17681 15589 17693 15592
rect 17727 15589 17739 15623
rect 17681 15583 17739 15589
rect 12912 15524 13676 15552
rect 13648 15493 13676 15524
rect 13357 15487 13415 15493
rect 13357 15484 13369 15487
rect 12728 15456 13369 15484
rect 8711 15453 8723 15456
rect 8665 15447 8723 15453
rect 13357 15453 13369 15456
rect 13403 15453 13415 15487
rect 13357 15447 13415 15453
rect 13449 15487 13507 15493
rect 13449 15453 13461 15487
rect 13495 15484 13507 15487
rect 13633 15487 13691 15493
rect 13495 15456 13584 15484
rect 13495 15453 13507 15456
rect 13449 15447 13507 15453
rect 1489 15419 1547 15425
rect 1489 15385 1501 15419
rect 1535 15416 1547 15419
rect 3234 15416 3240 15428
rect 1535 15388 3240 15416
rect 1535 15385 1547 15388
rect 1489 15379 1547 15385
rect 3234 15376 3240 15388
rect 3292 15376 3298 15428
rect 5626 15376 5632 15428
rect 5684 15376 5690 15428
rect 8754 15416 8760 15428
rect 8036 15388 8760 15416
rect 1578 15308 1584 15360
rect 1636 15308 1642 15360
rect 2038 15308 2044 15360
rect 2096 15308 2102 15360
rect 2774 15308 2780 15360
rect 2832 15348 2838 15360
rect 3145 15351 3203 15357
rect 3145 15348 3157 15351
rect 2832 15320 3157 15348
rect 2832 15308 2838 15320
rect 3145 15317 3157 15320
rect 3191 15348 3203 15351
rect 4062 15348 4068 15360
rect 3191 15320 4068 15348
rect 3191 15317 3203 15320
rect 3145 15311 3203 15317
rect 4062 15308 4068 15320
rect 4120 15308 4126 15360
rect 8036 15357 8064 15388
rect 8754 15376 8760 15388
rect 8812 15376 8818 15428
rect 10962 15376 10968 15428
rect 11020 15416 11026 15428
rect 11149 15419 11207 15425
rect 11149 15416 11161 15419
rect 11020 15388 11161 15416
rect 11020 15376 11026 15388
rect 11149 15385 11161 15388
rect 11195 15416 11207 15419
rect 11514 15416 11520 15428
rect 11195 15388 11520 15416
rect 11195 15385 11207 15388
rect 11149 15379 11207 15385
rect 11514 15376 11520 15388
rect 11572 15416 11578 15428
rect 12894 15416 12900 15428
rect 11572 15388 12900 15416
rect 11572 15376 11578 15388
rect 12894 15376 12900 15388
rect 12952 15416 12958 15428
rect 13556 15416 13584 15456
rect 13633 15453 13645 15487
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15484 13783 15487
rect 15212 15484 15240 15580
rect 17972 15552 18000 15648
rect 18782 15580 18788 15632
rect 18840 15580 18846 15632
rect 18892 15620 18920 15660
rect 20714 15648 20720 15700
rect 20772 15688 20778 15700
rect 22094 15688 22100 15700
rect 20772 15660 22100 15688
rect 20772 15648 20778 15660
rect 22094 15648 22100 15660
rect 22152 15648 22158 15700
rect 22738 15648 22744 15700
rect 22796 15688 22802 15700
rect 23842 15688 23848 15700
rect 22796 15660 23848 15688
rect 22796 15648 22802 15660
rect 23842 15648 23848 15660
rect 23900 15688 23906 15700
rect 25593 15691 25651 15697
rect 23900 15660 24348 15688
rect 23900 15648 23906 15660
rect 21450 15620 21456 15632
rect 18892 15592 21456 15620
rect 21450 15580 21456 15592
rect 21508 15580 21514 15632
rect 22756 15620 22784 15648
rect 21836 15592 22784 15620
rect 17972 15524 18276 15552
rect 13771 15456 15240 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 15286 15444 15292 15496
rect 15344 15444 15350 15496
rect 17037 15487 17095 15493
rect 17037 15453 17049 15487
rect 17083 15453 17095 15487
rect 17037 15447 17095 15453
rect 17313 15487 17371 15493
rect 17313 15453 17325 15487
rect 17359 15484 17371 15487
rect 17359 15456 17908 15484
rect 17359 15453 17371 15456
rect 17313 15447 17371 15453
rect 15304 15416 15332 15444
rect 15746 15416 15752 15428
rect 12952 15388 15332 15416
rect 15488 15388 15752 15416
rect 12952 15376 12958 15388
rect 8021 15351 8079 15357
rect 8021 15317 8033 15351
rect 8067 15317 8079 15351
rect 8021 15311 8079 15317
rect 8297 15351 8355 15357
rect 8297 15317 8309 15351
rect 8343 15348 8355 15351
rect 9950 15348 9956 15360
rect 8343 15320 9956 15348
rect 8343 15317 8355 15320
rect 8297 15311 8355 15317
rect 9950 15308 9956 15320
rect 10008 15308 10014 15360
rect 10778 15308 10784 15360
rect 10836 15308 10842 15360
rect 11054 15308 11060 15360
rect 11112 15348 11118 15360
rect 11241 15351 11299 15357
rect 11241 15348 11253 15351
rect 11112 15320 11253 15348
rect 11112 15308 11118 15320
rect 11241 15317 11253 15320
rect 11287 15317 11299 15351
rect 11241 15311 11299 15317
rect 13173 15351 13231 15357
rect 13173 15317 13185 15351
rect 13219 15348 13231 15351
rect 14274 15348 14280 15360
rect 13219 15320 14280 15348
rect 13219 15317 13231 15320
rect 13173 15311 13231 15317
rect 14274 15308 14280 15320
rect 14332 15308 14338 15360
rect 14458 15308 14464 15360
rect 14516 15348 14522 15360
rect 15488 15348 15516 15388
rect 15746 15376 15752 15388
rect 15804 15416 15810 15428
rect 17052 15416 17080 15447
rect 17880 15428 17908 15456
rect 18138 15444 18144 15496
rect 18196 15444 18202 15496
rect 18248 15484 18276 15524
rect 18443 15487 18501 15493
rect 18443 15484 18455 15487
rect 18248 15456 18455 15484
rect 18443 15453 18455 15456
rect 18489 15453 18501 15487
rect 18443 15447 18501 15453
rect 18601 15487 18659 15493
rect 18601 15453 18613 15487
rect 18647 15484 18659 15487
rect 18690 15484 18696 15496
rect 18647 15456 18696 15484
rect 18647 15453 18659 15456
rect 18601 15447 18659 15453
rect 18690 15444 18696 15456
rect 18748 15444 18754 15496
rect 15804 15388 16988 15416
rect 17052 15388 17356 15416
rect 15804 15376 15810 15388
rect 14516 15320 15516 15348
rect 14516 15308 14522 15320
rect 16850 15308 16856 15360
rect 16908 15308 16914 15360
rect 16960 15348 16988 15388
rect 17221 15351 17279 15357
rect 17221 15348 17233 15351
rect 16960 15320 17233 15348
rect 17221 15317 17233 15320
rect 17267 15317 17279 15351
rect 17328 15348 17356 15388
rect 17402 15376 17408 15428
rect 17460 15416 17466 15428
rect 17497 15419 17555 15425
rect 17497 15416 17509 15419
rect 17460 15388 17509 15416
rect 17460 15376 17466 15388
rect 17497 15385 17509 15388
rect 17543 15385 17555 15419
rect 17497 15379 17555 15385
rect 17862 15376 17868 15428
rect 17920 15376 17926 15428
rect 18233 15419 18291 15425
rect 18233 15385 18245 15419
rect 18279 15385 18291 15419
rect 18233 15379 18291 15385
rect 18325 15419 18383 15425
rect 18325 15385 18337 15419
rect 18371 15416 18383 15419
rect 18800 15416 18828 15580
rect 21174 15444 21180 15496
rect 21232 15484 21238 15496
rect 21269 15487 21327 15493
rect 21269 15484 21281 15487
rect 21232 15456 21281 15484
rect 21232 15444 21238 15456
rect 21269 15453 21281 15456
rect 21315 15453 21327 15487
rect 21269 15447 21327 15453
rect 21453 15487 21511 15493
rect 21453 15453 21465 15487
rect 21499 15484 21511 15487
rect 21634 15484 21640 15496
rect 21499 15456 21640 15484
rect 21499 15453 21511 15456
rect 21453 15447 21511 15453
rect 20714 15416 20720 15428
rect 18371 15388 20720 15416
rect 18371 15385 18383 15388
rect 18325 15379 18383 15385
rect 17957 15351 18015 15357
rect 17957 15348 17969 15351
rect 17328 15320 17969 15348
rect 17221 15311 17279 15317
rect 17957 15317 17969 15320
rect 18003 15317 18015 15351
rect 18248 15348 18276 15379
rect 20714 15376 20720 15388
rect 20772 15376 20778 15428
rect 21284 15416 21312 15447
rect 21634 15444 21640 15456
rect 21692 15444 21698 15496
rect 21836 15493 21864 15592
rect 24210 15580 24216 15632
rect 24268 15580 24274 15632
rect 24228 15552 24256 15580
rect 22020 15524 24256 15552
rect 24320 15552 24348 15660
rect 25593 15657 25605 15691
rect 25639 15688 25651 15691
rect 25682 15688 25688 15700
rect 25639 15660 25688 15688
rect 25639 15657 25651 15660
rect 25593 15651 25651 15657
rect 25682 15648 25688 15660
rect 25740 15648 25746 15700
rect 26878 15648 26884 15700
rect 26936 15648 26942 15700
rect 30098 15648 30104 15700
rect 30156 15648 30162 15700
rect 30282 15648 30288 15700
rect 30340 15648 30346 15700
rect 32214 15648 32220 15700
rect 32272 15688 32278 15700
rect 32861 15691 32919 15697
rect 32861 15688 32873 15691
rect 32272 15660 32873 15688
rect 32272 15648 32278 15660
rect 32861 15657 32873 15660
rect 32907 15657 32919 15691
rect 32861 15651 32919 15657
rect 35437 15691 35495 15697
rect 35437 15657 35449 15691
rect 35483 15688 35495 15691
rect 37458 15688 37464 15700
rect 35483 15660 37464 15688
rect 35483 15657 35495 15660
rect 35437 15651 35495 15657
rect 37458 15648 37464 15660
rect 37516 15648 37522 15700
rect 37921 15691 37979 15697
rect 37921 15657 37933 15691
rect 37967 15688 37979 15691
rect 39022 15688 39028 15700
rect 37967 15660 39028 15688
rect 37967 15657 37979 15660
rect 37921 15651 37979 15657
rect 39022 15648 39028 15660
rect 39080 15648 39086 15700
rect 39666 15648 39672 15700
rect 39724 15648 39730 15700
rect 39850 15648 39856 15700
rect 39908 15648 39914 15700
rect 40313 15691 40371 15697
rect 40313 15657 40325 15691
rect 40359 15688 40371 15691
rect 40586 15688 40592 15700
rect 40359 15660 40592 15688
rect 40359 15657 40371 15660
rect 40313 15651 40371 15657
rect 40586 15648 40592 15660
rect 40644 15648 40650 15700
rect 25700 15620 25728 15648
rect 25700 15592 26096 15620
rect 24320 15524 25820 15552
rect 22020 15493 22048 15524
rect 21821 15487 21879 15493
rect 21821 15453 21833 15487
rect 21867 15453 21879 15487
rect 21821 15447 21879 15453
rect 21913 15487 21971 15493
rect 21913 15453 21925 15487
rect 21959 15453 21971 15487
rect 21913 15447 21971 15453
rect 22005 15487 22063 15493
rect 22005 15453 22017 15487
rect 22051 15453 22063 15487
rect 22005 15447 22063 15453
rect 21928 15416 21956 15447
rect 22186 15444 22192 15496
rect 22244 15484 22250 15496
rect 22646 15484 22652 15496
rect 22244 15456 22652 15484
rect 22244 15444 22250 15456
rect 22646 15444 22652 15456
rect 22704 15444 22710 15496
rect 23845 15487 23903 15493
rect 23845 15453 23857 15487
rect 23891 15453 23903 15487
rect 23845 15447 23903 15453
rect 23937 15487 23995 15493
rect 23937 15453 23949 15487
rect 23983 15484 23995 15487
rect 24026 15484 24032 15496
rect 23983 15456 24032 15484
rect 23983 15453 23995 15456
rect 23937 15447 23995 15453
rect 23860 15416 23888 15447
rect 24026 15444 24032 15456
rect 24084 15444 24090 15496
rect 24121 15487 24179 15493
rect 24121 15453 24133 15487
rect 24167 15453 24179 15487
rect 24121 15447 24179 15453
rect 24213 15487 24271 15493
rect 24213 15453 24225 15487
rect 24259 15484 24271 15487
rect 24320 15484 24348 15524
rect 25792 15496 25820 15524
rect 24259 15456 24348 15484
rect 24259 15453 24271 15456
rect 24213 15447 24271 15453
rect 21284 15388 21956 15416
rect 22013 15388 23888 15416
rect 24136 15416 24164 15447
rect 24394 15444 24400 15496
rect 24452 15444 24458 15496
rect 25501 15487 25559 15493
rect 25501 15453 25513 15487
rect 25547 15453 25559 15487
rect 25501 15447 25559 15453
rect 24412 15416 24440 15444
rect 24136 15388 24440 15416
rect 25516 15416 25544 15447
rect 25774 15444 25780 15496
rect 25832 15444 25838 15496
rect 25869 15487 25927 15493
rect 25869 15453 25881 15487
rect 25915 15484 25927 15487
rect 25958 15484 25964 15496
rect 25915 15456 25964 15484
rect 25915 15453 25927 15456
rect 25869 15447 25927 15453
rect 25958 15444 25964 15456
rect 26016 15444 26022 15496
rect 26068 15493 26096 15592
rect 26142 15512 26148 15564
rect 26200 15512 26206 15564
rect 26234 15512 26240 15564
rect 26292 15552 26298 15564
rect 26292 15524 26924 15552
rect 26292 15512 26298 15524
rect 26344 15493 26372 15524
rect 26053 15487 26111 15493
rect 26053 15453 26065 15487
rect 26099 15453 26111 15487
rect 26053 15447 26111 15453
rect 26329 15487 26387 15493
rect 26329 15453 26341 15487
rect 26375 15453 26387 15487
rect 26329 15447 26387 15453
rect 26513 15487 26571 15493
rect 26513 15453 26525 15487
rect 26559 15484 26571 15487
rect 26602 15484 26608 15496
rect 26559 15456 26608 15484
rect 26559 15453 26571 15456
rect 26513 15447 26571 15453
rect 26602 15444 26608 15456
rect 26660 15444 26666 15496
rect 26697 15487 26755 15493
rect 26697 15453 26709 15487
rect 26743 15453 26755 15487
rect 26697 15447 26755 15453
rect 26142 15416 26148 15428
rect 25516 15388 26148 15416
rect 19150 15348 19156 15360
rect 18248 15320 19156 15348
rect 17957 15311 18015 15317
rect 19150 15308 19156 15320
rect 19208 15348 19214 15360
rect 19426 15348 19432 15360
rect 19208 15320 19432 15348
rect 19208 15308 19214 15320
rect 19426 15308 19432 15320
rect 19484 15308 19490 15360
rect 21174 15308 21180 15360
rect 21232 15348 21238 15360
rect 21361 15351 21419 15357
rect 21361 15348 21373 15351
rect 21232 15320 21373 15348
rect 21232 15308 21238 15320
rect 21361 15317 21373 15320
rect 21407 15317 21419 15351
rect 21361 15311 21419 15317
rect 21542 15308 21548 15360
rect 21600 15308 21606 15360
rect 21726 15308 21732 15360
rect 21784 15348 21790 15360
rect 22013 15348 22041 15388
rect 21784 15320 22041 15348
rect 21784 15308 21790 15320
rect 23658 15308 23664 15360
rect 23716 15308 23722 15360
rect 23860 15348 23888 15388
rect 26142 15376 26148 15388
rect 26200 15376 26206 15428
rect 26712 15416 26740 15447
rect 26786 15444 26792 15496
rect 26844 15444 26850 15496
rect 26896 15484 26924 15524
rect 26970 15512 26976 15564
rect 27028 15512 27034 15564
rect 30116 15552 30144 15648
rect 30190 15580 30196 15632
rect 30248 15580 30254 15632
rect 30377 15623 30435 15629
rect 30377 15589 30389 15623
rect 30423 15620 30435 15623
rect 34514 15620 34520 15632
rect 30423 15592 34520 15620
rect 30423 15589 30435 15592
rect 30377 15583 30435 15589
rect 34514 15580 34520 15592
rect 34572 15580 34578 15632
rect 36081 15555 36139 15561
rect 36081 15552 36093 15555
rect 30116 15524 36093 15552
rect 27246 15484 27252 15496
rect 26896 15456 27252 15484
rect 27246 15444 27252 15456
rect 27304 15444 27310 15496
rect 30098 15444 30104 15496
rect 30156 15484 30162 15496
rect 30374 15484 30380 15496
rect 30156 15456 30380 15484
rect 30156 15444 30162 15456
rect 30374 15444 30380 15456
rect 30432 15444 30438 15496
rect 30576 15493 30604 15524
rect 36081 15521 36093 15524
rect 36127 15521 36139 15555
rect 36081 15515 36139 15521
rect 37182 15512 37188 15564
rect 37240 15552 37246 15564
rect 37240 15524 37688 15552
rect 37240 15512 37246 15524
rect 30561 15487 30619 15493
rect 30561 15453 30573 15487
rect 30607 15484 30619 15487
rect 30607 15456 30641 15484
rect 30607 15453 30619 15456
rect 30561 15447 30619 15453
rect 30834 15444 30840 15496
rect 30892 15484 30898 15496
rect 31754 15484 31760 15496
rect 30892 15456 31760 15484
rect 30892 15444 30898 15456
rect 31754 15444 31760 15456
rect 31812 15444 31818 15496
rect 32582 15444 32588 15496
rect 32640 15444 32646 15496
rect 32677 15487 32735 15493
rect 32677 15453 32689 15487
rect 32723 15484 32735 15487
rect 33594 15484 33600 15496
rect 32723 15456 33600 15484
rect 32723 15453 32735 15456
rect 32677 15447 32735 15453
rect 33594 15444 33600 15456
rect 33652 15484 33658 15496
rect 33652 15456 35388 15484
rect 33652 15444 33658 15456
rect 35360 15428 35388 15456
rect 35618 15444 35624 15496
rect 35676 15484 35682 15496
rect 35676 15456 36216 15484
rect 35676 15444 35682 15456
rect 29825 15419 29883 15425
rect 29825 15416 29837 15419
rect 26712 15388 29837 15416
rect 29825 15385 29837 15388
rect 29871 15385 29883 15419
rect 29825 15379 29883 15385
rect 31202 15376 31208 15428
rect 31260 15416 31266 15428
rect 34054 15416 34060 15428
rect 31260 15388 34060 15416
rect 31260 15376 31266 15388
rect 34054 15376 34060 15388
rect 34112 15376 34118 15428
rect 35342 15376 35348 15428
rect 35400 15416 35406 15428
rect 35713 15419 35771 15425
rect 35713 15416 35725 15419
rect 35400 15388 35725 15416
rect 35400 15376 35406 15388
rect 35713 15385 35725 15388
rect 35759 15385 35771 15419
rect 35713 15379 35771 15385
rect 35805 15419 35863 15425
rect 35805 15385 35817 15419
rect 35851 15385 35863 15419
rect 35805 15379 35863 15385
rect 26326 15348 26332 15360
rect 23860 15320 26332 15348
rect 26326 15308 26332 15320
rect 26384 15308 26390 15360
rect 26878 15308 26884 15360
rect 26936 15348 26942 15360
rect 29730 15348 29736 15360
rect 26936 15320 29736 15348
rect 26936 15308 26942 15320
rect 29730 15308 29736 15320
rect 29788 15348 29794 15360
rect 30190 15348 30196 15360
rect 29788 15320 30196 15348
rect 29788 15308 29794 15320
rect 30190 15308 30196 15320
rect 30248 15308 30254 15360
rect 31662 15308 31668 15360
rect 31720 15348 31726 15360
rect 32306 15348 32312 15360
rect 31720 15320 32312 15348
rect 31720 15308 31726 15320
rect 32306 15308 32312 15320
rect 32364 15308 32370 15360
rect 34238 15308 34244 15360
rect 34296 15348 34302 15360
rect 34606 15348 34612 15360
rect 34296 15320 34612 15348
rect 34296 15308 34302 15320
rect 34606 15308 34612 15320
rect 34664 15308 34670 15360
rect 35618 15308 35624 15360
rect 35676 15348 35682 15360
rect 35820 15348 35848 15379
rect 35894 15376 35900 15428
rect 35952 15425 35958 15428
rect 35952 15419 36001 15425
rect 35952 15385 35955 15419
rect 35989 15416 36001 15419
rect 36078 15416 36084 15428
rect 35989 15388 36084 15416
rect 35989 15385 36001 15388
rect 35952 15379 36001 15385
rect 35952 15376 35958 15379
rect 36078 15376 36084 15388
rect 36136 15376 36142 15428
rect 36188 15416 36216 15456
rect 36998 15444 37004 15496
rect 37056 15484 37062 15496
rect 37458 15493 37464 15496
rect 37277 15487 37335 15493
rect 37277 15484 37289 15487
rect 37056 15456 37289 15484
rect 37056 15444 37062 15456
rect 37277 15453 37289 15456
rect 37323 15453 37335 15487
rect 37277 15447 37335 15453
rect 37425 15487 37464 15493
rect 37425 15453 37437 15487
rect 37425 15447 37464 15453
rect 37458 15444 37464 15447
rect 37516 15444 37522 15496
rect 37660 15493 37688 15524
rect 37645 15487 37703 15493
rect 37645 15453 37657 15487
rect 37691 15453 37703 15487
rect 37645 15447 37703 15453
rect 37783 15487 37841 15493
rect 37783 15453 37795 15487
rect 37829 15484 37841 15487
rect 38930 15484 38936 15496
rect 37829 15456 38936 15484
rect 37829 15453 37841 15456
rect 37783 15447 37841 15453
rect 38930 15444 38936 15456
rect 38988 15444 38994 15496
rect 39684 15484 39712 15648
rect 39758 15512 39764 15564
rect 39816 15552 39822 15564
rect 39945 15555 40003 15561
rect 39945 15552 39957 15555
rect 39816 15524 39957 15552
rect 39816 15512 39822 15524
rect 39945 15521 39957 15524
rect 39991 15521 40003 15555
rect 39945 15515 40003 15521
rect 39853 15487 39911 15493
rect 39853 15484 39865 15487
rect 39684 15456 39865 15484
rect 39853 15453 39865 15456
rect 39899 15453 39911 15487
rect 39853 15447 39911 15453
rect 40129 15487 40187 15493
rect 40129 15453 40141 15487
rect 40175 15453 40187 15487
rect 40129 15447 40187 15453
rect 37553 15419 37611 15425
rect 37553 15416 37565 15419
rect 36188 15388 37565 15416
rect 37553 15385 37565 15388
rect 37599 15416 37611 15419
rect 38378 15416 38384 15428
rect 37599 15388 38384 15416
rect 37599 15385 37611 15388
rect 37553 15379 37611 15385
rect 38378 15376 38384 15388
rect 38436 15376 38442 15428
rect 35676 15320 35848 15348
rect 35676 15308 35682 15320
rect 37182 15308 37188 15360
rect 37240 15348 37246 15360
rect 40144 15348 40172 15447
rect 37240 15320 40172 15348
rect 37240 15308 37246 15320
rect 1104 15258 41400 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 41400 15258
rect 1104 15184 41400 15206
rect 2038 15144 2044 15156
rect 1872 15116 2044 15144
rect 1872 15085 1900 15116
rect 2038 15104 2044 15116
rect 2096 15104 2102 15156
rect 3329 15147 3387 15153
rect 3329 15113 3341 15147
rect 3375 15144 3387 15147
rect 3694 15144 3700 15156
rect 3375 15116 3700 15144
rect 3375 15113 3387 15116
rect 3329 15107 3387 15113
rect 3694 15104 3700 15116
rect 3752 15104 3758 15156
rect 3970 15104 3976 15156
rect 4028 15144 4034 15156
rect 4028 15116 7972 15144
rect 4028 15104 4034 15116
rect 1857 15079 1915 15085
rect 1857 15045 1869 15079
rect 1903 15045 1915 15079
rect 3142 15076 3148 15088
rect 3082 15048 3148 15076
rect 1857 15039 1915 15045
rect 3142 15036 3148 15048
rect 3200 15076 3206 15088
rect 5626 15076 5632 15088
rect 3200 15048 5632 15076
rect 3200 15036 3206 15048
rect 5626 15036 5632 15048
rect 5684 15076 5690 15088
rect 7944 15076 7972 15116
rect 8018 15104 8024 15156
rect 8076 15144 8082 15156
rect 8113 15147 8171 15153
rect 8113 15144 8125 15147
rect 8076 15116 8125 15144
rect 8076 15104 8082 15116
rect 8113 15113 8125 15116
rect 8159 15113 8171 15147
rect 8113 15107 8171 15113
rect 10137 15147 10195 15153
rect 10137 15113 10149 15147
rect 10183 15144 10195 15147
rect 10778 15144 10784 15156
rect 10183 15116 10784 15144
rect 10183 15113 10195 15116
rect 10137 15107 10195 15113
rect 10778 15104 10784 15116
rect 10836 15104 10842 15156
rect 10962 15104 10968 15156
rect 11020 15104 11026 15156
rect 11422 15104 11428 15156
rect 11480 15104 11486 15156
rect 12069 15147 12127 15153
rect 12069 15113 12081 15147
rect 12115 15144 12127 15147
rect 12529 15147 12587 15153
rect 12529 15144 12541 15147
rect 12115 15116 12541 15144
rect 12115 15113 12127 15116
rect 12069 15107 12127 15113
rect 12529 15113 12541 15116
rect 12575 15113 12587 15147
rect 12529 15107 12587 15113
rect 12894 15104 12900 15156
rect 12952 15104 12958 15156
rect 15286 15104 15292 15156
rect 15344 15104 15350 15156
rect 15838 15104 15844 15156
rect 15896 15144 15902 15156
rect 19610 15144 19616 15156
rect 15896 15116 19616 15144
rect 15896 15104 15902 15116
rect 19610 15104 19616 15116
rect 19668 15104 19674 15156
rect 20162 15144 20168 15156
rect 19720 15116 20168 15144
rect 10229 15079 10287 15085
rect 5684 15048 7130 15076
rect 7944 15048 8248 15076
rect 5684 15036 5690 15048
rect 8220 15017 8248 15048
rect 10229 15045 10241 15079
rect 10275 15076 10287 15079
rect 11440 15076 11468 15104
rect 10275 15048 11468 15076
rect 12161 15079 12219 15085
rect 10275 15045 10287 15048
rect 10229 15039 10287 15045
rect 12161 15045 12173 15079
rect 12207 15076 12219 15079
rect 13630 15076 13636 15088
rect 12207 15048 13636 15076
rect 12207 15045 12219 15048
rect 12161 15039 12219 15045
rect 13630 15036 13636 15048
rect 13688 15036 13694 15088
rect 14645 15079 14703 15085
rect 14645 15045 14657 15079
rect 14691 15045 14703 15079
rect 14645 15039 14703 15045
rect 14737 15079 14795 15085
rect 14737 15045 14749 15079
rect 14783 15076 14795 15079
rect 15102 15076 15108 15088
rect 14783 15048 15108 15076
rect 14783 15045 14795 15048
rect 14737 15039 14795 15045
rect 8205 15011 8263 15017
rect 8205 14977 8217 15011
rect 8251 14977 8263 15011
rect 8205 14971 8263 14977
rect 8386 14968 8392 15020
rect 8444 14968 8450 15020
rect 8478 14968 8484 15020
rect 8536 14968 8542 15020
rect 8665 15011 8723 15017
rect 8665 14977 8677 15011
rect 8711 15008 8723 15011
rect 8711 14980 9674 15008
rect 8711 14977 8723 14980
rect 8665 14971 8723 14977
rect 1581 14943 1639 14949
rect 1581 14909 1593 14943
rect 1627 14909 1639 14943
rect 1581 14903 1639 14909
rect 1596 14816 1624 14903
rect 6270 14900 6276 14952
rect 6328 14940 6334 14952
rect 6365 14943 6423 14949
rect 6365 14940 6377 14943
rect 6328 14912 6377 14940
rect 6328 14900 6334 14912
rect 6365 14909 6377 14912
rect 6411 14909 6423 14943
rect 6365 14903 6423 14909
rect 6641 14943 6699 14949
rect 6641 14909 6653 14943
rect 6687 14940 6699 14943
rect 6730 14940 6736 14952
rect 6687 14912 6736 14940
rect 6687 14909 6699 14912
rect 6641 14903 6699 14909
rect 1578 14764 1584 14816
rect 1636 14764 1642 14816
rect 6380 14804 6408 14903
rect 6730 14900 6736 14912
rect 6788 14900 6794 14952
rect 8404 14940 8432 14968
rect 8680 14940 8708 14971
rect 8404 14912 8708 14940
rect 8297 14875 8355 14881
rect 8297 14841 8309 14875
rect 8343 14872 8355 14875
rect 9122 14872 9128 14884
rect 8343 14844 9128 14872
rect 8343 14841 8355 14844
rect 8297 14835 8355 14841
rect 9122 14832 9128 14844
rect 9180 14832 9186 14884
rect 9646 14872 9674 14980
rect 11054 14968 11060 15020
rect 11112 15008 11118 15020
rect 14458 15008 14464 15020
rect 11112 14980 13032 15008
rect 11112 14968 11118 14980
rect 10413 14943 10471 14949
rect 10413 14909 10425 14943
rect 10459 14940 10471 14943
rect 10778 14940 10784 14952
rect 10459 14912 10784 14940
rect 10459 14909 10471 14912
rect 10413 14903 10471 14909
rect 10778 14900 10784 14912
rect 10836 14900 10842 14952
rect 11146 14900 11152 14952
rect 11204 14900 11210 14952
rect 12345 14943 12403 14949
rect 12345 14909 12357 14943
rect 12391 14940 12403 14943
rect 12434 14940 12440 14952
rect 12391 14912 12440 14940
rect 12391 14909 12403 14912
rect 12345 14903 12403 14909
rect 12434 14900 12440 14912
rect 12492 14900 12498 14952
rect 13004 14949 13032 14980
rect 13924 14980 14464 15008
rect 12989 14943 13047 14949
rect 12989 14909 13001 14943
rect 13035 14940 13047 14943
rect 13173 14943 13231 14949
rect 13035 14912 13124 14940
rect 13035 14909 13047 14912
rect 12989 14903 13047 14909
rect 9646 14844 11100 14872
rect 11072 14816 11100 14844
rect 6638 14804 6644 14816
rect 6380 14776 6644 14804
rect 6638 14764 6644 14776
rect 6696 14764 6702 14816
rect 8570 14764 8576 14816
rect 8628 14764 8634 14816
rect 9398 14764 9404 14816
rect 9456 14804 9462 14816
rect 9769 14807 9827 14813
rect 9769 14804 9781 14807
rect 9456 14776 9781 14804
rect 9456 14764 9462 14776
rect 9769 14773 9781 14776
rect 9815 14773 9827 14807
rect 9769 14767 9827 14773
rect 10594 14764 10600 14816
rect 10652 14764 10658 14816
rect 11054 14764 11060 14816
rect 11112 14764 11118 14816
rect 11422 14764 11428 14816
rect 11480 14804 11486 14816
rect 11701 14807 11759 14813
rect 11701 14804 11713 14807
rect 11480 14776 11713 14804
rect 11480 14764 11486 14776
rect 11701 14773 11713 14776
rect 11747 14773 11759 14807
rect 11701 14767 11759 14773
rect 12894 14764 12900 14816
rect 12952 14804 12958 14816
rect 13096 14804 13124 14912
rect 13173 14909 13185 14943
rect 13219 14940 13231 14943
rect 13924 14940 13952 14980
rect 14458 14968 14464 14980
rect 14516 14968 14522 15020
rect 14660 15008 14688 15039
rect 15102 15036 15108 15048
rect 15160 15036 15166 15088
rect 16114 15036 16120 15088
rect 16172 15036 16178 15088
rect 16850 15036 16856 15088
rect 16908 15076 16914 15088
rect 16945 15079 17003 15085
rect 16945 15076 16957 15079
rect 16908 15048 16957 15076
rect 16908 15036 16914 15048
rect 16945 15045 16957 15048
rect 16991 15045 17003 15079
rect 16945 15039 17003 15045
rect 17218 15036 17224 15088
rect 17276 15076 17282 15088
rect 17276 15048 17434 15076
rect 17276 15036 17282 15048
rect 18322 15036 18328 15088
rect 18380 15076 18386 15088
rect 18782 15076 18788 15088
rect 18380 15048 18788 15076
rect 18380 15036 18386 15048
rect 18782 15036 18788 15048
rect 18840 15036 18846 15088
rect 19426 15076 19432 15088
rect 18984 15048 19432 15076
rect 15010 15008 15016 15020
rect 14660 14980 15016 15008
rect 15010 14968 15016 14980
rect 15068 14968 15074 15020
rect 16574 14968 16580 15020
rect 16632 15008 16638 15020
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 16632 14980 16681 15008
rect 16632 14968 16638 14980
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 13219 14912 13952 14940
rect 13219 14909 13231 14912
rect 13173 14903 13231 14909
rect 13998 14900 14004 14952
rect 14056 14940 14062 14952
rect 14167 14943 14225 14949
rect 14167 14940 14179 14943
rect 14056 14912 14179 14940
rect 14056 14900 14062 14912
rect 14167 14909 14179 14912
rect 14213 14909 14225 14943
rect 14167 14903 14225 14909
rect 14645 14943 14703 14949
rect 14645 14909 14657 14943
rect 14691 14940 14703 14943
rect 15381 14943 15439 14949
rect 14691 14912 14964 14940
rect 14691 14909 14703 14912
rect 14645 14903 14703 14909
rect 14936 14881 14964 14912
rect 15381 14909 15393 14943
rect 15427 14909 15439 14943
rect 15381 14903 15439 14909
rect 14921 14875 14979 14881
rect 14921 14841 14933 14875
rect 14967 14841 14979 14875
rect 14921 14835 14979 14841
rect 15396 14872 15424 14903
rect 15562 14900 15568 14952
rect 15620 14900 15626 14952
rect 16298 14900 16304 14952
rect 16356 14900 16362 14952
rect 16393 14943 16451 14949
rect 16393 14909 16405 14943
rect 16439 14940 16451 14943
rect 16942 14940 16948 14952
rect 16439 14912 16948 14940
rect 16439 14909 16451 14912
rect 16393 14903 16451 14909
rect 16942 14900 16948 14912
rect 17000 14900 17006 14952
rect 17310 14900 17316 14952
rect 17368 14940 17374 14952
rect 18984 14940 19012 15048
rect 19426 15036 19432 15048
rect 19484 15036 19490 15088
rect 19720 15085 19748 15116
rect 20162 15104 20168 15116
rect 20220 15104 20226 15156
rect 21177 15147 21235 15153
rect 21177 15113 21189 15147
rect 21223 15144 21235 15147
rect 21266 15144 21272 15156
rect 21223 15116 21272 15144
rect 21223 15113 21235 15116
rect 21177 15107 21235 15113
rect 21266 15104 21272 15116
rect 21324 15104 21330 15156
rect 22002 15144 22008 15156
rect 21744 15116 22008 15144
rect 19706 15079 19764 15085
rect 19706 15045 19718 15079
rect 19752 15045 19764 15079
rect 19706 15039 19764 15045
rect 19843 15079 19901 15085
rect 19843 15045 19855 15079
rect 19889 15076 19901 15079
rect 20346 15076 20352 15088
rect 19889 15048 20352 15076
rect 19889 15045 19901 15048
rect 19843 15039 19901 15045
rect 20346 15036 20352 15048
rect 20404 15036 20410 15088
rect 20898 15076 20904 15088
rect 20456 15048 20904 15076
rect 19518 14968 19524 15020
rect 19576 14968 19582 15020
rect 19614 15011 19672 15017
rect 19614 14977 19626 15011
rect 19660 14977 19672 15011
rect 19614 14971 19672 14977
rect 19981 15011 20039 15017
rect 19981 14977 19993 15011
rect 20027 15008 20039 15011
rect 20456 15008 20484 15048
rect 20898 15036 20904 15048
rect 20956 15036 20962 15088
rect 20027 14980 20484 15008
rect 20027 14977 20039 14980
rect 19981 14971 20039 14977
rect 19619 14940 19647 14971
rect 20806 14968 20812 15020
rect 20864 15008 20870 15020
rect 21085 15011 21143 15017
rect 21085 15008 21097 15011
rect 20864 14980 21097 15008
rect 20864 14968 20870 14980
rect 21085 14977 21097 14980
rect 21131 14977 21143 15011
rect 21085 14971 21143 14977
rect 21269 15011 21327 15017
rect 21269 14977 21281 15011
rect 21315 14977 21327 15011
rect 21269 14971 21327 14977
rect 21637 15011 21695 15017
rect 21637 14977 21649 15011
rect 21683 15008 21695 15011
rect 21744 15008 21772 15116
rect 22002 15104 22008 15116
rect 22060 15104 22066 15156
rect 22186 15104 22192 15156
rect 22244 15144 22250 15156
rect 22649 15147 22707 15153
rect 22649 15144 22661 15147
rect 22244 15116 22661 15144
rect 22244 15104 22250 15116
rect 22649 15113 22661 15116
rect 22695 15113 22707 15147
rect 22649 15107 22707 15113
rect 23658 15104 23664 15156
rect 23716 15104 23722 15156
rect 23845 15147 23903 15153
rect 23845 15113 23857 15147
rect 23891 15144 23903 15147
rect 26234 15144 26240 15156
rect 23891 15116 26240 15144
rect 23891 15113 23903 15116
rect 23845 15107 23903 15113
rect 26234 15104 26240 15116
rect 26292 15104 26298 15156
rect 26786 15104 26792 15156
rect 26844 15144 26850 15156
rect 26973 15147 27031 15153
rect 26973 15144 26985 15147
rect 26844 15116 26985 15144
rect 26844 15104 26850 15116
rect 26973 15113 26985 15116
rect 27019 15113 27031 15147
rect 26973 15107 27031 15113
rect 27062 15104 27068 15156
rect 27120 15104 27126 15156
rect 28442 15104 28448 15156
rect 28500 15104 28506 15156
rect 29270 15104 29276 15156
rect 29328 15104 29334 15156
rect 32214 15104 32220 15156
rect 32272 15104 32278 15156
rect 32398 15104 32404 15156
rect 32456 15144 32462 15156
rect 34057 15147 34115 15153
rect 32456 15116 33916 15144
rect 32456 15104 32462 15116
rect 21818 15036 21824 15088
rect 21876 15076 21882 15088
rect 23676 15076 23704 15104
rect 21876 15048 23612 15076
rect 23676 15048 24072 15076
rect 21876 15036 21882 15048
rect 21683 14980 21772 15008
rect 21683 14977 21695 14980
rect 21637 14971 21695 14977
rect 17368 14912 19012 14940
rect 19076 14912 19647 14940
rect 17368 14900 17374 14912
rect 16316 14872 16344 14900
rect 18417 14875 18475 14881
rect 18417 14872 18429 14875
rect 15396 14844 16344 14872
rect 17972 14844 18429 14872
rect 13354 14804 13360 14816
rect 12952 14776 13360 14804
rect 12952 14764 12958 14776
rect 13354 14764 13360 14776
rect 13412 14804 13418 14816
rect 15396 14804 15424 14844
rect 13412 14776 15424 14804
rect 13412 14764 13418 14776
rect 16482 14764 16488 14816
rect 16540 14804 16546 14816
rect 17310 14804 17316 14816
rect 16540 14776 17316 14804
rect 16540 14764 16546 14776
rect 17310 14764 17316 14776
rect 17368 14764 17374 14816
rect 17586 14764 17592 14816
rect 17644 14804 17650 14816
rect 17972 14804 18000 14844
rect 18417 14841 18429 14844
rect 18463 14872 18475 14875
rect 18690 14872 18696 14884
rect 18463 14844 18696 14872
rect 18463 14841 18475 14844
rect 18417 14835 18475 14841
rect 18690 14832 18696 14844
rect 18748 14832 18754 14884
rect 17644 14776 18000 14804
rect 17644 14764 17650 14776
rect 18322 14764 18328 14816
rect 18380 14804 18386 14816
rect 19076 14804 19104 14912
rect 19242 14832 19248 14884
rect 19300 14872 19306 14884
rect 21284 14872 21312 14971
rect 22002 14968 22008 15020
rect 22060 14968 22066 15020
rect 22373 15011 22431 15017
rect 22373 14977 22385 15011
rect 22419 15008 22431 15011
rect 22738 15008 22744 15020
rect 22419 14980 22744 15008
rect 22419 14977 22431 14980
rect 22373 14971 22431 14977
rect 22738 14968 22744 14980
rect 22796 14968 22802 15020
rect 22833 15011 22891 15017
rect 22833 14977 22845 15011
rect 22879 14977 22891 15011
rect 23584 15008 23612 15048
rect 23658 15008 23664 15020
rect 23584 14980 23664 15008
rect 22833 14971 22891 14977
rect 21913 14943 21971 14949
rect 21913 14940 21925 14943
rect 21468 14912 21925 14940
rect 21468 14881 21496 14912
rect 21913 14909 21925 14912
rect 21959 14940 21971 14943
rect 22848 14940 22876 14971
rect 23658 14968 23664 14980
rect 23716 14968 23722 15020
rect 23753 15011 23811 15017
rect 23753 14977 23765 15011
rect 23799 15008 23811 15011
rect 23934 15008 23940 15020
rect 23799 14980 23940 15008
rect 23799 14977 23811 14980
rect 23753 14971 23811 14977
rect 23934 14968 23940 14980
rect 23992 14968 23998 15020
rect 24044 15017 24072 15048
rect 25958 15036 25964 15088
rect 26016 15076 26022 15088
rect 27080 15076 27108 15104
rect 26016 15048 27108 15076
rect 27172 15048 28028 15076
rect 26016 15036 26022 15048
rect 24029 15011 24087 15017
rect 24029 14977 24041 15011
rect 24075 14977 24087 15011
rect 24029 14971 24087 14977
rect 24213 15011 24271 15017
rect 24213 14977 24225 15011
rect 24259 15008 24271 15011
rect 24302 15008 24308 15020
rect 24259 14980 24308 15008
rect 24259 14977 24271 14980
rect 24213 14971 24271 14977
rect 24302 14968 24308 14980
rect 24360 14968 24366 15020
rect 24394 14968 24400 15020
rect 24452 15008 24458 15020
rect 24489 15011 24547 15017
rect 24489 15008 24501 15011
rect 24452 14980 24501 15008
rect 24452 14968 24458 14980
rect 24489 14977 24501 14980
rect 24535 14977 24547 15011
rect 24489 14971 24547 14977
rect 26234 14968 26240 15020
rect 26292 15008 26298 15020
rect 27172 15017 27200 15048
rect 27157 15011 27215 15017
rect 27157 15008 27169 15011
rect 26292 14980 27169 15008
rect 26292 14968 26298 14980
rect 27157 14977 27169 14980
rect 27203 14977 27215 15011
rect 27157 14971 27215 14977
rect 27433 15011 27491 15017
rect 27433 14977 27445 15011
rect 27479 14977 27491 15011
rect 27433 14971 27491 14977
rect 27617 15011 27675 15017
rect 27617 14977 27629 15011
rect 27663 14977 27675 15011
rect 27617 14971 27675 14977
rect 24581 14943 24639 14949
rect 24581 14940 24593 14943
rect 21959 14912 22876 14940
rect 22940 14912 24593 14940
rect 21959 14909 21971 14912
rect 21913 14903 21971 14909
rect 19300 14844 21312 14872
rect 19300 14832 19306 14844
rect 18380 14776 19104 14804
rect 18380 14764 18386 14776
rect 19334 14764 19340 14816
rect 19392 14764 19398 14816
rect 19426 14764 19432 14816
rect 19484 14804 19490 14816
rect 20530 14804 20536 14816
rect 19484 14776 20536 14804
rect 19484 14764 19490 14776
rect 20530 14764 20536 14776
rect 20588 14764 20594 14816
rect 21284 14804 21312 14844
rect 21453 14875 21511 14881
rect 21453 14841 21465 14875
rect 21499 14841 21511 14875
rect 21453 14835 21511 14841
rect 21634 14832 21640 14884
rect 21692 14872 21698 14884
rect 22940 14872 22968 14912
rect 24581 14909 24593 14912
rect 24627 14909 24639 14943
rect 24581 14903 24639 14909
rect 25130 14900 25136 14952
rect 25188 14940 25194 14952
rect 25958 14940 25964 14952
rect 25188 14912 25964 14940
rect 25188 14900 25194 14912
rect 25958 14900 25964 14912
rect 26016 14900 26022 14952
rect 26510 14940 26516 14952
rect 26068 14912 26516 14940
rect 21692 14844 22968 14872
rect 23477 14875 23535 14881
rect 21692 14832 21698 14844
rect 23477 14841 23489 14875
rect 23523 14872 23535 14875
rect 24397 14875 24455 14881
rect 24397 14872 24409 14875
rect 23523 14844 24409 14872
rect 23523 14841 23535 14844
rect 23477 14835 23535 14841
rect 24397 14841 24409 14844
rect 24443 14841 24455 14875
rect 24397 14835 24455 14841
rect 24670 14832 24676 14884
rect 24728 14872 24734 14884
rect 26068 14872 26096 14912
rect 26510 14900 26516 14912
rect 26568 14940 26574 14952
rect 27448 14940 27476 14971
rect 26568 14912 27476 14940
rect 26568 14900 26574 14912
rect 27632 14884 27660 14971
rect 27890 14968 27896 15020
rect 27948 14968 27954 15020
rect 28000 15008 28028 15048
rect 28258 15036 28264 15088
rect 28316 15036 28322 15088
rect 29288 15076 29316 15104
rect 29822 15076 29828 15088
rect 29288 15048 29828 15076
rect 28902 15008 28908 15020
rect 28000 14980 28908 15008
rect 28902 14968 28908 14980
rect 28960 14968 28966 15020
rect 28997 15011 29055 15017
rect 28997 14977 29009 15011
rect 29043 15008 29055 15011
rect 29549 15011 29607 15017
rect 29549 15008 29561 15011
rect 29043 14980 29561 15008
rect 29043 14977 29055 14980
rect 28997 14971 29055 14977
rect 29549 14977 29561 14980
rect 29595 15008 29607 15011
rect 29638 15008 29644 15020
rect 29595 14980 29644 15008
rect 29595 14977 29607 14980
rect 29549 14971 29607 14977
rect 29638 14968 29644 14980
rect 29696 14968 29702 15020
rect 29748 15017 29776 15048
rect 29822 15036 29828 15048
rect 29880 15036 29886 15088
rect 29733 15011 29791 15017
rect 29733 14977 29745 15011
rect 29779 14977 29791 15011
rect 29733 14971 29791 14977
rect 31570 14968 31576 15020
rect 31628 15008 31634 15020
rect 31846 15008 31852 15020
rect 31628 14980 31852 15008
rect 31628 14968 31634 14980
rect 31846 14968 31852 14980
rect 31904 14968 31910 15020
rect 32232 15008 32260 15104
rect 33226 15036 33232 15088
rect 33284 15076 33290 15088
rect 33781 15079 33839 15085
rect 33781 15076 33793 15079
rect 33284 15048 33793 15076
rect 33284 15036 33290 15048
rect 33781 15045 33793 15048
rect 33827 15045 33839 15079
rect 33888 15076 33916 15116
rect 34057 15113 34069 15147
rect 34103 15144 34115 15147
rect 38654 15144 38660 15156
rect 34103 15116 38660 15144
rect 34103 15113 34115 15116
rect 34057 15107 34115 15113
rect 38654 15104 38660 15116
rect 38712 15104 38718 15156
rect 38746 15104 38752 15156
rect 38804 15144 38810 15156
rect 38841 15147 38899 15153
rect 38841 15144 38853 15147
rect 38804 15116 38853 15144
rect 38804 15104 38810 15116
rect 38841 15113 38853 15116
rect 38887 15113 38899 15147
rect 38841 15107 38899 15113
rect 34425 15079 34483 15085
rect 34425 15076 34437 15079
rect 33888 15048 34437 15076
rect 33781 15039 33839 15045
rect 34425 15045 34437 15048
rect 34471 15045 34483 15079
rect 34425 15039 34483 15045
rect 38120 15048 38332 15076
rect 38120 15020 38148 15048
rect 32309 15011 32367 15017
rect 32309 15008 32321 15011
rect 32232 14980 32321 15008
rect 32309 14977 32321 14980
rect 32355 14977 32367 15011
rect 32309 14971 32367 14977
rect 32401 15011 32459 15017
rect 32401 14977 32413 15011
rect 32447 14977 32459 15011
rect 32401 14971 32459 14977
rect 32493 15011 32551 15017
rect 32493 14977 32505 15011
rect 32539 14977 32551 15011
rect 32611 15011 32669 15017
rect 32611 15008 32623 15011
rect 32493 14971 32551 14977
rect 32600 14977 32623 15008
rect 32657 14977 32669 15011
rect 32600 14971 32669 14977
rect 28813 14943 28871 14949
rect 28813 14940 28825 14943
rect 27724 14912 28825 14940
rect 24728 14844 26096 14872
rect 24728 14832 24734 14844
rect 26142 14832 26148 14884
rect 26200 14872 26206 14884
rect 27154 14872 27160 14884
rect 26200 14844 27160 14872
rect 26200 14832 26206 14844
rect 27154 14832 27160 14844
rect 27212 14872 27218 14884
rect 27249 14875 27307 14881
rect 27249 14872 27261 14875
rect 27212 14844 27261 14872
rect 27212 14832 27218 14844
rect 27249 14841 27261 14844
rect 27295 14841 27307 14875
rect 27249 14835 27307 14841
rect 27338 14832 27344 14884
rect 27396 14832 27402 14884
rect 27614 14832 27620 14884
rect 27672 14832 27678 14884
rect 22002 14804 22008 14816
rect 21284 14776 22008 14804
rect 22002 14764 22008 14776
rect 22060 14764 22066 14816
rect 22278 14764 22284 14816
rect 22336 14764 22342 14816
rect 22554 14764 22560 14816
rect 22612 14764 22618 14816
rect 23290 14764 23296 14816
rect 23348 14764 23354 14816
rect 23566 14764 23572 14816
rect 23624 14764 23630 14816
rect 23658 14764 23664 14816
rect 23716 14764 23722 14816
rect 23750 14764 23756 14816
rect 23808 14804 23814 14816
rect 24118 14804 24124 14816
rect 23808 14776 24124 14804
rect 23808 14764 23814 14776
rect 24118 14764 24124 14776
rect 24176 14764 24182 14816
rect 24302 14764 24308 14816
rect 24360 14804 24366 14816
rect 27724 14804 27752 14912
rect 28813 14909 28825 14912
rect 28859 14909 28871 14943
rect 28813 14903 28871 14909
rect 29273 14943 29331 14949
rect 29273 14909 29285 14943
rect 29319 14940 29331 14943
rect 29454 14940 29460 14952
rect 29319 14912 29460 14940
rect 29319 14909 29331 14912
rect 29273 14903 29331 14909
rect 29454 14900 29460 14912
rect 29512 14900 29518 14952
rect 29825 14943 29883 14949
rect 29825 14909 29837 14943
rect 29871 14940 29883 14943
rect 29914 14940 29920 14952
rect 29871 14912 29920 14940
rect 29871 14909 29883 14912
rect 29825 14903 29883 14909
rect 29914 14900 29920 14912
rect 29972 14940 29978 14952
rect 30926 14940 30932 14952
rect 29972 14912 30932 14940
rect 29972 14900 29978 14912
rect 30926 14900 30932 14912
rect 30984 14900 30990 14952
rect 31864 14940 31892 14968
rect 32416 14940 32444 14971
rect 31864 14912 32444 14940
rect 29086 14872 29092 14884
rect 28276 14844 29092 14872
rect 28276 14813 28304 14844
rect 29086 14832 29092 14844
rect 29144 14832 29150 14884
rect 29178 14832 29184 14884
rect 29236 14872 29242 14884
rect 31662 14872 31668 14884
rect 29236 14844 31668 14872
rect 29236 14832 29242 14844
rect 31662 14832 31668 14844
rect 31720 14832 31726 14884
rect 31754 14832 31760 14884
rect 31812 14872 31818 14884
rect 32214 14872 32220 14884
rect 31812 14844 32220 14872
rect 31812 14832 31818 14844
rect 32214 14832 32220 14844
rect 32272 14872 32278 14884
rect 32508 14872 32536 14971
rect 32272 14844 32536 14872
rect 32600 14872 32628 14971
rect 32858 14968 32864 15020
rect 32916 15008 32922 15020
rect 33413 15011 33471 15017
rect 33413 15008 33425 15011
rect 32916 14980 33425 15008
rect 32916 14968 32922 14980
rect 33413 14977 33425 14980
rect 33459 14977 33471 15011
rect 33413 14971 33471 14977
rect 33506 15011 33564 15017
rect 33506 14977 33518 15011
rect 33552 14977 33564 15011
rect 33506 14971 33564 14977
rect 32766 14900 32772 14952
rect 32824 14900 32830 14952
rect 32674 14872 32680 14884
rect 32600 14844 32680 14872
rect 32272 14832 32278 14844
rect 32674 14832 32680 14844
rect 32732 14872 32738 14884
rect 33521 14872 33549 14971
rect 33594 14968 33600 15020
rect 33652 15008 33658 15020
rect 33689 15011 33747 15017
rect 33689 15008 33701 15011
rect 33652 14980 33701 15008
rect 33652 14968 33658 14980
rect 33689 14977 33701 14980
rect 33735 14977 33747 15011
rect 33689 14971 33747 14977
rect 33704 14940 33732 14971
rect 33870 14968 33876 15020
rect 33928 15017 33934 15020
rect 33928 15008 33936 15017
rect 34149 15011 34207 15017
rect 33928 14980 33973 15008
rect 33928 14971 33936 14980
rect 34149 14977 34161 15011
rect 34195 15008 34207 15011
rect 34238 15008 34244 15020
rect 34195 14980 34244 15008
rect 34195 14977 34207 14980
rect 34149 14971 34207 14977
rect 33928 14968 33934 14971
rect 34238 14968 34244 14980
rect 34296 14968 34302 15020
rect 34333 15011 34391 15017
rect 34333 14977 34345 15011
rect 34379 14977 34391 15011
rect 34517 15011 34575 15017
rect 34517 15008 34529 15011
rect 34333 14971 34391 14977
rect 34440 14980 34529 15008
rect 34348 14940 34376 14971
rect 34440 14952 34468 14980
rect 34517 14977 34529 14980
rect 34563 15008 34575 15011
rect 35250 15008 35256 15020
rect 34563 14980 35256 15008
rect 34563 14977 34575 14980
rect 34517 14971 34575 14977
rect 35250 14968 35256 14980
rect 35308 15008 35314 15020
rect 37642 15008 37648 15020
rect 35308 14980 37648 15008
rect 35308 14968 35314 14980
rect 37642 14968 37648 14980
rect 37700 14968 37706 15020
rect 38102 14968 38108 15020
rect 38160 14968 38166 15020
rect 38304 15017 38332 15048
rect 38378 15036 38384 15088
rect 38436 15076 38442 15088
rect 38473 15079 38531 15085
rect 38473 15076 38485 15079
rect 38436 15048 38485 15076
rect 38436 15036 38442 15048
rect 38473 15045 38485 15048
rect 38519 15045 38531 15079
rect 38473 15039 38531 15045
rect 38562 15036 38568 15088
rect 38620 15036 38626 15088
rect 38197 15011 38255 15017
rect 38197 14977 38209 15011
rect 38243 14977 38255 15011
rect 38197 14971 38255 14977
rect 38290 15011 38348 15017
rect 38290 14977 38302 15011
rect 38336 14977 38348 15011
rect 38290 14971 38348 14977
rect 38703 15011 38761 15017
rect 38703 14977 38715 15011
rect 38749 15008 38761 15011
rect 38930 15008 38936 15020
rect 38749 14980 38936 15008
rect 38749 14977 38761 14980
rect 38703 14971 38761 14977
rect 33704 14912 34376 14940
rect 34422 14900 34428 14952
rect 34480 14900 34486 14952
rect 35710 14900 35716 14952
rect 35768 14900 35774 14952
rect 38212 14940 38240 14971
rect 38930 14968 38936 14980
rect 38988 15008 38994 15020
rect 39390 15008 39396 15020
rect 38988 14980 39396 15008
rect 38988 14968 38994 14980
rect 39390 14968 39396 14980
rect 39448 14968 39454 15020
rect 38470 14940 38476 14952
rect 38212 14912 38476 14940
rect 38470 14900 38476 14912
rect 38528 14900 38534 14952
rect 35728 14872 35756 14900
rect 32732 14844 33272 14872
rect 33521 14844 35756 14872
rect 32732 14832 32738 14844
rect 24360 14776 27752 14804
rect 28261 14807 28319 14813
rect 24360 14764 24366 14776
rect 28261 14773 28273 14807
rect 28307 14773 28319 14807
rect 28261 14767 28319 14773
rect 28350 14764 28356 14816
rect 28408 14804 28414 14816
rect 29365 14807 29423 14813
rect 29365 14804 29377 14807
rect 28408 14776 29377 14804
rect 28408 14764 28414 14776
rect 29365 14773 29377 14776
rect 29411 14773 29423 14807
rect 29365 14767 29423 14773
rect 29914 14764 29920 14816
rect 29972 14804 29978 14816
rect 32030 14804 32036 14816
rect 29972 14776 32036 14804
rect 29972 14764 29978 14776
rect 32030 14764 32036 14776
rect 32088 14764 32094 14816
rect 32125 14807 32183 14813
rect 32125 14773 32137 14807
rect 32171 14804 32183 14807
rect 33134 14804 33140 14816
rect 32171 14776 33140 14804
rect 32171 14773 32183 14776
rect 32125 14767 32183 14773
rect 33134 14764 33140 14776
rect 33192 14764 33198 14816
rect 33244 14804 33272 14844
rect 34422 14804 34428 14816
rect 33244 14776 34428 14804
rect 34422 14764 34428 14776
rect 34480 14764 34486 14816
rect 34701 14807 34759 14813
rect 34701 14773 34713 14807
rect 34747 14804 34759 14807
rect 36998 14804 37004 14816
rect 34747 14776 37004 14804
rect 34747 14773 34759 14776
rect 34701 14767 34759 14773
rect 36998 14764 37004 14776
rect 37056 14764 37062 14816
rect 1104 14714 41400 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 41400 14714
rect 1104 14640 41400 14662
rect 4062 14560 4068 14612
rect 4120 14600 4126 14612
rect 8478 14600 8484 14612
rect 4120 14572 8484 14600
rect 4120 14560 4126 14572
rect 8478 14560 8484 14572
rect 8536 14560 8542 14612
rect 14829 14603 14887 14609
rect 12406 14572 14780 14600
rect 12406 14532 12434 14572
rect 3344 14504 12434 14532
rect 14185 14535 14243 14541
rect 3234 14424 3240 14476
rect 3292 14424 3298 14476
rect 3344 14473 3372 14504
rect 14185 14501 14197 14535
rect 14231 14532 14243 14535
rect 14642 14532 14648 14544
rect 14231 14504 14648 14532
rect 14231 14501 14243 14504
rect 14185 14495 14243 14501
rect 14642 14492 14648 14504
rect 14700 14492 14706 14544
rect 14752 14532 14780 14572
rect 14829 14569 14841 14603
rect 14875 14600 14887 14603
rect 14918 14600 14924 14612
rect 14875 14572 14924 14600
rect 14875 14569 14887 14572
rect 14829 14563 14887 14569
rect 14918 14560 14924 14572
rect 14976 14560 14982 14612
rect 16022 14560 16028 14612
rect 16080 14600 16086 14612
rect 16482 14600 16488 14612
rect 16080 14572 16488 14600
rect 16080 14560 16086 14572
rect 16482 14560 16488 14572
rect 16540 14560 16546 14612
rect 16942 14560 16948 14612
rect 17000 14600 17006 14612
rect 17678 14600 17684 14612
rect 17000 14572 17684 14600
rect 17000 14560 17006 14572
rect 17678 14560 17684 14572
rect 17736 14600 17742 14612
rect 17773 14603 17831 14609
rect 17773 14600 17785 14603
rect 17736 14572 17785 14600
rect 17736 14560 17742 14572
rect 17773 14569 17785 14572
rect 17819 14569 17831 14603
rect 17773 14563 17831 14569
rect 17954 14560 17960 14612
rect 18012 14600 18018 14612
rect 18138 14600 18144 14612
rect 18012 14572 18144 14600
rect 18012 14560 18018 14572
rect 18138 14560 18144 14572
rect 18196 14600 18202 14612
rect 18509 14603 18567 14609
rect 18509 14600 18521 14603
rect 18196 14572 18521 14600
rect 18196 14560 18202 14572
rect 18509 14569 18521 14572
rect 18555 14600 18567 14603
rect 18555 14572 19564 14600
rect 18555 14569 18567 14572
rect 18509 14563 18567 14569
rect 15562 14532 15568 14544
rect 14752 14504 15568 14532
rect 15562 14492 15568 14504
rect 15620 14532 15626 14544
rect 17494 14532 17500 14544
rect 15620 14504 17500 14532
rect 15620 14492 15626 14504
rect 17494 14492 17500 14504
rect 17552 14492 17558 14544
rect 19245 14535 19303 14541
rect 19245 14501 19257 14535
rect 19291 14532 19303 14535
rect 19426 14532 19432 14544
rect 19291 14504 19432 14532
rect 19291 14501 19303 14504
rect 19245 14495 19303 14501
rect 19426 14492 19432 14504
rect 19484 14492 19490 14544
rect 19536 14532 19564 14572
rect 19610 14560 19616 14612
rect 19668 14560 19674 14612
rect 20622 14600 20628 14612
rect 19721 14572 20628 14600
rect 19721 14532 19749 14572
rect 20622 14560 20628 14572
rect 20680 14560 20686 14612
rect 23658 14560 23664 14612
rect 23716 14600 23722 14612
rect 25317 14603 25375 14609
rect 25317 14600 25329 14603
rect 23716 14572 25329 14600
rect 23716 14560 23722 14572
rect 25317 14569 25329 14572
rect 25363 14569 25375 14603
rect 25317 14563 25375 14569
rect 25774 14560 25780 14612
rect 25832 14560 25838 14612
rect 26697 14603 26755 14609
rect 26697 14569 26709 14603
rect 26743 14600 26755 14603
rect 26878 14600 26884 14612
rect 26743 14572 26884 14600
rect 26743 14569 26755 14572
rect 26697 14563 26755 14569
rect 26878 14560 26884 14572
rect 26936 14560 26942 14612
rect 26973 14603 27031 14609
rect 26973 14569 26985 14603
rect 27019 14600 27031 14603
rect 27062 14600 27068 14612
rect 27019 14572 27068 14600
rect 27019 14569 27031 14572
rect 26973 14563 27031 14569
rect 19536 14504 19749 14532
rect 19794 14492 19800 14544
rect 19852 14532 19858 14544
rect 19889 14535 19947 14541
rect 19889 14532 19901 14535
rect 19852 14504 19901 14532
rect 19852 14492 19858 14504
rect 19889 14501 19901 14504
rect 19935 14501 19947 14535
rect 19889 14495 19947 14501
rect 19978 14492 19984 14544
rect 20036 14532 20042 14544
rect 20441 14535 20499 14541
rect 20441 14532 20453 14535
rect 20036 14504 20453 14532
rect 20036 14492 20042 14504
rect 20441 14501 20453 14504
rect 20487 14501 20499 14535
rect 20441 14495 20499 14501
rect 21266 14492 21272 14544
rect 21324 14532 21330 14544
rect 21729 14535 21787 14541
rect 21729 14532 21741 14535
rect 21324 14504 21741 14532
rect 21324 14492 21330 14504
rect 21729 14501 21741 14504
rect 21775 14501 21787 14535
rect 22554 14532 22560 14544
rect 21729 14495 21787 14501
rect 22066 14504 22560 14532
rect 3329 14467 3387 14473
rect 3329 14433 3341 14467
rect 3375 14433 3387 14467
rect 3329 14427 3387 14433
rect 3513 14467 3571 14473
rect 3513 14433 3525 14467
rect 3559 14464 3571 14467
rect 6270 14464 6276 14476
rect 3559 14436 6276 14464
rect 3559 14433 3571 14436
rect 3513 14427 3571 14433
rect 6270 14424 6276 14436
rect 6328 14424 6334 14476
rect 7101 14467 7159 14473
rect 7101 14433 7113 14467
rect 7147 14464 7159 14467
rect 7926 14464 7932 14476
rect 7147 14436 7932 14464
rect 7147 14433 7159 14436
rect 7101 14427 7159 14433
rect 7926 14424 7932 14436
rect 7984 14424 7990 14476
rect 9214 14424 9220 14476
rect 9272 14464 9278 14476
rect 9272 14436 10824 14464
rect 9272 14424 9278 14436
rect 3252 14396 3280 14424
rect 3789 14399 3847 14405
rect 3789 14396 3801 14399
rect 3252 14368 3801 14396
rect 3789 14365 3801 14368
rect 3835 14365 3847 14399
rect 3789 14359 3847 14365
rect 10594 14356 10600 14408
rect 10652 14396 10658 14408
rect 10689 14399 10747 14405
rect 10689 14396 10701 14399
rect 10652 14368 10701 14396
rect 10652 14356 10658 14368
rect 10689 14365 10701 14368
rect 10735 14365 10747 14399
rect 10796 14396 10824 14436
rect 10962 14424 10968 14476
rect 11020 14464 11026 14476
rect 12434 14464 12440 14476
rect 11020 14436 12440 14464
rect 11020 14424 11026 14436
rect 12434 14424 12440 14436
rect 12492 14424 12498 14476
rect 18969 14467 19027 14473
rect 14200 14436 15424 14464
rect 11793 14399 11851 14405
rect 11793 14396 11805 14399
rect 10796 14368 11805 14396
rect 10689 14359 10747 14365
rect 11793 14365 11805 14368
rect 11839 14365 11851 14399
rect 11793 14359 11851 14365
rect 11977 14399 12035 14405
rect 11977 14365 11989 14399
rect 12023 14365 12035 14399
rect 11977 14359 12035 14365
rect 3237 14331 3295 14337
rect 3237 14297 3249 14331
rect 3283 14328 3295 14331
rect 4433 14331 4491 14337
rect 4433 14328 4445 14331
rect 3283 14300 4445 14328
rect 3283 14297 3295 14300
rect 3237 14291 3295 14297
rect 4433 14297 4445 14300
rect 4479 14297 4491 14331
rect 4433 14291 4491 14297
rect 7834 14288 7840 14340
rect 7892 14328 7898 14340
rect 9858 14328 9864 14340
rect 7892 14300 9864 14328
rect 7892 14288 7898 14300
rect 9858 14288 9864 14300
rect 9916 14288 9922 14340
rect 10870 14288 10876 14340
rect 10928 14288 10934 14340
rect 11054 14288 11060 14340
rect 11112 14328 11118 14340
rect 11992 14328 12020 14359
rect 12250 14328 12256 14340
rect 11112 14300 12256 14328
rect 11112 14288 11118 14300
rect 12250 14288 12256 14300
rect 12308 14288 12314 14340
rect 14200 14337 14228 14436
rect 14274 14356 14280 14408
rect 14332 14396 14338 14408
rect 14461 14399 14519 14405
rect 14461 14396 14473 14399
rect 14332 14368 14473 14396
rect 14332 14356 14338 14368
rect 14461 14365 14473 14368
rect 14507 14365 14519 14399
rect 14461 14359 14519 14365
rect 14553 14399 14611 14405
rect 14553 14365 14565 14399
rect 14599 14396 14611 14399
rect 14918 14396 14924 14408
rect 14599 14368 14924 14396
rect 14599 14365 14611 14368
rect 14553 14359 14611 14365
rect 14185 14331 14243 14337
rect 14185 14328 14197 14331
rect 12406 14300 14197 14328
rect 2774 14220 2780 14272
rect 2832 14260 2838 14272
rect 2869 14263 2927 14269
rect 2869 14260 2881 14263
rect 2832 14232 2881 14260
rect 2832 14220 2838 14232
rect 2869 14229 2881 14232
rect 2915 14229 2927 14263
rect 2869 14223 2927 14229
rect 7650 14220 7656 14272
rect 7708 14220 7714 14272
rect 9030 14220 9036 14272
rect 9088 14260 9094 14272
rect 10321 14263 10379 14269
rect 10321 14260 10333 14263
rect 9088 14232 10333 14260
rect 9088 14220 9094 14232
rect 10321 14229 10333 14232
rect 10367 14229 10379 14263
rect 10321 14223 10379 14229
rect 10781 14263 10839 14269
rect 10781 14229 10793 14263
rect 10827 14260 10839 14263
rect 10888 14260 10916 14288
rect 10827 14232 10916 14260
rect 10827 14229 10839 14232
rect 10781 14223 10839 14229
rect 11974 14220 11980 14272
rect 12032 14260 12038 14272
rect 12406 14260 12434 14300
rect 14185 14297 14197 14300
rect 14231 14297 14243 14331
rect 14476 14328 14504 14359
rect 14918 14356 14924 14368
rect 14976 14356 14982 14408
rect 15396 14405 15424 14436
rect 17328 14436 18184 14464
rect 17328 14405 17356 14436
rect 15289 14399 15347 14405
rect 15289 14396 15301 14399
rect 15212 14368 15301 14396
rect 15105 14331 15163 14337
rect 15105 14328 15117 14331
rect 14476 14300 15117 14328
rect 14185 14291 14243 14297
rect 15105 14297 15117 14300
rect 15151 14297 15163 14331
rect 15105 14291 15163 14297
rect 12032 14232 12434 14260
rect 14369 14263 14427 14269
rect 12032 14220 12038 14232
rect 14369 14229 14381 14263
rect 14415 14260 14427 14263
rect 15013 14263 15071 14269
rect 15013 14260 15025 14263
rect 14415 14232 15025 14260
rect 14415 14229 14427 14232
rect 14369 14223 14427 14229
rect 15013 14229 15025 14232
rect 15059 14260 15071 14263
rect 15212 14260 15240 14368
rect 15289 14365 15301 14368
rect 15335 14365 15347 14399
rect 15289 14359 15347 14365
rect 15381 14399 15439 14405
rect 15381 14365 15393 14399
rect 15427 14365 15439 14399
rect 15381 14359 15439 14365
rect 17313 14399 17371 14405
rect 17313 14365 17325 14399
rect 17359 14365 17371 14399
rect 17313 14359 17371 14365
rect 17402 14356 17408 14408
rect 17460 14396 17466 14408
rect 17497 14399 17555 14405
rect 17497 14396 17509 14399
rect 17460 14368 17509 14396
rect 17460 14356 17466 14368
rect 17497 14365 17509 14368
rect 17543 14365 17555 14399
rect 17954 14396 17960 14408
rect 17497 14359 17555 14365
rect 17820 14368 17960 14396
rect 17586 14288 17592 14340
rect 17644 14288 17650 14340
rect 17820 14337 17848 14368
rect 17954 14356 17960 14368
rect 18012 14356 18018 14408
rect 18156 14337 18184 14436
rect 18969 14433 18981 14467
rect 19015 14464 19027 14467
rect 22066 14464 22094 14504
rect 22554 14492 22560 14504
rect 22612 14492 22618 14544
rect 23566 14492 23572 14544
rect 23624 14532 23630 14544
rect 24302 14532 24308 14544
rect 23624 14504 24308 14532
rect 23624 14492 23630 14504
rect 24302 14492 24308 14504
rect 24360 14492 24366 14544
rect 24394 14492 24400 14544
rect 24452 14492 24458 14544
rect 26237 14535 26295 14541
rect 26237 14532 26249 14535
rect 25792 14504 26249 14532
rect 23750 14464 23756 14476
rect 19015 14436 21680 14464
rect 19015 14433 19027 14436
rect 18969 14427 19027 14433
rect 18325 14399 18383 14405
rect 18325 14365 18337 14399
rect 18371 14396 18383 14399
rect 18414 14396 18420 14408
rect 18371 14368 18420 14396
rect 18371 14365 18383 14368
rect 18325 14359 18383 14365
rect 18414 14356 18420 14368
rect 18472 14356 18478 14408
rect 18785 14399 18843 14405
rect 18785 14365 18797 14399
rect 18831 14396 18843 14399
rect 18874 14396 18880 14408
rect 18831 14368 18880 14396
rect 18831 14365 18843 14368
rect 18785 14359 18843 14365
rect 18874 14356 18880 14368
rect 18932 14356 18938 14408
rect 19061 14399 19119 14405
rect 19061 14365 19073 14399
rect 19107 14396 19119 14399
rect 19242 14396 19248 14408
rect 19107 14368 19248 14396
rect 19107 14365 19119 14368
rect 19061 14359 19119 14365
rect 19242 14356 19248 14368
rect 19300 14356 19306 14408
rect 20042 14399 20100 14405
rect 19352 14368 19932 14396
rect 17805 14331 17863 14337
rect 17805 14297 17817 14331
rect 17851 14297 17863 14331
rect 17805 14291 17863 14297
rect 18141 14331 18199 14337
rect 18141 14297 18153 14331
rect 18187 14328 18199 14331
rect 19352 14328 19380 14368
rect 18187 14300 19380 14328
rect 18187 14297 18199 14300
rect 18141 14291 18199 14297
rect 19426 14288 19432 14340
rect 19484 14328 19490 14340
rect 19904 14328 19932 14368
rect 20042 14365 20054 14399
rect 20088 14396 20100 14399
rect 20346 14396 20352 14408
rect 20088 14368 20352 14396
rect 20088 14365 20100 14368
rect 20042 14359 20100 14365
rect 20346 14356 20352 14368
rect 20404 14356 20410 14408
rect 20530 14356 20536 14408
rect 20588 14356 20594 14408
rect 20139 14331 20197 14337
rect 19484 14300 19840 14328
rect 19904 14300 20085 14328
rect 19484 14288 19490 14300
rect 15059 14232 15240 14260
rect 15059 14229 15071 14232
rect 15013 14223 15071 14229
rect 15286 14220 15292 14272
rect 15344 14220 15350 14272
rect 17402 14220 17408 14272
rect 17460 14220 17466 14272
rect 17954 14220 17960 14272
rect 18012 14220 18018 14272
rect 18414 14220 18420 14272
rect 18472 14260 18478 14272
rect 18601 14263 18659 14269
rect 18601 14260 18613 14263
rect 18472 14232 18613 14260
rect 18472 14220 18478 14232
rect 18601 14229 18613 14232
rect 18647 14229 18659 14263
rect 18601 14223 18659 14229
rect 18690 14220 18696 14272
rect 18748 14260 18754 14272
rect 19058 14260 19064 14272
rect 18748 14232 19064 14260
rect 18748 14220 18754 14232
rect 19058 14220 19064 14232
rect 19116 14260 19122 14272
rect 19812 14269 19840 14300
rect 19613 14263 19671 14269
rect 19613 14260 19625 14263
rect 19116 14232 19625 14260
rect 19116 14220 19122 14232
rect 19613 14229 19625 14232
rect 19659 14229 19671 14263
rect 19613 14223 19671 14229
rect 19797 14263 19855 14269
rect 19797 14229 19809 14263
rect 19843 14229 19855 14263
rect 20057 14260 20085 14300
rect 20139 14297 20151 14331
rect 20185 14328 20197 14331
rect 20714 14328 20720 14340
rect 20185 14300 20720 14328
rect 20185 14297 20197 14300
rect 20139 14291 20197 14297
rect 20714 14288 20720 14300
rect 20772 14288 20778 14340
rect 21652 14328 21680 14436
rect 21744 14436 22094 14464
rect 23124 14436 23756 14464
rect 21744 14405 21772 14436
rect 21729 14399 21787 14405
rect 21729 14365 21741 14399
rect 21775 14365 21787 14399
rect 21729 14359 21787 14365
rect 21821 14399 21879 14405
rect 21821 14365 21833 14399
rect 21867 14396 21879 14399
rect 23124 14396 23152 14436
rect 23750 14424 23756 14436
rect 23808 14424 23814 14476
rect 24118 14424 24124 14476
rect 24176 14464 24182 14476
rect 24412 14464 24440 14492
rect 24176 14436 24440 14464
rect 24504 14436 25544 14464
rect 24176 14424 24182 14436
rect 21867 14368 23152 14396
rect 23201 14399 23259 14405
rect 21867 14365 21879 14368
rect 21821 14359 21879 14365
rect 23201 14365 23213 14399
rect 23247 14396 23259 14399
rect 23290 14396 23296 14408
rect 23247 14368 23296 14396
rect 23247 14365 23259 14368
rect 23201 14359 23259 14365
rect 23290 14356 23296 14368
rect 23348 14356 23354 14408
rect 24504 14396 24532 14436
rect 25516 14408 25544 14436
rect 25792 14408 25820 14504
rect 26237 14501 26249 14504
rect 26283 14501 26295 14535
rect 26237 14495 26295 14501
rect 26605 14535 26663 14541
rect 26605 14501 26617 14535
rect 26651 14532 26663 14535
rect 26988 14532 27016 14563
rect 27062 14560 27068 14572
rect 27120 14560 27126 14612
rect 27430 14560 27436 14612
rect 27488 14560 27494 14612
rect 27617 14603 27675 14609
rect 27617 14569 27629 14603
rect 27663 14600 27675 14603
rect 27890 14600 27896 14612
rect 27663 14572 27896 14600
rect 27663 14569 27675 14572
rect 27617 14563 27675 14569
rect 27890 14560 27896 14572
rect 27948 14560 27954 14612
rect 29178 14560 29184 14612
rect 29236 14560 29242 14612
rect 30650 14560 30656 14612
rect 30708 14600 30714 14612
rect 33413 14603 33471 14609
rect 30708 14572 31754 14600
rect 30708 14560 30714 14572
rect 26651 14504 27016 14532
rect 27448 14532 27476 14560
rect 28258 14532 28264 14544
rect 27448 14504 28264 14532
rect 26651 14501 26663 14504
rect 26605 14495 26663 14501
rect 23400 14368 24532 14396
rect 22005 14331 22063 14337
rect 22005 14328 22017 14331
rect 21652 14300 22017 14328
rect 22005 14297 22017 14300
rect 22051 14328 22063 14331
rect 22738 14328 22744 14340
rect 22051 14300 22744 14328
rect 22051 14297 22063 14300
rect 22005 14291 22063 14297
rect 22738 14288 22744 14300
rect 22796 14288 22802 14340
rect 23400 14328 23428 14368
rect 24670 14356 24676 14408
rect 24728 14356 24734 14408
rect 24946 14356 24952 14408
rect 25004 14396 25010 14408
rect 25004 14368 25452 14396
rect 25004 14356 25010 14368
rect 22848 14300 23428 14328
rect 24397 14331 24455 14337
rect 22848 14260 22876 14300
rect 24397 14297 24409 14331
rect 24443 14328 24455 14331
rect 24486 14328 24492 14340
rect 24443 14300 24492 14328
rect 24443 14297 24455 14300
rect 24397 14291 24455 14297
rect 24486 14288 24492 14300
rect 24544 14328 24550 14340
rect 24762 14328 24768 14340
rect 24544 14300 24768 14328
rect 24544 14288 24550 14300
rect 24762 14288 24768 14300
rect 24820 14288 24826 14340
rect 25222 14288 25228 14340
rect 25280 14328 25286 14340
rect 25317 14331 25375 14337
rect 25317 14328 25329 14331
rect 25280 14300 25329 14328
rect 25280 14288 25286 14300
rect 25317 14297 25329 14300
rect 25363 14297 25375 14331
rect 25424 14328 25452 14368
rect 25498 14356 25504 14408
rect 25556 14356 25562 14408
rect 25593 14399 25651 14405
rect 25593 14365 25605 14399
rect 25639 14365 25651 14399
rect 25593 14359 25651 14365
rect 25608 14328 25636 14359
rect 25774 14356 25780 14408
rect 25832 14356 25838 14408
rect 25958 14356 25964 14408
rect 26016 14356 26022 14408
rect 26252 14396 26280 14495
rect 28258 14492 28264 14504
rect 28316 14492 28322 14544
rect 26421 14467 26479 14473
rect 26421 14433 26433 14467
rect 26467 14464 26479 14467
rect 26789 14467 26847 14473
rect 26467 14436 26740 14464
rect 26467 14433 26479 14436
rect 26421 14427 26479 14433
rect 26513 14399 26571 14405
rect 26513 14396 26525 14399
rect 26252 14368 26525 14396
rect 26513 14365 26525 14368
rect 26559 14365 26571 14399
rect 26712 14396 26740 14436
rect 26789 14433 26801 14467
rect 26835 14464 26847 14467
rect 27157 14467 27215 14473
rect 27157 14464 27169 14467
rect 26835 14436 27169 14464
rect 26835 14433 26847 14436
rect 26789 14427 26847 14433
rect 27157 14433 27169 14436
rect 27203 14433 27215 14467
rect 27157 14427 27215 14433
rect 26881 14399 26939 14405
rect 26881 14396 26893 14399
rect 26712 14368 26893 14396
rect 26513 14359 26571 14365
rect 26881 14365 26893 14368
rect 26927 14365 26939 14399
rect 27172 14396 27200 14427
rect 27890 14424 27896 14476
rect 27948 14464 27954 14476
rect 28813 14467 28871 14473
rect 28813 14464 28825 14467
rect 27948 14436 28825 14464
rect 27948 14424 27954 14436
rect 28813 14433 28825 14436
rect 28859 14433 28871 14467
rect 28813 14427 28871 14433
rect 27706 14396 27712 14408
rect 27172 14368 27712 14396
rect 26881 14359 26939 14365
rect 27706 14356 27712 14368
rect 27764 14356 27770 14408
rect 28997 14399 29055 14405
rect 28997 14365 29009 14399
rect 29043 14396 29055 14399
rect 29196 14396 29224 14560
rect 31478 14492 31484 14544
rect 31536 14492 31542 14544
rect 31496 14464 31524 14492
rect 31726 14464 31754 14572
rect 33413 14569 33425 14603
rect 33459 14600 33471 14603
rect 33686 14600 33692 14612
rect 33459 14572 33692 14600
rect 33459 14569 33471 14572
rect 33413 14563 33471 14569
rect 33686 14560 33692 14572
rect 33744 14560 33750 14612
rect 35986 14560 35992 14612
rect 36044 14600 36050 14612
rect 36262 14600 36268 14612
rect 36044 14572 36268 14600
rect 36044 14560 36050 14572
rect 36262 14560 36268 14572
rect 36320 14560 36326 14612
rect 36633 14603 36691 14609
rect 36633 14569 36645 14603
rect 36679 14600 36691 14603
rect 37090 14600 37096 14612
rect 36679 14572 37096 14600
rect 36679 14569 36691 14572
rect 36633 14563 36691 14569
rect 37090 14560 37096 14572
rect 37148 14560 37154 14612
rect 38194 14560 38200 14612
rect 38252 14560 38258 14612
rect 38654 14560 38660 14612
rect 38712 14560 38718 14612
rect 39025 14603 39083 14609
rect 39025 14569 39037 14603
rect 39071 14600 39083 14603
rect 39758 14600 39764 14612
rect 39071 14572 39764 14600
rect 39071 14569 39083 14572
rect 39025 14563 39083 14569
rect 39758 14560 39764 14572
rect 39816 14560 39822 14612
rect 39853 14603 39911 14609
rect 39853 14569 39865 14603
rect 39899 14569 39911 14603
rect 39853 14563 39911 14569
rect 31938 14492 31944 14544
rect 31996 14492 32002 14544
rect 38212 14532 38240 14560
rect 39868 14532 39896 14563
rect 40310 14560 40316 14612
rect 40368 14560 40374 14612
rect 34624 14504 36860 14532
rect 38212 14504 39896 14532
rect 34624 14476 34652 14504
rect 34057 14467 34115 14473
rect 34057 14464 34069 14467
rect 31496 14436 31616 14464
rect 31726 14436 34069 14464
rect 31588 14408 31616 14436
rect 34057 14433 34069 14436
rect 34103 14433 34115 14467
rect 34330 14464 34336 14476
rect 34057 14427 34115 14433
rect 34169 14436 34336 14464
rect 29043 14368 29224 14396
rect 29043 14365 29055 14368
rect 28997 14359 29055 14365
rect 30374 14356 30380 14408
rect 30432 14396 30438 14408
rect 30653 14399 30711 14405
rect 30653 14396 30665 14399
rect 30432 14368 30665 14396
rect 30432 14356 30438 14368
rect 30653 14365 30665 14368
rect 30699 14365 30711 14399
rect 30653 14359 30711 14365
rect 30834 14356 30840 14408
rect 30892 14356 30898 14408
rect 30926 14356 30932 14408
rect 30984 14356 30990 14408
rect 31018 14356 31024 14408
rect 31076 14356 31082 14408
rect 31294 14356 31300 14408
rect 31352 14356 31358 14408
rect 31478 14405 31484 14408
rect 31445 14399 31484 14405
rect 31445 14365 31457 14399
rect 31445 14359 31484 14365
rect 31478 14356 31484 14359
rect 31536 14356 31542 14408
rect 31570 14356 31576 14408
rect 31628 14356 31634 14408
rect 31662 14356 31668 14408
rect 31720 14356 31726 14408
rect 31803 14399 31861 14405
rect 31803 14365 31815 14399
rect 31849 14396 31861 14399
rect 32398 14396 32404 14408
rect 31849 14368 32404 14396
rect 31849 14365 31861 14368
rect 31803 14359 31861 14365
rect 32398 14356 32404 14368
rect 32456 14356 32462 14408
rect 32490 14356 32496 14408
rect 32548 14356 32554 14408
rect 33410 14356 33416 14408
rect 33468 14396 33474 14408
rect 33597 14399 33655 14405
rect 33597 14396 33609 14399
rect 33468 14368 33609 14396
rect 33468 14356 33474 14368
rect 33597 14365 33609 14368
rect 33643 14365 33655 14399
rect 33597 14359 33655 14365
rect 33919 14399 33977 14405
rect 33919 14365 33931 14399
rect 33965 14396 33977 14399
rect 34169 14396 34197 14436
rect 34330 14424 34336 14436
rect 34388 14424 34394 14476
rect 34606 14424 34612 14476
rect 34664 14424 34670 14476
rect 34900 14436 35572 14464
rect 33965 14368 34197 14396
rect 33965 14365 33977 14368
rect 33919 14359 33977 14365
rect 34238 14356 34244 14408
rect 34296 14396 34302 14408
rect 34900 14405 34928 14436
rect 34885 14399 34943 14405
rect 34296 14368 34744 14396
rect 34296 14356 34302 14368
rect 26694 14328 26700 14340
rect 25424 14300 26700 14328
rect 25317 14291 25375 14297
rect 26694 14288 26700 14300
rect 26752 14288 26758 14340
rect 27280 14331 27338 14337
rect 27280 14328 27292 14331
rect 26804 14300 27292 14328
rect 20057 14232 22876 14260
rect 19797 14223 19855 14229
rect 23014 14220 23020 14272
rect 23072 14220 23078 14272
rect 24581 14263 24639 14269
rect 24581 14229 24593 14263
rect 24627 14260 24639 14263
rect 25406 14260 25412 14272
rect 24627 14232 25412 14260
rect 24627 14229 24639 14232
rect 24581 14223 24639 14229
rect 25406 14220 25412 14232
rect 25464 14220 25470 14272
rect 25866 14220 25872 14272
rect 25924 14260 25930 14272
rect 26804 14260 26832 14300
rect 27280 14297 27292 14300
rect 27326 14328 27338 14331
rect 27326 14300 27660 14328
rect 27326 14297 27338 14300
rect 27280 14291 27338 14297
rect 25924 14232 26832 14260
rect 27157 14263 27215 14269
rect 25924 14220 25930 14232
rect 27157 14229 27169 14263
rect 27203 14260 27215 14263
rect 27430 14260 27436 14272
rect 27203 14232 27436 14260
rect 27203 14229 27215 14232
rect 27157 14223 27215 14229
rect 27430 14220 27436 14232
rect 27488 14220 27494 14272
rect 27632 14260 27660 14300
rect 27798 14288 27804 14340
rect 27856 14328 27862 14340
rect 29181 14331 29239 14337
rect 29181 14328 29193 14331
rect 27856 14300 29193 14328
rect 27856 14288 27862 14300
rect 29181 14297 29193 14300
rect 29227 14297 29239 14331
rect 29181 14291 29239 14297
rect 30558 14288 30564 14340
rect 30616 14328 30622 14340
rect 32508 14328 32536 14356
rect 33686 14328 33692 14340
rect 30616 14300 33692 14328
rect 30616 14288 30622 14300
rect 33686 14288 33692 14300
rect 33744 14288 33750 14340
rect 33781 14331 33839 14337
rect 33781 14297 33793 14331
rect 33827 14328 33839 14331
rect 34422 14328 34428 14340
rect 33827 14300 34428 14328
rect 33827 14297 33839 14300
rect 33781 14291 33839 14297
rect 33980 14272 34008 14300
rect 34422 14288 34428 14300
rect 34480 14288 34486 14340
rect 34716 14328 34744 14368
rect 34885 14365 34897 14399
rect 34931 14365 34943 14399
rect 34885 14359 34943 14365
rect 35345 14399 35403 14405
rect 35345 14365 35357 14399
rect 35391 14396 35403 14399
rect 35434 14396 35440 14408
rect 35391 14368 35440 14396
rect 35391 14365 35403 14368
rect 35345 14359 35403 14365
rect 35434 14356 35440 14368
rect 35492 14356 35498 14408
rect 35544 14340 35572 14436
rect 36832 14405 36860 14504
rect 38746 14424 38752 14476
rect 38804 14424 38810 14476
rect 39942 14424 39948 14476
rect 40000 14424 40006 14476
rect 36817 14399 36875 14405
rect 36817 14365 36829 14399
rect 36863 14365 36875 14399
rect 36817 14359 36875 14365
rect 36906 14356 36912 14408
rect 36964 14356 36970 14408
rect 36998 14356 37004 14408
rect 37056 14396 37062 14408
rect 37093 14399 37151 14405
rect 37093 14396 37105 14399
rect 37056 14368 37105 14396
rect 37056 14356 37062 14368
rect 37093 14365 37105 14368
rect 37139 14365 37151 14399
rect 37093 14359 37151 14365
rect 37185 14399 37243 14405
rect 37185 14365 37197 14399
rect 37231 14396 37243 14399
rect 37826 14396 37832 14408
rect 37231 14368 37832 14396
rect 37231 14365 37243 14368
rect 37185 14359 37243 14365
rect 37826 14356 37832 14368
rect 37884 14396 37890 14408
rect 38565 14399 38623 14405
rect 38565 14396 38577 14399
rect 37884 14368 38577 14396
rect 37884 14356 37890 14368
rect 38565 14365 38577 14368
rect 38611 14365 38623 14399
rect 38565 14359 38623 14365
rect 38838 14356 38844 14408
rect 38896 14396 38902 14408
rect 39206 14396 39212 14408
rect 38896 14368 39212 14396
rect 38896 14356 38902 14368
rect 39206 14356 39212 14368
rect 39264 14356 39270 14408
rect 40034 14356 40040 14408
rect 40092 14396 40098 14408
rect 40129 14399 40187 14405
rect 40129 14396 40141 14399
rect 40092 14368 40141 14396
rect 40092 14356 40098 14368
rect 40129 14365 40141 14368
rect 40175 14365 40187 14399
rect 40129 14359 40187 14365
rect 34977 14331 35035 14337
rect 34977 14328 34989 14331
rect 34716 14300 34989 14328
rect 34977 14297 34989 14300
rect 35023 14297 35035 14331
rect 34977 14291 35035 14297
rect 35066 14288 35072 14340
rect 35124 14288 35130 14340
rect 35158 14288 35164 14340
rect 35216 14337 35222 14340
rect 35216 14331 35245 14337
rect 35233 14297 35245 14331
rect 35216 14291 35245 14297
rect 35216 14288 35222 14291
rect 35526 14288 35532 14340
rect 35584 14288 35590 14340
rect 35618 14288 35624 14340
rect 35676 14328 35682 14340
rect 35986 14328 35992 14340
rect 35676 14300 35992 14328
rect 35676 14288 35682 14300
rect 35986 14288 35992 14300
rect 36044 14288 36050 14340
rect 39853 14331 39911 14337
rect 39853 14297 39865 14331
rect 39899 14297 39911 14331
rect 39853 14291 39911 14297
rect 28166 14260 28172 14272
rect 27632 14232 28172 14260
rect 28166 14220 28172 14232
rect 28224 14220 28230 14272
rect 28534 14220 28540 14272
rect 28592 14260 28598 14272
rect 28902 14260 28908 14272
rect 28592 14232 28908 14260
rect 28592 14220 28598 14232
rect 28902 14220 28908 14232
rect 28960 14260 28966 14272
rect 30190 14260 30196 14272
rect 28960 14232 30196 14260
rect 28960 14220 28966 14232
rect 30190 14220 30196 14232
rect 30248 14220 30254 14272
rect 31205 14263 31263 14269
rect 31205 14229 31217 14263
rect 31251 14260 31263 14263
rect 31294 14260 31300 14272
rect 31251 14232 31300 14260
rect 31251 14229 31263 14232
rect 31205 14223 31263 14229
rect 31294 14220 31300 14232
rect 31352 14260 31358 14272
rect 32122 14260 32128 14272
rect 31352 14232 32128 14260
rect 31352 14220 31358 14232
rect 32122 14220 32128 14232
rect 32180 14220 32186 14272
rect 32766 14220 32772 14272
rect 32824 14260 32830 14272
rect 33594 14260 33600 14272
rect 32824 14232 33600 14260
rect 32824 14220 32830 14232
rect 33594 14220 33600 14232
rect 33652 14220 33658 14272
rect 33962 14220 33968 14272
rect 34020 14220 34026 14272
rect 34698 14220 34704 14272
rect 34756 14260 34762 14272
rect 39868 14260 39896 14291
rect 34756 14232 39896 14260
rect 34756 14220 34762 14232
rect 1104 14170 41400 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 41400 14170
rect 1104 14096 41400 14118
rect 1578 14056 1584 14068
rect 1504 14028 1584 14056
rect 1504 13929 1532 14028
rect 1578 14016 1584 14028
rect 1636 14056 1642 14068
rect 3510 14056 3516 14068
rect 1636 14028 3516 14056
rect 1636 14016 1642 14028
rect 3510 14016 3516 14028
rect 3568 14016 3574 14068
rect 6730 14016 6736 14068
rect 6788 14056 6794 14068
rect 6917 14059 6975 14065
rect 6917 14056 6929 14059
rect 6788 14028 6929 14056
rect 6788 14016 6794 14028
rect 6917 14025 6929 14028
rect 6963 14025 6975 14059
rect 6917 14019 6975 14025
rect 7650 14016 7656 14068
rect 7708 14016 7714 14068
rect 9493 14059 9551 14065
rect 7944 14028 9444 14056
rect 3142 13988 3148 14000
rect 2990 13960 3148 13988
rect 3142 13948 3148 13960
rect 3200 13948 3206 14000
rect 3234 13948 3240 14000
rect 3292 13948 3298 14000
rect 3528 13988 3556 14016
rect 5626 13988 5632 14000
rect 3436 13960 3556 13988
rect 4922 13960 5632 13988
rect 1489 13923 1547 13929
rect 1489 13889 1501 13923
rect 1535 13889 1547 13923
rect 1489 13883 1547 13889
rect 1762 13812 1768 13864
rect 1820 13812 1826 13864
rect 3252 13861 3280 13948
rect 3436 13929 3464 13960
rect 5626 13948 5632 13960
rect 5684 13948 5690 14000
rect 6641 13991 6699 13997
rect 6641 13957 6653 13991
rect 6687 13988 6699 13991
rect 7668 13988 7696 14016
rect 6687 13960 7696 13988
rect 6687 13957 6699 13960
rect 6641 13951 6699 13957
rect 7944 13932 7972 14028
rect 8021 13991 8079 13997
rect 8021 13957 8033 13991
rect 8067 13988 8079 13991
rect 8067 13960 8708 13988
rect 8067 13957 8079 13960
rect 8021 13951 8079 13957
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13889 3479 13923
rect 3421 13883 3479 13889
rect 5350 13880 5356 13932
rect 5408 13880 5414 13932
rect 6365 13923 6423 13929
rect 6365 13889 6377 13923
rect 6411 13889 6423 13923
rect 6365 13883 6423 13889
rect 3237 13855 3295 13861
rect 3237 13821 3249 13855
rect 3283 13821 3295 13855
rect 3237 13815 3295 13821
rect 3694 13812 3700 13864
rect 3752 13812 3758 13864
rect 5169 13855 5227 13861
rect 5169 13821 5181 13855
rect 5215 13852 5227 13855
rect 5368 13852 5396 13880
rect 5215 13824 5396 13852
rect 6380 13852 6408 13883
rect 6546 13880 6552 13932
rect 6604 13880 6610 13932
rect 6730 13880 6736 13932
rect 6788 13880 6794 13932
rect 7745 13923 7803 13929
rect 7745 13889 7757 13923
rect 7791 13920 7803 13923
rect 7834 13920 7840 13932
rect 7791 13892 7840 13920
rect 7791 13889 7803 13892
rect 7745 13883 7803 13889
rect 7834 13880 7840 13892
rect 7892 13880 7898 13932
rect 7926 13880 7932 13932
rect 7984 13880 7990 13932
rect 8680 13929 8708 13960
rect 8846 13948 8852 14000
rect 8904 13948 8910 14000
rect 9030 13948 9036 14000
rect 9088 13948 9094 14000
rect 9416 13988 9444 14028
rect 9493 14025 9505 14059
rect 9539 14056 9551 14059
rect 9858 14056 9864 14068
rect 9539 14028 9864 14056
rect 9539 14025 9551 14028
rect 9493 14019 9551 14025
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 12253 14059 12311 14065
rect 12253 14025 12265 14059
rect 12299 14056 12311 14059
rect 12299 14028 18552 14056
rect 12299 14025 12311 14028
rect 12253 14019 12311 14025
rect 10045 13991 10103 13997
rect 10045 13988 10057 13991
rect 9416 13960 10057 13988
rect 10045 13957 10057 13960
rect 10091 13988 10103 13991
rect 12342 13988 12348 14000
rect 10091 13960 12348 13988
rect 10091 13957 10103 13960
rect 10045 13951 10103 13957
rect 12342 13948 12348 13960
rect 12400 13988 12406 14000
rect 13170 13988 13176 14000
rect 12400 13960 13176 13988
rect 12400 13948 12406 13960
rect 13170 13948 13176 13960
rect 13228 13948 13234 14000
rect 16574 13948 16580 14000
rect 16632 13988 16638 14000
rect 17405 13991 17463 13997
rect 17405 13988 17417 13991
rect 16632 13960 17417 13988
rect 16632 13948 16638 13960
rect 17405 13957 17417 13960
rect 17451 13957 17463 13991
rect 17405 13951 17463 13957
rect 17696 13960 18460 13988
rect 8205 13923 8263 13929
rect 8205 13889 8217 13923
rect 8251 13920 8263 13923
rect 8665 13923 8723 13929
rect 8251 13892 8524 13920
rect 8251 13889 8263 13892
rect 8205 13883 8263 13889
rect 7098 13852 7104 13864
rect 6380 13824 7104 13852
rect 5215 13821 5227 13824
rect 5169 13815 5227 13821
rect 7098 13812 7104 13824
rect 7156 13812 7162 13864
rect 8496 13861 8524 13892
rect 8665 13889 8677 13923
rect 8711 13920 8723 13923
rect 9048 13920 9076 13948
rect 17696 13932 17724 13960
rect 8711 13892 9076 13920
rect 8711 13889 8723 13892
rect 8665 13883 8723 13889
rect 9122 13880 9128 13932
rect 9180 13920 9186 13932
rect 9309 13923 9367 13929
rect 9309 13920 9321 13923
rect 9180 13892 9321 13920
rect 9180 13880 9186 13892
rect 9309 13889 9321 13892
rect 9355 13889 9367 13923
rect 9309 13883 9367 13889
rect 8481 13855 8539 13861
rect 8481 13821 8493 13855
rect 8527 13852 8539 13855
rect 8570 13852 8576 13864
rect 8527 13824 8576 13852
rect 8527 13821 8539 13824
rect 8481 13815 8539 13821
rect 8570 13812 8576 13824
rect 8628 13852 8634 13864
rect 9214 13852 9220 13864
rect 8628 13824 9220 13852
rect 8628 13812 8634 13824
rect 9214 13812 9220 13824
rect 9272 13812 9278 13864
rect 9324 13852 9352 13883
rect 9398 13880 9404 13932
rect 9456 13920 9462 13932
rect 9861 13923 9919 13929
rect 9861 13920 9873 13923
rect 9456 13892 9873 13920
rect 9456 13880 9462 13892
rect 9861 13889 9873 13892
rect 9907 13889 9919 13923
rect 9861 13883 9919 13889
rect 12158 13880 12164 13932
rect 12216 13920 12222 13932
rect 12216 13892 12756 13920
rect 12216 13880 12222 13892
rect 9490 13852 9496 13864
rect 9324 13824 9496 13852
rect 9490 13812 9496 13824
rect 9548 13852 9554 13864
rect 12728 13861 12756 13892
rect 12802 13880 12808 13932
rect 12860 13880 12866 13932
rect 12986 13880 12992 13932
rect 13044 13880 13050 13932
rect 16669 13923 16727 13929
rect 16669 13889 16681 13923
rect 16715 13920 16727 13923
rect 16758 13920 16764 13932
rect 16715 13892 16764 13920
rect 16715 13889 16727 13892
rect 16669 13883 16727 13889
rect 16758 13880 16764 13892
rect 16816 13880 16822 13932
rect 17678 13880 17684 13932
rect 17736 13880 17742 13932
rect 17788 13892 18000 13920
rect 9677 13855 9735 13861
rect 9677 13852 9689 13855
rect 9548 13824 9689 13852
rect 9548 13812 9554 13824
rect 9677 13821 9689 13824
rect 9723 13821 9735 13855
rect 9677 13815 9735 13821
rect 12713 13855 12771 13861
rect 12713 13821 12725 13855
rect 12759 13852 12771 13855
rect 13078 13852 13084 13864
rect 12759 13824 13084 13852
rect 12759 13821 12771 13824
rect 12713 13815 12771 13821
rect 13078 13812 13084 13824
rect 13136 13812 13142 13864
rect 17788 13852 17816 13892
rect 16776 13824 17816 13852
rect 17865 13855 17923 13861
rect 5534 13744 5540 13796
rect 5592 13784 5598 13796
rect 5592 13756 6868 13784
rect 5592 13744 5598 13756
rect 6840 13728 6868 13756
rect 7282 13744 7288 13796
rect 7340 13784 7346 13796
rect 7745 13787 7803 13793
rect 7745 13784 7757 13787
rect 7340 13756 7757 13784
rect 7340 13744 7346 13756
rect 7745 13753 7757 13756
rect 7791 13784 7803 13787
rect 7791 13756 8616 13784
rect 7791 13753 7803 13756
rect 7745 13747 7803 13753
rect 5994 13676 6000 13728
rect 6052 13676 6058 13728
rect 6822 13676 6828 13728
rect 6880 13676 6886 13728
rect 7006 13676 7012 13728
rect 7064 13716 7070 13728
rect 8297 13719 8355 13725
rect 8297 13716 8309 13719
rect 7064 13688 8309 13716
rect 7064 13676 7070 13688
rect 8297 13685 8309 13688
rect 8343 13716 8355 13719
rect 8478 13716 8484 13728
rect 8343 13688 8484 13716
rect 8343 13685 8355 13688
rect 8297 13679 8355 13685
rect 8478 13676 8484 13688
rect 8536 13676 8542 13728
rect 8588 13716 8616 13756
rect 8662 13744 8668 13796
rect 8720 13784 8726 13796
rect 12066 13784 12072 13796
rect 8720 13756 12072 13784
rect 8720 13744 8726 13756
rect 12066 13744 12072 13756
rect 12124 13744 12130 13796
rect 12529 13787 12587 13793
rect 12529 13753 12541 13787
rect 12575 13784 12587 13787
rect 16776 13784 16804 13824
rect 17865 13821 17877 13855
rect 17911 13821 17923 13855
rect 17972 13852 18000 13892
rect 18138 13880 18144 13932
rect 18196 13920 18202 13932
rect 18432 13929 18460 13960
rect 18524 13929 18552 14028
rect 19334 14016 19340 14068
rect 19392 14016 19398 14068
rect 20441 14059 20499 14065
rect 20441 14025 20453 14059
rect 20487 14056 20499 14059
rect 20714 14056 20720 14068
rect 20487 14028 20720 14056
rect 20487 14025 20499 14028
rect 20441 14019 20499 14025
rect 19352 13988 19380 14016
rect 20456 13988 20484 14019
rect 20714 14016 20720 14028
rect 20772 14016 20778 14068
rect 22002 14016 22008 14068
rect 22060 14056 22066 14068
rect 24946 14056 24952 14068
rect 22060 14028 24952 14056
rect 22060 14016 22066 14028
rect 24946 14016 24952 14028
rect 25004 14016 25010 14068
rect 25774 14016 25780 14068
rect 25832 14016 25838 14068
rect 27338 14056 27344 14068
rect 26436 14028 27344 14056
rect 22830 13988 22836 14000
rect 18892 13960 19380 13988
rect 19444 13960 20484 13988
rect 20640 13960 22836 13988
rect 18892 13929 18920 13960
rect 19444 13929 19472 13960
rect 18233 13923 18291 13929
rect 18233 13920 18245 13923
rect 18196 13892 18245 13920
rect 18196 13880 18202 13892
rect 18233 13889 18245 13892
rect 18279 13889 18291 13923
rect 18233 13883 18291 13889
rect 18417 13923 18475 13929
rect 18417 13889 18429 13923
rect 18463 13889 18475 13923
rect 18417 13883 18475 13889
rect 18509 13923 18567 13929
rect 18509 13889 18521 13923
rect 18555 13889 18567 13923
rect 18509 13883 18567 13889
rect 18877 13923 18935 13929
rect 18877 13889 18889 13923
rect 18923 13889 18935 13923
rect 18877 13883 18935 13889
rect 19429 13923 19487 13929
rect 19429 13889 19441 13923
rect 19475 13889 19487 13923
rect 19429 13883 19487 13889
rect 19794 13880 19800 13932
rect 19852 13880 19858 13932
rect 19978 13880 19984 13932
rect 20036 13880 20042 13932
rect 20640 13929 20668 13960
rect 22830 13948 22836 13960
rect 22888 13948 22894 14000
rect 25038 13948 25044 14000
rect 25096 13988 25102 14000
rect 25096 13960 25820 13988
rect 25096 13948 25102 13960
rect 25792 13932 25820 13960
rect 20625 13923 20683 13929
rect 20625 13889 20637 13923
rect 20671 13889 20683 13923
rect 20625 13883 20683 13889
rect 20809 13923 20867 13929
rect 20809 13889 20821 13923
rect 20855 13889 20867 13923
rect 20809 13883 20867 13889
rect 18322 13852 18328 13864
rect 17972 13824 18328 13852
rect 17865 13815 17923 13821
rect 12575 13756 16804 13784
rect 12575 13753 12587 13756
rect 12529 13747 12587 13753
rect 17310 13744 17316 13796
rect 17368 13784 17374 13796
rect 17880 13784 17908 13815
rect 18322 13812 18328 13824
rect 18380 13812 18386 13864
rect 19521 13855 19579 13861
rect 19521 13821 19533 13855
rect 19567 13852 19579 13855
rect 19702 13852 19708 13864
rect 19567 13824 19708 13852
rect 19567 13821 19579 13824
rect 19521 13815 19579 13821
rect 19702 13812 19708 13824
rect 19760 13812 19766 13864
rect 19996 13852 20024 13880
rect 20824 13852 20852 13883
rect 25590 13880 25596 13932
rect 25648 13920 25654 13932
rect 25685 13923 25743 13929
rect 25685 13920 25697 13923
rect 25648 13892 25697 13920
rect 25648 13880 25654 13892
rect 25685 13889 25697 13892
rect 25731 13889 25743 13923
rect 25685 13883 25743 13889
rect 25774 13880 25780 13932
rect 25832 13920 25838 13932
rect 26436 13929 26464 14028
rect 27338 14016 27344 14028
rect 27396 14016 27402 14068
rect 27706 14016 27712 14068
rect 27764 14016 27770 14068
rect 27798 14016 27804 14068
rect 27856 14056 27862 14068
rect 27856 14028 28028 14056
rect 27856 14016 27862 14028
rect 28000 13997 28028 14028
rect 28074 14016 28080 14068
rect 28132 14056 28138 14068
rect 28353 14059 28411 14065
rect 28353 14056 28365 14059
rect 28132 14028 28365 14056
rect 28132 14016 28138 14028
rect 28353 14025 28365 14028
rect 28399 14025 28411 14059
rect 28353 14019 28411 14025
rect 28442 14016 28448 14068
rect 28500 14056 28506 14068
rect 28629 14059 28687 14065
rect 28629 14056 28641 14059
rect 28500 14028 28641 14056
rect 28500 14016 28506 14028
rect 28629 14025 28641 14028
rect 28675 14025 28687 14059
rect 28629 14019 28687 14025
rect 29362 14016 29368 14068
rect 29420 14016 29426 14068
rect 29549 14059 29607 14065
rect 29549 14025 29561 14059
rect 29595 14025 29607 14059
rect 29549 14019 29607 14025
rect 26789 13991 26847 13997
rect 26789 13957 26801 13991
rect 26835 13988 26847 13991
rect 27985 13991 28043 13997
rect 26835 13960 27108 13988
rect 26835 13957 26847 13960
rect 26789 13951 26847 13957
rect 27080 13932 27108 13960
rect 27985 13957 27997 13991
rect 28031 13957 28043 13991
rect 29380 13988 29408 14016
rect 27985 13951 28043 13957
rect 28828 13960 29408 13988
rect 29564 13988 29592 14019
rect 29914 14016 29920 14068
rect 29972 14016 29978 14068
rect 30466 14016 30472 14068
rect 30524 14056 30530 14068
rect 30524 14028 31248 14056
rect 30524 14016 30530 14028
rect 31220 13997 31248 14028
rect 31386 14016 31392 14068
rect 31444 14056 31450 14068
rect 31573 14059 31631 14065
rect 31573 14056 31585 14059
rect 31444 14028 31585 14056
rect 31444 14016 31450 14028
rect 31573 14025 31585 14028
rect 31619 14056 31631 14059
rect 31619 14028 32168 14056
rect 31619 14025 31631 14028
rect 31573 14019 31631 14025
rect 31205 13991 31263 13997
rect 29564 13960 31156 13988
rect 25869 13923 25927 13929
rect 25869 13920 25881 13923
rect 25832 13892 25881 13920
rect 25832 13880 25838 13892
rect 25869 13889 25881 13892
rect 25915 13889 25927 13923
rect 25869 13883 25927 13889
rect 26421 13923 26479 13929
rect 26421 13889 26433 13923
rect 26467 13920 26479 13923
rect 26510 13920 26516 13932
rect 26467 13892 26516 13920
rect 26467 13889 26479 13892
rect 26421 13883 26479 13889
rect 26510 13880 26516 13892
rect 26568 13880 26574 13932
rect 26970 13880 26976 13932
rect 27028 13880 27034 13932
rect 27062 13880 27068 13932
rect 27120 13880 27126 13932
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13920 27215 13923
rect 27258 13923 27316 13929
rect 27203 13889 27228 13920
rect 27157 13883 27228 13889
rect 27258 13889 27270 13923
rect 27304 13920 27316 13923
rect 27525 13923 27583 13929
rect 27304 13892 27476 13920
rect 27304 13889 27316 13892
rect 27258 13883 27316 13889
rect 19996 13824 20852 13852
rect 26329 13855 26387 13861
rect 26329 13821 26341 13855
rect 26375 13821 26387 13855
rect 27200 13852 27228 13883
rect 26329 13815 26387 13821
rect 26620 13824 27228 13852
rect 27341 13855 27399 13861
rect 18690 13784 18696 13796
rect 17368 13756 18696 13784
rect 17368 13744 17374 13756
rect 18690 13744 18696 13756
rect 18748 13744 18754 13796
rect 18892 13756 19472 13784
rect 10226 13716 10232 13728
rect 8588 13688 10232 13716
rect 10226 13676 10232 13688
rect 10284 13676 10290 13728
rect 12621 13719 12679 13725
rect 12621 13685 12633 13719
rect 12667 13716 12679 13719
rect 13538 13716 13544 13728
rect 12667 13688 13544 13716
rect 12667 13685 12679 13688
rect 12621 13679 12679 13685
rect 13538 13676 13544 13688
rect 13596 13676 13602 13728
rect 14826 13676 14832 13728
rect 14884 13716 14890 13728
rect 18046 13716 18052 13728
rect 14884 13688 18052 13716
rect 14884 13676 14890 13688
rect 18046 13676 18052 13688
rect 18104 13676 18110 13728
rect 18892 13725 18920 13756
rect 19444 13728 19472 13756
rect 20806 13744 20812 13796
rect 20864 13784 20870 13796
rect 25222 13784 25228 13796
rect 20864 13756 25228 13784
rect 20864 13744 20870 13756
rect 25222 13744 25228 13756
rect 25280 13744 25286 13796
rect 18877 13719 18935 13725
rect 18877 13685 18889 13719
rect 18923 13685 18935 13719
rect 18877 13679 18935 13685
rect 19058 13676 19064 13728
rect 19116 13676 19122 13728
rect 19426 13676 19432 13728
rect 19484 13676 19490 13728
rect 26344 13716 26372 13815
rect 26620 13796 26648 13824
rect 27341 13821 27353 13855
rect 27387 13821 27399 13855
rect 27448 13852 27476 13892
rect 27525 13889 27537 13923
rect 27571 13920 27583 13923
rect 27801 13923 27859 13929
rect 27801 13920 27813 13923
rect 27571 13892 27813 13920
rect 27571 13889 27583 13892
rect 27525 13883 27583 13889
rect 27724 13864 27752 13892
rect 27801 13889 27813 13892
rect 27847 13889 27859 13923
rect 27801 13883 27859 13889
rect 28069 13923 28127 13929
rect 28069 13889 28081 13923
rect 28115 13889 28127 13923
rect 28069 13883 28127 13889
rect 27614 13852 27620 13864
rect 27448 13824 27620 13852
rect 27341 13815 27399 13821
rect 26418 13744 26424 13796
rect 26476 13744 26482 13796
rect 26602 13744 26608 13796
rect 26660 13744 26666 13796
rect 26786 13744 26792 13796
rect 26844 13784 26850 13796
rect 27356 13784 27384 13815
rect 27614 13812 27620 13824
rect 27672 13812 27678 13864
rect 27706 13812 27712 13864
rect 27764 13812 27770 13864
rect 26844 13756 27384 13784
rect 28092 13784 28120 13883
rect 28166 13880 28172 13932
rect 28224 13880 28230 13932
rect 28828 13929 28856 13960
rect 28813 13923 28871 13929
rect 28813 13889 28825 13923
rect 28859 13889 28871 13923
rect 28813 13883 28871 13889
rect 28902 13880 28908 13932
rect 28960 13920 28966 13932
rect 28997 13923 29055 13929
rect 28997 13920 29009 13923
rect 28960 13892 29009 13920
rect 28960 13880 28966 13892
rect 28997 13889 29009 13892
rect 29043 13889 29055 13923
rect 28997 13883 29055 13889
rect 29089 13923 29147 13929
rect 29089 13889 29101 13923
rect 29135 13920 29147 13923
rect 29730 13920 29736 13932
rect 29135 13892 29736 13920
rect 29135 13889 29147 13892
rect 29089 13883 29147 13889
rect 29730 13880 29736 13892
rect 29788 13880 29794 13932
rect 29914 13880 29920 13932
rect 29972 13880 29978 13932
rect 31018 13880 31024 13932
rect 31076 13880 31082 13932
rect 29932 13852 29960 13880
rect 28966 13824 29960 13852
rect 28966 13784 28994 13824
rect 30006 13812 30012 13864
rect 30064 13812 30070 13864
rect 30193 13855 30251 13861
rect 30193 13821 30205 13855
rect 30239 13821 30251 13855
rect 31128 13852 31156 13960
rect 31205 13957 31217 13991
rect 31251 13957 31263 13991
rect 31205 13951 31263 13957
rect 31297 13991 31355 13997
rect 31297 13957 31309 13991
rect 31343 13988 31355 13991
rect 32030 13988 32036 14000
rect 31343 13960 32036 13988
rect 31343 13957 31355 13960
rect 31297 13951 31355 13957
rect 32030 13948 32036 13960
rect 32088 13948 32094 14000
rect 32140 13997 32168 14028
rect 32582 14016 32588 14068
rect 32640 14016 32646 14068
rect 34698 14056 34704 14068
rect 34532 14028 34704 14056
rect 32125 13991 32183 13997
rect 32125 13957 32137 13991
rect 32171 13957 32183 13991
rect 32125 13951 32183 13957
rect 33778 13948 33784 14000
rect 33836 13988 33842 14000
rect 34241 13991 34299 13997
rect 34241 13988 34253 13991
rect 33836 13960 34253 13988
rect 33836 13948 33842 13960
rect 34241 13957 34253 13960
rect 34287 13957 34299 13991
rect 34532 13988 34560 14028
rect 34698 14016 34704 14028
rect 34756 14016 34762 14068
rect 37182 14056 37188 14068
rect 34808 14028 37188 14056
rect 34241 13951 34299 13957
rect 34440 13960 34560 13988
rect 31389 13923 31447 13929
rect 31389 13889 31401 13923
rect 31435 13920 31447 13923
rect 31754 13920 31760 13932
rect 31435 13892 31760 13920
rect 31435 13889 31447 13892
rect 31389 13883 31447 13889
rect 31754 13880 31760 13892
rect 31812 13880 31818 13932
rect 32401 13923 32459 13929
rect 32401 13889 32413 13923
rect 32447 13920 32459 13923
rect 32674 13920 32680 13932
rect 32447 13892 32680 13920
rect 32447 13889 32459 13892
rect 32401 13883 32459 13889
rect 32674 13880 32680 13892
rect 32732 13880 32738 13932
rect 33134 13880 33140 13932
rect 33192 13880 33198 13932
rect 34440 13929 34468 13960
rect 34425 13923 34483 13929
rect 34425 13889 34437 13923
rect 34471 13889 34483 13923
rect 34425 13883 34483 13889
rect 34517 13923 34575 13929
rect 34517 13889 34529 13923
rect 34563 13889 34575 13923
rect 34517 13883 34575 13889
rect 32217 13855 32275 13861
rect 32217 13852 32229 13855
rect 31128 13824 32229 13852
rect 30193 13815 30251 13821
rect 32217 13821 32229 13824
rect 32263 13852 32275 13855
rect 32858 13852 32864 13864
rect 32263 13824 32864 13852
rect 32263 13821 32275 13824
rect 32217 13815 32275 13821
rect 28092 13756 28994 13784
rect 26844 13744 26850 13756
rect 28092 13716 28120 13756
rect 30098 13744 30104 13796
rect 30156 13744 30162 13796
rect 30208 13784 30236 13815
rect 32858 13812 32864 13824
rect 32916 13812 32922 13864
rect 33152 13852 33180 13880
rect 34532 13852 34560 13883
rect 34808 13852 34836 14028
rect 37182 14016 37188 14028
rect 37240 14016 37246 14068
rect 37476 14028 37688 14056
rect 37476 13988 37504 14028
rect 35176 13960 37504 13988
rect 35176 13932 35204 13960
rect 37550 13948 37556 14000
rect 37608 13948 37614 14000
rect 35158 13880 35164 13932
rect 35216 13880 35222 13932
rect 35805 13923 35863 13929
rect 35805 13920 35817 13923
rect 35728 13892 35817 13920
rect 35728 13864 35756 13892
rect 35805 13889 35817 13892
rect 35851 13889 35863 13923
rect 35805 13883 35863 13889
rect 35897 13923 35955 13929
rect 35897 13889 35909 13923
rect 35943 13889 35955 13923
rect 35897 13883 35955 13889
rect 33152 13824 34560 13852
rect 34716 13824 34836 13852
rect 32490 13784 32496 13796
rect 30208 13756 32496 13784
rect 32490 13744 32496 13756
rect 32548 13744 32554 13796
rect 33226 13744 33232 13796
rect 33284 13784 33290 13796
rect 34146 13784 34152 13796
rect 33284 13756 34152 13784
rect 33284 13744 33290 13756
rect 34146 13744 34152 13756
rect 34204 13744 34210 13796
rect 34422 13744 34428 13796
rect 34480 13784 34486 13796
rect 34716 13793 34744 13824
rect 35710 13812 35716 13864
rect 35768 13812 35774 13864
rect 35912 13852 35940 13883
rect 35986 13880 35992 13932
rect 36044 13880 36050 13932
rect 36078 13880 36084 13932
rect 36136 13929 36142 13932
rect 36136 13923 36165 13929
rect 36153 13889 36165 13923
rect 36136 13883 36165 13889
rect 36136 13880 36142 13883
rect 36262 13880 36268 13932
rect 36320 13880 36326 13932
rect 36906 13880 36912 13932
rect 36964 13880 36970 13932
rect 37274 13880 37280 13932
rect 37332 13880 37338 13932
rect 37660 13929 37688 14028
rect 37826 14016 37832 14068
rect 37884 14016 37890 14068
rect 37461 13923 37519 13929
rect 37461 13889 37473 13923
rect 37507 13889 37519 13923
rect 37461 13883 37519 13889
rect 37645 13923 37703 13929
rect 37645 13889 37657 13923
rect 37691 13920 37703 13923
rect 39482 13920 39488 13932
rect 37691 13892 39488 13920
rect 37691 13889 37703 13892
rect 37645 13883 37703 13889
rect 36924 13852 36952 13880
rect 35912 13824 36952 13852
rect 37476 13852 37504 13883
rect 39482 13880 39488 13892
rect 39540 13880 39546 13932
rect 38930 13852 38936 13864
rect 37476 13824 38936 13852
rect 38930 13812 38936 13824
rect 38988 13852 38994 13864
rect 39114 13852 39120 13864
rect 38988 13824 39120 13852
rect 38988 13812 38994 13824
rect 39114 13812 39120 13824
rect 39172 13812 39178 13864
rect 34701 13787 34759 13793
rect 34480 13756 34652 13784
rect 34480 13744 34486 13756
rect 26344 13688 28120 13716
rect 28166 13676 28172 13728
rect 28224 13716 28230 13728
rect 30116 13716 30144 13744
rect 28224 13688 30144 13716
rect 28224 13676 28230 13688
rect 32122 13676 32128 13728
rect 32180 13676 32186 13728
rect 34514 13676 34520 13728
rect 34572 13676 34578 13728
rect 34624 13716 34652 13756
rect 34701 13753 34713 13787
rect 34747 13753 34759 13787
rect 36446 13784 36452 13796
rect 34701 13747 34759 13753
rect 34808 13756 36452 13784
rect 34808 13716 34836 13756
rect 36446 13744 36452 13756
rect 36504 13744 36510 13796
rect 36722 13744 36728 13796
rect 36780 13784 36786 13796
rect 36998 13784 37004 13796
rect 36780 13756 37004 13784
rect 36780 13744 36786 13756
rect 36998 13744 37004 13756
rect 37056 13744 37062 13796
rect 34624 13688 34836 13716
rect 35618 13676 35624 13728
rect 35676 13676 35682 13728
rect 1104 13626 41400 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 41400 13626
rect 1104 13552 41400 13574
rect 1762 13472 1768 13524
rect 1820 13512 1826 13524
rect 2225 13515 2283 13521
rect 2225 13512 2237 13515
rect 1820 13484 2237 13512
rect 1820 13472 1826 13484
rect 2225 13481 2237 13484
rect 2271 13481 2283 13515
rect 2225 13475 2283 13481
rect 3694 13472 3700 13524
rect 3752 13512 3758 13524
rect 4709 13515 4767 13521
rect 4709 13512 4721 13515
rect 3752 13484 4721 13512
rect 3752 13472 3758 13484
rect 4709 13481 4721 13484
rect 4755 13481 4767 13515
rect 4709 13475 4767 13481
rect 5537 13515 5595 13521
rect 5537 13481 5549 13515
rect 5583 13512 5595 13515
rect 6546 13512 6552 13524
rect 5583 13484 6552 13512
rect 5583 13481 5595 13484
rect 5537 13475 5595 13481
rect 6546 13472 6552 13484
rect 6604 13472 6610 13524
rect 6822 13472 6828 13524
rect 6880 13512 6886 13524
rect 7377 13515 7435 13521
rect 7377 13512 7389 13515
rect 6880 13484 7389 13512
rect 6880 13472 6886 13484
rect 7377 13481 7389 13484
rect 7423 13481 7435 13515
rect 7377 13475 7435 13481
rect 8294 13472 8300 13524
rect 8352 13512 8358 13524
rect 10778 13512 10784 13524
rect 8352 13484 10784 13512
rect 8352 13472 8358 13484
rect 10778 13472 10784 13484
rect 10836 13472 10842 13524
rect 14642 13472 14648 13524
rect 14700 13512 14706 13524
rect 14829 13515 14887 13521
rect 14829 13512 14841 13515
rect 14700 13484 14841 13512
rect 14700 13472 14706 13484
rect 14829 13481 14841 13484
rect 14875 13481 14887 13515
rect 15657 13515 15715 13521
rect 15657 13512 15669 13515
rect 14829 13475 14887 13481
rect 14936 13484 15669 13512
rect 6086 13444 6092 13456
rect 4908 13416 6092 13444
rect 2409 13311 2467 13317
rect 2409 13277 2421 13311
rect 2455 13308 2467 13311
rect 2774 13308 2780 13320
rect 2455 13280 2780 13308
rect 2455 13277 2467 13280
rect 2409 13271 2467 13277
rect 2774 13268 2780 13280
rect 2832 13268 2838 13320
rect 4908 13317 4936 13416
rect 6086 13404 6092 13416
rect 6144 13444 6150 13456
rect 6730 13444 6736 13456
rect 6144 13416 6736 13444
rect 6144 13404 6150 13416
rect 6730 13404 6736 13416
rect 6788 13404 6794 13456
rect 7926 13444 7932 13456
rect 7576 13416 7932 13444
rect 5000 13348 6040 13376
rect 5000 13317 5028 13348
rect 6012 13320 6040 13348
rect 4893 13311 4951 13317
rect 4893 13277 4905 13311
rect 4939 13277 4951 13311
rect 4893 13271 4951 13277
rect 4985 13311 5043 13317
rect 4985 13277 4997 13311
rect 5031 13277 5043 13311
rect 4985 13271 5043 13277
rect 5169 13311 5227 13317
rect 5169 13277 5181 13311
rect 5215 13277 5227 13311
rect 5169 13271 5227 13277
rect 5184 13240 5212 13271
rect 5258 13268 5264 13320
rect 5316 13268 5322 13320
rect 5442 13268 5448 13320
rect 5500 13268 5506 13320
rect 5534 13268 5540 13320
rect 5592 13268 5598 13320
rect 5629 13311 5687 13317
rect 5629 13277 5641 13311
rect 5675 13277 5687 13311
rect 5629 13271 5687 13277
rect 5552 13240 5580 13268
rect 5184 13212 5580 13240
rect 5644 13240 5672 13271
rect 5994 13268 6000 13320
rect 6052 13268 6058 13320
rect 6454 13268 6460 13320
rect 6512 13308 6518 13320
rect 6549 13311 6607 13317
rect 6549 13308 6561 13311
rect 6512 13280 6561 13308
rect 6512 13268 6518 13280
rect 6549 13277 6561 13280
rect 6595 13277 6607 13311
rect 6549 13271 6607 13277
rect 6733 13311 6791 13317
rect 6733 13277 6745 13311
rect 6779 13308 6791 13311
rect 7006 13308 7012 13320
rect 6779 13280 7012 13308
rect 6779 13277 6791 13280
rect 6733 13271 6791 13277
rect 7006 13268 7012 13280
rect 7064 13268 7070 13320
rect 7101 13311 7159 13317
rect 7101 13277 7113 13311
rect 7147 13308 7159 13311
rect 7576 13308 7604 13416
rect 7926 13404 7932 13416
rect 7984 13404 7990 13456
rect 8110 13404 8116 13456
rect 8168 13444 8174 13456
rect 9677 13447 9735 13453
rect 9677 13444 9689 13447
rect 8168 13416 9689 13444
rect 8168 13404 8174 13416
rect 9677 13413 9689 13416
rect 9723 13413 9735 13447
rect 9677 13407 9735 13413
rect 10410 13404 10416 13456
rect 10468 13444 10474 13456
rect 11241 13447 11299 13453
rect 11241 13444 11253 13447
rect 10468 13416 11253 13444
rect 10468 13404 10474 13416
rect 11241 13413 11253 13416
rect 11287 13413 11299 13447
rect 12437 13447 12495 13453
rect 12437 13444 12449 13447
rect 11241 13407 11299 13413
rect 11348 13416 12449 13444
rect 8846 13376 8852 13388
rect 7944 13348 8852 13376
rect 7147 13280 7604 13308
rect 7147 13277 7159 13280
rect 7101 13271 7159 13277
rect 7650 13268 7656 13320
rect 7708 13268 7714 13320
rect 7944 13317 7972 13348
rect 8846 13336 8852 13348
rect 8904 13376 8910 13388
rect 9309 13379 9367 13385
rect 8904 13348 9168 13376
rect 8904 13336 8910 13348
rect 7929 13311 7987 13317
rect 7929 13277 7941 13311
rect 7975 13277 7987 13311
rect 7929 13271 7987 13277
rect 8110 13268 8116 13320
rect 8168 13306 8174 13320
rect 8205 13311 8263 13317
rect 8205 13306 8217 13311
rect 8168 13278 8217 13306
rect 8168 13268 8174 13278
rect 8205 13277 8217 13278
rect 8251 13277 8263 13311
rect 8205 13271 8263 13277
rect 8573 13311 8631 13317
rect 8573 13277 8585 13311
rect 8619 13308 8631 13311
rect 8662 13308 8668 13320
rect 8619 13280 8668 13308
rect 8619 13277 8631 13280
rect 8573 13271 8631 13277
rect 8662 13268 8668 13280
rect 8720 13268 8726 13320
rect 8938 13268 8944 13320
rect 8996 13268 9002 13320
rect 9140 13317 9168 13348
rect 9309 13345 9321 13379
rect 9355 13376 9367 13379
rect 9398 13376 9404 13388
rect 9355 13348 9404 13376
rect 9355 13345 9367 13348
rect 9309 13339 9367 13345
rect 9398 13336 9404 13348
rect 9456 13336 9462 13388
rect 10594 13336 10600 13388
rect 10652 13336 10658 13388
rect 11348 13376 11376 13416
rect 12437 13413 12449 13416
rect 12483 13444 12495 13447
rect 12805 13447 12863 13453
rect 12483 13416 12664 13444
rect 12483 13413 12495 13416
rect 12437 13407 12495 13413
rect 10980 13348 11376 13376
rect 11716 13348 12480 13376
rect 9125 13311 9183 13317
rect 9125 13277 9137 13311
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 9217 13311 9275 13317
rect 9217 13277 9229 13311
rect 9263 13284 9275 13311
rect 9504 13311 9562 13317
rect 9263 13277 9352 13284
rect 9217 13271 9352 13277
rect 9504 13277 9516 13311
rect 9550 13308 9562 13311
rect 9550 13280 9628 13308
rect 9550 13277 9562 13280
rect 9504 13271 9562 13277
rect 9232 13256 9352 13271
rect 7374 13240 7380 13252
rect 5644 13212 7380 13240
rect 7374 13200 7380 13212
rect 7432 13200 7438 13252
rect 7561 13243 7619 13249
rect 7561 13209 7573 13243
rect 7607 13240 7619 13243
rect 7607 13212 8156 13240
rect 7607 13209 7619 13212
rect 7561 13203 7619 13209
rect 6730 13132 6736 13184
rect 6788 13132 6794 13184
rect 7190 13132 7196 13184
rect 7248 13132 7254 13184
rect 8018 13132 8024 13184
rect 8076 13132 8082 13184
rect 8128 13172 8156 13212
rect 8386 13200 8392 13252
rect 8444 13200 8450 13252
rect 8478 13200 8484 13252
rect 8536 13240 8542 13252
rect 9324 13240 9352 13256
rect 9398 13240 9404 13252
rect 8536 13212 9076 13240
rect 9324 13212 9404 13240
rect 8536 13200 8542 13212
rect 9048 13184 9076 13212
rect 9398 13200 9404 13212
rect 9456 13200 9462 13252
rect 9600 13240 9628 13280
rect 9858 13268 9864 13320
rect 9916 13308 9922 13320
rect 10413 13311 10471 13317
rect 10413 13308 10425 13311
rect 9916 13280 10425 13308
rect 9916 13268 9922 13280
rect 10413 13277 10425 13280
rect 10459 13308 10471 13311
rect 10980 13308 11008 13348
rect 10459 13280 11008 13308
rect 10459 13277 10471 13280
rect 10413 13271 10471 13277
rect 11054 13268 11060 13320
rect 11112 13268 11118 13320
rect 11146 13268 11152 13320
rect 11204 13308 11210 13320
rect 11333 13311 11391 13317
rect 11333 13308 11345 13311
rect 11204 13280 11345 13308
rect 11204 13268 11210 13280
rect 11333 13277 11345 13280
rect 11379 13308 11391 13311
rect 11716 13308 11744 13348
rect 11379 13280 11744 13308
rect 11793 13311 11851 13317
rect 11379 13277 11391 13280
rect 11333 13271 11391 13277
rect 11793 13277 11805 13311
rect 11839 13308 11851 13311
rect 11882 13308 11888 13320
rect 11839 13280 11888 13308
rect 11839 13277 11851 13280
rect 11793 13271 11851 13277
rect 11808 13240 11836 13271
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 11974 13268 11980 13320
rect 12032 13268 12038 13320
rect 12158 13268 12164 13320
rect 12216 13308 12222 13320
rect 12253 13311 12311 13317
rect 12253 13308 12265 13311
rect 12216 13280 12265 13308
rect 12216 13268 12222 13280
rect 12253 13277 12265 13280
rect 12299 13277 12311 13311
rect 12253 13271 12311 13277
rect 12345 13311 12403 13317
rect 12345 13277 12357 13311
rect 12391 13277 12403 13311
rect 12345 13271 12403 13277
rect 9600 13212 11836 13240
rect 8757 13175 8815 13181
rect 8757 13172 8769 13175
rect 8128 13144 8769 13172
rect 8757 13141 8769 13144
rect 8803 13141 8815 13175
rect 8757 13135 8815 13141
rect 9030 13132 9036 13184
rect 9088 13132 9094 13184
rect 9490 13132 9496 13184
rect 9548 13172 9554 13184
rect 9600 13172 9628 13212
rect 9548 13144 9628 13172
rect 9548 13132 9554 13144
rect 9674 13132 9680 13184
rect 9732 13172 9738 13184
rect 10045 13175 10103 13181
rect 10045 13172 10057 13175
rect 9732 13144 10057 13172
rect 9732 13132 9738 13144
rect 10045 13141 10057 13144
rect 10091 13141 10103 13175
rect 10045 13135 10103 13141
rect 10502 13132 10508 13184
rect 10560 13132 10566 13184
rect 10594 13132 10600 13184
rect 10652 13172 10658 13184
rect 10873 13175 10931 13181
rect 10873 13172 10885 13175
rect 10652 13144 10885 13172
rect 10652 13132 10658 13144
rect 10873 13141 10885 13144
rect 10919 13141 10931 13175
rect 10873 13135 10931 13141
rect 11885 13175 11943 13181
rect 11885 13141 11897 13175
rect 11931 13172 11943 13175
rect 11974 13172 11980 13184
rect 11931 13144 11980 13172
rect 11931 13141 11943 13144
rect 11885 13135 11943 13141
rect 11974 13132 11980 13144
rect 12032 13132 12038 13184
rect 12069 13175 12127 13181
rect 12069 13141 12081 13175
rect 12115 13172 12127 13175
rect 12158 13172 12164 13184
rect 12115 13144 12164 13172
rect 12115 13141 12127 13144
rect 12069 13135 12127 13141
rect 12158 13132 12164 13144
rect 12216 13132 12222 13184
rect 12360 13172 12388 13271
rect 12452 13240 12480 13348
rect 12526 13268 12532 13320
rect 12584 13268 12590 13320
rect 12636 13318 12664 13416
rect 12805 13413 12817 13447
rect 12851 13444 12863 13447
rect 12986 13444 12992 13456
rect 12851 13416 12992 13444
rect 12851 13413 12863 13416
rect 12805 13407 12863 13413
rect 12986 13404 12992 13416
rect 13044 13404 13050 13456
rect 14936 13444 14964 13484
rect 15657 13481 15669 13484
rect 15703 13512 15715 13515
rect 16022 13512 16028 13524
rect 15703 13484 16028 13512
rect 15703 13481 15715 13484
rect 15657 13475 15715 13481
rect 16022 13472 16028 13484
rect 16080 13472 16086 13524
rect 16390 13472 16396 13524
rect 16448 13472 16454 13524
rect 17218 13512 17224 13524
rect 16500 13484 17224 13512
rect 14108 13416 14964 13444
rect 13078 13336 13084 13388
rect 13136 13336 13142 13388
rect 12705 13321 12763 13327
rect 12705 13318 12717 13321
rect 12636 13290 12717 13318
rect 12705 13287 12717 13290
rect 12751 13287 12763 13321
rect 12705 13281 12763 13287
rect 12989 13311 13047 13317
rect 12989 13277 13001 13311
rect 13035 13277 13047 13311
rect 12989 13271 13047 13277
rect 12802 13240 12808 13252
rect 12452 13212 12808 13240
rect 12802 13200 12808 13212
rect 12860 13240 12866 13252
rect 13004 13240 13032 13271
rect 13170 13268 13176 13320
rect 13228 13268 13234 13320
rect 14108 13252 14136 13416
rect 15286 13404 15292 13456
rect 15344 13404 15350 13456
rect 15304 13376 15332 13404
rect 16500 13376 16528 13484
rect 17218 13472 17224 13484
rect 17276 13472 17282 13524
rect 23014 13512 23020 13524
rect 20916 13484 21956 13512
rect 16577 13447 16635 13453
rect 16577 13413 16589 13447
rect 16623 13444 16635 13447
rect 20806 13444 20812 13456
rect 16623 13416 16712 13444
rect 16623 13413 16635 13416
rect 16577 13407 16635 13413
rect 16684 13388 16712 13416
rect 16868 13416 20812 13444
rect 14752 13348 15332 13376
rect 15396 13348 16528 13376
rect 14752 13317 14780 13348
rect 14737 13311 14795 13317
rect 14737 13277 14749 13311
rect 14783 13277 14795 13311
rect 15289 13311 15347 13317
rect 15289 13308 15301 13311
rect 14737 13271 14795 13277
rect 14844 13280 15301 13308
rect 12860 13212 13032 13240
rect 12860 13200 12866 13212
rect 13630 13200 13636 13252
rect 13688 13240 13694 13252
rect 13998 13240 14004 13252
rect 13688 13212 14004 13240
rect 13688 13200 13694 13212
rect 13998 13200 14004 13212
rect 14056 13200 14062 13252
rect 14090 13200 14096 13252
rect 14148 13200 14154 13252
rect 14182 13200 14188 13252
rect 14240 13240 14246 13252
rect 14844 13240 14872 13280
rect 15289 13277 15301 13280
rect 15335 13308 15347 13311
rect 15396 13308 15424 13348
rect 16666 13336 16672 13388
rect 16724 13336 16730 13388
rect 15335 13280 15424 13308
rect 15473 13311 15531 13317
rect 15335 13277 15347 13280
rect 15289 13271 15347 13277
rect 15473 13277 15485 13311
rect 15519 13277 15531 13311
rect 15473 13271 15531 13277
rect 15488 13240 15516 13271
rect 15654 13268 15660 13320
rect 15712 13268 15718 13320
rect 15841 13311 15899 13317
rect 15841 13277 15853 13311
rect 15887 13308 15899 13311
rect 16117 13311 16175 13317
rect 16117 13308 16129 13311
rect 15887 13280 16129 13308
rect 15887 13277 15899 13280
rect 15841 13271 15899 13277
rect 16117 13277 16129 13280
rect 16163 13277 16175 13311
rect 16117 13271 16175 13277
rect 16209 13311 16267 13317
rect 16209 13277 16221 13311
rect 16255 13308 16267 13311
rect 16761 13311 16819 13317
rect 16761 13308 16773 13311
rect 16255 13280 16773 13308
rect 16255 13277 16267 13280
rect 16209 13271 16267 13277
rect 16761 13277 16773 13280
rect 16807 13308 16819 13311
rect 16868 13308 16896 13416
rect 20806 13404 20812 13416
rect 20864 13404 20870 13456
rect 17402 13336 17408 13388
rect 17460 13376 17466 13388
rect 17957 13379 18015 13385
rect 17957 13376 17969 13379
rect 17460 13348 17969 13376
rect 17460 13336 17466 13348
rect 17957 13345 17969 13348
rect 18003 13345 18015 13379
rect 17957 13339 18015 13345
rect 18049 13379 18107 13385
rect 18049 13345 18061 13379
rect 18095 13376 18107 13379
rect 19978 13376 19984 13388
rect 18095 13348 19984 13376
rect 18095 13345 18107 13348
rect 18049 13339 18107 13345
rect 19978 13336 19984 13348
rect 20036 13336 20042 13388
rect 16807 13280 16896 13308
rect 17221 13311 17279 13317
rect 16807 13277 16819 13280
rect 16761 13271 16819 13277
rect 17221 13277 17233 13311
rect 17267 13277 17279 13311
rect 17221 13271 17279 13277
rect 17497 13311 17555 13317
rect 17497 13277 17509 13311
rect 17543 13308 17555 13311
rect 17586 13308 17592 13320
rect 17543 13280 17592 13308
rect 17543 13277 17555 13280
rect 17497 13271 17555 13277
rect 14240 13212 14872 13240
rect 15212 13212 15516 13240
rect 14240 13200 14246 13212
rect 12618 13172 12624 13184
rect 12360 13144 12624 13172
rect 12618 13132 12624 13144
rect 12676 13132 12682 13184
rect 14274 13132 14280 13184
rect 14332 13172 14338 13184
rect 15212 13181 15240 13212
rect 15197 13175 15255 13181
rect 15197 13172 15209 13175
rect 14332 13144 15209 13172
rect 14332 13132 14338 13144
rect 15197 13141 15209 13144
rect 15243 13141 15255 13175
rect 15197 13135 15255 13141
rect 15378 13132 15384 13184
rect 15436 13132 15442 13184
rect 15672 13172 15700 13268
rect 16132 13240 16160 13271
rect 17236 13240 17264 13271
rect 17586 13268 17592 13280
rect 17644 13268 17650 13320
rect 17678 13268 17684 13320
rect 17736 13268 17742 13320
rect 18138 13268 18144 13320
rect 18196 13308 18202 13320
rect 19702 13308 19708 13320
rect 18196 13280 19708 13308
rect 18196 13268 18202 13280
rect 19702 13268 19708 13280
rect 19760 13268 19766 13320
rect 17696 13240 17724 13268
rect 16132 13212 17724 13240
rect 20806 13200 20812 13252
rect 20864 13200 20870 13252
rect 15838 13172 15844 13184
rect 15672 13144 15844 13172
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 17678 13132 17684 13184
rect 17736 13132 17742 13184
rect 20916 13172 20944 13484
rect 21928 13444 21956 13484
rect 22296 13484 23020 13512
rect 22186 13444 22192 13456
rect 21008 13416 21864 13444
rect 21928 13416 22192 13444
rect 21008 13317 21036 13416
rect 21836 13376 21864 13416
rect 22186 13404 22192 13416
rect 22244 13404 22250 13456
rect 22296 13376 22324 13484
rect 23014 13472 23020 13484
rect 23072 13472 23078 13524
rect 26970 13472 26976 13524
rect 27028 13472 27034 13524
rect 27706 13472 27712 13524
rect 27764 13512 27770 13524
rect 28166 13512 28172 13524
rect 27764 13484 28172 13512
rect 27764 13472 27770 13484
rect 28166 13472 28172 13484
rect 28224 13472 28230 13524
rect 29362 13472 29368 13524
rect 29420 13512 29426 13524
rect 29733 13515 29791 13521
rect 29733 13512 29745 13515
rect 29420 13484 29745 13512
rect 29420 13472 29426 13484
rect 29733 13481 29745 13484
rect 29779 13481 29791 13515
rect 29733 13475 29791 13481
rect 32858 13472 32864 13524
rect 32916 13512 32922 13524
rect 34606 13512 34612 13524
rect 32916 13484 34612 13512
rect 32916 13472 32922 13484
rect 34606 13472 34612 13484
rect 34664 13472 34670 13524
rect 35802 13472 35808 13524
rect 35860 13472 35866 13524
rect 37829 13515 37887 13521
rect 37829 13481 37841 13515
rect 37875 13512 37887 13515
rect 37918 13512 37924 13524
rect 37875 13484 37924 13512
rect 37875 13481 37887 13484
rect 37829 13475 37887 13481
rect 37918 13472 37924 13484
rect 37976 13472 37982 13524
rect 39850 13472 39856 13524
rect 39908 13472 39914 13524
rect 40034 13472 40040 13524
rect 40092 13512 40098 13524
rect 40221 13515 40279 13521
rect 40221 13512 40233 13515
rect 40092 13484 40233 13512
rect 40092 13472 40098 13484
rect 40221 13481 40233 13484
rect 40267 13481 40279 13515
rect 40221 13475 40279 13481
rect 26786 13404 26792 13456
rect 26844 13444 26850 13456
rect 26881 13447 26939 13453
rect 26881 13444 26893 13447
rect 26844 13416 26893 13444
rect 26844 13404 26850 13416
rect 26881 13413 26893 13416
rect 26927 13413 26939 13447
rect 26881 13407 26939 13413
rect 21192 13348 21680 13376
rect 21836 13348 22324 13376
rect 26988 13376 27016 13472
rect 31478 13404 31484 13456
rect 31536 13444 31542 13456
rect 33226 13444 33232 13456
rect 31536 13416 33232 13444
rect 31536 13404 31542 13416
rect 33226 13404 33232 13416
rect 33284 13404 33290 13456
rect 35268 13416 36308 13444
rect 35268 13388 35296 13416
rect 27065 13379 27123 13385
rect 27065 13376 27077 13379
rect 26988 13348 27077 13376
rect 20993 13311 21051 13317
rect 20993 13277 21005 13311
rect 21039 13277 21051 13311
rect 20993 13271 21051 13277
rect 21192 13184 21220 13348
rect 21266 13268 21272 13320
rect 21324 13308 21330 13320
rect 21453 13311 21511 13317
rect 21453 13308 21465 13311
rect 21324 13280 21465 13308
rect 21324 13268 21330 13280
rect 21453 13277 21465 13280
rect 21499 13277 21511 13311
rect 21652 13308 21680 13348
rect 27065 13345 27077 13348
rect 27111 13376 27123 13379
rect 27249 13379 27307 13385
rect 27249 13376 27261 13379
rect 27111 13348 27261 13376
rect 27111 13345 27123 13348
rect 27065 13339 27123 13345
rect 27249 13345 27261 13348
rect 27295 13345 27307 13379
rect 27249 13339 27307 13345
rect 30469 13379 30527 13385
rect 30469 13345 30481 13379
rect 30515 13376 30527 13379
rect 32674 13376 32680 13388
rect 30515 13348 32680 13376
rect 30515 13345 30527 13348
rect 30469 13339 30527 13345
rect 32674 13336 32680 13348
rect 32732 13336 32738 13388
rect 33870 13336 33876 13388
rect 33928 13376 33934 13388
rect 33928 13348 34376 13376
rect 33928 13336 33934 13348
rect 21713 13311 21771 13317
rect 21713 13308 21725 13311
rect 21652 13280 21725 13308
rect 21453 13271 21511 13277
rect 21713 13277 21725 13280
rect 21759 13277 21771 13311
rect 21713 13271 21771 13277
rect 21821 13311 21879 13317
rect 21821 13277 21833 13311
rect 21867 13308 21879 13311
rect 22649 13311 22707 13317
rect 21867 13280 22324 13308
rect 21867 13277 21879 13280
rect 21821 13271 21879 13277
rect 21361 13243 21419 13249
rect 21361 13209 21373 13243
rect 21407 13240 21419 13243
rect 22186 13240 22192 13252
rect 21407 13212 22192 13240
rect 21407 13209 21419 13212
rect 21361 13203 21419 13209
rect 22186 13200 22192 13212
rect 22244 13200 22250 13252
rect 21085 13175 21143 13181
rect 21085 13172 21097 13175
rect 20916 13144 21097 13172
rect 21085 13141 21097 13144
rect 21131 13141 21143 13175
rect 21085 13135 21143 13141
rect 21174 13132 21180 13184
rect 21232 13132 21238 13184
rect 22296 13172 22324 13280
rect 22649 13277 22661 13311
rect 22695 13308 22707 13311
rect 22738 13308 22744 13320
rect 22695 13280 22744 13308
rect 22695 13277 22707 13280
rect 22649 13271 22707 13277
rect 22738 13268 22744 13280
rect 22796 13268 22802 13320
rect 22925 13311 22983 13317
rect 22925 13277 22937 13311
rect 22971 13277 22983 13311
rect 22925 13271 22983 13277
rect 22370 13200 22376 13252
rect 22428 13240 22434 13252
rect 22940 13240 22968 13271
rect 26234 13268 26240 13320
rect 26292 13308 26298 13320
rect 26789 13311 26847 13317
rect 26789 13308 26801 13311
rect 26292 13280 26801 13308
rect 26292 13268 26298 13280
rect 26789 13277 26801 13280
rect 26835 13277 26847 13311
rect 26789 13271 26847 13277
rect 27157 13311 27215 13317
rect 27157 13277 27169 13311
rect 27203 13308 27215 13311
rect 27341 13311 27399 13317
rect 27203 13280 27292 13308
rect 27203 13277 27215 13280
rect 27157 13271 27215 13277
rect 27264 13252 27292 13280
rect 27341 13277 27353 13311
rect 27387 13308 27399 13311
rect 27430 13308 27436 13320
rect 27387 13280 27436 13308
rect 27387 13277 27399 13280
rect 27341 13271 27399 13277
rect 27430 13268 27436 13280
rect 27488 13308 27494 13320
rect 27890 13308 27896 13320
rect 27488 13280 27896 13308
rect 27488 13268 27494 13280
rect 27890 13268 27896 13280
rect 27948 13308 27954 13320
rect 29641 13311 29699 13317
rect 29641 13308 29653 13311
rect 27948 13280 29653 13308
rect 27948 13268 27954 13280
rect 29641 13277 29653 13280
rect 29687 13277 29699 13311
rect 29641 13271 29699 13277
rect 29730 13268 29736 13320
rect 29788 13308 29794 13320
rect 30377 13311 30435 13317
rect 30377 13308 30389 13311
rect 29788 13280 30389 13308
rect 29788 13268 29794 13280
rect 30377 13277 30389 13280
rect 30423 13277 30435 13311
rect 30377 13271 30435 13277
rect 33962 13268 33968 13320
rect 34020 13268 34026 13320
rect 34054 13268 34060 13320
rect 34112 13308 34118 13320
rect 34348 13317 34376 13348
rect 35250 13336 35256 13388
rect 35308 13336 35314 13388
rect 36280 13385 36308 13416
rect 36354 13404 36360 13456
rect 36412 13444 36418 13456
rect 36412 13416 39988 13444
rect 36412 13404 36418 13416
rect 36173 13379 36231 13385
rect 36173 13376 36185 13379
rect 35729 13348 36185 13376
rect 34241 13311 34299 13317
rect 34241 13308 34253 13311
rect 34112 13280 34253 13308
rect 34112 13268 34118 13280
rect 34241 13277 34253 13280
rect 34287 13277 34299 13311
rect 34241 13271 34299 13277
rect 34333 13311 34391 13317
rect 34333 13277 34345 13311
rect 34379 13308 34391 13311
rect 35434 13308 35440 13320
rect 34379 13280 35440 13308
rect 34379 13277 34391 13280
rect 34333 13271 34391 13277
rect 35434 13268 35440 13280
rect 35492 13268 35498 13320
rect 22428 13212 22968 13240
rect 22428 13200 22434 13212
rect 27062 13200 27068 13252
rect 27120 13200 27126 13252
rect 27246 13200 27252 13252
rect 27304 13240 27310 13252
rect 27522 13240 27528 13252
rect 27304 13212 27528 13240
rect 27304 13200 27310 13212
rect 27522 13200 27528 13212
rect 27580 13200 27586 13252
rect 32306 13200 32312 13252
rect 32364 13200 32370 13252
rect 33318 13200 33324 13252
rect 33376 13240 33382 13252
rect 34149 13243 34207 13249
rect 34149 13240 34161 13243
rect 33376 13212 34161 13240
rect 33376 13200 33382 13212
rect 34149 13209 34161 13212
rect 34195 13209 34207 13243
rect 34149 13203 34207 13209
rect 34882 13200 34888 13252
rect 34940 13240 34946 13252
rect 35729 13240 35757 13348
rect 36173 13345 36185 13348
rect 36219 13345 36231 13379
rect 36173 13339 36231 13345
rect 36265 13379 36323 13385
rect 36265 13345 36277 13379
rect 36311 13376 36323 13379
rect 38838 13376 38844 13388
rect 36311 13348 36768 13376
rect 36311 13345 36323 13348
rect 36265 13339 36323 13345
rect 35802 13268 35808 13320
rect 35860 13308 35866 13320
rect 35989 13311 36047 13317
rect 35989 13308 36001 13311
rect 35860 13280 36001 13308
rect 35860 13268 35866 13280
rect 35989 13277 36001 13280
rect 36035 13277 36047 13311
rect 35989 13271 36047 13277
rect 36081 13311 36139 13317
rect 36081 13277 36093 13311
rect 36127 13308 36139 13311
rect 36280 13308 36400 13310
rect 36446 13308 36452 13320
rect 36127 13282 36452 13308
rect 36127 13280 36308 13282
rect 36372 13280 36452 13282
rect 36127 13277 36139 13280
rect 36081 13271 36139 13277
rect 36446 13268 36452 13280
rect 36504 13268 36510 13320
rect 36541 13243 36599 13249
rect 36541 13240 36553 13243
rect 34940 13212 36553 13240
rect 34940 13200 34946 13212
rect 36004 13184 36032 13212
rect 36541 13209 36553 13212
rect 36587 13209 36599 13243
rect 36541 13203 36599 13209
rect 22741 13175 22799 13181
rect 22741 13172 22753 13175
rect 22296 13144 22753 13172
rect 22741 13141 22753 13144
rect 22787 13141 22799 13175
rect 22741 13135 22799 13141
rect 22830 13132 22836 13184
rect 22888 13172 22894 13184
rect 28074 13172 28080 13184
rect 22888 13144 28080 13172
rect 22888 13132 22894 13144
rect 28074 13132 28080 13144
rect 28132 13132 28138 13184
rect 31846 13132 31852 13184
rect 31904 13172 31910 13184
rect 32214 13172 32220 13184
rect 31904 13144 32220 13172
rect 31904 13132 31910 13144
rect 32214 13132 32220 13144
rect 32272 13172 32278 13184
rect 32401 13175 32459 13181
rect 32401 13172 32413 13175
rect 32272 13144 32413 13172
rect 32272 13132 32278 13144
rect 32401 13141 32413 13144
rect 32447 13172 32459 13175
rect 33778 13172 33784 13184
rect 32447 13144 33784 13172
rect 32447 13141 32459 13144
rect 32401 13135 32459 13141
rect 33778 13132 33784 13144
rect 33836 13132 33842 13184
rect 34514 13132 34520 13184
rect 34572 13132 34578 13184
rect 35986 13132 35992 13184
rect 36044 13132 36050 13184
rect 36630 13132 36636 13184
rect 36688 13132 36694 13184
rect 36740 13172 36768 13348
rect 37292 13348 38844 13376
rect 37292 13320 37320 13348
rect 38838 13336 38844 13348
rect 38896 13336 38902 13388
rect 39482 13376 39488 13388
rect 39132 13348 39488 13376
rect 37274 13268 37280 13320
rect 37332 13268 37338 13320
rect 37553 13311 37611 13317
rect 37553 13277 37565 13311
rect 37599 13277 37611 13311
rect 37553 13271 37611 13277
rect 37182 13200 37188 13252
rect 37240 13240 37246 13252
rect 37461 13243 37519 13249
rect 37461 13240 37473 13243
rect 37240 13212 37473 13240
rect 37240 13200 37246 13212
rect 37461 13209 37473 13212
rect 37507 13209 37519 13243
rect 37568 13240 37596 13271
rect 37642 13268 37648 13320
rect 37700 13268 37706 13320
rect 37826 13268 37832 13320
rect 37884 13268 37890 13320
rect 38102 13268 38108 13320
rect 38160 13308 38166 13320
rect 38749 13311 38807 13317
rect 38749 13308 38761 13311
rect 38160 13280 38761 13308
rect 38160 13268 38166 13280
rect 38749 13277 38761 13280
rect 38795 13277 38807 13311
rect 38749 13271 38807 13277
rect 39022 13268 39028 13320
rect 39080 13268 39086 13320
rect 39132 13317 39160 13348
rect 39482 13336 39488 13348
rect 39540 13336 39546 13388
rect 39960 13385 39988 13416
rect 39945 13379 40003 13385
rect 39945 13345 39957 13379
rect 39991 13345 40003 13379
rect 39945 13339 40003 13345
rect 39117 13311 39175 13317
rect 39117 13277 39129 13311
rect 39163 13277 39175 13311
rect 39853 13311 39911 13317
rect 39853 13308 39865 13311
rect 39117 13271 39175 13277
rect 39316 13280 39865 13308
rect 37844 13240 37872 13268
rect 37568 13212 37872 13240
rect 37461 13203 37519 13209
rect 38654 13200 38660 13252
rect 38712 13200 38718 13252
rect 38838 13200 38844 13252
rect 38896 13240 38902 13252
rect 38933 13243 38991 13249
rect 38933 13240 38945 13243
rect 38896 13212 38945 13240
rect 38896 13200 38902 13212
rect 38933 13209 38945 13212
rect 38979 13209 38991 13243
rect 38933 13203 38991 13209
rect 38672 13172 38700 13200
rect 39316 13181 39344 13280
rect 39853 13277 39865 13280
rect 39899 13277 39911 13311
rect 39853 13271 39911 13277
rect 36740 13144 38700 13172
rect 39301 13175 39359 13181
rect 39301 13141 39313 13175
rect 39347 13141 39359 13175
rect 39301 13135 39359 13141
rect 1104 13082 41400 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 41400 13082
rect 1104 13008 41400 13030
rect 6549 12971 6607 12977
rect 6549 12937 6561 12971
rect 6595 12968 6607 12971
rect 7006 12968 7012 12980
rect 6595 12940 7012 12968
rect 6595 12937 6607 12940
rect 6549 12931 6607 12937
rect 7006 12928 7012 12940
rect 7064 12928 7070 12980
rect 7190 12928 7196 12980
rect 7248 12968 7254 12980
rect 7745 12971 7803 12977
rect 7745 12968 7757 12971
rect 7248 12940 7757 12968
rect 7248 12928 7254 12940
rect 7745 12937 7757 12940
rect 7791 12937 7803 12971
rect 7745 12931 7803 12937
rect 8386 12928 8392 12980
rect 8444 12968 8450 12980
rect 8757 12971 8815 12977
rect 8757 12968 8769 12971
rect 8444 12940 8769 12968
rect 8444 12928 8450 12940
rect 8757 12937 8769 12940
rect 8803 12937 8815 12971
rect 9122 12968 9128 12980
rect 8757 12931 8815 12937
rect 8864 12940 9128 12968
rect 6454 12860 6460 12912
rect 6512 12900 6518 12912
rect 8864 12900 8892 12940
rect 9122 12928 9128 12940
rect 9180 12928 9186 12980
rect 9858 12928 9864 12980
rect 9916 12968 9922 12980
rect 10229 12971 10287 12977
rect 10229 12968 10241 12971
rect 9916 12940 10241 12968
rect 9916 12928 9922 12940
rect 10229 12937 10241 12940
rect 10275 12937 10287 12971
rect 10229 12931 10287 12937
rect 10410 12928 10416 12980
rect 10468 12928 10474 12980
rect 10502 12928 10508 12980
rect 10560 12968 10566 12980
rect 10597 12971 10655 12977
rect 10597 12968 10609 12971
rect 10560 12940 10609 12968
rect 10560 12928 10566 12940
rect 10597 12937 10609 12940
rect 10643 12937 10655 12971
rect 10597 12931 10655 12937
rect 11057 12971 11115 12977
rect 11057 12937 11069 12971
rect 11103 12968 11115 12971
rect 12345 12971 12403 12977
rect 12345 12968 12357 12971
rect 11103 12940 12357 12968
rect 11103 12937 11115 12940
rect 11057 12931 11115 12937
rect 12345 12937 12357 12940
rect 12391 12937 12403 12971
rect 12345 12931 12403 12937
rect 12618 12928 12624 12980
rect 12676 12968 12682 12980
rect 13998 12968 14004 12980
rect 12676 12940 14004 12968
rect 12676 12928 12682 12940
rect 13998 12928 14004 12940
rect 14056 12968 14062 12980
rect 16945 12971 17003 12977
rect 16945 12968 16957 12971
rect 14056 12940 16957 12968
rect 14056 12928 14062 12940
rect 16945 12937 16957 12940
rect 16991 12937 17003 12971
rect 16945 12931 17003 12937
rect 17494 12928 17500 12980
rect 17552 12968 17558 12980
rect 17773 12971 17831 12977
rect 17773 12968 17785 12971
rect 17552 12940 17785 12968
rect 17552 12928 17558 12940
rect 17773 12937 17785 12940
rect 17819 12937 17831 12971
rect 17773 12931 17831 12937
rect 22278 12928 22284 12980
rect 22336 12928 22342 12980
rect 24302 12928 24308 12980
rect 24360 12928 24366 12980
rect 26421 12971 26479 12977
rect 24688 12940 26372 12968
rect 6512 12872 6684 12900
rect 6512 12860 6518 12872
rect 6362 12792 6368 12844
rect 6420 12792 6426 12844
rect 6656 12841 6684 12872
rect 6748 12872 7880 12900
rect 6748 12844 6776 12872
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12801 6699 12835
rect 6641 12795 6699 12801
rect 6730 12792 6736 12844
rect 6788 12792 6794 12844
rect 6917 12835 6975 12841
rect 6917 12801 6929 12835
rect 6963 12832 6975 12835
rect 7190 12832 7196 12844
rect 6963 12804 7196 12832
rect 6963 12801 6975 12804
rect 6917 12795 6975 12801
rect 7190 12792 7196 12804
rect 7248 12792 7254 12844
rect 7285 12835 7343 12841
rect 7285 12801 7297 12835
rect 7331 12832 7343 12835
rect 7561 12835 7619 12841
rect 7561 12832 7573 12835
rect 7331 12804 7573 12832
rect 7331 12801 7343 12804
rect 7285 12795 7343 12801
rect 7561 12801 7573 12804
rect 7607 12832 7619 12835
rect 7742 12832 7748 12844
rect 7607 12804 7748 12832
rect 7607 12801 7619 12804
rect 7561 12795 7619 12801
rect 7742 12792 7748 12804
rect 7800 12792 7806 12844
rect 7852 12841 7880 12872
rect 8772 12872 8892 12900
rect 7837 12835 7895 12841
rect 7837 12801 7849 12835
rect 7883 12801 7895 12835
rect 7837 12795 7895 12801
rect 8294 12792 8300 12844
rect 8352 12832 8358 12844
rect 8389 12835 8447 12841
rect 8389 12832 8401 12835
rect 8352 12804 8401 12832
rect 8352 12792 8358 12804
rect 8389 12801 8401 12804
rect 8435 12801 8447 12835
rect 8389 12795 8447 12801
rect 8570 12792 8576 12844
rect 8628 12841 8634 12844
rect 8628 12832 8639 12841
rect 8628 12804 8708 12832
rect 8628 12795 8639 12804
rect 8628 12792 8634 12795
rect 7098 12724 7104 12776
rect 7156 12764 7162 12776
rect 8680 12764 8708 12804
rect 8772 12830 8800 12872
rect 9214 12860 9220 12912
rect 9272 12900 9278 12912
rect 9272 12872 10088 12900
rect 9272 12860 9278 12872
rect 10060 12844 10088 12872
rect 10778 12860 10784 12912
rect 10836 12900 10842 12912
rect 10836 12872 14228 12900
rect 10836 12860 10842 12872
rect 8849 12835 8907 12841
rect 8849 12830 8861 12835
rect 8772 12802 8861 12830
rect 8849 12801 8861 12802
rect 8895 12801 8907 12835
rect 8849 12795 8907 12801
rect 9030 12792 9036 12844
rect 9088 12792 9094 12844
rect 9674 12792 9680 12844
rect 9732 12832 9738 12844
rect 9861 12835 9919 12841
rect 9861 12832 9873 12835
rect 9732 12804 9873 12832
rect 9732 12792 9738 12804
rect 9861 12801 9873 12804
rect 9907 12801 9919 12835
rect 9861 12795 9919 12801
rect 10042 12792 10048 12844
rect 10100 12792 10106 12844
rect 10226 12792 10232 12844
rect 10284 12832 10290 12844
rect 10321 12835 10379 12841
rect 10321 12832 10333 12835
rect 10284 12804 10333 12832
rect 10284 12792 10290 12804
rect 10321 12801 10333 12804
rect 10367 12832 10379 12835
rect 10965 12835 11023 12841
rect 10965 12832 10977 12835
rect 10367 12804 10977 12832
rect 10367 12801 10379 12804
rect 10321 12795 10379 12801
rect 10965 12801 10977 12804
rect 11011 12801 11023 12835
rect 10965 12795 11023 12801
rect 8941 12767 8999 12773
rect 8941 12764 8953 12767
rect 7156 12736 7328 12764
rect 8680 12736 8953 12764
rect 7156 12724 7162 12736
rect 4614 12656 4620 12708
rect 4672 12696 4678 12708
rect 7193 12699 7251 12705
rect 7193 12696 7205 12699
rect 4672 12668 7205 12696
rect 4672 12656 4678 12668
rect 7193 12665 7205 12668
rect 7239 12665 7251 12699
rect 7193 12659 7251 12665
rect 6365 12631 6423 12637
rect 6365 12597 6377 12631
rect 6411 12628 6423 12631
rect 6730 12628 6736 12640
rect 6411 12600 6736 12628
rect 6411 12597 6423 12600
rect 6365 12591 6423 12597
rect 6730 12588 6736 12600
rect 6788 12588 6794 12640
rect 7300 12628 7328 12736
rect 8941 12733 8953 12736
rect 8987 12733 8999 12767
rect 8941 12727 8999 12733
rect 9048 12736 10456 12764
rect 7374 12656 7380 12708
rect 7432 12696 7438 12708
rect 9048 12696 9076 12736
rect 7432 12668 9076 12696
rect 7432 12656 7438 12668
rect 9858 12628 9864 12640
rect 7300 12600 9864 12628
rect 9858 12588 9864 12600
rect 9916 12588 9922 12640
rect 10045 12631 10103 12637
rect 10045 12597 10057 12631
rect 10091 12628 10103 12631
rect 10226 12628 10232 12640
rect 10091 12600 10232 12628
rect 10091 12597 10103 12600
rect 10045 12591 10103 12597
rect 10226 12588 10232 12600
rect 10284 12588 10290 12640
rect 10428 12628 10456 12736
rect 10502 12724 10508 12776
rect 10560 12764 10566 12776
rect 10778 12764 10784 12776
rect 10560 12736 10784 12764
rect 10560 12724 10566 12736
rect 10778 12724 10784 12736
rect 10836 12724 10842 12776
rect 11256 12773 11284 12872
rect 14200 12844 14228 12872
rect 14476 12872 15240 12900
rect 11790 12792 11796 12844
rect 11848 12792 11854 12844
rect 12158 12792 12164 12844
rect 12216 12832 12222 12844
rect 12253 12835 12311 12841
rect 12253 12832 12265 12835
rect 12216 12804 12265 12832
rect 12216 12792 12222 12804
rect 12253 12801 12265 12804
rect 12299 12801 12311 12835
rect 12253 12795 12311 12801
rect 12342 12792 12348 12844
rect 12400 12832 12406 12844
rect 12529 12835 12587 12841
rect 12529 12832 12541 12835
rect 12400 12804 12541 12832
rect 12400 12792 12406 12804
rect 12529 12801 12541 12804
rect 12575 12801 12587 12835
rect 12529 12795 12587 12801
rect 12621 12835 12679 12841
rect 12621 12801 12633 12835
rect 12667 12832 12679 12835
rect 14090 12832 14096 12844
rect 12667 12804 14096 12832
rect 12667 12801 12679 12804
rect 12621 12795 12679 12801
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 14182 12792 14188 12844
rect 14240 12792 14246 12844
rect 14274 12792 14280 12844
rect 14332 12792 14338 12844
rect 14476 12832 14504 12872
rect 14384 12804 14504 12832
rect 11241 12767 11299 12773
rect 11241 12733 11253 12767
rect 11287 12733 11299 12767
rect 11241 12727 11299 12733
rect 11330 12724 11336 12776
rect 11388 12764 11394 12776
rect 11885 12767 11943 12773
rect 11885 12764 11897 12767
rect 11388 12736 11897 12764
rect 11388 12724 11394 12736
rect 11885 12733 11897 12736
rect 11931 12733 11943 12767
rect 11885 12727 11943 12733
rect 11977 12767 12035 12773
rect 11977 12733 11989 12767
rect 12023 12733 12035 12767
rect 11977 12727 12035 12733
rect 11606 12656 11612 12708
rect 11664 12656 11670 12708
rect 11992 12628 12020 12727
rect 12066 12724 12072 12776
rect 12124 12724 12130 12776
rect 14384 12773 14412 12804
rect 14642 12792 14648 12844
rect 14700 12832 14706 12844
rect 15010 12832 15016 12844
rect 14700 12804 15016 12832
rect 14700 12792 14706 12804
rect 15010 12792 15016 12804
rect 15068 12832 15074 12844
rect 15105 12835 15163 12841
rect 15105 12832 15117 12835
rect 15068 12804 15117 12832
rect 15068 12792 15074 12804
rect 15105 12801 15117 12804
rect 15151 12801 15163 12835
rect 15212 12832 15240 12872
rect 15286 12860 15292 12912
rect 15344 12900 15350 12912
rect 15841 12903 15899 12909
rect 15344 12872 15700 12900
rect 15344 12860 15350 12872
rect 15381 12835 15439 12841
rect 15381 12832 15393 12835
rect 15212 12804 15393 12832
rect 15105 12795 15163 12801
rect 15381 12801 15393 12804
rect 15427 12832 15439 12835
rect 15562 12832 15568 12844
rect 15427 12804 15568 12832
rect 15427 12801 15439 12804
rect 15381 12795 15439 12801
rect 15562 12792 15568 12804
rect 15620 12792 15626 12844
rect 15672 12841 15700 12872
rect 15841 12869 15853 12903
rect 15887 12900 15899 12903
rect 15887 12872 16712 12900
rect 15887 12869 15899 12872
rect 15841 12863 15899 12869
rect 15657 12835 15715 12841
rect 15657 12801 15669 12835
rect 15703 12801 15715 12835
rect 15657 12795 15715 12801
rect 15749 12835 15807 12841
rect 15749 12801 15761 12835
rect 15795 12832 15807 12835
rect 15795 12804 15884 12832
rect 15795 12801 15807 12804
rect 15749 12795 15807 12801
rect 15856 12776 15884 12804
rect 15930 12792 15936 12844
rect 15988 12841 15994 12844
rect 15988 12835 16017 12841
rect 16005 12801 16017 12835
rect 15988 12795 16017 12801
rect 15988 12792 15994 12795
rect 16114 12792 16120 12844
rect 16172 12792 16178 12844
rect 12897 12767 12955 12773
rect 12897 12733 12909 12767
rect 12943 12733 12955 12767
rect 12897 12727 12955 12733
rect 12989 12767 13047 12773
rect 12989 12733 13001 12767
rect 13035 12764 13047 12767
rect 14369 12767 14427 12773
rect 14369 12764 14381 12767
rect 13035 12736 14381 12764
rect 13035 12733 13047 12736
rect 12989 12727 13047 12733
rect 14369 12733 14381 12736
rect 14415 12733 14427 12767
rect 14369 12727 14427 12733
rect 14476 12736 15608 12764
rect 12912 12696 12940 12727
rect 14476 12696 14504 12736
rect 12912 12668 14504 12696
rect 13004 12640 13032 12668
rect 15102 12656 15108 12708
rect 15160 12696 15166 12708
rect 15580 12696 15608 12736
rect 15838 12724 15844 12776
rect 15896 12724 15902 12776
rect 16132 12696 16160 12792
rect 16684 12764 16712 12872
rect 16776 12872 18000 12900
rect 16776 12841 16804 12872
rect 17972 12844 18000 12872
rect 18064 12872 18736 12900
rect 18064 12844 18092 12872
rect 18708 12844 18736 12872
rect 18782 12860 18788 12912
rect 18840 12900 18846 12912
rect 22373 12903 22431 12909
rect 18840 12872 19334 12900
rect 18840 12860 18846 12872
rect 16761 12835 16819 12841
rect 16761 12801 16773 12835
rect 16807 12801 16819 12835
rect 16761 12795 16819 12801
rect 17405 12835 17463 12841
rect 17405 12801 17417 12835
rect 17451 12832 17463 12835
rect 17494 12832 17500 12844
rect 17451 12804 17500 12832
rect 17451 12801 17463 12804
rect 17405 12795 17463 12801
rect 17494 12792 17500 12804
rect 17552 12792 17558 12844
rect 17589 12835 17647 12841
rect 17589 12801 17601 12835
rect 17635 12801 17647 12835
rect 17589 12795 17647 12801
rect 17310 12764 17316 12776
rect 16684 12736 17316 12764
rect 17310 12724 17316 12736
rect 17368 12724 17374 12776
rect 17604 12764 17632 12795
rect 17862 12792 17868 12844
rect 17920 12792 17926 12844
rect 17954 12792 17960 12844
rect 18012 12792 18018 12844
rect 18046 12792 18052 12844
rect 18104 12792 18110 12844
rect 18598 12792 18604 12844
rect 18656 12792 18662 12844
rect 18690 12792 18696 12844
rect 18748 12792 18754 12844
rect 19306 12832 19334 12872
rect 22373 12869 22385 12903
rect 22419 12900 22431 12903
rect 22462 12900 22468 12912
rect 22419 12872 22468 12900
rect 22419 12869 22431 12872
rect 22373 12863 22431 12869
rect 22462 12860 22468 12872
rect 22520 12860 22526 12912
rect 23934 12860 23940 12912
rect 23992 12860 23998 12912
rect 24026 12860 24032 12912
rect 24084 12900 24090 12912
rect 24137 12903 24195 12909
rect 24137 12900 24149 12903
rect 24084 12872 24149 12900
rect 24084 12860 24090 12872
rect 24137 12869 24149 12872
rect 24183 12869 24195 12903
rect 24578 12900 24584 12912
rect 24137 12863 24195 12869
rect 24320 12872 24584 12900
rect 21358 12832 21364 12844
rect 19306 12804 21364 12832
rect 21358 12792 21364 12804
rect 21416 12792 21422 12844
rect 22097 12835 22155 12841
rect 22097 12801 22109 12835
rect 22143 12832 22155 12835
rect 22186 12832 22192 12844
rect 22143 12804 22192 12832
rect 22143 12801 22155 12804
rect 22097 12795 22155 12801
rect 22186 12792 22192 12804
rect 22244 12832 22250 12844
rect 22244 12804 23520 12832
rect 22244 12792 22250 12804
rect 23492 12776 23520 12804
rect 18325 12767 18383 12773
rect 18325 12764 18337 12767
rect 17604 12736 18337 12764
rect 18325 12733 18337 12736
rect 18371 12733 18383 12767
rect 18325 12727 18383 12733
rect 18509 12767 18567 12773
rect 18509 12733 18521 12767
rect 18555 12733 18567 12767
rect 18509 12727 18567 12733
rect 18785 12767 18843 12773
rect 18785 12733 18797 12767
rect 18831 12764 18843 12767
rect 19610 12764 19616 12776
rect 18831 12736 19616 12764
rect 18831 12733 18843 12736
rect 18785 12727 18843 12733
rect 15160 12668 15516 12696
rect 15580 12668 16160 12696
rect 15160 12656 15166 12668
rect 10428 12600 12020 12628
rect 12986 12588 12992 12640
rect 13044 12588 13050 12640
rect 14366 12588 14372 12640
rect 14424 12628 14430 12640
rect 14645 12631 14703 12637
rect 14645 12628 14657 12631
rect 14424 12600 14657 12628
rect 14424 12588 14430 12600
rect 14645 12597 14657 12600
rect 14691 12597 14703 12631
rect 14645 12591 14703 12597
rect 14921 12631 14979 12637
rect 14921 12597 14933 12631
rect 14967 12628 14979 12631
rect 15286 12628 15292 12640
rect 14967 12600 15292 12628
rect 14967 12597 14979 12600
rect 14921 12591 14979 12597
rect 15286 12588 15292 12600
rect 15344 12588 15350 12640
rect 15488 12637 15516 12668
rect 15473 12631 15531 12637
rect 15473 12597 15485 12631
rect 15519 12597 15531 12631
rect 17328 12628 17356 12724
rect 18524 12696 18552 12727
rect 19610 12724 19616 12736
rect 19668 12724 19674 12776
rect 23474 12724 23480 12776
rect 23532 12724 23538 12776
rect 18966 12696 18972 12708
rect 18524 12668 18972 12696
rect 18966 12656 18972 12668
rect 19024 12656 19030 12708
rect 24320 12696 24348 12872
rect 24578 12860 24584 12872
rect 24636 12860 24642 12912
rect 24688 12909 24716 12940
rect 24673 12903 24731 12909
rect 24673 12869 24685 12903
rect 24719 12869 24731 12903
rect 24673 12863 24731 12869
rect 25869 12903 25927 12909
rect 25869 12869 25881 12903
rect 25915 12900 25927 12903
rect 26344 12900 26372 12940
rect 26421 12937 26433 12971
rect 26467 12968 26479 12971
rect 26602 12968 26608 12980
rect 26467 12940 26608 12968
rect 26467 12937 26479 12940
rect 26421 12931 26479 12937
rect 26602 12928 26608 12940
rect 26660 12928 26666 12980
rect 29641 12971 29699 12977
rect 26804 12940 29316 12968
rect 26804 12900 26832 12940
rect 25915 12872 26280 12900
rect 26344 12872 26832 12900
rect 25915 12869 25927 12872
rect 25869 12863 25927 12869
rect 26252 12844 26280 12872
rect 27890 12860 27896 12912
rect 27948 12900 27954 12912
rect 29288 12909 29316 12940
rect 29641 12937 29653 12971
rect 29687 12968 29699 12971
rect 29730 12968 29736 12980
rect 29687 12940 29736 12968
rect 29687 12937 29699 12940
rect 29641 12931 29699 12937
rect 29730 12928 29736 12940
rect 29788 12928 29794 12980
rect 29825 12971 29883 12977
rect 29825 12937 29837 12971
rect 29871 12968 29883 12971
rect 30282 12968 30288 12980
rect 29871 12940 30288 12968
rect 29871 12937 29883 12940
rect 29825 12931 29883 12937
rect 30282 12928 30288 12940
rect 30340 12928 30346 12980
rect 31754 12928 31760 12980
rect 31812 12968 31818 12980
rect 32122 12968 32128 12980
rect 31812 12940 32128 12968
rect 31812 12928 31818 12940
rect 32122 12928 32128 12940
rect 32180 12968 32186 12980
rect 32401 12971 32459 12977
rect 32401 12968 32413 12971
rect 32180 12940 32413 12968
rect 32180 12928 32186 12940
rect 32401 12937 32413 12940
rect 32447 12968 32459 12971
rect 32582 12968 32588 12980
rect 32447 12940 32588 12968
rect 32447 12937 32459 12940
rect 32401 12931 32459 12937
rect 32582 12928 32588 12940
rect 32640 12928 32646 12980
rect 32769 12971 32827 12977
rect 32769 12937 32781 12971
rect 32815 12968 32827 12971
rect 32950 12968 32956 12980
rect 32815 12940 32956 12968
rect 32815 12937 32827 12940
rect 32769 12931 32827 12937
rect 32950 12928 32956 12940
rect 33008 12928 33014 12980
rect 33042 12928 33048 12980
rect 33100 12968 33106 12980
rect 33100 12940 34744 12968
rect 33100 12928 33106 12940
rect 28905 12903 28963 12909
rect 28905 12900 28917 12903
rect 27948 12872 28917 12900
rect 27948 12860 27954 12872
rect 28905 12869 28917 12872
rect 28951 12869 28963 12903
rect 28905 12863 28963 12869
rect 29273 12903 29331 12909
rect 29273 12869 29285 12903
rect 29319 12900 29331 12903
rect 30098 12900 30104 12912
rect 29319 12872 30104 12900
rect 29319 12869 29331 12872
rect 29273 12863 29331 12869
rect 30098 12860 30104 12872
rect 30156 12860 30162 12912
rect 31662 12860 31668 12912
rect 31720 12900 31726 12912
rect 32217 12903 32275 12909
rect 32217 12900 32229 12903
rect 31720 12872 32229 12900
rect 31720 12860 31726 12872
rect 32217 12869 32229 12872
rect 32263 12900 32275 12903
rect 32490 12900 32496 12912
rect 32263 12872 32496 12900
rect 32263 12869 32275 12872
rect 32217 12863 32275 12869
rect 32490 12860 32496 12872
rect 32548 12860 32554 12912
rect 32674 12860 32680 12912
rect 32732 12900 32738 12912
rect 32732 12872 34376 12900
rect 32732 12860 32738 12872
rect 24397 12835 24455 12841
rect 24397 12801 24409 12835
rect 24443 12801 24455 12835
rect 24397 12795 24455 12801
rect 24765 12835 24823 12841
rect 24765 12801 24777 12835
rect 24811 12832 24823 12835
rect 24854 12832 24860 12844
rect 24811 12804 24860 12832
rect 24811 12801 24823 12804
rect 24765 12795 24823 12801
rect 24412 12764 24440 12795
rect 24854 12792 24860 12804
rect 24912 12792 24918 12844
rect 25130 12792 25136 12844
rect 25188 12792 25194 12844
rect 26053 12835 26111 12841
rect 26053 12801 26065 12835
rect 26099 12801 26111 12835
rect 26053 12795 26111 12801
rect 25148 12764 25176 12792
rect 24412 12736 25176 12764
rect 25866 12724 25872 12776
rect 25924 12764 25930 12776
rect 26068 12764 26096 12795
rect 26234 12792 26240 12844
rect 26292 12832 26298 12844
rect 26329 12835 26387 12841
rect 26329 12832 26341 12835
rect 26292 12804 26341 12832
rect 26292 12792 26298 12804
rect 26329 12801 26341 12804
rect 26375 12801 26387 12835
rect 26329 12795 26387 12801
rect 26513 12835 26571 12841
rect 26513 12801 26525 12835
rect 26559 12832 26571 12835
rect 27706 12832 27712 12844
rect 26559 12804 27712 12832
rect 26559 12801 26571 12804
rect 26513 12795 26571 12801
rect 26528 12764 26556 12795
rect 27706 12792 27712 12804
rect 27764 12792 27770 12844
rect 29086 12792 29092 12844
rect 29144 12792 29150 12844
rect 29822 12832 29828 12844
rect 29783 12804 29828 12832
rect 29822 12792 29828 12804
rect 29880 12792 29886 12844
rect 32858 12832 32864 12844
rect 32600 12804 32864 12832
rect 25924 12736 26556 12764
rect 25924 12724 25930 12736
rect 26694 12724 26700 12776
rect 26752 12764 26758 12776
rect 27614 12764 27620 12776
rect 26752 12736 27620 12764
rect 26752 12724 26758 12736
rect 27614 12724 27620 12736
rect 27672 12724 27678 12776
rect 29104 12764 29132 12792
rect 30098 12764 30104 12776
rect 29104 12736 30104 12764
rect 30098 12724 30104 12736
rect 30156 12764 30162 12776
rect 30193 12767 30251 12773
rect 30193 12764 30205 12767
rect 30156 12736 30205 12764
rect 30156 12724 30162 12736
rect 30193 12733 30205 12736
rect 30239 12733 30251 12767
rect 30193 12727 30251 12733
rect 30285 12767 30343 12773
rect 30285 12733 30297 12767
rect 30331 12764 30343 12767
rect 31294 12764 31300 12776
rect 30331 12736 31300 12764
rect 30331 12733 30343 12736
rect 30285 12727 30343 12733
rect 31294 12724 31300 12736
rect 31352 12724 31358 12776
rect 32600 12705 32628 12804
rect 32858 12792 32864 12804
rect 32916 12832 32922 12844
rect 32953 12835 33011 12841
rect 32953 12832 32965 12835
rect 32916 12804 32965 12832
rect 32916 12792 32922 12804
rect 32953 12801 32965 12804
rect 32999 12801 33011 12835
rect 32953 12795 33011 12801
rect 33045 12835 33103 12841
rect 33045 12801 33057 12835
rect 33091 12801 33103 12835
rect 33045 12795 33103 12801
rect 32674 12724 32680 12776
rect 32732 12764 32738 12776
rect 33060 12764 33088 12795
rect 33134 12792 33140 12844
rect 33192 12832 33198 12844
rect 33229 12835 33287 12841
rect 33229 12832 33241 12835
rect 33192 12804 33241 12832
rect 33192 12792 33198 12804
rect 33229 12801 33241 12804
rect 33275 12801 33287 12835
rect 33229 12795 33287 12801
rect 33321 12835 33379 12841
rect 33321 12801 33333 12835
rect 33367 12801 33379 12835
rect 33321 12795 33379 12801
rect 32732 12736 33088 12764
rect 32732 12724 32738 12736
rect 23768 12668 24348 12696
rect 32585 12699 32643 12705
rect 19058 12628 19064 12640
rect 17328 12600 19064 12628
rect 15473 12591 15531 12597
rect 19058 12588 19064 12600
rect 19116 12588 19122 12640
rect 21910 12588 21916 12640
rect 21968 12588 21974 12640
rect 23290 12588 23296 12640
rect 23348 12628 23354 12640
rect 23768 12628 23796 12668
rect 32585 12665 32597 12699
rect 32631 12665 32643 12699
rect 32585 12659 32643 12665
rect 32950 12656 32956 12708
rect 33008 12696 33014 12708
rect 33336 12696 33364 12795
rect 33778 12792 33784 12844
rect 33836 12792 33842 12844
rect 33929 12835 33987 12841
rect 33929 12801 33941 12835
rect 33975 12801 33987 12835
rect 33929 12795 33987 12801
rect 33944 12764 33972 12795
rect 34054 12792 34060 12844
rect 34112 12792 34118 12844
rect 34146 12792 34152 12844
rect 34204 12792 34210 12844
rect 34246 12835 34304 12841
rect 34246 12801 34258 12835
rect 34292 12801 34304 12835
rect 34246 12795 34304 12801
rect 33944 12736 34192 12764
rect 34164 12708 34192 12736
rect 33008 12668 33364 12696
rect 33008 12656 33014 12668
rect 34146 12656 34152 12708
rect 34204 12656 34210 12708
rect 23348 12600 23796 12628
rect 23348 12588 23354 12600
rect 23842 12588 23848 12640
rect 23900 12628 23906 12640
rect 24118 12628 24124 12640
rect 23900 12600 24124 12628
rect 23900 12588 23906 12600
rect 24118 12588 24124 12600
rect 24176 12588 24182 12640
rect 24946 12588 24952 12640
rect 25004 12588 25010 12640
rect 25406 12588 25412 12640
rect 25464 12628 25470 12640
rect 26145 12631 26203 12637
rect 26145 12628 26157 12631
rect 25464 12600 26157 12628
rect 25464 12588 25470 12600
rect 26145 12597 26157 12600
rect 26191 12597 26203 12631
rect 26145 12591 26203 12597
rect 32306 12588 32312 12640
rect 32364 12628 32370 12640
rect 32401 12631 32459 12637
rect 32401 12628 32413 12631
rect 32364 12600 32413 12628
rect 32364 12588 32370 12600
rect 32401 12597 32413 12600
rect 32447 12597 32459 12631
rect 32401 12591 32459 12597
rect 33870 12588 33876 12640
rect 33928 12628 33934 12640
rect 34261 12628 34289 12795
rect 33928 12600 34289 12628
rect 34348 12628 34376 12872
rect 34716 12841 34744 12940
rect 34882 12928 34888 12980
rect 34940 12928 34946 12980
rect 35618 12928 35624 12980
rect 35676 12928 35682 12980
rect 35894 12928 35900 12980
rect 35952 12968 35958 12980
rect 36170 12968 36176 12980
rect 35952 12940 36176 12968
rect 35952 12928 35958 12940
rect 36170 12928 36176 12940
rect 36228 12928 36234 12980
rect 36725 12971 36783 12977
rect 36725 12937 36737 12971
rect 36771 12968 36783 12971
rect 38194 12968 38200 12980
rect 36771 12940 38200 12968
rect 36771 12937 36783 12940
rect 36725 12931 36783 12937
rect 38194 12928 38200 12940
rect 38252 12928 38258 12980
rect 39393 12971 39451 12977
rect 39393 12937 39405 12971
rect 39439 12968 39451 12971
rect 39850 12968 39856 12980
rect 39439 12940 39856 12968
rect 39439 12937 39451 12940
rect 39393 12931 39451 12937
rect 39850 12928 39856 12940
rect 39908 12928 39914 12980
rect 34701 12835 34759 12841
rect 34701 12801 34713 12835
rect 34747 12801 34759 12835
rect 35636 12832 35664 12928
rect 38930 12860 38936 12912
rect 38988 12900 38994 12912
rect 39025 12903 39083 12909
rect 39025 12900 39037 12903
rect 38988 12872 39037 12900
rect 38988 12860 38994 12872
rect 39025 12869 39037 12872
rect 39071 12869 39083 12903
rect 39025 12863 39083 12869
rect 39114 12860 39120 12912
rect 39172 12860 39178 12912
rect 36357 12835 36415 12841
rect 36357 12832 36369 12835
rect 35636 12804 36369 12832
rect 34701 12795 34759 12801
rect 36357 12801 36369 12804
rect 36403 12801 36415 12835
rect 36357 12795 36415 12801
rect 36538 12792 36544 12844
rect 36596 12792 36602 12844
rect 38838 12792 38844 12844
rect 38896 12792 38902 12844
rect 39209 12835 39267 12841
rect 39209 12801 39221 12835
rect 39255 12832 39267 12835
rect 39390 12832 39396 12844
rect 39255 12804 39396 12832
rect 39255 12801 39267 12804
rect 39209 12795 39267 12801
rect 34514 12724 34520 12776
rect 34572 12724 34578 12776
rect 38654 12724 38660 12776
rect 38712 12764 38718 12776
rect 39224 12764 39252 12795
rect 39390 12792 39396 12804
rect 39448 12792 39454 12844
rect 38712 12736 39252 12764
rect 38712 12724 38718 12736
rect 34425 12699 34483 12705
rect 34425 12665 34437 12699
rect 34471 12696 34483 12699
rect 35250 12696 35256 12708
rect 34471 12668 35256 12696
rect 34471 12665 34483 12668
rect 34425 12659 34483 12665
rect 35250 12656 35256 12668
rect 35308 12656 35314 12708
rect 38930 12656 38936 12708
rect 38988 12696 38994 12708
rect 39482 12696 39488 12708
rect 38988 12668 39488 12696
rect 38988 12656 38994 12668
rect 39482 12656 39488 12668
rect 39540 12656 39546 12708
rect 36357 12631 36415 12637
rect 36357 12628 36369 12631
rect 34348 12600 36369 12628
rect 33928 12588 33934 12600
rect 36357 12597 36369 12600
rect 36403 12597 36415 12631
rect 36357 12591 36415 12597
rect 1104 12538 41400 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 41400 12538
rect 1104 12464 41400 12486
rect 4341 12427 4399 12433
rect 4341 12393 4353 12427
rect 4387 12424 4399 12427
rect 5261 12427 5319 12433
rect 5261 12424 5273 12427
rect 4387 12396 5273 12424
rect 4387 12393 4399 12396
rect 4341 12387 4399 12393
rect 5261 12393 5273 12396
rect 5307 12393 5319 12427
rect 5261 12387 5319 12393
rect 6454 12384 6460 12436
rect 6512 12424 6518 12436
rect 7101 12427 7159 12433
rect 7101 12424 7113 12427
rect 6512 12396 7113 12424
rect 6512 12384 6518 12396
rect 7101 12393 7113 12396
rect 7147 12393 7159 12427
rect 7101 12387 7159 12393
rect 8202 12384 8208 12436
rect 8260 12384 8266 12436
rect 10413 12427 10471 12433
rect 10413 12393 10425 12427
rect 10459 12424 10471 12427
rect 11054 12424 11060 12436
rect 10459 12396 11060 12424
rect 10459 12393 10471 12396
rect 10413 12387 10471 12393
rect 11054 12384 11060 12396
rect 11112 12384 11118 12436
rect 14921 12427 14979 12433
rect 11164 12396 14872 12424
rect 4890 12356 4896 12368
rect 4448 12328 4896 12356
rect 3973 12223 4031 12229
rect 3973 12189 3985 12223
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 4065 12223 4123 12229
rect 4065 12189 4077 12223
rect 4111 12220 4123 12223
rect 4338 12220 4344 12232
rect 4111 12192 4344 12220
rect 4111 12189 4123 12192
rect 4065 12183 4123 12189
rect 3988 12096 4016 12183
rect 4338 12180 4344 12192
rect 4396 12180 4402 12232
rect 4448 12229 4476 12328
rect 4890 12316 4896 12328
rect 4948 12316 4954 12368
rect 5629 12359 5687 12365
rect 5629 12325 5641 12359
rect 5675 12356 5687 12359
rect 7374 12356 7380 12368
rect 5675 12328 7380 12356
rect 5675 12325 5687 12328
rect 5629 12319 5687 12325
rect 7374 12316 7380 12328
rect 7432 12316 7438 12368
rect 8220 12356 8248 12384
rect 11164 12356 11192 12396
rect 14844 12368 14872 12396
rect 14921 12393 14933 12427
rect 14967 12424 14979 12427
rect 15102 12424 15108 12436
rect 14967 12396 15108 12424
rect 14967 12393 14979 12396
rect 14921 12387 14979 12393
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 15378 12384 15384 12436
rect 15436 12384 15442 12436
rect 17218 12384 17224 12436
rect 17276 12424 17282 12436
rect 18138 12424 18144 12436
rect 17276 12396 18144 12424
rect 17276 12384 17282 12396
rect 18138 12384 18144 12396
rect 18196 12384 18202 12436
rect 18966 12384 18972 12436
rect 19024 12384 19030 12436
rect 19334 12384 19340 12436
rect 19392 12424 19398 12436
rect 19429 12427 19487 12433
rect 19429 12424 19441 12427
rect 19392 12396 19441 12424
rect 19392 12384 19398 12396
rect 19429 12393 19441 12396
rect 19475 12393 19487 12427
rect 19429 12387 19487 12393
rect 8220 12328 11192 12356
rect 14369 12359 14427 12365
rect 14369 12325 14381 12359
rect 14415 12356 14427 12359
rect 14734 12356 14740 12368
rect 14415 12328 14740 12356
rect 14415 12325 14427 12328
rect 14369 12319 14427 12325
rect 14734 12316 14740 12328
rect 14792 12316 14798 12368
rect 14826 12316 14832 12368
rect 14884 12316 14890 12368
rect 15013 12359 15071 12365
rect 15013 12325 15025 12359
rect 15059 12356 15071 12359
rect 15396 12356 15424 12384
rect 15059 12328 15424 12356
rect 15059 12325 15071 12328
rect 15013 12319 15071 12325
rect 5258 12288 5264 12300
rect 4724 12260 5264 12288
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12189 4491 12223
rect 4433 12183 4491 12189
rect 4724 12152 4752 12260
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 6362 12248 6368 12300
rect 6420 12288 6426 12300
rect 7282 12288 7288 12300
rect 6420 12260 7288 12288
rect 6420 12248 6426 12260
rect 7282 12248 7288 12260
rect 7340 12248 7346 12300
rect 11146 12288 11152 12300
rect 10612 12260 11152 12288
rect 4798 12180 4804 12232
rect 4856 12180 4862 12232
rect 4890 12180 4896 12232
rect 4948 12180 4954 12232
rect 4982 12180 4988 12232
rect 5040 12180 5046 12232
rect 5077 12223 5135 12229
rect 5077 12189 5089 12223
rect 5123 12189 5135 12223
rect 5077 12183 5135 12189
rect 4448 12124 4752 12152
rect 5092 12152 5120 12183
rect 5350 12180 5356 12232
rect 5408 12220 5414 12232
rect 5445 12223 5503 12229
rect 5445 12220 5457 12223
rect 5408 12192 5457 12220
rect 5408 12180 5414 12192
rect 5445 12189 5457 12192
rect 5491 12189 5503 12223
rect 5445 12183 5503 12189
rect 5537 12223 5595 12229
rect 5537 12189 5549 12223
rect 5583 12189 5595 12223
rect 5537 12183 5595 12189
rect 5721 12223 5779 12229
rect 5721 12189 5733 12223
rect 5767 12189 5779 12223
rect 5721 12183 5779 12189
rect 5552 12152 5580 12183
rect 5092 12124 5580 12152
rect 3970 12044 3976 12096
rect 4028 12044 4034 12096
rect 4157 12087 4215 12093
rect 4157 12053 4169 12087
rect 4203 12084 4215 12087
rect 4338 12084 4344 12096
rect 4203 12056 4344 12084
rect 4203 12053 4215 12056
rect 4157 12047 4215 12053
rect 4338 12044 4344 12056
rect 4396 12044 4402 12096
rect 4448 12093 4476 12124
rect 4433 12087 4491 12093
rect 4433 12053 4445 12087
rect 4479 12053 4491 12087
rect 4433 12047 4491 12053
rect 4617 12087 4675 12093
rect 4617 12053 4629 12087
rect 4663 12084 4675 12087
rect 5442 12084 5448 12096
rect 4663 12056 5448 12084
rect 4663 12053 4675 12056
rect 4617 12047 4675 12053
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 5552 12084 5580 12124
rect 5626 12112 5632 12164
rect 5684 12152 5690 12164
rect 5736 12152 5764 12183
rect 5902 12180 5908 12232
rect 5960 12180 5966 12232
rect 5684 12124 6408 12152
rect 5684 12112 5690 12124
rect 6380 12096 6408 12124
rect 6638 12112 6644 12164
rect 6696 12112 6702 12164
rect 6917 12155 6975 12161
rect 6917 12121 6929 12155
rect 6963 12152 6975 12155
rect 7006 12152 7012 12164
rect 6963 12124 7012 12152
rect 6963 12121 6975 12124
rect 6917 12115 6975 12121
rect 7006 12112 7012 12124
rect 7064 12112 7070 12164
rect 7133 12155 7191 12161
rect 7133 12121 7145 12155
rect 7179 12152 7191 12155
rect 7300 12152 7328 12248
rect 9030 12180 9036 12232
rect 9088 12180 9094 12232
rect 9122 12180 9128 12232
rect 9180 12180 9186 12232
rect 10612 12229 10640 12260
rect 11146 12248 11152 12260
rect 11204 12248 11210 12300
rect 12161 12291 12219 12297
rect 12161 12257 12173 12291
rect 12207 12288 12219 12291
rect 16574 12288 16580 12300
rect 12207 12260 16580 12288
rect 12207 12257 12219 12260
rect 12161 12251 12219 12257
rect 16574 12248 16580 12260
rect 16632 12248 16638 12300
rect 18984 12288 19012 12384
rect 19444 12356 19472 12387
rect 19610 12384 19616 12436
rect 19668 12424 19674 12436
rect 20070 12424 20076 12436
rect 19668 12396 20076 12424
rect 19668 12384 19674 12396
rect 20070 12384 20076 12396
rect 20128 12384 20134 12436
rect 23474 12384 23480 12436
rect 23532 12384 23538 12436
rect 23934 12424 23940 12436
rect 23584 12396 23940 12424
rect 23293 12359 23351 12365
rect 19444 12328 19886 12356
rect 18984 12260 19748 12288
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12220 9367 12223
rect 10597 12223 10655 12229
rect 10597 12220 10609 12223
rect 9355 12192 10609 12220
rect 9355 12189 9367 12192
rect 9309 12183 9367 12189
rect 10597 12189 10609 12192
rect 10643 12189 10655 12223
rect 10597 12183 10655 12189
rect 10686 12180 10692 12232
rect 10744 12180 10750 12232
rect 14274 12180 14280 12232
rect 14332 12180 14338 12232
rect 14458 12180 14464 12232
rect 14516 12220 14522 12232
rect 14829 12223 14887 12229
rect 14829 12220 14841 12223
rect 14516 12192 14841 12220
rect 14516 12180 14522 12192
rect 14829 12189 14841 12192
rect 14875 12189 14887 12223
rect 14829 12183 14887 12189
rect 15102 12180 15108 12232
rect 15160 12180 15166 12232
rect 15289 12223 15347 12229
rect 15289 12189 15301 12223
rect 15335 12220 15347 12223
rect 15746 12220 15752 12232
rect 15335 12192 15752 12220
rect 15335 12189 15347 12192
rect 15289 12183 15347 12189
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 17126 12180 17132 12232
rect 17184 12220 17190 12232
rect 17310 12220 17316 12232
rect 17184 12192 17316 12220
rect 17184 12180 17190 12192
rect 17310 12180 17316 12192
rect 17368 12180 17374 12232
rect 17494 12180 17500 12232
rect 17552 12180 17558 12232
rect 18782 12180 18788 12232
rect 18840 12180 18846 12232
rect 18877 12223 18935 12229
rect 18877 12189 18889 12223
rect 18923 12189 18935 12223
rect 18877 12183 18935 12189
rect 7179 12124 7328 12152
rect 10413 12155 10471 12161
rect 7179 12121 7191 12124
rect 7133 12115 7191 12121
rect 10413 12121 10425 12155
rect 10459 12152 10471 12155
rect 11146 12152 11152 12164
rect 10459 12124 11152 12152
rect 10459 12121 10471 12124
rect 10413 12115 10471 12121
rect 11146 12112 11152 12124
rect 11204 12112 11210 12164
rect 12437 12155 12495 12161
rect 12437 12121 12449 12155
rect 12483 12152 12495 12155
rect 12710 12152 12716 12164
rect 12483 12124 12716 12152
rect 12483 12121 12495 12124
rect 12437 12115 12495 12121
rect 12710 12112 12716 12124
rect 12768 12112 12774 12164
rect 13078 12112 13084 12164
rect 13136 12112 13142 12164
rect 13722 12112 13728 12164
rect 13780 12152 13786 12164
rect 13780 12124 14044 12152
rect 13780 12112 13786 12124
rect 5810 12084 5816 12096
rect 5552 12056 5816 12084
rect 5810 12044 5816 12056
rect 5868 12044 5874 12096
rect 6362 12044 6368 12096
rect 6420 12044 6426 12096
rect 7282 12044 7288 12096
rect 7340 12044 7346 12096
rect 13814 12044 13820 12096
rect 13872 12084 13878 12096
rect 13909 12087 13967 12093
rect 13909 12084 13921 12087
rect 13872 12056 13921 12084
rect 13872 12044 13878 12056
rect 13909 12053 13921 12056
rect 13955 12053 13967 12087
rect 14016 12084 14044 12124
rect 14090 12112 14096 12164
rect 14148 12152 14154 12164
rect 14553 12155 14611 12161
rect 14553 12152 14565 12155
rect 14148 12124 14565 12152
rect 14148 12112 14154 12124
rect 14553 12121 14565 12124
rect 14599 12121 14611 12155
rect 14553 12115 14611 12121
rect 17405 12087 17463 12093
rect 17405 12084 17417 12087
rect 14016 12056 17417 12084
rect 13909 12047 13967 12053
rect 17405 12053 17417 12056
rect 17451 12053 17463 12087
rect 17405 12047 17463 12053
rect 18598 12044 18604 12096
rect 18656 12044 18662 12096
rect 18892 12084 18920 12183
rect 19058 12180 19064 12232
rect 19116 12180 19122 12232
rect 19720 12229 19748 12260
rect 19858 12229 19886 12328
rect 21100 12328 21956 12356
rect 21100 12300 21128 12328
rect 21928 12300 21956 12328
rect 23293 12325 23305 12359
rect 23339 12356 23351 12359
rect 23584 12356 23612 12396
rect 23934 12384 23940 12396
rect 23992 12384 23998 12436
rect 24854 12384 24860 12436
rect 24912 12424 24918 12436
rect 24949 12427 25007 12433
rect 24949 12424 24961 12427
rect 24912 12396 24961 12424
rect 24912 12384 24918 12396
rect 24949 12393 24961 12396
rect 24995 12393 25007 12427
rect 24949 12387 25007 12393
rect 25590 12384 25596 12436
rect 25648 12384 25654 12436
rect 25866 12384 25872 12436
rect 25924 12384 25930 12436
rect 26050 12384 26056 12436
rect 26108 12384 26114 12436
rect 26145 12427 26203 12433
rect 26145 12393 26157 12427
rect 26191 12393 26203 12427
rect 26145 12387 26203 12393
rect 25608 12356 25636 12384
rect 26160 12356 26188 12387
rect 26602 12384 26608 12436
rect 26660 12384 26666 12436
rect 26697 12427 26755 12433
rect 26697 12393 26709 12427
rect 26743 12424 26755 12427
rect 26878 12424 26884 12436
rect 26743 12396 26884 12424
rect 26743 12393 26755 12396
rect 26697 12387 26755 12393
rect 26878 12384 26884 12396
rect 26936 12384 26942 12436
rect 31570 12424 31576 12436
rect 30300 12396 31576 12424
rect 23339 12328 23612 12356
rect 23768 12328 24072 12356
rect 25608 12328 26188 12356
rect 23339 12325 23351 12328
rect 23293 12319 23351 12325
rect 21082 12248 21088 12300
rect 21140 12248 21146 12300
rect 21358 12248 21364 12300
rect 21416 12248 21422 12300
rect 21542 12248 21548 12300
rect 21600 12248 21606 12300
rect 21910 12248 21916 12300
rect 21968 12248 21974 12300
rect 23474 12248 23480 12300
rect 23532 12248 23538 12300
rect 23768 12297 23796 12328
rect 24044 12300 24072 12328
rect 23753 12291 23811 12297
rect 23753 12257 23765 12291
rect 23799 12257 23811 12291
rect 23753 12251 23811 12257
rect 23842 12248 23848 12300
rect 23900 12248 23906 12300
rect 24026 12248 24032 12300
rect 24084 12248 24090 12300
rect 24596 12260 25636 12288
rect 19705 12223 19763 12229
rect 19705 12189 19717 12223
rect 19751 12189 19763 12223
rect 19705 12183 19763 12189
rect 19843 12223 19901 12229
rect 19843 12189 19855 12223
rect 19889 12189 19901 12223
rect 19843 12183 19901 12189
rect 20254 12180 20260 12232
rect 20312 12180 20318 12232
rect 21729 12223 21787 12229
rect 21729 12189 21741 12223
rect 21775 12189 21787 12223
rect 21729 12183 21787 12189
rect 23201 12223 23259 12229
rect 23201 12189 23213 12223
rect 23247 12220 23259 12223
rect 23290 12220 23296 12232
rect 23247 12192 23296 12220
rect 23247 12189 23259 12192
rect 23201 12183 23259 12189
rect 19076 12152 19104 12180
rect 19245 12155 19303 12161
rect 19245 12152 19257 12155
rect 19076 12124 19257 12152
rect 19245 12121 19257 12124
rect 19291 12121 19303 12155
rect 19461 12155 19519 12161
rect 19461 12152 19473 12155
rect 19245 12115 19303 12121
rect 19352 12124 19473 12152
rect 19352 12084 19380 12124
rect 19461 12121 19473 12124
rect 19507 12152 19519 12155
rect 20272 12152 20300 12180
rect 19507 12124 20300 12152
rect 21744 12152 21772 12183
rect 23290 12180 23296 12192
rect 23348 12180 23354 12232
rect 23385 12223 23443 12229
rect 23385 12189 23397 12223
rect 23431 12220 23443 12223
rect 23492 12220 23520 12248
rect 23431 12192 23520 12220
rect 23431 12189 23443 12192
rect 23385 12183 23443 12189
rect 23658 12180 23664 12232
rect 23716 12180 23722 12232
rect 23937 12223 23995 12229
rect 23937 12189 23949 12223
rect 23983 12220 23995 12223
rect 24394 12220 24400 12232
rect 23983 12192 24400 12220
rect 23983 12189 23995 12192
rect 23937 12183 23995 12189
rect 23952 12152 23980 12183
rect 24394 12180 24400 12192
rect 24452 12180 24458 12232
rect 24596 12161 24624 12260
rect 25608 12232 25636 12260
rect 24765 12223 24823 12229
rect 24765 12189 24777 12223
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 21744 12124 23980 12152
rect 24581 12155 24639 12161
rect 19507 12121 19519 12124
rect 19461 12115 19519 12121
rect 24581 12121 24593 12155
rect 24627 12121 24639 12155
rect 24780 12152 24808 12183
rect 25590 12180 25596 12232
rect 25648 12180 25654 12232
rect 25701 12220 25729 12328
rect 25777 12291 25835 12297
rect 25777 12257 25789 12291
rect 25823 12288 25835 12291
rect 26050 12288 26056 12300
rect 25823 12260 26056 12288
rect 25823 12257 25835 12260
rect 25777 12251 25835 12257
rect 26050 12248 26056 12260
rect 26108 12248 26114 12300
rect 26252 12260 27292 12288
rect 25866 12220 25872 12232
rect 25701 12192 25872 12220
rect 25866 12180 25872 12192
rect 25924 12180 25930 12232
rect 25682 12152 25688 12164
rect 24780 12124 25688 12152
rect 24581 12115 24639 12121
rect 18892 12056 19380 12084
rect 19978 12044 19984 12096
rect 20036 12084 20042 12096
rect 20073 12087 20131 12093
rect 20073 12084 20085 12087
rect 20036 12056 20085 12084
rect 20036 12044 20042 12056
rect 20073 12053 20085 12056
rect 20119 12053 20131 12087
rect 20073 12047 20131 12053
rect 20898 12044 20904 12096
rect 20956 12044 20962 12096
rect 21269 12087 21327 12093
rect 21269 12053 21281 12087
rect 21315 12084 21327 12087
rect 21358 12084 21364 12096
rect 21315 12056 21364 12084
rect 21315 12053 21327 12056
rect 21269 12047 21327 12053
rect 21358 12044 21364 12056
rect 21416 12044 21422 12096
rect 23106 12044 23112 12096
rect 23164 12084 23170 12096
rect 24596 12084 24624 12115
rect 25682 12112 25688 12124
rect 25740 12152 25746 12164
rect 26050 12152 26056 12164
rect 25740 12124 26056 12152
rect 25740 12112 25746 12124
rect 26050 12112 26056 12124
rect 26108 12112 26114 12164
rect 26145 12155 26203 12161
rect 26145 12121 26157 12155
rect 26191 12152 26203 12155
rect 26252 12152 26280 12260
rect 26326 12180 26332 12232
rect 26384 12180 26390 12232
rect 26421 12223 26479 12229
rect 26421 12189 26433 12223
rect 26467 12220 26479 12223
rect 26602 12220 26608 12232
rect 26467 12192 26608 12220
rect 26467 12189 26479 12192
rect 26421 12183 26479 12189
rect 26602 12180 26608 12192
rect 26660 12180 26666 12232
rect 26881 12223 26939 12229
rect 26881 12189 26893 12223
rect 26927 12189 26939 12223
rect 26881 12183 26939 12189
rect 26191 12124 26280 12152
rect 26896 12152 26924 12183
rect 26970 12180 26976 12232
rect 27028 12180 27034 12232
rect 27062 12180 27068 12232
rect 27120 12220 27126 12232
rect 27264 12229 27292 12260
rect 28626 12248 28632 12300
rect 28684 12288 28690 12300
rect 28684 12260 28994 12288
rect 28684 12248 28690 12260
rect 27157 12223 27215 12229
rect 27157 12220 27169 12223
rect 27120 12192 27169 12220
rect 27120 12180 27126 12192
rect 27157 12189 27169 12192
rect 27203 12189 27215 12223
rect 27157 12183 27215 12189
rect 27249 12223 27307 12229
rect 27249 12189 27261 12223
rect 27295 12220 27307 12223
rect 27295 12192 27472 12220
rect 27295 12189 27307 12192
rect 27249 12183 27307 12189
rect 27341 12155 27399 12161
rect 27341 12152 27353 12155
rect 26896 12124 27353 12152
rect 26191 12121 26203 12124
rect 26145 12115 26203 12121
rect 27341 12121 27353 12124
rect 27387 12121 27399 12155
rect 27444 12152 27472 12192
rect 27522 12180 27528 12232
rect 27580 12180 27586 12232
rect 27614 12180 27620 12232
rect 27672 12180 27678 12232
rect 27706 12180 27712 12232
rect 27764 12220 27770 12232
rect 27801 12223 27859 12229
rect 27801 12220 27813 12223
rect 27764 12192 27813 12220
rect 27764 12180 27770 12192
rect 27801 12189 27813 12192
rect 27847 12189 27859 12223
rect 27801 12183 27859 12189
rect 27893 12223 27951 12229
rect 27893 12189 27905 12223
rect 27939 12220 27951 12223
rect 28074 12220 28080 12232
rect 27939 12192 28080 12220
rect 27939 12189 27951 12192
rect 27893 12183 27951 12189
rect 28074 12180 28080 12192
rect 28132 12180 28138 12232
rect 28966 12152 28994 12260
rect 29380 12260 29868 12288
rect 29380 12232 29408 12260
rect 29362 12180 29368 12232
rect 29420 12180 29426 12232
rect 29840 12229 29868 12260
rect 29549 12223 29607 12229
rect 29549 12189 29561 12223
rect 29595 12189 29607 12223
rect 29549 12183 29607 12189
rect 29825 12223 29883 12229
rect 29825 12189 29837 12223
rect 29871 12189 29883 12223
rect 29825 12183 29883 12189
rect 29564 12152 29592 12183
rect 29914 12180 29920 12232
rect 29972 12220 29978 12232
rect 30009 12223 30067 12229
rect 30009 12220 30021 12223
rect 29972 12192 30021 12220
rect 29972 12180 29978 12192
rect 30009 12189 30021 12192
rect 30055 12189 30067 12223
rect 30009 12183 30067 12189
rect 30193 12223 30251 12229
rect 30193 12189 30205 12223
rect 30239 12189 30251 12223
rect 30300 12220 30328 12396
rect 31570 12384 31576 12396
rect 31628 12424 31634 12436
rect 32217 12427 32275 12433
rect 31628 12396 32076 12424
rect 31628 12384 31634 12396
rect 31018 12316 31024 12368
rect 31076 12316 31082 12368
rect 32048 12356 32076 12396
rect 32217 12393 32229 12427
rect 32263 12424 32275 12427
rect 32306 12424 32312 12436
rect 32263 12396 32312 12424
rect 32263 12393 32275 12396
rect 32217 12387 32275 12393
rect 32306 12384 32312 12396
rect 32364 12424 32370 12436
rect 33042 12424 33048 12436
rect 32364 12396 33048 12424
rect 32364 12384 32370 12396
rect 33042 12384 33048 12396
rect 33100 12424 33106 12436
rect 33413 12427 33471 12433
rect 33413 12424 33425 12427
rect 33100 12396 33425 12424
rect 33100 12384 33106 12396
rect 33413 12393 33425 12396
rect 33459 12393 33471 12427
rect 33413 12387 33471 12393
rect 33502 12384 33508 12436
rect 33560 12424 33566 12436
rect 33597 12427 33655 12433
rect 33597 12424 33609 12427
rect 33560 12396 33609 12424
rect 33560 12384 33566 12396
rect 33597 12393 33609 12396
rect 33643 12393 33655 12427
rect 33597 12387 33655 12393
rect 34241 12427 34299 12433
rect 34241 12393 34253 12427
rect 34287 12424 34299 12427
rect 37182 12424 37188 12436
rect 34287 12396 37188 12424
rect 34287 12393 34299 12396
rect 34241 12387 34299 12393
rect 37182 12384 37188 12396
rect 37240 12424 37246 12436
rect 38102 12424 38108 12436
rect 37240 12396 38108 12424
rect 37240 12384 37246 12396
rect 38102 12384 38108 12396
rect 38160 12384 38166 12436
rect 32048 12328 33088 12356
rect 30374 12248 30380 12300
rect 30432 12248 30438 12300
rect 31297 12291 31355 12297
rect 31297 12257 31309 12291
rect 31343 12288 31355 12291
rect 31343 12260 32168 12288
rect 31343 12257 31355 12260
rect 31297 12251 31355 12257
rect 30466 12220 30472 12232
rect 30300 12192 30472 12220
rect 30193 12183 30251 12189
rect 29730 12152 29736 12164
rect 27444 12124 27936 12152
rect 28966 12124 29736 12152
rect 27341 12115 27399 12121
rect 23164 12056 24624 12084
rect 23164 12044 23170 12056
rect 24670 12044 24676 12096
rect 24728 12084 24734 12096
rect 26160 12084 26188 12115
rect 27908 12096 27936 12124
rect 29730 12112 29736 12124
rect 29788 12112 29794 12164
rect 24728 12056 26188 12084
rect 24728 12044 24734 12056
rect 26510 12044 26516 12096
rect 26568 12084 26574 12096
rect 27062 12084 27068 12096
rect 26568 12056 27068 12084
rect 26568 12044 26574 12056
rect 27062 12044 27068 12056
rect 27120 12044 27126 12096
rect 27890 12044 27896 12096
rect 27948 12044 27954 12096
rect 30208 12084 30236 12183
rect 30466 12180 30472 12192
rect 30524 12180 30530 12232
rect 30653 12223 30711 12229
rect 30653 12189 30665 12223
rect 30699 12220 30711 12223
rect 31312 12220 31340 12251
rect 30699 12192 31340 12220
rect 30699 12189 30711 12192
rect 30653 12183 30711 12189
rect 31570 12180 31576 12232
rect 31628 12180 31634 12232
rect 32140 12229 32168 12260
rect 32306 12248 32312 12300
rect 32364 12248 32370 12300
rect 32033 12223 32091 12229
rect 32033 12189 32045 12223
rect 32079 12189 32091 12223
rect 32033 12183 32091 12189
rect 32125 12223 32183 12229
rect 32125 12189 32137 12223
rect 32171 12220 32183 12223
rect 32582 12220 32588 12232
rect 32171 12192 32588 12220
rect 32171 12189 32183 12192
rect 32125 12183 32183 12189
rect 30282 12112 30288 12164
rect 30340 12152 30346 12164
rect 30837 12155 30895 12161
rect 30837 12152 30849 12155
rect 30340 12124 30849 12152
rect 30340 12112 30346 12124
rect 30837 12121 30849 12124
rect 30883 12152 30895 12155
rect 31202 12152 31208 12164
rect 30883 12124 31208 12152
rect 30883 12121 30895 12124
rect 30837 12115 30895 12121
rect 31202 12112 31208 12124
rect 31260 12112 31266 12164
rect 31386 12112 31392 12164
rect 31444 12152 31450 12164
rect 31665 12155 31723 12161
rect 31665 12152 31677 12155
rect 31444 12124 31677 12152
rect 31444 12112 31450 12124
rect 31665 12121 31677 12124
rect 31711 12121 31723 12155
rect 31665 12115 31723 12121
rect 31782 12155 31840 12161
rect 31782 12121 31794 12155
rect 31828 12152 31840 12155
rect 32048 12152 32076 12183
rect 32582 12180 32588 12192
rect 32640 12180 32646 12232
rect 33060 12220 33088 12328
rect 33134 12316 33140 12368
rect 33192 12356 33198 12368
rect 39022 12356 39028 12368
rect 33192 12328 39028 12356
rect 33192 12316 33198 12328
rect 39022 12316 39028 12328
rect 39080 12316 39086 12368
rect 33686 12248 33692 12300
rect 33744 12288 33750 12300
rect 35250 12288 35256 12300
rect 33744 12260 35256 12288
rect 33744 12248 33750 12260
rect 35250 12248 35256 12260
rect 35308 12248 35314 12300
rect 36446 12248 36452 12300
rect 36504 12288 36510 12300
rect 36998 12288 37004 12300
rect 36504 12260 37004 12288
rect 36504 12248 36510 12260
rect 36998 12248 37004 12260
rect 37056 12248 37062 12300
rect 32692 12192 32904 12220
rect 33060 12192 33472 12220
rect 31828 12124 32076 12152
rect 31828 12121 31840 12124
rect 31782 12115 31840 12121
rect 30374 12084 30380 12096
rect 30208 12056 30380 12084
rect 30374 12044 30380 12056
rect 30432 12044 30438 12096
rect 30650 12044 30656 12096
rect 30708 12044 30714 12096
rect 30926 12044 30932 12096
rect 30984 12084 30990 12096
rect 31797 12084 31825 12115
rect 32490 12112 32496 12164
rect 32548 12152 32554 12164
rect 32692 12152 32720 12192
rect 32548 12124 32720 12152
rect 32548 12112 32554 12124
rect 32766 12112 32772 12164
rect 32824 12112 32830 12164
rect 30984 12056 31825 12084
rect 31941 12087 31999 12093
rect 30984 12044 30990 12056
rect 31941 12053 31953 12087
rect 31987 12084 31999 12087
rect 32784 12084 32812 12112
rect 31987 12056 32812 12084
rect 32876 12084 32904 12192
rect 33134 12112 33140 12164
rect 33192 12112 33198 12164
rect 33444 12161 33472 12192
rect 34054 12180 34060 12232
rect 34112 12180 34118 12232
rect 34330 12180 34336 12232
rect 34388 12220 34394 12232
rect 35802 12220 35808 12232
rect 34388 12192 35808 12220
rect 34388 12180 34394 12192
rect 35802 12180 35808 12192
rect 35860 12180 35866 12232
rect 36262 12180 36268 12232
rect 36320 12180 36326 12232
rect 33229 12155 33287 12161
rect 33229 12121 33241 12155
rect 33275 12121 33287 12155
rect 33229 12115 33287 12121
rect 33429 12155 33487 12161
rect 33429 12121 33441 12155
rect 33475 12121 33487 12155
rect 33429 12115 33487 12121
rect 33244 12084 33272 12115
rect 33594 12112 33600 12164
rect 33652 12152 33658 12164
rect 36280 12152 36308 12180
rect 37182 12152 37188 12164
rect 33652 12124 37188 12152
rect 33652 12112 33658 12124
rect 37182 12112 37188 12124
rect 37240 12112 37246 12164
rect 34514 12084 34520 12096
rect 32876 12056 34520 12084
rect 31987 12053 31999 12056
rect 31941 12047 31999 12053
rect 34514 12044 34520 12056
rect 34572 12044 34578 12096
rect 36262 12044 36268 12096
rect 36320 12084 36326 12096
rect 36814 12084 36820 12096
rect 36320 12056 36820 12084
rect 36320 12044 36326 12056
rect 36814 12044 36820 12056
rect 36872 12044 36878 12096
rect 1104 11994 41400 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 41400 11994
rect 1104 11920 41400 11942
rect 3970 11840 3976 11892
rect 4028 11880 4034 11892
rect 4065 11883 4123 11889
rect 4065 11880 4077 11883
rect 4028 11852 4077 11880
rect 4028 11840 4034 11852
rect 4065 11849 4077 11852
rect 4111 11849 4123 11883
rect 4065 11843 4123 11849
rect 4798 11840 4804 11892
rect 4856 11880 4862 11892
rect 4893 11883 4951 11889
rect 4893 11880 4905 11883
rect 4856 11852 4905 11880
rect 4856 11840 4862 11852
rect 4893 11849 4905 11852
rect 4939 11849 4951 11883
rect 4893 11843 4951 11849
rect 5810 11840 5816 11892
rect 5868 11840 5874 11892
rect 6730 11840 6736 11892
rect 6788 11840 6794 11892
rect 7282 11840 7288 11892
rect 7340 11840 7346 11892
rect 8110 11840 8116 11892
rect 8168 11840 8174 11892
rect 9122 11840 9128 11892
rect 9180 11840 9186 11892
rect 10226 11840 10232 11892
rect 10284 11880 10290 11892
rect 11330 11880 11336 11892
rect 10284 11852 11336 11880
rect 10284 11840 10290 11852
rect 11330 11840 11336 11852
rect 11388 11840 11394 11892
rect 12710 11840 12716 11892
rect 12768 11880 12774 11892
rect 14553 11883 14611 11889
rect 14553 11880 14565 11883
rect 12768 11852 14565 11880
rect 12768 11840 12774 11852
rect 14553 11849 14565 11852
rect 14599 11849 14611 11883
rect 14553 11843 14611 11849
rect 18598 11840 18604 11892
rect 18656 11880 18662 11892
rect 18656 11852 18736 11880
rect 18656 11840 18662 11852
rect 6748 11812 6776 11840
rect 3068 11784 4752 11812
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 3068 11753 3096 11784
rect 4724 11753 4752 11784
rect 6104 11784 6776 11812
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 992 11716 1409 11744
rect 992 11704 998 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 3053 11747 3111 11753
rect 3053 11713 3065 11747
rect 3099 11713 3111 11747
rect 3053 11707 3111 11713
rect 3697 11747 3755 11753
rect 3697 11713 3709 11747
rect 3743 11744 3755 11747
rect 4341 11747 4399 11753
rect 4341 11744 4353 11747
rect 3743 11716 4353 11744
rect 3743 11713 3755 11716
rect 3697 11707 3755 11713
rect 4341 11713 4353 11716
rect 4387 11713 4399 11747
rect 4341 11707 4399 11713
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11744 4767 11747
rect 5626 11744 5632 11756
rect 4755 11716 5632 11744
rect 4755 11713 4767 11716
rect 4709 11707 4767 11713
rect 1670 11636 1676 11688
rect 1728 11636 1734 11688
rect 3145 11679 3203 11685
rect 3145 11645 3157 11679
rect 3191 11676 3203 11679
rect 3605 11679 3663 11685
rect 3605 11676 3617 11679
rect 3191 11648 3372 11676
rect 3191 11645 3203 11648
rect 3145 11639 3203 11645
rect 3344 11540 3372 11648
rect 3436 11648 3617 11676
rect 3436 11617 3464 11648
rect 3605 11645 3617 11648
rect 3651 11645 3663 11679
rect 3605 11639 3663 11645
rect 3421 11611 3479 11617
rect 3421 11577 3433 11611
rect 3467 11577 3479 11611
rect 4356 11608 4384 11707
rect 5626 11704 5632 11716
rect 5684 11704 5690 11756
rect 5721 11747 5779 11753
rect 5721 11713 5733 11747
rect 5767 11713 5779 11747
rect 5721 11707 5779 11713
rect 5905 11747 5963 11753
rect 5905 11713 5917 11747
rect 5951 11742 5963 11747
rect 6104 11744 6132 11784
rect 6012 11742 6132 11744
rect 5951 11716 6132 11742
rect 5951 11714 6040 11716
rect 5951 11713 5963 11714
rect 5905 11707 5963 11713
rect 4430 11636 4436 11688
rect 4488 11676 4494 11688
rect 4798 11676 4804 11688
rect 4488 11648 4804 11676
rect 4488 11636 4494 11648
rect 4798 11636 4804 11648
rect 4856 11676 4862 11688
rect 5736 11676 5764 11707
rect 6178 11704 6184 11756
rect 6236 11744 6242 11756
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 6236 11716 6561 11744
rect 6236 11704 6242 11716
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 6733 11747 6791 11753
rect 6733 11713 6745 11747
rect 6779 11744 6791 11747
rect 7300 11744 7328 11840
rect 8294 11812 8300 11824
rect 8128 11784 8300 11812
rect 6779 11716 7328 11744
rect 8021 11747 8079 11753
rect 6779 11713 6791 11716
rect 6733 11707 6791 11713
rect 8021 11713 8033 11747
rect 8067 11742 8079 11747
rect 8128 11742 8156 11784
rect 8294 11772 8300 11784
rect 8352 11812 8358 11824
rect 9140 11812 9168 11840
rect 12526 11812 12532 11824
rect 8352 11784 9168 11812
rect 9232 11784 12532 11812
rect 8352 11772 8358 11784
rect 8067 11714 8156 11742
rect 8067 11713 8079 11714
rect 8021 11707 8079 11713
rect 6748 11676 6776 11707
rect 8202 11704 8208 11756
rect 8260 11704 8266 11756
rect 4856 11648 5488 11676
rect 5736 11648 6776 11676
rect 4856 11636 4862 11648
rect 5350 11608 5356 11620
rect 4356 11580 5356 11608
rect 3421 11571 3479 11577
rect 5350 11568 5356 11580
rect 5408 11568 5414 11620
rect 4709 11543 4767 11549
rect 4709 11540 4721 11543
rect 3344 11512 4721 11540
rect 4709 11509 4721 11512
rect 4755 11540 4767 11543
rect 5258 11540 5264 11552
rect 4755 11512 5264 11540
rect 4755 11509 4767 11512
rect 4709 11503 4767 11509
rect 5258 11500 5264 11512
rect 5316 11500 5322 11552
rect 5460 11540 5488 11648
rect 6822 11636 6828 11688
rect 6880 11636 6886 11688
rect 7558 11636 7564 11688
rect 7616 11676 7622 11688
rect 9232 11676 9260 11784
rect 12526 11772 12532 11784
rect 12584 11772 12590 11824
rect 14090 11772 14096 11824
rect 14148 11772 14154 11824
rect 14185 11815 14243 11821
rect 14185 11781 14197 11815
rect 14231 11812 14243 11815
rect 14734 11812 14740 11824
rect 14231 11784 14740 11812
rect 14231 11781 14243 11784
rect 14185 11775 14243 11781
rect 14734 11772 14740 11784
rect 14792 11772 14798 11824
rect 18708 11821 18736 11852
rect 20898 11840 20904 11892
rect 20956 11840 20962 11892
rect 23658 11840 23664 11892
rect 23716 11880 23722 11892
rect 23753 11883 23811 11889
rect 23753 11880 23765 11883
rect 23716 11852 23765 11880
rect 23716 11840 23722 11852
rect 23753 11849 23765 11852
rect 23799 11849 23811 11883
rect 25774 11880 25780 11892
rect 23753 11843 23811 11849
rect 24136 11852 25780 11880
rect 18693 11815 18751 11821
rect 18693 11781 18705 11815
rect 18739 11781 18751 11815
rect 18693 11775 18751 11781
rect 19334 11772 19340 11824
rect 19392 11772 19398 11824
rect 20162 11772 20168 11824
rect 20220 11812 20226 11824
rect 20441 11815 20499 11821
rect 20441 11812 20453 11815
rect 20220 11784 20453 11812
rect 20220 11772 20226 11784
rect 20441 11781 20453 11784
rect 20487 11781 20499 11815
rect 20441 11775 20499 11781
rect 10870 11704 10876 11756
rect 10928 11704 10934 11756
rect 11054 11704 11060 11756
rect 11112 11704 11118 11756
rect 13357 11747 13415 11753
rect 13357 11713 13369 11747
rect 13403 11744 13415 11747
rect 13814 11744 13820 11756
rect 13403 11716 13820 11744
rect 13403 11713 13415 11716
rect 13357 11707 13415 11713
rect 13814 11704 13820 11716
rect 13872 11704 13878 11756
rect 14001 11747 14059 11753
rect 14001 11713 14013 11747
rect 14047 11744 14059 11747
rect 14108 11744 14136 11772
rect 14047 11716 14136 11744
rect 14277 11747 14335 11753
rect 14047 11713 14059 11716
rect 14001 11707 14059 11713
rect 14277 11713 14289 11747
rect 14323 11713 14335 11747
rect 14277 11707 14335 11713
rect 14369 11747 14427 11753
rect 14369 11713 14381 11747
rect 14415 11744 14427 11747
rect 15102 11744 15108 11756
rect 14415 11716 15108 11744
rect 14415 11713 14427 11716
rect 14369 11707 14427 11713
rect 7616 11648 9260 11676
rect 13909 11679 13967 11685
rect 7616 11636 7622 11648
rect 13909 11645 13921 11679
rect 13955 11676 13967 11679
rect 14292 11676 14320 11707
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 16574 11704 16580 11756
rect 16632 11744 16638 11756
rect 17402 11744 17408 11756
rect 16632 11716 17408 11744
rect 16632 11704 16638 11716
rect 17402 11704 17408 11716
rect 17460 11744 17466 11756
rect 20916 11753 20944 11840
rect 24136 11821 24164 11852
rect 25774 11840 25780 11852
rect 25832 11880 25838 11892
rect 26697 11883 26755 11889
rect 25832 11852 26464 11880
rect 25832 11840 25838 11852
rect 24121 11815 24179 11821
rect 23768 11784 24072 11812
rect 23768 11756 23796 11784
rect 18417 11747 18475 11753
rect 18417 11744 18429 11747
rect 17460 11716 18429 11744
rect 17460 11704 17466 11716
rect 18417 11713 18429 11716
rect 18463 11713 18475 11747
rect 18417 11707 18475 11713
rect 20901 11747 20959 11753
rect 20901 11713 20913 11747
rect 20947 11713 20959 11747
rect 20901 11707 20959 11713
rect 23661 11747 23719 11753
rect 23661 11713 23673 11747
rect 23707 11744 23719 11747
rect 23750 11744 23756 11756
rect 23707 11716 23756 11744
rect 23707 11713 23719 11716
rect 23661 11707 23719 11713
rect 23750 11704 23756 11716
rect 23808 11704 23814 11756
rect 23845 11747 23903 11753
rect 23845 11713 23857 11747
rect 23891 11713 23903 11747
rect 23845 11707 23903 11713
rect 23937 11747 23995 11753
rect 23937 11713 23949 11747
rect 23983 11713 23995 11747
rect 24044 11744 24072 11784
rect 24121 11781 24133 11815
rect 24167 11781 24179 11815
rect 24121 11775 24179 11781
rect 25590 11772 25596 11824
rect 25648 11812 25654 11824
rect 25961 11815 26019 11821
rect 25648 11784 25912 11812
rect 25648 11772 25654 11784
rect 24213 11747 24271 11753
rect 24213 11744 24225 11747
rect 24044 11716 24225 11744
rect 23937 11707 23995 11713
rect 24213 11713 24225 11716
rect 24259 11713 24271 11747
rect 24213 11707 24271 11713
rect 13955 11648 14320 11676
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 14826 11636 14832 11688
rect 14884 11676 14890 11688
rect 14884 11648 22094 11676
rect 14884 11636 14890 11648
rect 5534 11568 5540 11620
rect 5592 11608 5598 11620
rect 13722 11608 13728 11620
rect 5592 11580 13728 11608
rect 5592 11568 5598 11580
rect 13722 11568 13728 11580
rect 13780 11568 13786 11620
rect 15562 11568 15568 11620
rect 15620 11608 15626 11620
rect 16298 11608 16304 11620
rect 15620 11580 16304 11608
rect 15620 11568 15626 11580
rect 16298 11568 16304 11580
rect 16356 11568 16362 11620
rect 16850 11568 16856 11620
rect 16908 11608 16914 11620
rect 18322 11608 18328 11620
rect 16908 11580 18328 11608
rect 16908 11568 16914 11580
rect 18322 11568 18328 11580
rect 18380 11568 18386 11620
rect 21818 11608 21824 11620
rect 19720 11580 21824 11608
rect 6365 11543 6423 11549
rect 6365 11540 6377 11543
rect 5460 11512 6377 11540
rect 6365 11509 6377 11512
rect 6411 11540 6423 11543
rect 10226 11540 10232 11552
rect 6411 11512 10232 11540
rect 6411 11509 6423 11512
rect 6365 11503 6423 11509
rect 10226 11500 10232 11512
rect 10284 11500 10290 11552
rect 10318 11500 10324 11552
rect 10376 11540 10382 11552
rect 11241 11543 11299 11549
rect 11241 11540 11253 11543
rect 10376 11512 11253 11540
rect 10376 11500 10382 11512
rect 11241 11509 11253 11512
rect 11287 11509 11299 11543
rect 11241 11503 11299 11509
rect 16390 11500 16396 11552
rect 16448 11540 16454 11552
rect 17494 11540 17500 11552
rect 16448 11512 17500 11540
rect 16448 11500 16454 11512
rect 17494 11500 17500 11512
rect 17552 11540 17558 11552
rect 19720 11540 19748 11580
rect 21818 11568 21824 11580
rect 21876 11568 21882 11620
rect 17552 11512 19748 11540
rect 17552 11500 17558 11512
rect 20254 11500 20260 11552
rect 20312 11540 20318 11552
rect 20717 11543 20775 11549
rect 20717 11540 20729 11543
rect 20312 11512 20729 11540
rect 20312 11500 20318 11512
rect 20717 11509 20729 11512
rect 20763 11509 20775 11543
rect 22066 11540 22094 11648
rect 23474 11636 23480 11688
rect 23532 11676 23538 11688
rect 23860 11676 23888 11707
rect 23532 11648 23888 11676
rect 23952 11676 23980 11707
rect 24946 11704 24952 11756
rect 25004 11704 25010 11756
rect 25777 11747 25835 11753
rect 25777 11713 25789 11747
rect 25823 11713 25835 11747
rect 25884 11744 25912 11784
rect 25961 11781 25973 11815
rect 26007 11812 26019 11815
rect 26007 11784 26372 11812
rect 26007 11781 26019 11784
rect 25961 11775 26019 11781
rect 26145 11747 26203 11753
rect 26145 11744 26157 11747
rect 25884 11716 26157 11744
rect 25777 11707 25835 11713
rect 26145 11713 26157 11716
rect 26191 11713 26203 11747
rect 26145 11707 26203 11713
rect 26237 11747 26295 11753
rect 26237 11713 26249 11747
rect 26283 11713 26295 11747
rect 26237 11707 26295 11713
rect 24964 11676 24992 11704
rect 23952 11648 24992 11676
rect 23532 11636 23538 11648
rect 23937 11611 23995 11617
rect 23937 11577 23949 11611
rect 23983 11608 23995 11611
rect 24026 11608 24032 11620
rect 23983 11580 24032 11608
rect 23983 11577 23995 11580
rect 23937 11571 23995 11577
rect 24026 11568 24032 11580
rect 24084 11568 24090 11620
rect 25792 11608 25820 11707
rect 25958 11636 25964 11688
rect 26016 11676 26022 11688
rect 26252 11676 26280 11707
rect 26016 11648 26280 11676
rect 26344 11676 26372 11784
rect 26436 11756 26464 11852
rect 26697 11849 26709 11883
rect 26743 11880 26755 11883
rect 26786 11880 26792 11892
rect 26743 11852 26792 11880
rect 26743 11849 26755 11852
rect 26697 11843 26755 11849
rect 26786 11840 26792 11852
rect 26844 11840 26850 11892
rect 26878 11840 26884 11892
rect 26936 11880 26942 11892
rect 27433 11883 27491 11889
rect 27433 11880 27445 11883
rect 26936 11852 27445 11880
rect 26936 11840 26942 11852
rect 27433 11849 27445 11852
rect 27479 11849 27491 11883
rect 27433 11843 27491 11849
rect 29641 11883 29699 11889
rect 29641 11849 29653 11883
rect 29687 11880 29699 11883
rect 30558 11880 30564 11892
rect 29687 11852 30564 11880
rect 29687 11849 29699 11852
rect 29641 11843 29699 11849
rect 30558 11840 30564 11852
rect 30616 11840 30622 11892
rect 30650 11840 30656 11892
rect 30708 11840 30714 11892
rect 31202 11840 31208 11892
rect 31260 11840 31266 11892
rect 31294 11840 31300 11892
rect 31352 11840 31358 11892
rect 31386 11840 31392 11892
rect 31444 11880 31450 11892
rect 32306 11880 32312 11892
rect 31444 11852 32312 11880
rect 31444 11840 31450 11852
rect 32306 11840 32312 11852
rect 32364 11840 32370 11892
rect 36265 11883 36323 11889
rect 34716 11852 35112 11880
rect 26602 11772 26608 11824
rect 26660 11812 26666 11824
rect 26973 11815 27031 11821
rect 26973 11812 26985 11815
rect 26660 11784 26985 11812
rect 26660 11772 26666 11784
rect 26973 11781 26985 11784
rect 27019 11812 27031 11815
rect 27019 11784 27384 11812
rect 27019 11781 27031 11784
rect 26973 11775 27031 11781
rect 26418 11704 26424 11756
rect 26476 11704 26482 11756
rect 26510 11676 26516 11688
rect 26344 11648 26516 11676
rect 26016 11636 26022 11648
rect 26390 11617 26418 11648
rect 26510 11636 26516 11648
rect 26568 11636 26574 11688
rect 26375 11611 26433 11617
rect 25792 11580 26004 11608
rect 25866 11540 25872 11552
rect 22066 11512 25872 11540
rect 20717 11503 20775 11509
rect 25866 11500 25872 11512
rect 25924 11500 25930 11552
rect 25976 11540 26004 11580
rect 26375 11577 26387 11611
rect 26421 11577 26433 11611
rect 26375 11571 26433 11577
rect 26513 11543 26571 11549
rect 26513 11540 26525 11543
rect 25976 11512 26525 11540
rect 26513 11509 26525 11512
rect 26559 11540 26571 11543
rect 26620 11540 26648 11772
rect 27356 11756 27384 11784
rect 29730 11772 29736 11824
rect 29788 11812 29794 11824
rect 30193 11815 30251 11821
rect 30193 11812 30205 11815
rect 29788 11784 30205 11812
rect 29788 11772 29794 11784
rect 30193 11781 30205 11784
rect 30239 11781 30251 11815
rect 30193 11775 30251 11781
rect 26694 11704 26700 11756
rect 26752 11704 26758 11756
rect 27246 11704 27252 11756
rect 27304 11704 27310 11756
rect 27338 11704 27344 11756
rect 27396 11704 27402 11756
rect 28994 11704 29000 11756
rect 29052 11744 29058 11756
rect 29362 11744 29368 11756
rect 29052 11716 29368 11744
rect 29052 11704 29058 11716
rect 29362 11704 29368 11716
rect 29420 11704 29426 11756
rect 29549 11747 29607 11753
rect 29549 11713 29561 11747
rect 29595 11713 29607 11747
rect 29549 11707 29607 11713
rect 30009 11747 30067 11753
rect 30009 11713 30021 11747
rect 30055 11744 30067 11747
rect 30098 11744 30104 11756
rect 30055 11716 30104 11744
rect 30055 11713 30067 11716
rect 30009 11707 30067 11713
rect 26786 11636 26792 11688
rect 26844 11676 26850 11688
rect 27065 11679 27123 11685
rect 27065 11676 27077 11679
rect 26844 11648 27077 11676
rect 26844 11636 26850 11648
rect 27065 11645 27077 11648
rect 27111 11645 27123 11679
rect 27065 11639 27123 11645
rect 29270 11636 29276 11688
rect 29328 11636 29334 11688
rect 29564 11676 29592 11707
rect 30098 11704 30104 11716
rect 30156 11704 30162 11756
rect 30208 11744 30236 11775
rect 30282 11772 30288 11824
rect 30340 11812 30346 11824
rect 30377 11815 30435 11821
rect 30377 11812 30389 11815
rect 30340 11784 30389 11812
rect 30340 11772 30346 11784
rect 30377 11781 30389 11784
rect 30423 11781 30435 11815
rect 30668 11812 30696 11840
rect 30668 11784 30972 11812
rect 30377 11775 30435 11781
rect 30469 11747 30527 11753
rect 30469 11744 30481 11747
rect 30208 11716 30481 11744
rect 30469 11713 30481 11716
rect 30515 11744 30527 11747
rect 30558 11744 30564 11756
rect 30515 11716 30564 11744
rect 30515 11713 30527 11716
rect 30469 11707 30527 11713
rect 30558 11704 30564 11716
rect 30616 11704 30622 11756
rect 30653 11747 30711 11753
rect 30653 11713 30665 11747
rect 30699 11713 30711 11747
rect 30653 11707 30711 11713
rect 29914 11676 29920 11688
rect 29564 11648 29920 11676
rect 29914 11636 29920 11648
rect 29972 11636 29978 11688
rect 30116 11676 30144 11704
rect 30668 11676 30696 11707
rect 30742 11704 30748 11756
rect 30800 11744 30806 11756
rect 30944 11753 30972 11784
rect 30929 11747 30987 11753
rect 30800 11716 30880 11744
rect 30800 11704 30806 11716
rect 30116 11648 30696 11676
rect 30852 11676 30880 11716
rect 30929 11713 30941 11747
rect 30975 11713 30987 11747
rect 31220 11744 31248 11840
rect 32030 11772 32036 11824
rect 32088 11812 32094 11824
rect 34716 11812 34744 11852
rect 35084 11824 35112 11852
rect 35912 11852 36216 11880
rect 32088 11784 34744 11812
rect 32088 11772 32094 11784
rect 34882 11772 34888 11824
rect 34940 11812 34946 11824
rect 34977 11815 35035 11821
rect 34977 11812 34989 11815
rect 34940 11784 34989 11812
rect 34940 11772 34946 11784
rect 34977 11781 34989 11784
rect 35023 11781 35035 11815
rect 34977 11775 35035 11781
rect 35066 11772 35072 11824
rect 35124 11772 35130 11824
rect 35250 11772 35256 11824
rect 35308 11812 35314 11824
rect 35912 11821 35940 11852
rect 35897 11815 35955 11821
rect 35897 11812 35909 11815
rect 35308 11784 35909 11812
rect 35308 11772 35314 11784
rect 35897 11781 35909 11784
rect 35943 11781 35955 11815
rect 35897 11775 35955 11781
rect 35986 11772 35992 11824
rect 36044 11772 36050 11824
rect 33870 11744 33876 11756
rect 31220 11716 33876 11744
rect 30929 11707 30987 11713
rect 33870 11704 33876 11716
rect 33928 11744 33934 11756
rect 34057 11747 34115 11753
rect 34057 11744 34069 11747
rect 33928 11716 34069 11744
rect 33928 11704 33934 11716
rect 34057 11713 34069 11716
rect 34103 11744 34115 11747
rect 34793 11747 34851 11753
rect 34793 11744 34805 11747
rect 34103 11716 34805 11744
rect 34103 11713 34115 11716
rect 34057 11707 34115 11713
rect 34793 11713 34805 11716
rect 34839 11713 34851 11747
rect 34793 11707 34851 11713
rect 35161 11747 35219 11753
rect 35161 11713 35173 11747
rect 35207 11713 35219 11747
rect 35161 11707 35219 11713
rect 35621 11747 35679 11753
rect 35621 11713 35633 11747
rect 35667 11713 35679 11747
rect 35621 11707 35679 11713
rect 31021 11679 31079 11685
rect 31021 11676 31033 11679
rect 30852 11648 31033 11676
rect 29730 11568 29736 11620
rect 29788 11608 29794 11620
rect 30116 11608 30144 11648
rect 31021 11645 31033 11648
rect 31067 11645 31079 11679
rect 31021 11639 31079 11645
rect 31570 11636 31576 11688
rect 31628 11636 31634 11688
rect 33778 11636 33784 11688
rect 33836 11676 33842 11688
rect 34146 11676 34152 11688
rect 33836 11648 34152 11676
rect 33836 11636 33842 11648
rect 34146 11636 34152 11648
rect 34204 11636 34210 11688
rect 34422 11636 34428 11688
rect 34480 11676 34486 11688
rect 35176 11676 35204 11707
rect 35636 11676 35664 11707
rect 35710 11704 35716 11756
rect 35768 11704 35774 11756
rect 36078 11704 36084 11756
rect 36136 11753 36142 11756
rect 36136 11707 36144 11753
rect 36188 11744 36216 11852
rect 36265 11849 36277 11883
rect 36311 11880 36323 11883
rect 36630 11880 36636 11892
rect 36311 11852 36636 11880
rect 36311 11849 36323 11852
rect 36265 11843 36323 11849
rect 36630 11840 36636 11852
rect 36688 11840 36694 11892
rect 36814 11840 36820 11892
rect 36872 11880 36878 11892
rect 37458 11880 37464 11892
rect 36872 11852 37464 11880
rect 36872 11840 36878 11852
rect 37458 11840 37464 11852
rect 37516 11840 37522 11892
rect 40313 11883 40371 11889
rect 38488 11852 39804 11880
rect 38488 11812 38516 11852
rect 36924 11784 38516 11812
rect 36630 11744 36636 11756
rect 36188 11716 36636 11744
rect 36136 11704 36142 11707
rect 36630 11704 36636 11716
rect 36688 11704 36694 11756
rect 36924 11676 36952 11784
rect 39390 11775 39396 11824
rect 39385 11772 39396 11775
rect 39448 11772 39454 11824
rect 39385 11769 39443 11772
rect 39385 11735 39397 11769
rect 39431 11735 39443 11769
rect 39385 11729 39443 11735
rect 39485 11747 39543 11753
rect 39485 11713 39497 11747
rect 39531 11713 39543 11747
rect 39485 11707 39543 11713
rect 34480 11648 35204 11676
rect 34480 11636 34486 11648
rect 29788 11580 30144 11608
rect 30745 11611 30803 11617
rect 29788 11568 29794 11580
rect 30745 11577 30757 11611
rect 30791 11608 30803 11611
rect 31588 11608 31616 11636
rect 30791 11580 31616 11608
rect 30791 11577 30803 11580
rect 30745 11571 30803 11577
rect 32398 11568 32404 11620
rect 32456 11608 32462 11620
rect 33134 11608 33140 11620
rect 32456 11580 33140 11608
rect 32456 11568 32462 11580
rect 33134 11568 33140 11580
rect 33192 11568 33198 11620
rect 26559 11512 26648 11540
rect 26559 11509 26571 11512
rect 26513 11503 26571 11509
rect 27154 11500 27160 11552
rect 27212 11500 27218 11552
rect 27614 11500 27620 11552
rect 27672 11540 27678 11552
rect 29362 11540 29368 11552
rect 27672 11512 29368 11540
rect 27672 11500 27678 11512
rect 29362 11500 29368 11512
rect 29420 11500 29426 11552
rect 30374 11500 30380 11552
rect 30432 11540 30438 11552
rect 30650 11540 30656 11552
rect 30432 11512 30656 11540
rect 30432 11500 30438 11512
rect 30650 11500 30656 11512
rect 30708 11540 30714 11552
rect 30929 11543 30987 11549
rect 30929 11540 30941 11543
rect 30708 11512 30941 11540
rect 30708 11500 30714 11512
rect 30929 11509 30941 11512
rect 30975 11509 30987 11543
rect 30929 11503 30987 11509
rect 34054 11500 34060 11552
rect 34112 11540 34118 11552
rect 34149 11543 34207 11549
rect 34149 11540 34161 11543
rect 34112 11512 34161 11540
rect 34112 11500 34118 11512
rect 34149 11509 34161 11512
rect 34195 11540 34207 11543
rect 34514 11540 34520 11552
rect 34195 11512 34520 11540
rect 34195 11509 34207 11512
rect 34149 11503 34207 11509
rect 34514 11500 34520 11512
rect 34572 11500 34578 11552
rect 35176 11540 35204 11648
rect 35360 11648 36952 11676
rect 35360 11617 35388 11648
rect 37734 11636 37740 11688
rect 37792 11676 37798 11688
rect 37792 11648 38976 11676
rect 37792 11636 37798 11648
rect 35345 11611 35403 11617
rect 35345 11577 35357 11611
rect 35391 11577 35403 11611
rect 38838 11608 38844 11620
rect 35345 11571 35403 11577
rect 36280 11580 38844 11608
rect 36280 11540 36308 11580
rect 38838 11568 38844 11580
rect 38896 11568 38902 11620
rect 38948 11608 38976 11648
rect 39114 11636 39120 11688
rect 39172 11676 39178 11688
rect 39209 11679 39267 11685
rect 39209 11676 39221 11679
rect 39172 11648 39221 11676
rect 39172 11636 39178 11648
rect 39209 11645 39221 11648
rect 39255 11645 39267 11679
rect 39209 11639 39267 11645
rect 39500 11608 39528 11707
rect 39666 11704 39672 11756
rect 39724 11704 39730 11756
rect 39776 11753 39804 11852
rect 40313 11849 40325 11883
rect 40359 11880 40371 11883
rect 41230 11880 41236 11892
rect 40359 11852 41236 11880
rect 40359 11849 40371 11852
rect 40313 11843 40371 11849
rect 41230 11840 41236 11852
rect 41288 11840 41294 11892
rect 39761 11747 39819 11753
rect 39761 11713 39773 11747
rect 39807 11713 39819 11747
rect 39761 11707 39819 11713
rect 39850 11704 39856 11756
rect 39908 11704 39914 11756
rect 40126 11704 40132 11756
rect 40184 11704 40190 11756
rect 40034 11636 40040 11688
rect 40092 11636 40098 11688
rect 38948 11580 39528 11608
rect 35176 11512 36308 11540
rect 36354 11500 36360 11552
rect 36412 11540 36418 11552
rect 39206 11540 39212 11552
rect 36412 11512 39212 11540
rect 36412 11500 36418 11512
rect 39206 11500 39212 11512
rect 39264 11540 39270 11552
rect 39853 11543 39911 11549
rect 39853 11540 39865 11543
rect 39264 11512 39865 11540
rect 39264 11500 39270 11512
rect 39853 11509 39865 11512
rect 39899 11509 39911 11543
rect 39853 11503 39911 11509
rect 1104 11450 41400 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 41400 11450
rect 1104 11376 41400 11398
rect 1670 11296 1676 11348
rect 1728 11336 1734 11348
rect 1728 11308 2774 11336
rect 1728 11296 1734 11308
rect 2746 11268 2774 11308
rect 4982 11296 4988 11348
rect 5040 11336 5046 11348
rect 6178 11336 6184 11348
rect 5040 11308 6184 11336
rect 5040 11296 5046 11308
rect 6178 11296 6184 11308
rect 6236 11296 6242 11348
rect 6362 11296 6368 11348
rect 6420 11296 6426 11348
rect 7561 11339 7619 11345
rect 7561 11305 7573 11339
rect 7607 11336 7619 11339
rect 7650 11336 7656 11348
rect 7607 11308 7656 11336
rect 7607 11305 7619 11308
rect 7561 11299 7619 11305
rect 7650 11296 7656 11308
rect 7708 11296 7714 11348
rect 8110 11296 8116 11348
rect 8168 11296 8174 11348
rect 8205 11339 8263 11345
rect 8205 11305 8217 11339
rect 8251 11336 8263 11339
rect 8294 11336 8300 11348
rect 8251 11308 8300 11336
rect 8251 11305 8263 11308
rect 8205 11299 8263 11305
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 12250 11296 12256 11348
rect 12308 11336 12314 11348
rect 12308 11308 13308 11336
rect 12308 11296 12314 11308
rect 7926 11268 7932 11280
rect 2746 11240 7932 11268
rect 7926 11228 7932 11240
rect 7984 11228 7990 11280
rect 5905 11203 5963 11209
rect 5905 11169 5917 11203
rect 5951 11200 5963 11203
rect 7837 11203 7895 11209
rect 7837 11200 7849 11203
rect 5951 11172 6500 11200
rect 5951 11169 5963 11172
rect 5905 11163 5963 11169
rect 6472 11144 6500 11172
rect 7576 11172 7849 11200
rect 5997 11135 6055 11141
rect 5997 11101 6009 11135
rect 6043 11132 6055 11135
rect 6273 11135 6331 11141
rect 6273 11132 6285 11135
rect 6043 11104 6285 11132
rect 6043 11101 6055 11104
rect 5997 11095 6055 11101
rect 6273 11101 6285 11104
rect 6319 11101 6331 11135
rect 6273 11095 6331 11101
rect 5537 11067 5595 11073
rect 5537 11064 5549 11067
rect 5276 11036 5549 11064
rect 5276 11008 5304 11036
rect 5537 11033 5549 11036
rect 5583 11033 5595 11067
rect 6288 11064 6316 11095
rect 6454 11092 6460 11144
rect 6512 11092 6518 11144
rect 6288 11036 7144 11064
rect 5537 11027 5595 11033
rect 7116 11008 7144 11036
rect 5258 10956 5264 11008
rect 5316 10956 5322 11008
rect 7098 10956 7104 11008
rect 7156 10956 7162 11008
rect 7190 10956 7196 11008
rect 7248 10996 7254 11008
rect 7576 10996 7604 11172
rect 7837 11169 7849 11172
rect 7883 11169 7895 11203
rect 7837 11163 7895 11169
rect 8021 11203 8079 11209
rect 8021 11169 8033 11203
rect 8067 11200 8079 11203
rect 8128 11200 8156 11296
rect 12894 11268 12900 11280
rect 11716 11240 12900 11268
rect 8067 11172 8156 11200
rect 9585 11203 9643 11209
rect 8067 11169 8079 11172
rect 8021 11163 8079 11169
rect 9585 11169 9597 11203
rect 9631 11200 9643 11203
rect 10134 11200 10140 11212
rect 9631 11172 10140 11200
rect 9631 11169 9643 11172
rect 9585 11163 9643 11169
rect 10134 11160 10140 11172
rect 10192 11160 10198 11212
rect 10686 11160 10692 11212
rect 10744 11200 10750 11212
rect 10962 11200 10968 11212
rect 10744 11172 10968 11200
rect 10744 11160 10750 11172
rect 10962 11160 10968 11172
rect 11020 11160 11026 11212
rect 11716 11209 11744 11240
rect 12894 11228 12900 11240
rect 12952 11228 12958 11280
rect 11701 11203 11759 11209
rect 11701 11169 11713 11203
rect 11747 11169 11759 11203
rect 11701 11163 11759 11169
rect 11885 11203 11943 11209
rect 11885 11169 11897 11203
rect 11931 11200 11943 11203
rect 12158 11200 12164 11212
rect 11931 11172 12164 11200
rect 11931 11169 11943 11172
rect 11885 11163 11943 11169
rect 7745 11135 7803 11141
rect 7745 11101 7757 11135
rect 7791 11101 7803 11135
rect 7745 11095 7803 11101
rect 7650 11024 7656 11076
rect 7708 11064 7714 11076
rect 7760 11064 7788 11095
rect 7926 11092 7932 11144
rect 7984 11132 7990 11144
rect 8389 11135 8447 11141
rect 8389 11132 8401 11135
rect 7984 11104 8401 11132
rect 7984 11092 7990 11104
rect 8389 11101 8401 11104
rect 8435 11132 8447 11135
rect 8570 11132 8576 11144
rect 8435 11104 8576 11132
rect 8435 11101 8447 11104
rect 8389 11095 8447 11101
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 8665 11135 8723 11141
rect 8665 11101 8677 11135
rect 8711 11101 8723 11135
rect 8665 11095 8723 11101
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11101 9551 11135
rect 9493 11095 9551 11101
rect 9769 11135 9827 11141
rect 9769 11101 9781 11135
rect 9815 11132 9827 11135
rect 9950 11132 9956 11144
rect 9815 11104 9956 11132
rect 9815 11101 9827 11104
rect 9769 11095 9827 11101
rect 8680 11064 8708 11095
rect 9508 11064 9536 11095
rect 9950 11092 9956 11104
rect 10008 11092 10014 11144
rect 10318 11092 10324 11144
rect 10376 11092 10382 11144
rect 10873 11135 10931 11141
rect 10873 11101 10885 11135
rect 10919 11132 10931 11135
rect 11716 11132 11744 11163
rect 12158 11160 12164 11172
rect 12216 11160 12222 11212
rect 12250 11160 12256 11212
rect 12308 11160 12314 11212
rect 13280 11200 13308 11308
rect 14550 11296 14556 11348
rect 14608 11336 14614 11348
rect 15841 11339 15899 11345
rect 14608 11308 15700 11336
rect 14608 11296 14614 11308
rect 15473 11203 15531 11209
rect 15473 11200 15485 11203
rect 13096 11172 15485 11200
rect 10919 11104 11744 11132
rect 10919 11101 10931 11104
rect 10873 11095 10931 11101
rect 12434 11092 12440 11144
rect 12492 11092 12498 11144
rect 12526 11092 12532 11144
rect 12584 11132 12590 11144
rect 13096 11141 13124 11172
rect 15473 11169 15485 11172
rect 15519 11200 15531 11203
rect 15562 11200 15568 11212
rect 15519 11172 15568 11200
rect 15519 11169 15531 11172
rect 15473 11163 15531 11169
rect 15562 11160 15568 11172
rect 15620 11160 15626 11212
rect 15672 11141 15700 11308
rect 15841 11305 15853 11339
rect 15887 11336 15899 11339
rect 15930 11336 15936 11348
rect 15887 11308 15936 11336
rect 15887 11305 15899 11308
rect 15841 11299 15899 11305
rect 15930 11296 15936 11308
rect 15988 11296 15994 11348
rect 16114 11296 16120 11348
rect 16172 11296 16178 11348
rect 21358 11296 21364 11348
rect 21416 11296 21422 11348
rect 26050 11296 26056 11348
rect 26108 11336 26114 11348
rect 26697 11339 26755 11345
rect 26697 11336 26709 11339
rect 26108 11308 26709 11336
rect 26108 11296 26114 11308
rect 26697 11305 26709 11308
rect 26743 11336 26755 11339
rect 26786 11336 26792 11348
rect 26743 11308 26792 11336
rect 26743 11305 26755 11308
rect 26697 11299 26755 11305
rect 26786 11296 26792 11308
rect 26844 11296 26850 11348
rect 27522 11296 27528 11348
rect 27580 11336 27586 11348
rect 27580 11308 30972 11336
rect 27580 11296 27586 11308
rect 16132 11200 16160 11296
rect 22094 11228 22100 11280
rect 22152 11268 22158 11280
rect 22373 11271 22431 11277
rect 22373 11268 22385 11271
rect 22152 11240 22385 11268
rect 22152 11228 22158 11240
rect 22373 11237 22385 11240
rect 22419 11237 22431 11271
rect 28994 11268 29000 11280
rect 22373 11231 22431 11237
rect 25204 11240 29000 11268
rect 16132 11172 16528 11200
rect 12897 11135 12955 11141
rect 12897 11132 12909 11135
rect 12584 11104 12909 11132
rect 12584 11092 12590 11104
rect 12897 11101 12909 11104
rect 12943 11101 12955 11135
rect 12897 11095 12955 11101
rect 13081 11135 13139 11141
rect 13081 11101 13093 11135
rect 13127 11101 13139 11135
rect 15657 11135 15715 11141
rect 13081 11095 13139 11101
rect 13188 11104 14872 11132
rect 10336 11064 10364 11092
rect 7708 11036 8708 11064
rect 8772 11036 9444 11064
rect 9508 11036 10364 11064
rect 10781 11067 10839 11073
rect 7708 11024 7714 11036
rect 8110 10996 8116 11008
rect 7248 10968 8116 10996
rect 7248 10956 7254 10968
rect 8110 10956 8116 10968
rect 8168 10996 8174 11008
rect 8573 10999 8631 11005
rect 8573 10996 8585 10999
rect 8168 10968 8585 10996
rect 8168 10956 8174 10968
rect 8573 10965 8585 10968
rect 8619 10996 8631 10999
rect 8772 10996 8800 11036
rect 8619 10968 8800 10996
rect 9416 10996 9444 11036
rect 10781 11033 10793 11067
rect 10827 11064 10839 11067
rect 11606 11064 11612 11076
rect 10827 11036 11612 11064
rect 10827 11033 10839 11036
rect 10781 11027 10839 11033
rect 11606 11024 11612 11036
rect 11664 11024 11670 11076
rect 11882 11024 11888 11076
rect 11940 11064 11946 11076
rect 13188 11064 13216 11104
rect 11940 11036 13216 11064
rect 13265 11067 13323 11073
rect 11940 11024 11946 11036
rect 13265 11033 13277 11067
rect 13311 11033 13323 11067
rect 14844 11064 14872 11104
rect 15657 11101 15669 11135
rect 15703 11132 15715 11135
rect 16209 11135 16267 11141
rect 16209 11132 16221 11135
rect 15703 11104 16221 11132
rect 15703 11101 15715 11104
rect 15657 11095 15715 11101
rect 16209 11101 16221 11104
rect 16255 11101 16267 11135
rect 16209 11095 16267 11101
rect 16298 11092 16304 11144
rect 16356 11132 16362 11144
rect 16500 11141 16528 11172
rect 17402 11160 17408 11212
rect 17460 11160 17466 11212
rect 17494 11160 17500 11212
rect 17552 11160 17558 11212
rect 17681 11203 17739 11209
rect 17681 11169 17693 11203
rect 17727 11200 17739 11203
rect 17770 11200 17776 11212
rect 17727 11172 17776 11200
rect 17727 11169 17739 11172
rect 17681 11163 17739 11169
rect 17770 11160 17776 11172
rect 17828 11200 17834 11212
rect 18598 11200 18604 11212
rect 17828 11172 18604 11200
rect 17828 11160 17834 11172
rect 18598 11160 18604 11172
rect 18656 11160 18662 11212
rect 19889 11203 19947 11209
rect 19889 11169 19901 11203
rect 19935 11200 19947 11203
rect 20254 11200 20260 11212
rect 19935 11172 20260 11200
rect 19935 11169 19947 11172
rect 19889 11163 19947 11169
rect 20254 11160 20260 11172
rect 20312 11160 20318 11212
rect 21913 11203 21971 11209
rect 21913 11169 21925 11203
rect 21959 11200 21971 11203
rect 25204 11200 25232 11240
rect 28994 11228 29000 11240
rect 29052 11228 29058 11280
rect 30834 11228 30840 11280
rect 30892 11228 30898 11280
rect 30944 11268 30972 11308
rect 31018 11296 31024 11348
rect 31076 11296 31082 11348
rect 36078 11336 36084 11348
rect 31128 11308 36084 11336
rect 31128 11268 31156 11308
rect 36078 11296 36084 11308
rect 36136 11296 36142 11348
rect 36170 11296 36176 11348
rect 36228 11336 36234 11348
rect 38473 11339 38531 11345
rect 38473 11336 38485 11339
rect 36228 11308 38485 11336
rect 36228 11296 36234 11308
rect 38473 11305 38485 11308
rect 38519 11336 38531 11339
rect 38654 11336 38660 11348
rect 38519 11308 38660 11336
rect 38519 11305 38531 11308
rect 38473 11299 38531 11305
rect 38654 11296 38660 11308
rect 38712 11336 38718 11348
rect 39114 11336 39120 11348
rect 38712 11308 39120 11336
rect 38712 11296 38718 11308
rect 39114 11296 39120 11308
rect 39172 11296 39178 11348
rect 39298 11296 39304 11348
rect 39356 11296 39362 11348
rect 30944 11240 31156 11268
rect 32125 11271 32183 11277
rect 32125 11237 32137 11271
rect 32171 11268 32183 11271
rect 33502 11268 33508 11280
rect 32171 11240 33508 11268
rect 32171 11237 32183 11240
rect 32125 11231 32183 11237
rect 33502 11228 33508 11240
rect 33560 11228 33566 11280
rect 33781 11271 33839 11277
rect 33781 11268 33793 11271
rect 33612 11240 33793 11268
rect 21959 11172 25232 11200
rect 21959 11169 21971 11172
rect 21913 11163 21971 11169
rect 25866 11160 25872 11212
rect 25924 11200 25930 11212
rect 25924 11172 29224 11200
rect 25924 11160 25930 11172
rect 16393 11135 16451 11141
rect 16393 11132 16405 11135
rect 16356 11104 16405 11132
rect 16356 11092 16362 11104
rect 16393 11101 16405 11104
rect 16439 11101 16451 11135
rect 16393 11095 16451 11101
rect 16485 11135 16543 11141
rect 16485 11101 16497 11135
rect 16531 11101 16543 11135
rect 17420 11132 17448 11160
rect 19613 11135 19671 11141
rect 19613 11132 19625 11135
rect 17420 11104 19625 11132
rect 16485 11095 16543 11101
rect 19613 11101 19625 11104
rect 19659 11101 19671 11135
rect 19613 11095 19671 11101
rect 22005 11135 22063 11141
rect 22005 11101 22017 11135
rect 22051 11132 22063 11135
rect 22370 11132 22376 11144
rect 22051 11104 22376 11132
rect 22051 11101 22063 11104
rect 22005 11095 22063 11101
rect 22370 11092 22376 11104
rect 22428 11092 22434 11144
rect 22646 11092 22652 11144
rect 22704 11092 22710 11144
rect 23106 11092 23112 11144
rect 23164 11092 23170 11144
rect 29089 11135 29147 11141
rect 29089 11132 29101 11135
rect 23216 11104 29101 11132
rect 16577 11067 16635 11073
rect 16577 11064 16589 11067
rect 14844 11036 16589 11064
rect 13265 11027 13323 11033
rect 16577 11033 16589 11036
rect 16623 11064 16635 11067
rect 17126 11064 17132 11076
rect 16623 11036 17132 11064
rect 16623 11033 16635 11036
rect 16577 11027 16635 11033
rect 9858 10996 9864 11008
rect 9416 10968 9864 10996
rect 8619 10965 8631 10968
rect 8573 10959 8631 10965
rect 9858 10956 9864 10968
rect 9916 10996 9922 11008
rect 9953 10999 10011 11005
rect 9953 10996 9965 10999
rect 9916 10968 9965 10996
rect 9916 10956 9922 10968
rect 9953 10965 9965 10968
rect 9999 10965 10011 10999
rect 9953 10959 10011 10965
rect 10410 10956 10416 11008
rect 10468 10956 10474 11008
rect 11238 10956 11244 11008
rect 11296 10956 11302 11008
rect 12618 10956 12624 11008
rect 12676 10956 12682 11008
rect 13280 10996 13308 11027
rect 17126 11024 17132 11036
rect 17184 11024 17190 11076
rect 22462 11064 22468 11076
rect 21114 11036 22468 11064
rect 22462 11024 22468 11036
rect 22520 11024 22526 11076
rect 13814 10996 13820 11008
rect 13280 10968 13820 10996
rect 13814 10956 13820 10968
rect 13872 10956 13878 11008
rect 16298 10956 16304 11008
rect 16356 10956 16362 11008
rect 17034 10956 17040 11008
rect 17092 10956 17098 11008
rect 17310 10956 17316 11008
rect 17368 10996 17374 11008
rect 17405 10999 17463 11005
rect 17405 10996 17417 10999
rect 17368 10968 17417 10996
rect 17368 10956 17374 10968
rect 17405 10965 17417 10968
rect 17451 10965 17463 10999
rect 17405 10959 17463 10965
rect 21450 10956 21456 11008
rect 21508 10996 21514 11008
rect 23216 10996 23244 11104
rect 29089 11101 29101 11104
rect 29135 11101 29147 11135
rect 29196 11132 29224 11172
rect 31036 11172 31892 11200
rect 31036 11132 31064 11172
rect 29196 11104 31064 11132
rect 29089 11095 29147 11101
rect 25958 11024 25964 11076
rect 26016 11064 26022 11076
rect 26605 11067 26663 11073
rect 26605 11064 26617 11067
rect 26016 11036 26617 11064
rect 26016 11024 26022 11036
rect 26605 11033 26617 11036
rect 26651 11033 26663 11067
rect 26605 11027 26663 11033
rect 26694 11024 26700 11076
rect 26752 11064 26758 11076
rect 27154 11064 27160 11076
rect 26752 11036 27160 11064
rect 26752 11024 26758 11036
rect 27154 11024 27160 11036
rect 27212 11024 27218 11076
rect 29104 11064 29132 11095
rect 31478 11092 31484 11144
rect 31536 11132 31542 11144
rect 31864 11141 31892 11172
rect 32950 11160 32956 11212
rect 33008 11160 33014 11212
rect 33612 11200 33640 11240
rect 33781 11237 33793 11240
rect 33827 11237 33839 11271
rect 33781 11231 33839 11237
rect 36354 11228 36360 11280
rect 36412 11228 36418 11280
rect 36630 11228 36636 11280
rect 36688 11228 36694 11280
rect 37642 11228 37648 11280
rect 37700 11228 37706 11280
rect 38013 11271 38071 11277
rect 38013 11237 38025 11271
rect 38059 11237 38071 11271
rect 39942 11268 39948 11280
rect 38013 11231 38071 11237
rect 39040 11240 39948 11268
rect 33870 11200 33876 11212
rect 33152 11172 33640 11200
rect 33704 11172 33876 11200
rect 31849 11135 31907 11141
rect 31536 11104 31800 11132
rect 31536 11092 31542 11104
rect 30190 11064 30196 11076
rect 29104 11036 30196 11064
rect 30190 11024 30196 11036
rect 30248 11024 30254 11076
rect 30558 11024 30564 11076
rect 30616 11064 30622 11076
rect 31573 11067 31631 11073
rect 31573 11064 31585 11067
rect 30616 11036 31585 11064
rect 30616 11024 30622 11036
rect 31573 11033 31585 11036
rect 31619 11064 31631 11067
rect 31662 11064 31668 11076
rect 31619 11036 31668 11064
rect 31619 11033 31631 11036
rect 31573 11027 31631 11033
rect 31662 11024 31668 11036
rect 31720 11024 31726 11076
rect 31772 11064 31800 11104
rect 31849 11101 31861 11135
rect 31895 11132 31907 11135
rect 32030 11132 32036 11144
rect 31895 11104 32036 11132
rect 31895 11101 31907 11104
rect 31849 11095 31907 11101
rect 32030 11092 32036 11104
rect 32088 11092 32094 11144
rect 33152 11141 33180 11172
rect 33137 11135 33195 11141
rect 33137 11101 33149 11135
rect 33183 11101 33195 11135
rect 33137 11095 33195 11101
rect 33594 11092 33600 11144
rect 33652 11092 33658 11144
rect 33704 11143 33732 11172
rect 33870 11160 33876 11172
rect 33928 11160 33934 11212
rect 35434 11160 35440 11212
rect 35492 11200 35498 11212
rect 35492 11172 36216 11200
rect 35492 11160 35498 11172
rect 36188 11144 36216 11172
rect 33689 11137 33747 11143
rect 33689 11103 33701 11137
rect 33735 11103 33747 11137
rect 34054 11132 34060 11144
rect 33689 11097 33747 11103
rect 33796 11104 34060 11132
rect 31941 11067 31999 11073
rect 31941 11064 31953 11067
rect 31772 11036 31953 11064
rect 31941 11033 31953 11036
rect 31987 11033 31999 11067
rect 31941 11027 31999 11033
rect 33229 11067 33287 11073
rect 33229 11033 33241 11067
rect 33275 11033 33287 11067
rect 33229 11027 33287 11033
rect 21508 10968 23244 10996
rect 21508 10956 21514 10968
rect 25130 10956 25136 11008
rect 25188 10996 25194 11008
rect 29178 10996 29184 11008
rect 25188 10968 29184 10996
rect 25188 10956 25194 10968
rect 29178 10956 29184 10968
rect 29236 10956 29242 11008
rect 29273 10999 29331 11005
rect 29273 10965 29285 10999
rect 29319 10996 29331 10999
rect 29546 10996 29552 11008
rect 29319 10968 29552 10996
rect 29319 10965 29331 10968
rect 29273 10959 29331 10965
rect 29546 10956 29552 10968
rect 29604 10956 29610 11008
rect 31202 10956 31208 11008
rect 31260 10996 31266 11008
rect 31757 10999 31815 11005
rect 31757 10996 31769 10999
rect 31260 10968 31769 10996
rect 31260 10956 31266 10968
rect 31757 10965 31769 10968
rect 31803 10965 31815 10999
rect 31956 10996 31984 11027
rect 32950 10996 32956 11008
rect 31956 10968 32956 10996
rect 31757 10959 31815 10965
rect 32950 10956 32956 10968
rect 33008 10956 33014 11008
rect 33134 10956 33140 11008
rect 33192 10996 33198 11008
rect 33244 10996 33272 11027
rect 33318 11024 33324 11076
rect 33376 11024 33382 11076
rect 33439 11067 33497 11073
rect 33439 11033 33451 11067
rect 33485 11064 33497 11067
rect 33796 11064 33824 11104
rect 34054 11092 34060 11104
rect 34112 11092 34118 11144
rect 35158 11092 35164 11144
rect 35216 11132 35222 11144
rect 35805 11135 35863 11141
rect 35805 11132 35817 11135
rect 35216 11104 35817 11132
rect 35216 11092 35222 11104
rect 35805 11101 35817 11104
rect 35851 11101 35863 11135
rect 35805 11095 35863 11101
rect 36078 11092 36084 11144
rect 36136 11092 36142 11144
rect 36170 11092 36176 11144
rect 36228 11092 36234 11144
rect 36354 11092 36360 11144
rect 36412 11132 36418 11144
rect 36648 11141 36676 11228
rect 37660 11200 37688 11228
rect 36832 11172 37596 11200
rect 37660 11172 37872 11200
rect 36832 11144 36860 11172
rect 37568 11144 37596 11172
rect 36449 11135 36507 11141
rect 36449 11132 36461 11135
rect 36412 11104 36461 11132
rect 36412 11092 36418 11104
rect 36449 11101 36461 11104
rect 36495 11101 36507 11135
rect 36449 11095 36507 11101
rect 36633 11135 36691 11141
rect 36633 11101 36645 11135
rect 36679 11101 36691 11135
rect 36633 11095 36691 11101
rect 36814 11092 36820 11144
rect 36872 11092 36878 11144
rect 37461 11135 37519 11141
rect 37461 11101 37473 11135
rect 37507 11101 37519 11135
rect 37461 11095 37519 11101
rect 35986 11064 35992 11076
rect 33485 11036 33824 11064
rect 34716 11036 35992 11064
rect 33485 11033 33497 11036
rect 33439 11027 33497 11033
rect 33192 10968 33272 10996
rect 33336 10996 33364 11024
rect 34716 10996 34744 11036
rect 35986 11024 35992 11036
rect 36044 11064 36050 11076
rect 36044 11036 36216 11064
rect 36044 11024 36050 11036
rect 33336 10968 34744 10996
rect 36188 10996 36216 11036
rect 37182 11024 37188 11076
rect 37240 11064 37246 11076
rect 37476 11064 37504 11095
rect 37550 11092 37556 11144
rect 37608 11132 37614 11144
rect 37844 11141 37872 11172
rect 37645 11135 37703 11141
rect 37645 11132 37657 11135
rect 37608 11104 37657 11132
rect 37608 11092 37614 11104
rect 37645 11101 37657 11104
rect 37691 11101 37703 11135
rect 37645 11095 37703 11101
rect 37829 11135 37887 11141
rect 37829 11101 37841 11135
rect 37875 11101 37887 11135
rect 38028 11132 38056 11231
rect 38378 11132 38384 11144
rect 38028 11104 38384 11132
rect 37829 11095 37887 11101
rect 37240 11036 37504 11064
rect 37737 11067 37795 11073
rect 37240 11024 37246 11036
rect 37737 11033 37749 11067
rect 37783 11033 37795 11067
rect 37844 11064 37872 11095
rect 38378 11092 38384 11104
rect 38436 11132 38442 11144
rect 38657 11135 38715 11141
rect 38657 11132 38669 11135
rect 38436 11104 38669 11132
rect 38436 11092 38442 11104
rect 38657 11101 38669 11104
rect 38703 11101 38715 11135
rect 38657 11095 38715 11101
rect 38746 11092 38752 11144
rect 38804 11092 38810 11144
rect 39040 11141 39068 11240
rect 39942 11228 39948 11240
rect 40000 11228 40006 11280
rect 39025 11135 39083 11141
rect 39025 11101 39037 11135
rect 39071 11101 39083 11135
rect 39025 11095 39083 11101
rect 39114 11092 39120 11144
rect 39172 11141 39178 11144
rect 39172 11132 39180 11141
rect 39172 11104 39217 11132
rect 39172 11095 39180 11104
rect 39172 11092 39178 11095
rect 38197 11067 38255 11073
rect 38197 11064 38209 11067
rect 37844 11036 38209 11064
rect 37737 11027 37795 11033
rect 38197 11033 38209 11036
rect 38243 11033 38255 11067
rect 38197 11027 38255 11033
rect 38933 11067 38991 11073
rect 38933 11033 38945 11067
rect 38979 11064 38991 11067
rect 38979 11036 39068 11064
rect 38979 11033 38991 11036
rect 38933 11027 38991 11033
rect 36630 10996 36636 11008
rect 36188 10968 36636 10996
rect 33192 10956 33198 10968
rect 36630 10956 36636 10968
rect 36688 10956 36694 11008
rect 36814 10956 36820 11008
rect 36872 10956 36878 11008
rect 37090 10956 37096 11008
rect 37148 10996 37154 11008
rect 37752 10996 37780 11027
rect 39040 11008 39068 11036
rect 37148 10968 37780 10996
rect 37148 10956 37154 10968
rect 39022 10956 39028 11008
rect 39080 10956 39086 11008
rect 1104 10906 41400 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 41400 10906
rect 1104 10832 41400 10854
rect 6454 10752 6460 10804
rect 6512 10752 6518 10804
rect 7098 10752 7104 10804
rect 7156 10752 7162 10804
rect 7926 10752 7932 10804
rect 7984 10752 7990 10804
rect 11238 10752 11244 10804
rect 11296 10792 11302 10804
rect 11885 10795 11943 10801
rect 11885 10792 11897 10795
rect 11296 10764 11897 10792
rect 11296 10752 11302 10764
rect 11885 10761 11897 10764
rect 11931 10761 11943 10795
rect 11885 10755 11943 10761
rect 11974 10752 11980 10804
rect 12032 10752 12038 10804
rect 12158 10752 12164 10804
rect 12216 10792 12222 10804
rect 16482 10792 16488 10804
rect 12216 10764 16488 10792
rect 12216 10752 12222 10764
rect 16482 10752 16488 10764
rect 16540 10792 16546 10804
rect 17954 10792 17960 10804
rect 16540 10764 17960 10792
rect 16540 10752 16546 10764
rect 17954 10752 17960 10764
rect 18012 10752 18018 10804
rect 19334 10792 19340 10804
rect 18984 10764 19340 10792
rect 7944 10724 7972 10752
rect 18984 10736 19012 10764
rect 19334 10752 19340 10764
rect 19392 10792 19398 10804
rect 20257 10795 20315 10801
rect 20257 10792 20269 10795
rect 19392 10764 20269 10792
rect 19392 10752 19398 10764
rect 20257 10761 20269 10764
rect 20303 10761 20315 10795
rect 20257 10755 20315 10761
rect 20898 10752 20904 10804
rect 20956 10792 20962 10804
rect 30101 10795 30159 10801
rect 30101 10792 30113 10795
rect 20956 10764 26924 10792
rect 20956 10752 20962 10764
rect 9677 10727 9735 10733
rect 9677 10724 9689 10727
rect 6656 10696 7972 10724
rect 8588 10696 9689 10724
rect 6656 10665 6684 10696
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10625 6699 10659
rect 6641 10619 6699 10625
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10625 6883 10659
rect 6825 10619 6883 10625
rect 6840 10588 6868 10619
rect 6914 10616 6920 10668
rect 6972 10656 6978 10668
rect 7009 10659 7067 10665
rect 7009 10656 7021 10659
rect 6972 10628 7021 10656
rect 6972 10616 6978 10628
rect 7009 10625 7021 10628
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 7190 10616 7196 10668
rect 7248 10616 7254 10668
rect 7300 10665 7328 10696
rect 7285 10659 7343 10665
rect 7285 10625 7297 10659
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 7929 10659 7987 10665
rect 7929 10625 7941 10659
rect 7975 10625 7987 10659
rect 7929 10619 7987 10625
rect 8113 10659 8171 10665
rect 8113 10625 8125 10659
rect 8159 10656 8171 10659
rect 8478 10656 8484 10668
rect 8159 10628 8484 10656
rect 8159 10625 8171 10628
rect 8113 10619 8171 10625
rect 7208 10588 7236 10616
rect 6840 10560 7236 10588
rect 7944 10520 7972 10619
rect 8478 10616 8484 10628
rect 8536 10616 8542 10668
rect 8588 10665 8616 10696
rect 9677 10693 9689 10696
rect 9723 10693 9735 10727
rect 9677 10687 9735 10693
rect 10505 10727 10563 10733
rect 10505 10693 10517 10727
rect 10551 10724 10563 10727
rect 10870 10724 10876 10736
rect 10551 10696 10876 10724
rect 10551 10693 10563 10696
rect 10505 10687 10563 10693
rect 10870 10684 10876 10696
rect 10928 10724 10934 10736
rect 16301 10727 16359 10733
rect 10928 10696 12112 10724
rect 10928 10684 10934 10696
rect 8573 10659 8631 10665
rect 8573 10625 8585 10659
rect 8619 10625 8631 10659
rect 8573 10619 8631 10625
rect 8662 10616 8668 10668
rect 8720 10656 8726 10668
rect 8757 10659 8815 10665
rect 8757 10656 8769 10659
rect 8720 10628 8769 10656
rect 8720 10616 8726 10628
rect 8757 10625 8769 10628
rect 8803 10625 8815 10659
rect 8757 10619 8815 10625
rect 8938 10616 8944 10668
rect 8996 10616 9002 10668
rect 9125 10659 9183 10665
rect 9125 10625 9137 10659
rect 9171 10625 9183 10659
rect 9125 10619 9183 10625
rect 8202 10548 8208 10600
rect 8260 10588 8266 10600
rect 8297 10591 8355 10597
rect 8297 10588 8309 10591
rect 8260 10560 8309 10588
rect 8260 10548 8266 10560
rect 8297 10557 8309 10560
rect 8343 10588 8355 10591
rect 8849 10591 8907 10597
rect 8849 10588 8861 10591
rect 8343 10560 8861 10588
rect 8343 10557 8355 10560
rect 8297 10551 8355 10557
rect 8849 10557 8861 10560
rect 8895 10557 8907 10591
rect 8849 10551 8907 10557
rect 9140 10520 9168 10619
rect 9306 10616 9312 10668
rect 9364 10616 9370 10668
rect 9398 10616 9404 10668
rect 9456 10616 9462 10668
rect 9490 10616 9496 10668
rect 9548 10616 9554 10668
rect 9950 10616 9956 10668
rect 10008 10616 10014 10668
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 10229 10659 10287 10665
rect 10229 10656 10241 10659
rect 10192 10628 10241 10656
rect 10192 10616 10198 10628
rect 10229 10625 10241 10628
rect 10275 10656 10287 10659
rect 10275 10628 11008 10656
rect 10275 10625 10287 10628
rect 10229 10619 10287 10625
rect 9217 10591 9275 10597
rect 9217 10557 9229 10591
rect 9263 10588 9275 10591
rect 9416 10588 9444 10616
rect 9263 10560 9444 10588
rect 9263 10557 9275 10560
rect 9217 10551 9275 10557
rect 10318 10548 10324 10600
rect 10376 10548 10382 10600
rect 10980 10597 11008 10628
rect 12084 10597 12112 10696
rect 16301 10693 16313 10727
rect 16347 10724 16359 10727
rect 16850 10724 16856 10736
rect 16347 10696 16856 10724
rect 16347 10693 16359 10696
rect 16301 10687 16359 10693
rect 16850 10684 16856 10696
rect 16908 10684 16914 10736
rect 17034 10684 17040 10736
rect 17092 10684 17098 10736
rect 17678 10684 17684 10736
rect 17736 10684 17742 10736
rect 18966 10724 18972 10736
rect 18906 10696 18972 10724
rect 18966 10684 18972 10696
rect 19024 10684 19030 10736
rect 19058 10684 19064 10736
rect 19116 10724 19122 10736
rect 20165 10727 20223 10733
rect 20165 10724 20177 10727
rect 19116 10696 20177 10724
rect 19116 10684 19122 10696
rect 20165 10693 20177 10696
rect 20211 10724 20223 10727
rect 20714 10724 20720 10736
rect 20211 10696 20720 10724
rect 20211 10693 20223 10696
rect 20165 10687 20223 10693
rect 20714 10684 20720 10696
rect 20772 10684 20778 10736
rect 25501 10727 25559 10733
rect 25501 10693 25513 10727
rect 25547 10724 25559 10727
rect 25547 10696 26832 10724
rect 25547 10693 25559 10696
rect 25501 10687 25559 10693
rect 12805 10659 12863 10665
rect 12805 10625 12817 10659
rect 12851 10625 12863 10659
rect 12805 10619 12863 10625
rect 10965 10591 11023 10597
rect 10965 10557 10977 10591
rect 11011 10557 11023 10591
rect 10965 10551 11023 10557
rect 12069 10591 12127 10597
rect 12069 10557 12081 10591
rect 12115 10557 12127 10591
rect 12069 10551 12127 10557
rect 9769 10523 9827 10529
rect 9769 10520 9781 10523
rect 7944 10492 9781 10520
rect 9769 10489 9781 10492
rect 9815 10489 9827 10523
rect 9769 10483 9827 10489
rect 10137 10523 10195 10529
rect 10137 10489 10149 10523
rect 10183 10520 10195 10523
rect 10336 10520 10364 10548
rect 10183 10492 10364 10520
rect 10183 10489 10195 10492
rect 10137 10483 10195 10489
rect 10410 10480 10416 10532
rect 10468 10520 10474 10532
rect 10781 10523 10839 10529
rect 10781 10520 10793 10523
rect 10468 10492 10793 10520
rect 10468 10480 10474 10492
rect 10781 10489 10793 10492
rect 10827 10489 10839 10523
rect 12084 10520 12112 10551
rect 12618 10548 12624 10600
rect 12676 10588 12682 10600
rect 12820 10588 12848 10619
rect 12986 10616 12992 10668
rect 13044 10616 13050 10668
rect 16117 10659 16175 10665
rect 16117 10625 16129 10659
rect 16163 10656 16175 10659
rect 17052 10656 17080 10684
rect 16163 10628 17080 10656
rect 16163 10625 16175 10628
rect 16117 10619 16175 10625
rect 17402 10616 17408 10668
rect 17460 10616 17466 10668
rect 18690 10616 18696 10668
rect 18748 10616 18754 10668
rect 19797 10659 19855 10665
rect 19797 10625 19809 10659
rect 19843 10656 19855 10659
rect 19978 10656 19984 10668
rect 19843 10628 19984 10656
rect 19843 10625 19855 10628
rect 19797 10619 19855 10625
rect 19978 10616 19984 10628
rect 20036 10616 20042 10668
rect 26053 10659 26111 10665
rect 26053 10625 26065 10659
rect 26099 10656 26111 10659
rect 26234 10656 26240 10668
rect 26099 10628 26240 10656
rect 26099 10625 26111 10628
rect 26053 10619 26111 10625
rect 26234 10616 26240 10628
rect 26292 10656 26298 10668
rect 26694 10656 26700 10668
rect 26292 10628 26700 10656
rect 26292 10616 26298 10628
rect 26694 10616 26700 10628
rect 26752 10616 26758 10668
rect 12676 10560 12848 10588
rect 16393 10591 16451 10597
rect 12676 10548 12682 10560
rect 16393 10557 16405 10591
rect 16439 10557 16451 10591
rect 18708 10588 18736 10616
rect 19150 10588 19156 10600
rect 18708 10560 19156 10588
rect 16393 10551 16451 10557
rect 15654 10520 15660 10532
rect 12084 10492 15660 10520
rect 10781 10483 10839 10489
rect 15654 10480 15660 10492
rect 15712 10520 15718 10532
rect 16408 10520 16436 10551
rect 19150 10548 19156 10560
rect 19208 10548 19214 10600
rect 19334 10548 19340 10600
rect 19392 10548 19398 10600
rect 19705 10591 19763 10597
rect 19705 10557 19717 10591
rect 19751 10557 19763 10591
rect 19996 10588 20024 10616
rect 20254 10588 20260 10600
rect 19996 10560 20260 10588
rect 19705 10551 19763 10557
rect 15712 10492 16436 10520
rect 19720 10520 19748 10551
rect 20254 10548 20260 10560
rect 20312 10548 20318 10600
rect 23293 10591 23351 10597
rect 23293 10557 23305 10591
rect 23339 10588 23351 10591
rect 23566 10588 23572 10600
rect 23339 10560 23572 10588
rect 23339 10557 23351 10560
rect 23293 10551 23351 10557
rect 23566 10548 23572 10560
rect 23624 10548 23630 10600
rect 21450 10520 21456 10532
rect 19720 10492 21456 10520
rect 15712 10480 15718 10492
rect 21450 10480 21456 10492
rect 21508 10480 21514 10532
rect 4798 10412 4804 10464
rect 4856 10452 4862 10464
rect 5350 10452 5356 10464
rect 4856 10424 5356 10452
rect 4856 10412 4862 10424
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 8386 10412 8392 10464
rect 8444 10412 8450 10464
rect 10226 10412 10232 10464
rect 10284 10452 10290 10464
rect 11517 10455 11575 10461
rect 11517 10452 11529 10455
rect 10284 10424 11529 10452
rect 10284 10412 10290 10424
rect 11517 10421 11529 10424
rect 11563 10421 11575 10455
rect 11517 10415 11575 10421
rect 12894 10412 12900 10464
rect 12952 10412 12958 10464
rect 15841 10455 15899 10461
rect 15841 10421 15853 10455
rect 15887 10452 15899 10455
rect 16114 10452 16120 10464
rect 15887 10424 16120 10452
rect 15887 10421 15899 10424
rect 15841 10415 15899 10421
rect 16114 10412 16120 10424
rect 16172 10412 16178 10464
rect 19978 10412 19984 10464
rect 20036 10412 20042 10464
rect 21634 10412 21640 10464
rect 21692 10452 21698 10464
rect 23750 10452 23756 10464
rect 21692 10424 23756 10452
rect 21692 10412 21698 10424
rect 23750 10412 23756 10424
rect 23808 10412 23814 10464
rect 23842 10412 23848 10464
rect 23900 10412 23906 10464
rect 25130 10412 25136 10464
rect 25188 10452 25194 10464
rect 25593 10455 25651 10461
rect 25593 10452 25605 10455
rect 25188 10424 25605 10452
rect 25188 10412 25194 10424
rect 25593 10421 25605 10424
rect 25639 10421 25651 10455
rect 25593 10415 25651 10421
rect 26329 10455 26387 10461
rect 26329 10421 26341 10455
rect 26375 10452 26387 10455
rect 26418 10452 26424 10464
rect 26375 10424 26424 10452
rect 26375 10421 26387 10424
rect 26329 10415 26387 10421
rect 26418 10412 26424 10424
rect 26476 10412 26482 10464
rect 26804 10452 26832 10696
rect 26896 10588 26924 10764
rect 27724 10764 30113 10792
rect 27724 10733 27752 10764
rect 30101 10761 30113 10764
rect 30147 10761 30159 10795
rect 30101 10755 30159 10761
rect 30466 10752 30472 10804
rect 30524 10792 30530 10804
rect 30561 10795 30619 10801
rect 30561 10792 30573 10795
rect 30524 10764 30573 10792
rect 30524 10752 30530 10764
rect 30561 10761 30573 10764
rect 30607 10761 30619 10795
rect 30561 10755 30619 10761
rect 31754 10752 31760 10804
rect 31812 10752 31818 10804
rect 32953 10795 33011 10801
rect 31864 10764 32904 10792
rect 27709 10727 27767 10733
rect 27709 10693 27721 10727
rect 27755 10693 27767 10727
rect 31864 10724 31892 10764
rect 27709 10687 27767 10693
rect 29104 10696 31892 10724
rect 27430 10616 27436 10668
rect 27488 10616 27494 10668
rect 28718 10616 28724 10668
rect 28776 10656 28782 10668
rect 28776 10628 28842 10656
rect 28776 10616 28782 10628
rect 29104 10588 29132 10696
rect 32398 10684 32404 10736
rect 32456 10724 32462 10736
rect 32585 10727 32643 10733
rect 32585 10724 32597 10727
rect 32456 10696 32597 10724
rect 32456 10684 32462 10696
rect 32585 10693 32597 10696
rect 32631 10693 32643 10727
rect 32585 10687 32643 10693
rect 32766 10684 32772 10736
rect 32824 10733 32830 10736
rect 32824 10727 32843 10733
rect 32831 10693 32843 10727
rect 32876 10724 32904 10764
rect 32953 10761 32965 10795
rect 32999 10792 33011 10795
rect 33042 10792 33048 10804
rect 32999 10764 33048 10792
rect 32999 10761 33011 10764
rect 32953 10755 33011 10761
rect 33042 10752 33048 10764
rect 33100 10752 33106 10804
rect 33137 10795 33195 10801
rect 33137 10761 33149 10795
rect 33183 10792 33195 10795
rect 34422 10792 34428 10804
rect 33183 10764 34428 10792
rect 33183 10761 33195 10764
rect 33137 10755 33195 10761
rect 34422 10752 34428 10764
rect 34480 10752 34486 10804
rect 40954 10792 40960 10804
rect 34532 10764 40960 10792
rect 34532 10724 34560 10764
rect 40954 10752 40960 10764
rect 41012 10752 41018 10804
rect 32876 10696 34560 10724
rect 32824 10687 32843 10693
rect 32824 10684 32830 10687
rect 35894 10684 35900 10736
rect 35952 10724 35958 10736
rect 37553 10727 37611 10733
rect 37553 10724 37565 10727
rect 35952 10696 37565 10724
rect 35952 10684 35958 10696
rect 37553 10693 37565 10696
rect 37599 10693 37611 10727
rect 37553 10687 37611 10693
rect 29178 10616 29184 10668
rect 29236 10656 29242 10668
rect 29457 10659 29515 10665
rect 29457 10656 29469 10659
rect 29236 10628 29469 10656
rect 29236 10616 29242 10628
rect 29457 10625 29469 10628
rect 29503 10625 29515 10659
rect 29457 10619 29515 10625
rect 26896 10560 29132 10588
rect 29472 10588 29500 10619
rect 29546 10616 29552 10668
rect 29604 10616 29610 10668
rect 29638 10616 29644 10668
rect 29696 10656 29702 10668
rect 29733 10659 29791 10665
rect 29733 10656 29745 10659
rect 29696 10628 29745 10656
rect 29696 10616 29702 10628
rect 29733 10625 29745 10628
rect 29779 10625 29791 10659
rect 29733 10619 29791 10625
rect 29825 10659 29883 10665
rect 29825 10625 29837 10659
rect 29871 10625 29883 10659
rect 29825 10619 29883 10625
rect 29917 10659 29975 10665
rect 29917 10625 29929 10659
rect 29963 10656 29975 10659
rect 30098 10656 30104 10668
rect 29963 10628 30104 10656
rect 29963 10625 29975 10628
rect 29917 10619 29975 10625
rect 29840 10588 29868 10619
rect 30098 10616 30104 10628
rect 30156 10616 30162 10668
rect 30190 10616 30196 10668
rect 30248 10616 30254 10668
rect 30377 10659 30435 10665
rect 30377 10625 30389 10659
rect 30423 10656 30435 10659
rect 30834 10656 30840 10668
rect 30423 10628 30840 10656
rect 30423 10625 30435 10628
rect 30377 10619 30435 10625
rect 30834 10616 30840 10628
rect 30892 10656 30898 10668
rect 30892 10628 31064 10656
rect 30892 10616 30898 10628
rect 29472 10560 29868 10588
rect 31036 10532 31064 10628
rect 31478 10616 31484 10668
rect 31536 10616 31542 10668
rect 31665 10659 31723 10665
rect 31665 10625 31677 10659
rect 31711 10625 31723 10659
rect 31665 10619 31723 10625
rect 31849 10659 31907 10665
rect 31849 10625 31861 10659
rect 31895 10656 31907 10659
rect 32030 10656 32036 10668
rect 31895 10628 32036 10656
rect 31895 10625 31907 10628
rect 31849 10619 31907 10625
rect 31113 10591 31171 10597
rect 31113 10557 31125 10591
rect 31159 10588 31171 10591
rect 31202 10588 31208 10600
rect 31159 10560 31208 10588
rect 31159 10557 31171 10560
rect 31113 10551 31171 10557
rect 31202 10548 31208 10560
rect 31260 10548 31266 10600
rect 31297 10591 31355 10597
rect 31297 10557 31309 10591
rect 31343 10557 31355 10591
rect 31496 10588 31524 10616
rect 31680 10588 31708 10619
rect 32030 10616 32036 10628
rect 32088 10616 32094 10668
rect 32950 10616 32956 10668
rect 33008 10616 33014 10668
rect 33229 10659 33287 10665
rect 33229 10625 33241 10659
rect 33275 10656 33287 10659
rect 33502 10656 33508 10668
rect 33275 10628 33508 10656
rect 33275 10625 33287 10628
rect 33229 10619 33287 10625
rect 33502 10616 33508 10628
rect 33560 10616 33566 10668
rect 33778 10616 33784 10668
rect 33836 10616 33842 10668
rect 36078 10616 36084 10668
rect 36136 10656 36142 10668
rect 37277 10659 37335 10665
rect 37277 10656 37289 10659
rect 36136 10628 37289 10656
rect 36136 10616 36142 10628
rect 37277 10625 37289 10628
rect 37323 10625 37335 10659
rect 37277 10619 37335 10625
rect 37461 10659 37519 10665
rect 37461 10625 37473 10659
rect 37507 10656 37519 10659
rect 37507 10628 37596 10656
rect 37507 10625 37519 10628
rect 37461 10619 37519 10625
rect 31496 10560 31708 10588
rect 32968 10588 32996 10616
rect 37568 10600 37596 10628
rect 37642 10616 37648 10668
rect 37700 10616 37706 10668
rect 33873 10591 33931 10597
rect 33873 10588 33885 10591
rect 32968 10560 33885 10588
rect 31297 10551 31355 10557
rect 33873 10557 33885 10560
rect 33919 10588 33931 10591
rect 34054 10588 34060 10600
rect 33919 10560 34060 10588
rect 33919 10557 33931 10560
rect 33873 10551 33931 10557
rect 31018 10480 31024 10532
rect 31076 10480 31082 10532
rect 31312 10520 31340 10551
rect 34054 10548 34060 10560
rect 34112 10548 34118 10600
rect 35434 10548 35440 10600
rect 35492 10588 35498 10600
rect 36354 10588 36360 10600
rect 35492 10560 36360 10588
rect 35492 10548 35498 10560
rect 36354 10548 36360 10560
rect 36412 10548 36418 10600
rect 37550 10548 37556 10600
rect 37608 10548 37614 10600
rect 32122 10520 32128 10532
rect 31312 10492 32128 10520
rect 32122 10480 32128 10492
rect 32180 10480 32186 10532
rect 28442 10452 28448 10464
rect 26804 10424 28448 10452
rect 28442 10412 28448 10424
rect 28500 10412 28506 10464
rect 29546 10412 29552 10464
rect 29604 10452 29610 10464
rect 29914 10452 29920 10464
rect 29604 10424 29920 10452
rect 29604 10412 29610 10424
rect 29914 10412 29920 10424
rect 29972 10452 29978 10464
rect 30558 10452 30564 10464
rect 29972 10424 30564 10452
rect 29972 10412 29978 10424
rect 30558 10412 30564 10424
rect 30616 10412 30622 10464
rect 32674 10412 32680 10464
rect 32732 10452 32738 10464
rect 32769 10455 32827 10461
rect 32769 10452 32781 10455
rect 32732 10424 32781 10452
rect 32732 10412 32738 10424
rect 32769 10421 32781 10424
rect 32815 10421 32827 10455
rect 32769 10415 32827 10421
rect 37826 10412 37832 10464
rect 37884 10412 37890 10464
rect 1104 10362 41400 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 41400 10362
rect 1104 10288 41400 10310
rect 4798 10208 4804 10260
rect 4856 10248 4862 10260
rect 4893 10251 4951 10257
rect 4893 10248 4905 10251
rect 4856 10220 4905 10248
rect 4856 10208 4862 10220
rect 4893 10217 4905 10220
rect 4939 10217 4951 10251
rect 4893 10211 4951 10217
rect 5169 10251 5227 10257
rect 5169 10217 5181 10251
rect 5215 10248 5227 10251
rect 5813 10251 5871 10257
rect 5813 10248 5825 10251
rect 5215 10220 5825 10248
rect 5215 10217 5227 10220
rect 5169 10211 5227 10217
rect 5813 10217 5825 10220
rect 5859 10217 5871 10251
rect 5813 10211 5871 10217
rect 8386 10208 8392 10260
rect 8444 10208 8450 10260
rect 8478 10208 8484 10260
rect 8536 10248 8542 10260
rect 9769 10251 9827 10257
rect 9769 10248 9781 10251
rect 8536 10220 9781 10248
rect 8536 10208 8542 10220
rect 9769 10217 9781 10220
rect 9815 10217 9827 10251
rect 9769 10211 9827 10217
rect 11422 10208 11428 10260
rect 11480 10248 11486 10260
rect 17494 10248 17500 10260
rect 11480 10220 17500 10248
rect 11480 10208 11486 10220
rect 17494 10208 17500 10220
rect 17552 10208 17558 10260
rect 19334 10208 19340 10260
rect 19392 10248 19398 10260
rect 20073 10251 20131 10257
rect 20073 10248 20085 10251
rect 19392 10220 20085 10248
rect 19392 10208 19398 10220
rect 20073 10217 20085 10220
rect 20119 10217 20131 10251
rect 20073 10211 20131 10217
rect 20438 10208 20444 10260
rect 20496 10248 20502 10260
rect 20806 10248 20812 10260
rect 20496 10220 20812 10248
rect 20496 10208 20502 10220
rect 20806 10208 20812 10220
rect 20864 10208 20870 10260
rect 21450 10208 21456 10260
rect 21508 10208 21514 10260
rect 22186 10208 22192 10260
rect 22244 10248 22250 10260
rect 22370 10248 22376 10260
rect 22244 10220 22376 10248
rect 22244 10208 22250 10220
rect 22370 10208 22376 10220
rect 22428 10208 22434 10260
rect 22554 10208 22560 10260
rect 22612 10208 22618 10260
rect 23842 10208 23848 10260
rect 23900 10208 23906 10260
rect 24486 10208 24492 10260
rect 24544 10208 24550 10260
rect 26145 10251 26203 10257
rect 26145 10217 26157 10251
rect 26191 10248 26203 10251
rect 26234 10248 26240 10260
rect 26191 10220 26240 10248
rect 26191 10217 26203 10220
rect 26145 10211 26203 10217
rect 26234 10208 26240 10220
rect 26292 10208 26298 10260
rect 26510 10208 26516 10260
rect 26568 10248 26574 10260
rect 26970 10248 26976 10260
rect 26568 10220 26976 10248
rect 26568 10208 26574 10220
rect 26970 10208 26976 10220
rect 27028 10208 27034 10260
rect 27430 10208 27436 10260
rect 27488 10248 27494 10260
rect 28718 10248 28724 10260
rect 27488 10220 28724 10248
rect 27488 10208 27494 10220
rect 28718 10208 28724 10220
rect 28776 10248 28782 10260
rect 28813 10251 28871 10257
rect 28813 10248 28825 10251
rect 28776 10220 28825 10248
rect 28776 10208 28782 10220
rect 28813 10217 28825 10220
rect 28859 10217 28871 10251
rect 28813 10211 28871 10217
rect 30190 10208 30196 10260
rect 30248 10248 30254 10260
rect 31478 10248 31484 10260
rect 30248 10220 31484 10248
rect 30248 10208 30254 10220
rect 31478 10208 31484 10220
rect 31536 10208 31542 10260
rect 32674 10208 32680 10260
rect 32732 10208 32738 10260
rect 37826 10208 37832 10260
rect 37884 10248 37890 10260
rect 38105 10251 38163 10257
rect 38105 10248 38117 10251
rect 37884 10220 38117 10248
rect 37884 10208 37890 10220
rect 38105 10217 38117 10220
rect 38151 10217 38163 10251
rect 38105 10211 38163 10217
rect 38565 10251 38623 10257
rect 38565 10217 38577 10251
rect 38611 10248 38623 10251
rect 39850 10248 39856 10260
rect 38611 10220 39856 10248
rect 38611 10217 38623 10220
rect 38565 10211 38623 10217
rect 39850 10208 39856 10220
rect 39908 10208 39914 10260
rect 5077 10183 5135 10189
rect 5077 10149 5089 10183
rect 5123 10149 5135 10183
rect 5077 10143 5135 10149
rect 5092 10112 5120 10143
rect 7742 10140 7748 10192
rect 7800 10180 7806 10192
rect 7929 10183 7987 10189
rect 7929 10180 7941 10183
rect 7800 10152 7941 10180
rect 7800 10140 7806 10152
rect 7929 10149 7941 10152
rect 7975 10149 7987 10183
rect 7929 10143 7987 10149
rect 5905 10115 5963 10121
rect 5092 10084 5856 10112
rect 5828 10053 5856 10084
rect 5905 10081 5917 10115
rect 5951 10112 5963 10115
rect 5994 10112 6000 10124
rect 5951 10084 6000 10112
rect 5951 10081 5963 10084
rect 5905 10075 5963 10081
rect 5994 10072 6000 10084
rect 6052 10072 6058 10124
rect 8404 10112 8432 10208
rect 8754 10140 8760 10192
rect 8812 10140 8818 10192
rect 13630 10140 13636 10192
rect 13688 10140 13694 10192
rect 16022 10140 16028 10192
rect 16080 10140 16086 10192
rect 22094 10140 22100 10192
rect 22152 10140 22158 10192
rect 22572 10180 22600 10208
rect 22204 10152 22600 10180
rect 7944 10084 8432 10112
rect 8772 10112 8800 10140
rect 9306 10112 9312 10124
rect 8772 10084 9312 10112
rect 7944 10053 7972 10084
rect 5445 10047 5503 10053
rect 5445 10044 5457 10047
rect 5000 10016 5457 10044
rect 4709 9979 4767 9985
rect 4709 9945 4721 9979
rect 4755 9945 4767 9979
rect 4709 9939 4767 9945
rect 4724 9908 4752 9939
rect 4890 9936 4896 9988
rect 4948 9985 4954 9988
rect 4948 9979 4972 9985
rect 4960 9976 4972 9979
rect 5000 9976 5028 10016
rect 5445 10013 5457 10016
rect 5491 10013 5503 10047
rect 5445 10007 5503 10013
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10013 5871 10047
rect 5813 10007 5871 10013
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 8110 10004 8116 10056
rect 8168 10004 8174 10056
rect 8205 10047 8263 10053
rect 8205 10013 8217 10047
rect 8251 10044 8263 10047
rect 8772 10044 8800 10084
rect 9306 10072 9312 10084
rect 9364 10072 9370 10124
rect 9766 10112 9772 10124
rect 9416 10084 9772 10112
rect 8251 10016 8800 10044
rect 8251 10013 8263 10016
rect 8205 10007 8263 10013
rect 8846 10004 8852 10056
rect 8904 10044 8910 10056
rect 9416 10053 9444 10084
rect 9766 10072 9772 10084
rect 9824 10112 9830 10124
rect 10226 10112 10232 10124
rect 9824 10084 10232 10112
rect 9824 10072 9830 10084
rect 10226 10072 10232 10084
rect 10284 10072 10290 10124
rect 13648 10112 13676 10140
rect 16298 10112 16304 10124
rect 13648 10084 14136 10112
rect 9217 10047 9275 10053
rect 9217 10044 9229 10047
rect 8904 10016 9229 10044
rect 8904 10004 8910 10016
rect 9217 10013 9229 10016
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10013 9459 10047
rect 9401 10007 9459 10013
rect 9677 10047 9735 10053
rect 9677 10013 9689 10047
rect 9723 10044 9735 10047
rect 9858 10044 9864 10056
rect 9723 10016 9864 10044
rect 9723 10013 9735 10016
rect 9677 10007 9735 10013
rect 4960 9948 5028 9976
rect 5169 9979 5227 9985
rect 4960 9945 4972 9948
rect 4948 9939 4972 9945
rect 5169 9945 5181 9979
rect 5215 9976 5227 9979
rect 5258 9976 5264 9988
rect 5215 9948 5264 9976
rect 5215 9945 5227 9948
rect 5169 9939 5227 9945
rect 4948 9936 4954 9939
rect 5184 9908 5212 9939
rect 5258 9936 5264 9948
rect 5316 9936 5322 9988
rect 5350 9936 5356 9988
rect 5408 9936 5414 9988
rect 9232 9976 9260 10007
rect 9858 10004 9864 10016
rect 9916 10004 9922 10056
rect 12069 10047 12127 10053
rect 12069 10013 12081 10047
rect 12115 10044 12127 10047
rect 12618 10044 12624 10056
rect 12115 10016 12624 10044
rect 12115 10013 12127 10016
rect 12069 10007 12127 10013
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 13740 10053 13768 10084
rect 14108 10053 14136 10084
rect 16040 10084 16304 10112
rect 13633 10047 13691 10053
rect 13633 10013 13645 10047
rect 13679 10013 13691 10047
rect 13633 10007 13691 10013
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10044 13783 10047
rect 14093 10047 14151 10053
rect 13771 10016 13805 10044
rect 13771 10013 13783 10016
rect 13725 10007 13783 10013
rect 14093 10013 14105 10047
rect 14139 10044 14151 10047
rect 14182 10044 14188 10056
rect 14139 10016 14188 10044
rect 14139 10013 14151 10016
rect 14093 10007 14151 10013
rect 13648 9976 13676 10007
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 15749 10047 15807 10053
rect 15749 10013 15761 10047
rect 15795 10044 15807 10047
rect 15795 10016 15976 10044
rect 15795 10013 15807 10016
rect 15749 10007 15807 10013
rect 15948 9988 15976 10016
rect 13814 9976 13820 9988
rect 9232 9948 9904 9976
rect 13648 9948 13820 9976
rect 9876 9920 9904 9948
rect 13814 9936 13820 9948
rect 13872 9976 13878 9988
rect 14277 9979 14335 9985
rect 14277 9976 14289 9979
rect 13872 9948 14289 9976
rect 13872 9936 13878 9948
rect 14277 9945 14289 9948
rect 14323 9945 14335 9979
rect 14277 9939 14335 9945
rect 15930 9936 15936 9988
rect 15988 9936 15994 9988
rect 4724 9880 5212 9908
rect 5718 9868 5724 9920
rect 5776 9908 5782 9920
rect 6181 9911 6239 9917
rect 6181 9908 6193 9911
rect 5776 9880 6193 9908
rect 5776 9868 5782 9880
rect 6181 9877 6193 9880
rect 6227 9877 6239 9911
rect 6181 9871 6239 9877
rect 9582 9868 9588 9920
rect 9640 9868 9646 9920
rect 9858 9868 9864 9920
rect 9916 9868 9922 9920
rect 12158 9868 12164 9920
rect 12216 9868 12222 9920
rect 13906 9868 13912 9920
rect 13964 9868 13970 9920
rect 13998 9868 14004 9920
rect 14056 9908 14062 9920
rect 14461 9911 14519 9917
rect 14461 9908 14473 9911
rect 14056 9880 14473 9908
rect 14056 9868 14062 9880
rect 14461 9877 14473 9880
rect 14507 9877 14519 9911
rect 14461 9871 14519 9877
rect 15838 9868 15844 9920
rect 15896 9908 15902 9920
rect 16040 9908 16068 10084
rect 16298 10072 16304 10084
rect 16356 10112 16362 10124
rect 16356 10084 16804 10112
rect 16356 10072 16362 10084
rect 16114 10004 16120 10056
rect 16172 10004 16178 10056
rect 16776 10053 16804 10084
rect 16850 10072 16856 10124
rect 16908 10112 16914 10124
rect 20162 10112 20168 10124
rect 16908 10084 20168 10112
rect 16908 10072 16914 10084
rect 20162 10072 20168 10084
rect 20220 10072 20226 10124
rect 20990 10112 20996 10124
rect 20272 10084 20996 10112
rect 16761 10047 16819 10053
rect 16761 10013 16773 10047
rect 16807 10013 16819 10047
rect 16761 10007 16819 10013
rect 16945 10047 17003 10053
rect 16945 10013 16957 10047
rect 16991 10013 17003 10047
rect 16945 10007 17003 10013
rect 16132 9976 16160 10004
rect 16960 9976 16988 10007
rect 19150 10004 19156 10056
rect 19208 10044 19214 10056
rect 20272 10053 20300 10084
rect 20990 10072 20996 10084
rect 21048 10072 21054 10124
rect 20257 10047 20315 10053
rect 20257 10044 20269 10047
rect 19208 10016 20269 10044
rect 19208 10004 19214 10016
rect 20257 10013 20269 10016
rect 20303 10013 20315 10047
rect 20257 10007 20315 10013
rect 20441 10047 20499 10053
rect 20441 10013 20453 10047
rect 20487 10044 20499 10047
rect 20809 10047 20867 10053
rect 20809 10044 20821 10047
rect 20487 10016 20821 10044
rect 20487 10013 20499 10016
rect 20441 10007 20499 10013
rect 20809 10013 20821 10016
rect 20855 10044 20867 10047
rect 21174 10044 21180 10056
rect 20855 10016 21180 10044
rect 20855 10013 20867 10016
rect 20809 10007 20867 10013
rect 21174 10004 21180 10016
rect 21232 10004 21238 10056
rect 21545 10047 21603 10053
rect 21545 10013 21557 10047
rect 21591 10044 21603 10047
rect 21634 10044 21640 10056
rect 21591 10016 21640 10044
rect 21591 10013 21603 10016
rect 21545 10007 21603 10013
rect 21634 10004 21640 10016
rect 21692 10004 21698 10056
rect 21913 10047 21971 10053
rect 21913 10013 21925 10047
rect 21959 10044 21971 10047
rect 22002 10044 22008 10056
rect 21959 10016 22008 10044
rect 21959 10013 21971 10016
rect 21913 10007 21971 10013
rect 22002 10004 22008 10016
rect 22060 10044 22066 10056
rect 22204 10044 22232 10152
rect 23382 10140 23388 10192
rect 23440 10140 23446 10192
rect 23860 10112 23888 10208
rect 22296 10084 23888 10112
rect 24397 10115 24455 10121
rect 22296 10053 22324 10084
rect 24397 10081 24409 10115
rect 24443 10112 24455 10115
rect 24504 10112 24532 10208
rect 30101 10183 30159 10189
rect 30101 10180 30113 10183
rect 26896 10152 30113 10180
rect 25222 10112 25228 10124
rect 24443 10084 25228 10112
rect 24443 10081 24455 10084
rect 24397 10075 24455 10081
rect 25222 10072 25228 10084
rect 25280 10072 25286 10124
rect 26896 10121 26924 10152
rect 30101 10149 30113 10152
rect 30147 10149 30159 10183
rect 31846 10180 31852 10192
rect 30101 10143 30159 10149
rect 30392 10152 31852 10180
rect 26881 10115 26939 10121
rect 26881 10081 26893 10115
rect 26927 10081 26939 10115
rect 26881 10075 26939 10081
rect 27062 10072 27068 10124
rect 27120 10072 27126 10124
rect 28534 10072 28540 10124
rect 28592 10112 28598 10124
rect 29270 10112 29276 10124
rect 28592 10084 29276 10112
rect 28592 10072 28598 10084
rect 29270 10072 29276 10084
rect 29328 10072 29334 10124
rect 30392 10112 30420 10152
rect 31846 10140 31852 10152
rect 31904 10180 31910 10192
rect 32490 10180 32496 10192
rect 31904 10152 32496 10180
rect 31904 10140 31910 10152
rect 32490 10140 32496 10152
rect 32548 10140 32554 10192
rect 32692 10180 32720 10208
rect 32692 10152 33180 10180
rect 30300 10084 30420 10112
rect 22060 10016 22232 10044
rect 22281 10047 22339 10053
rect 22060 10004 22066 10016
rect 22281 10013 22293 10047
rect 22327 10013 22339 10047
rect 22281 10007 22339 10013
rect 22554 10004 22560 10056
rect 22612 10004 22618 10056
rect 23106 10004 23112 10056
rect 23164 10044 23170 10056
rect 23385 10047 23443 10053
rect 23385 10044 23397 10047
rect 23164 10016 23397 10044
rect 23164 10004 23170 10016
rect 23385 10013 23397 10016
rect 23431 10013 23443 10047
rect 23385 10007 23443 10013
rect 23566 10004 23572 10056
rect 23624 10044 23630 10056
rect 23624 10016 24118 10044
rect 23624 10004 23630 10016
rect 16132 9948 16988 9976
rect 19797 9979 19855 9985
rect 19797 9945 19809 9979
rect 19843 9976 19855 9979
rect 20717 9979 20775 9985
rect 20717 9976 20729 9979
rect 19843 9948 20729 9976
rect 19843 9945 19855 9948
rect 19797 9939 19855 9945
rect 20717 9945 20729 9948
rect 20763 9976 20775 9979
rect 20898 9976 20904 9988
rect 20763 9948 20904 9976
rect 20763 9945 20775 9948
rect 20717 9939 20775 9945
rect 20898 9936 20904 9948
rect 20956 9936 20962 9988
rect 21266 9936 21272 9988
rect 21324 9976 21330 9988
rect 21729 9979 21787 9985
rect 21729 9976 21741 9979
rect 21324 9948 21741 9976
rect 21324 9936 21330 9948
rect 21729 9945 21741 9948
rect 21775 9945 21787 9979
rect 21729 9939 21787 9945
rect 21821 9979 21879 9985
rect 21821 9945 21833 9979
rect 21867 9976 21879 9979
rect 23584 9976 23612 10004
rect 21867 9948 23612 9976
rect 21867 9945 21879 9948
rect 21821 9939 21879 9945
rect 24090 9920 24118 10016
rect 26786 10004 26792 10056
rect 26844 10004 26850 10056
rect 27614 10004 27620 10056
rect 27672 10044 27678 10056
rect 28077 10047 28135 10053
rect 28077 10044 28089 10047
rect 27672 10016 28089 10044
rect 27672 10004 27678 10016
rect 28077 10013 28089 10016
rect 28123 10013 28135 10047
rect 28077 10007 28135 10013
rect 28237 10047 28295 10053
rect 28237 10013 28249 10047
rect 28283 10044 28295 10047
rect 29730 10044 29736 10056
rect 28283 10013 28304 10044
rect 28237 10007 28304 10013
rect 24673 9979 24731 9985
rect 24673 9945 24685 9979
rect 24719 9976 24731 9979
rect 24946 9976 24952 9988
rect 24719 9948 24952 9976
rect 24719 9945 24731 9948
rect 24673 9939 24731 9945
rect 24946 9936 24952 9948
rect 25004 9936 25010 9988
rect 25130 9936 25136 9988
rect 25188 9936 25194 9988
rect 28276 9976 28304 10007
rect 28460 10016 29736 10044
rect 28460 9976 28488 10016
rect 29730 10004 29736 10016
rect 29788 10004 29794 10056
rect 30300 10053 30328 10084
rect 30466 10072 30472 10124
rect 30524 10072 30530 10124
rect 31018 10072 31024 10124
rect 31076 10112 31082 10124
rect 31665 10115 31723 10121
rect 31665 10112 31677 10115
rect 31076 10084 31677 10112
rect 31076 10072 31082 10084
rect 31665 10081 31677 10084
rect 31711 10112 31723 10115
rect 32398 10112 32404 10124
rect 31711 10084 32404 10112
rect 31711 10081 31723 10084
rect 31665 10075 31723 10081
rect 32398 10072 32404 10084
rect 32456 10112 32462 10124
rect 32456 10084 32996 10112
rect 32456 10072 32462 10084
rect 30285 10047 30343 10053
rect 30285 10013 30297 10047
rect 30331 10013 30343 10047
rect 30285 10007 30343 10013
rect 30377 10047 30435 10053
rect 30377 10013 30389 10047
rect 30423 10044 30435 10047
rect 30484 10044 30512 10072
rect 30423 10016 30512 10044
rect 30423 10013 30435 10016
rect 30377 10007 30435 10013
rect 31294 10004 31300 10056
rect 31352 10004 31358 10056
rect 31570 10004 31576 10056
rect 31628 10004 31634 10056
rect 31757 10047 31815 10053
rect 31757 10013 31769 10047
rect 31803 10013 31815 10047
rect 31757 10007 31815 10013
rect 25976 9948 28304 9976
rect 28368 9948 28488 9976
rect 28721 9979 28779 9985
rect 15896 9880 16068 9908
rect 15896 9868 15902 9880
rect 16942 9868 16948 9920
rect 17000 9908 17006 9920
rect 17129 9911 17187 9917
rect 17129 9908 17141 9911
rect 17000 9880 17141 9908
rect 17000 9868 17006 9880
rect 17129 9877 17141 9880
rect 17175 9877 17187 9911
rect 24090 9880 24124 9920
rect 17129 9871 17187 9877
rect 24118 9868 24124 9880
rect 24176 9908 24182 9920
rect 25976 9908 26004 9948
rect 24176 9880 26004 9908
rect 24176 9868 24182 9880
rect 26418 9868 26424 9920
rect 26476 9868 26482 9920
rect 27062 9868 27068 9920
rect 27120 9908 27126 9920
rect 27982 9908 27988 9920
rect 27120 9880 27988 9908
rect 27120 9868 27126 9880
rect 27982 9868 27988 9880
rect 28040 9868 28046 9920
rect 28074 9868 28080 9920
rect 28132 9908 28138 9920
rect 28169 9911 28227 9917
rect 28169 9908 28181 9911
rect 28132 9880 28181 9908
rect 28132 9868 28138 9880
rect 28169 9877 28181 9880
rect 28215 9908 28227 9911
rect 28368 9908 28396 9948
rect 28721 9945 28733 9979
rect 28767 9945 28779 9979
rect 28721 9939 28779 9945
rect 30101 9979 30159 9985
rect 30101 9945 30113 9979
rect 30147 9976 30159 9979
rect 31312 9976 31340 10004
rect 31772 9976 31800 10007
rect 32122 10004 32128 10056
rect 32180 10044 32186 10056
rect 32968 10053 32996 10084
rect 33152 10053 33180 10152
rect 38194 10072 38200 10124
rect 38252 10072 38258 10124
rect 32769 10047 32827 10053
rect 32769 10044 32781 10047
rect 32180 10016 32781 10044
rect 32180 10004 32186 10016
rect 32769 10013 32781 10016
rect 32815 10013 32827 10047
rect 32769 10007 32827 10013
rect 32953 10047 33011 10053
rect 32953 10013 32965 10047
rect 32999 10013 33011 10047
rect 32953 10007 33011 10013
rect 33137 10047 33195 10053
rect 33137 10013 33149 10047
rect 33183 10013 33195 10047
rect 33137 10007 33195 10013
rect 33502 10004 33508 10056
rect 33560 10004 33566 10056
rect 38102 10004 38108 10056
rect 38160 10004 38166 10056
rect 38378 10004 38384 10056
rect 38436 10004 38442 10056
rect 30147 9948 30328 9976
rect 31312 9948 31800 9976
rect 32861 9979 32919 9985
rect 30147 9945 30159 9948
rect 30101 9939 30159 9945
rect 28215 9880 28396 9908
rect 28215 9877 28227 9880
rect 28169 9871 28227 9877
rect 28442 9868 28448 9920
rect 28500 9908 28506 9920
rect 28736 9908 28764 9939
rect 30300 9920 30328 9948
rect 32861 9945 32873 9979
rect 32907 9976 32919 9979
rect 33321 9979 33379 9985
rect 33321 9976 33333 9979
rect 32907 9948 33333 9976
rect 32907 9945 32919 9948
rect 32861 9939 32919 9945
rect 33321 9945 33333 9948
rect 33367 9945 33379 9979
rect 33321 9939 33379 9945
rect 33413 9979 33471 9985
rect 33413 9945 33425 9979
rect 33459 9945 33471 9979
rect 33413 9939 33471 9945
rect 28994 9908 29000 9920
rect 28500 9880 29000 9908
rect 28500 9868 28506 9880
rect 28994 9868 29000 9880
rect 29052 9868 29058 9920
rect 30282 9868 30288 9920
rect 30340 9868 30346 9920
rect 31846 9868 31852 9920
rect 31904 9908 31910 9920
rect 32030 9908 32036 9920
rect 31904 9880 32036 9908
rect 31904 9868 31910 9880
rect 32030 9868 32036 9880
rect 32088 9908 32094 9920
rect 32306 9908 32312 9920
rect 32088 9880 32312 9908
rect 32088 9868 32094 9880
rect 32306 9868 32312 9880
rect 32364 9868 32370 9920
rect 33134 9868 33140 9920
rect 33192 9908 33198 9920
rect 33428 9908 33456 9939
rect 33192 9880 33456 9908
rect 33192 9868 33198 9880
rect 33686 9868 33692 9920
rect 33744 9868 33750 9920
rect 1104 9818 41400 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 41400 9818
rect 1104 9744 41400 9766
rect 7193 9707 7251 9713
rect 7193 9673 7205 9707
rect 7239 9673 7251 9707
rect 7193 9667 7251 9673
rect 5537 9639 5595 9645
rect 5537 9605 5549 9639
rect 5583 9636 5595 9639
rect 5905 9639 5963 9645
rect 5905 9636 5917 9639
rect 5583 9608 5917 9636
rect 5583 9605 5595 9608
rect 5537 9599 5595 9605
rect 5905 9605 5917 9608
rect 5951 9605 5963 9639
rect 7208 9636 7236 9667
rect 8662 9664 8668 9716
rect 8720 9704 8726 9716
rect 9398 9704 9404 9716
rect 8720 9676 9404 9704
rect 8720 9664 8726 9676
rect 9398 9664 9404 9676
rect 9456 9664 9462 9716
rect 11256 9676 11836 9704
rect 5905 9599 5963 9605
rect 6104 9608 7236 9636
rect 7469 9639 7527 9645
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9568 5043 9571
rect 5074 9568 5080 9580
rect 5031 9540 5080 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 5074 9528 5080 9540
rect 5132 9568 5138 9580
rect 5442 9568 5448 9580
rect 5132 9540 5448 9568
rect 5132 9528 5138 9540
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9568 5687 9571
rect 5718 9568 5724 9580
rect 5675 9540 5724 9568
rect 5675 9537 5687 9540
rect 5629 9531 5687 9537
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9537 5871 9571
rect 5813 9531 5871 9537
rect 5828 9500 5856 9531
rect 5994 9528 6000 9580
rect 6052 9528 6058 9580
rect 6104 9500 6132 9608
rect 7469 9605 7481 9639
rect 7515 9636 7527 9639
rect 7650 9636 7656 9648
rect 7515 9608 7656 9636
rect 7515 9605 7527 9608
rect 7469 9599 7527 9605
rect 7650 9596 7656 9608
rect 7708 9596 7714 9648
rect 7834 9596 7840 9648
rect 7892 9596 7898 9648
rect 8938 9596 8944 9648
rect 8996 9596 9002 9648
rect 9122 9636 9128 9648
rect 9048 9608 9128 9636
rect 7835 9593 7893 9596
rect 6546 9528 6552 9580
rect 6604 9528 6610 9580
rect 6733 9571 6791 9577
rect 6733 9537 6745 9571
rect 6779 9568 6791 9571
rect 6914 9568 6920 9580
rect 6779 9540 6920 9568
rect 6779 9537 6791 9540
rect 6733 9531 6791 9537
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 7377 9571 7435 9577
rect 7377 9537 7389 9571
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 5828 9472 6132 9500
rect 7392 9500 7420 9531
rect 7558 9528 7564 9580
rect 7616 9528 7622 9580
rect 7742 9528 7748 9580
rect 7800 9528 7806 9580
rect 7835 9559 7847 9593
rect 7881 9559 7893 9593
rect 7835 9553 7893 9559
rect 8849 9571 8907 9577
rect 8849 9537 8861 9571
rect 8895 9568 8907 9571
rect 8956 9568 8984 9596
rect 9048 9577 9076 9608
rect 9122 9596 9128 9608
rect 9180 9636 9186 9648
rect 9582 9636 9588 9648
rect 9180 9608 9588 9636
rect 9180 9596 9186 9608
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 9677 9639 9735 9645
rect 9677 9605 9689 9639
rect 9723 9636 9735 9639
rect 9766 9636 9772 9648
rect 9723 9608 9772 9636
rect 9723 9605 9735 9608
rect 9677 9599 9735 9605
rect 9766 9596 9772 9608
rect 9824 9596 9830 9648
rect 9858 9596 9864 9648
rect 9916 9636 9922 9648
rect 11256 9636 11284 9676
rect 9916 9608 11284 9636
rect 11333 9639 11391 9645
rect 9916 9596 9922 9608
rect 11333 9605 11345 9639
rect 11379 9636 11391 9639
rect 11379 9608 11744 9636
rect 11379 9605 11391 9608
rect 11333 9599 11391 9605
rect 8895 9540 8984 9568
rect 9033 9571 9091 9577
rect 8895 9537 8907 9540
rect 8849 9531 8907 9537
rect 9033 9537 9045 9571
rect 9079 9537 9091 9571
rect 9033 9531 9091 9537
rect 9401 9571 9459 9577
rect 9401 9537 9413 9571
rect 9447 9568 9459 9571
rect 9490 9568 9496 9580
rect 9447 9540 9496 9568
rect 9447 9537 9459 9540
rect 9401 9531 9459 9537
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 9950 9528 9956 9580
rect 10008 9528 10014 9580
rect 11716 9577 11744 9608
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9568 11207 9571
rect 11517 9571 11575 9577
rect 11195 9540 11284 9568
rect 11195 9537 11207 9540
rect 11149 9531 11207 9537
rect 9125 9503 9183 9509
rect 7392 9472 8064 9500
rect 5258 9392 5264 9444
rect 5316 9432 5322 9444
rect 6549 9435 6607 9441
rect 6549 9432 6561 9435
rect 5316 9404 6561 9432
rect 5316 9392 5322 9404
rect 6549 9401 6561 9404
rect 6595 9401 6607 9435
rect 6549 9395 6607 9401
rect 7558 9392 7564 9444
rect 7616 9432 7622 9444
rect 7926 9432 7932 9444
rect 7616 9404 7932 9432
rect 7616 9392 7622 9404
rect 7926 9392 7932 9404
rect 7984 9392 7990 9444
rect 8036 9376 8064 9472
rect 9125 9469 9137 9503
rect 9171 9469 9183 9503
rect 9125 9463 9183 9469
rect 9217 9503 9275 9509
rect 9217 9469 9229 9503
rect 9263 9500 9275 9503
rect 9968 9500 9996 9528
rect 11256 9512 11284 9540
rect 11517 9537 11529 9571
rect 11563 9537 11575 9571
rect 11517 9531 11575 9537
rect 11701 9571 11759 9577
rect 11701 9537 11713 9571
rect 11747 9537 11759 9571
rect 11808 9568 11836 9676
rect 12894 9664 12900 9716
rect 12952 9664 12958 9716
rect 16114 9704 16120 9716
rect 15304 9676 16120 9704
rect 11882 9596 11888 9648
rect 11940 9636 11946 9648
rect 12912 9636 12940 9664
rect 11940 9608 12112 9636
rect 11940 9596 11946 9608
rect 12084 9577 12112 9608
rect 12452 9608 12940 9636
rect 13004 9608 13952 9636
rect 12452 9577 12480 9608
rect 12069 9571 12127 9577
rect 11808 9540 11928 9568
rect 11701 9531 11759 9537
rect 9263 9472 9996 9500
rect 10965 9503 11023 9509
rect 9263 9469 9275 9472
rect 9217 9463 9275 9469
rect 10965 9469 10977 9503
rect 11011 9500 11023 9503
rect 11054 9500 11060 9512
rect 11011 9472 11060 9500
rect 11011 9469 11023 9472
rect 10965 9463 11023 9469
rect 9140 9432 9168 9463
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 11238 9460 11244 9512
rect 11296 9460 11302 9512
rect 11330 9460 11336 9512
rect 11388 9500 11394 9512
rect 11532 9500 11560 9531
rect 11900 9509 11928 9540
rect 12069 9537 12081 9571
rect 12115 9537 12127 9571
rect 12069 9531 12127 9537
rect 12437 9571 12495 9577
rect 12437 9537 12449 9571
rect 12483 9537 12495 9571
rect 12437 9531 12495 9537
rect 12526 9528 12532 9580
rect 12584 9568 12590 9580
rect 12621 9571 12679 9577
rect 12621 9568 12633 9571
rect 12584 9540 12633 9568
rect 12584 9528 12590 9540
rect 12621 9537 12633 9540
rect 12667 9537 12679 9571
rect 12621 9531 12679 9537
rect 12710 9528 12716 9580
rect 12768 9528 12774 9580
rect 13004 9577 13032 9608
rect 13924 9580 13952 9608
rect 12989 9571 13047 9577
rect 12989 9537 13001 9571
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 13814 9528 13820 9580
rect 13872 9528 13878 9580
rect 13906 9528 13912 9580
rect 13964 9528 13970 9580
rect 14182 9528 14188 9580
rect 14240 9568 14246 9580
rect 15304 9577 15332 9676
rect 16114 9664 16120 9676
rect 16172 9664 16178 9716
rect 20714 9664 20720 9716
rect 20772 9704 20778 9716
rect 23106 9704 23112 9716
rect 20772 9676 21036 9704
rect 20772 9664 20778 9676
rect 19337 9639 19395 9645
rect 16040 9608 16988 9636
rect 14369 9571 14427 9577
rect 14369 9568 14381 9571
rect 14240 9540 14381 9568
rect 14240 9528 14246 9540
rect 14369 9537 14381 9540
rect 14415 9537 14427 9571
rect 14369 9531 14427 9537
rect 15289 9571 15347 9577
rect 15289 9537 15301 9571
rect 15335 9537 15347 9571
rect 15289 9531 15347 9537
rect 15473 9571 15531 9577
rect 15473 9537 15485 9571
rect 15519 9568 15531 9571
rect 15838 9568 15844 9580
rect 15519 9540 15844 9568
rect 15519 9537 15531 9540
rect 15473 9531 15531 9537
rect 15838 9528 15844 9540
rect 15896 9528 15902 9580
rect 16040 9577 16068 9608
rect 16960 9580 16988 9608
rect 19337 9605 19349 9639
rect 19383 9636 19395 9639
rect 19426 9636 19432 9648
rect 19383 9608 19432 9636
rect 19383 9605 19395 9608
rect 19337 9599 19395 9605
rect 19426 9596 19432 9608
rect 19484 9636 19490 9648
rect 19794 9636 19800 9648
rect 19484 9608 19800 9636
rect 19484 9596 19490 9608
rect 19794 9596 19800 9608
rect 19852 9596 19858 9648
rect 19889 9639 19947 9645
rect 19889 9605 19901 9639
rect 19935 9636 19947 9639
rect 19978 9636 19984 9648
rect 19935 9608 19984 9636
rect 19935 9605 19947 9608
rect 19889 9599 19947 9605
rect 19978 9596 19984 9608
rect 20036 9596 20042 9648
rect 16025 9571 16083 9577
rect 16025 9537 16037 9571
rect 16071 9537 16083 9571
rect 16025 9531 16083 9537
rect 16114 9528 16120 9580
rect 16172 9528 16178 9580
rect 16209 9571 16267 9577
rect 16209 9537 16221 9571
rect 16255 9568 16267 9571
rect 16393 9571 16451 9577
rect 16255 9540 16344 9568
rect 16255 9537 16267 9540
rect 16209 9531 16267 9537
rect 11388 9472 11560 9500
rect 11793 9503 11851 9509
rect 11388 9460 11394 9472
rect 11793 9469 11805 9503
rect 11839 9469 11851 9503
rect 11793 9463 11851 9469
rect 11885 9503 11943 9509
rect 11885 9469 11897 9503
rect 11931 9469 11943 9503
rect 12805 9503 12863 9509
rect 12805 9500 12817 9503
rect 11885 9463 11943 9469
rect 12406 9472 12817 9500
rect 9140 9404 9260 9432
rect 9232 9376 9260 9404
rect 9582 9392 9588 9444
rect 9640 9392 9646 9444
rect 9858 9392 9864 9444
rect 9916 9432 9922 9444
rect 10045 9435 10103 9441
rect 10045 9432 10057 9435
rect 9916 9404 10057 9432
rect 9916 9392 9922 9404
rect 10045 9401 10057 9404
rect 10091 9401 10103 9435
rect 11808 9432 11836 9463
rect 12406 9432 12434 9472
rect 12805 9469 12817 9472
rect 12851 9500 12863 9503
rect 16316 9500 16344 9540
rect 16393 9537 16405 9571
rect 16439 9570 16451 9571
rect 16439 9568 16528 9570
rect 16439 9542 16712 9568
rect 16439 9537 16451 9542
rect 16500 9540 16712 9542
rect 16393 9531 16451 9537
rect 16574 9500 16580 9512
rect 12851 9472 13308 9500
rect 16316 9472 16580 9500
rect 12851 9469 12863 9472
rect 12805 9463 12863 9469
rect 10045 9395 10103 9401
rect 11072 9404 12434 9432
rect 6178 9324 6184 9376
rect 6236 9324 6242 9376
rect 8018 9324 8024 9376
rect 8076 9324 8082 9376
rect 9214 9324 9220 9376
rect 9272 9364 9278 9376
rect 11072 9364 11100 9404
rect 9272 9336 11100 9364
rect 9272 9324 9278 9336
rect 11422 9324 11428 9376
rect 11480 9364 11486 9376
rect 12158 9364 12164 9376
rect 11480 9336 12164 9364
rect 11480 9324 11486 9336
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 12250 9324 12256 9376
rect 12308 9324 12314 9376
rect 13170 9324 13176 9376
rect 13228 9324 13234 9376
rect 13280 9364 13308 9472
rect 16574 9460 16580 9472
rect 16632 9460 16638 9512
rect 16684 9509 16712 9540
rect 16850 9528 16856 9580
rect 16908 9528 16914 9580
rect 16942 9528 16948 9580
rect 17000 9528 17006 9580
rect 17126 9528 17132 9580
rect 17184 9528 17190 9580
rect 17313 9571 17371 9577
rect 17313 9537 17325 9571
rect 17359 9537 17371 9571
rect 17313 9531 17371 9537
rect 16669 9503 16727 9509
rect 16669 9469 16681 9503
rect 16715 9469 16727 9503
rect 16669 9463 16727 9469
rect 13722 9392 13728 9444
rect 13780 9432 13786 9444
rect 14553 9435 14611 9441
rect 14553 9432 14565 9435
rect 13780 9404 14565 9432
rect 13780 9392 13786 9404
rect 14553 9401 14565 9404
rect 14599 9401 14611 9435
rect 14553 9395 14611 9401
rect 15289 9435 15347 9441
rect 15289 9401 15301 9435
rect 15335 9432 15347 9435
rect 16868 9432 16896 9528
rect 17037 9503 17095 9509
rect 17037 9500 17049 9503
rect 16960 9472 17049 9500
rect 16960 9444 16988 9472
rect 17037 9469 17049 9472
rect 17083 9469 17095 9503
rect 17037 9463 17095 9469
rect 15335 9404 16896 9432
rect 15335 9401 15347 9404
rect 15289 9395 15347 9401
rect 16942 9392 16948 9444
rect 17000 9392 17006 9444
rect 15194 9364 15200 9376
rect 13280 9336 15200 9364
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 15749 9367 15807 9373
rect 15749 9333 15761 9367
rect 15795 9364 15807 9367
rect 16390 9364 16396 9376
rect 15795 9336 16396 9364
rect 15795 9333 15807 9336
rect 15749 9327 15807 9333
rect 16390 9324 16396 9336
rect 16448 9324 16454 9376
rect 16482 9324 16488 9376
rect 16540 9364 16546 9376
rect 17328 9364 17356 9531
rect 19150 9528 19156 9580
rect 19208 9528 19214 9580
rect 21008 9554 21036 9676
rect 21652 9676 23112 9704
rect 21174 9596 21180 9648
rect 21232 9636 21238 9648
rect 21652 9645 21680 9676
rect 23106 9664 23112 9676
rect 23164 9664 23170 9716
rect 24854 9664 24860 9716
rect 24912 9704 24918 9716
rect 25130 9704 25136 9716
rect 24912 9676 25136 9704
rect 24912 9664 24918 9676
rect 25130 9664 25136 9676
rect 25188 9664 25194 9716
rect 25958 9664 25964 9716
rect 26016 9664 26022 9716
rect 26252 9676 26464 9704
rect 21637 9639 21695 9645
rect 21637 9636 21649 9639
rect 21232 9608 21649 9636
rect 21232 9596 21238 9608
rect 21637 9605 21649 9608
rect 21683 9605 21695 9639
rect 21637 9599 21695 9605
rect 22097 9639 22155 9645
rect 22097 9605 22109 9639
rect 22143 9636 22155 9639
rect 24872 9636 24900 9664
rect 26252 9645 26280 9676
rect 26237 9639 26295 9645
rect 22143 9608 22416 9636
rect 22143 9605 22155 9608
rect 22097 9599 22155 9605
rect 22002 9528 22008 9580
rect 22060 9528 22066 9580
rect 22186 9528 22192 9580
rect 22244 9528 22250 9580
rect 22388 9568 22416 9608
rect 22649 9571 22707 9577
rect 22649 9568 22661 9571
rect 22388 9540 22661 9568
rect 22649 9537 22661 9540
rect 22695 9537 22707 9571
rect 22649 9531 22707 9537
rect 23400 9568 23428 9622
rect 24136 9608 24978 9636
rect 25792 9608 26188 9636
rect 24136 9568 24164 9608
rect 25792 9568 25820 9608
rect 23400 9540 24164 9568
rect 25700 9540 25820 9568
rect 19613 9503 19671 9509
rect 19613 9469 19625 9503
rect 19659 9500 19671 9503
rect 19659 9472 19748 9500
rect 19659 9469 19671 9472
rect 19613 9463 19671 9469
rect 19720 9376 19748 9472
rect 21818 9460 21824 9512
rect 21876 9500 21882 9512
rect 22281 9503 22339 9509
rect 21876 9472 22094 9500
rect 21876 9460 21882 9472
rect 16540 9336 17356 9364
rect 16540 9324 16546 9336
rect 19426 9324 19432 9376
rect 19484 9364 19490 9376
rect 19521 9367 19579 9373
rect 19521 9364 19533 9367
rect 19484 9336 19533 9364
rect 19484 9324 19490 9336
rect 19521 9333 19533 9336
rect 19567 9333 19579 9367
rect 19521 9327 19579 9333
rect 19702 9324 19708 9376
rect 19760 9364 19766 9376
rect 21836 9364 21864 9460
rect 22066 9432 22094 9472
rect 22281 9469 22293 9503
rect 22327 9469 22339 9503
rect 22281 9463 22339 9469
rect 22296 9432 22324 9463
rect 22554 9460 22560 9512
rect 22612 9500 22618 9512
rect 23400 9500 23428 9540
rect 24118 9509 24124 9512
rect 22612 9472 23428 9500
rect 24075 9503 24124 9509
rect 22612 9460 22618 9472
rect 24075 9469 24087 9503
rect 24121 9469 24124 9503
rect 24075 9463 24124 9469
rect 24118 9460 24124 9463
rect 24176 9460 24182 9512
rect 24210 9460 24216 9512
rect 24268 9460 24274 9512
rect 24486 9460 24492 9512
rect 24544 9460 24550 9512
rect 24946 9460 24952 9512
rect 25004 9500 25010 9512
rect 25700 9500 25728 9540
rect 26050 9528 26056 9580
rect 26108 9528 26114 9580
rect 25004 9472 25728 9500
rect 25004 9460 25010 9472
rect 22066 9404 22324 9432
rect 26160 9432 26188 9608
rect 26237 9605 26249 9639
rect 26283 9605 26295 9639
rect 26237 9599 26295 9605
rect 26326 9596 26332 9648
rect 26384 9596 26390 9648
rect 26436 9636 26464 9676
rect 27264 9676 28488 9704
rect 27264 9636 27292 9676
rect 26436 9608 27292 9636
rect 27341 9639 27399 9645
rect 27341 9605 27353 9639
rect 27387 9636 27399 9639
rect 28353 9639 28411 9645
rect 28353 9636 28365 9639
rect 27387 9608 28365 9636
rect 27387 9605 27399 9608
rect 27341 9599 27399 9605
rect 28353 9605 28365 9608
rect 28399 9605 28411 9639
rect 28460 9636 28488 9676
rect 31478 9664 31484 9716
rect 31536 9704 31542 9716
rect 33134 9704 33140 9716
rect 31536 9676 33140 9704
rect 31536 9664 31542 9676
rect 33134 9664 33140 9676
rect 33192 9664 33198 9716
rect 33594 9664 33600 9716
rect 33652 9704 33658 9716
rect 35161 9707 35219 9713
rect 33652 9676 34100 9704
rect 33652 9664 33658 9676
rect 30374 9636 30380 9648
rect 28460 9608 30380 9636
rect 28353 9599 28411 9605
rect 30374 9596 30380 9608
rect 30432 9596 30438 9648
rect 31389 9639 31447 9645
rect 31389 9605 31401 9639
rect 31435 9636 31447 9639
rect 31570 9636 31576 9648
rect 31435 9608 31576 9636
rect 31435 9605 31447 9608
rect 31389 9599 31447 9605
rect 31570 9596 31576 9608
rect 31628 9636 31634 9648
rect 32493 9639 32551 9645
rect 31628 9608 32352 9636
rect 31628 9596 31634 9608
rect 26421 9571 26479 9577
rect 26421 9537 26433 9571
rect 26467 9537 26479 9571
rect 26421 9531 26479 9537
rect 27065 9571 27123 9577
rect 27065 9537 27077 9571
rect 27111 9568 27123 9571
rect 27154 9568 27160 9580
rect 27111 9540 27160 9568
rect 27111 9537 27123 9540
rect 27065 9531 27123 9537
rect 26436 9500 26464 9531
rect 27154 9528 27160 9540
rect 27212 9528 27218 9580
rect 27246 9528 27252 9580
rect 27304 9528 27310 9580
rect 27433 9571 27491 9577
rect 27433 9537 27445 9571
rect 27479 9568 27491 9571
rect 30098 9568 30104 9580
rect 27479 9540 30104 9568
rect 27479 9537 27491 9540
rect 27433 9531 27491 9537
rect 27448 9500 27476 9531
rect 28368 9512 28396 9540
rect 30098 9528 30104 9540
rect 30156 9528 30162 9580
rect 31297 9571 31355 9577
rect 31297 9537 31309 9571
rect 31343 9537 31355 9571
rect 31297 9531 31355 9537
rect 31481 9571 31539 9577
rect 31481 9537 31493 9571
rect 31527 9568 31539 9571
rect 31846 9568 31852 9580
rect 31527 9540 31852 9568
rect 31527 9537 31539 9540
rect 31481 9531 31539 9537
rect 27522 9500 27528 9512
rect 26436 9472 27528 9500
rect 27522 9460 27528 9472
rect 27580 9460 27586 9512
rect 27801 9503 27859 9509
rect 27801 9469 27813 9503
rect 27847 9500 27859 9503
rect 27847 9472 27936 9500
rect 27847 9469 27859 9472
rect 27801 9463 27859 9469
rect 26605 9435 26663 9441
rect 26605 9432 26617 9435
rect 26160 9404 26617 9432
rect 26605 9401 26617 9404
rect 26651 9401 26663 9435
rect 26605 9395 26663 9401
rect 27338 9392 27344 9444
rect 27396 9432 27402 9444
rect 27908 9432 27936 9472
rect 28350 9460 28356 9512
rect 28408 9460 28414 9512
rect 29638 9460 29644 9512
rect 29696 9500 29702 9512
rect 31312 9500 31340 9531
rect 31846 9528 31852 9540
rect 31904 9528 31910 9580
rect 32324 9577 32352 9608
rect 32493 9605 32505 9639
rect 32539 9636 32551 9639
rect 33502 9636 33508 9648
rect 32539 9608 33508 9636
rect 32539 9605 32551 9608
rect 32493 9599 32551 9605
rect 33502 9596 33508 9608
rect 33560 9596 33566 9648
rect 33962 9596 33968 9648
rect 34020 9596 34026 9648
rect 32125 9571 32183 9577
rect 32125 9537 32137 9571
rect 32171 9537 32183 9571
rect 32125 9531 32183 9537
rect 32309 9571 32367 9577
rect 32309 9537 32321 9571
rect 32355 9537 32367 9571
rect 32309 9531 32367 9537
rect 31386 9500 31392 9512
rect 29696 9472 31392 9500
rect 29696 9460 29702 9472
rect 31386 9460 31392 9472
rect 31444 9460 31450 9512
rect 27396 9404 27936 9432
rect 27396 9392 27402 9404
rect 27908 9376 27936 9404
rect 19760 9336 21864 9364
rect 19760 9324 19766 9336
rect 27614 9324 27620 9376
rect 27672 9324 27678 9376
rect 27890 9324 27896 9376
rect 27948 9324 27954 9376
rect 32030 9324 32036 9376
rect 32088 9364 32094 9376
rect 32146 9364 32174 9531
rect 33410 9528 33416 9580
rect 33468 9568 33474 9580
rect 33597 9571 33655 9577
rect 33597 9568 33609 9571
rect 33468 9540 33609 9568
rect 33468 9528 33474 9540
rect 33597 9537 33609 9540
rect 33643 9537 33655 9571
rect 33597 9531 33655 9537
rect 33781 9571 33839 9577
rect 33781 9537 33793 9571
rect 33827 9537 33839 9571
rect 33781 9531 33839 9537
rect 32766 9460 32772 9512
rect 32824 9500 32830 9512
rect 33796 9500 33824 9531
rect 33870 9528 33876 9580
rect 33928 9528 33934 9580
rect 34072 9574 34100 9676
rect 35161 9673 35173 9707
rect 35207 9704 35219 9707
rect 35207 9676 35756 9704
rect 35207 9673 35219 9676
rect 35161 9667 35219 9673
rect 35728 9648 35756 9676
rect 34238 9596 34244 9648
rect 34296 9636 34302 9648
rect 34514 9636 34520 9648
rect 34296 9608 34520 9636
rect 34296 9596 34302 9608
rect 34514 9596 34520 9608
rect 34572 9596 34578 9648
rect 35621 9639 35679 9645
rect 35621 9636 35633 9639
rect 34624 9608 35633 9636
rect 34149 9574 34207 9577
rect 34072 9571 34207 9574
rect 34072 9546 34161 9571
rect 34149 9537 34161 9546
rect 34195 9537 34207 9571
rect 34149 9531 34207 9537
rect 34422 9528 34428 9580
rect 34480 9528 34486 9580
rect 34624 9577 34652 9608
rect 35621 9605 35633 9608
rect 35667 9605 35679 9639
rect 35621 9599 35679 9605
rect 35710 9596 35716 9648
rect 35768 9596 35774 9648
rect 38930 9596 38936 9648
rect 38988 9636 38994 9648
rect 39025 9639 39083 9645
rect 39025 9636 39037 9639
rect 38988 9608 39037 9636
rect 38988 9596 38994 9608
rect 39025 9605 39037 9608
rect 39071 9605 39083 9639
rect 39025 9599 39083 9605
rect 39393 9639 39451 9645
rect 39393 9605 39405 9639
rect 39439 9636 39451 9639
rect 39574 9636 39580 9648
rect 39439 9608 39580 9636
rect 39439 9605 39451 9608
rect 39393 9599 39451 9605
rect 39574 9596 39580 9608
rect 39632 9596 39638 9648
rect 34609 9571 34667 9577
rect 34609 9537 34621 9571
rect 34655 9537 34667 9571
rect 34609 9531 34667 9537
rect 35069 9571 35127 9577
rect 35069 9537 35081 9571
rect 35115 9568 35127 9571
rect 35529 9571 35587 9577
rect 35529 9568 35541 9571
rect 35115 9540 35541 9568
rect 35115 9537 35127 9540
rect 35069 9531 35127 9537
rect 35529 9537 35541 9540
rect 35575 9568 35587 9571
rect 35575 9540 36032 9568
rect 35575 9537 35587 9540
rect 35529 9531 35587 9537
rect 32824 9472 33824 9500
rect 34333 9503 34391 9509
rect 32824 9460 32830 9472
rect 34333 9469 34345 9503
rect 34379 9469 34391 9503
rect 34333 9463 34391 9469
rect 32306 9392 32312 9444
rect 32364 9432 32370 9444
rect 33502 9432 33508 9444
rect 32364 9404 33508 9432
rect 32364 9392 32370 9404
rect 33502 9392 33508 9404
rect 33560 9392 33566 9444
rect 33597 9435 33655 9441
rect 33597 9401 33609 9435
rect 33643 9432 33655 9435
rect 33962 9432 33968 9444
rect 33643 9404 33968 9432
rect 33643 9401 33655 9404
rect 33597 9395 33655 9401
rect 33962 9392 33968 9404
rect 34020 9392 34026 9444
rect 34238 9432 34244 9444
rect 34072 9404 34244 9432
rect 34072 9364 34100 9404
rect 34238 9392 34244 9404
rect 34296 9392 34302 9444
rect 34348 9432 34376 9463
rect 35250 9460 35256 9512
rect 35308 9460 35314 9512
rect 35342 9460 35348 9512
rect 35400 9500 35406 9512
rect 35437 9503 35495 9509
rect 35437 9500 35449 9503
rect 35400 9472 35449 9500
rect 35400 9460 35406 9472
rect 35437 9469 35449 9472
rect 35483 9469 35495 9503
rect 35437 9463 35495 9469
rect 34606 9432 34612 9444
rect 34348 9404 34612 9432
rect 34606 9392 34612 9404
rect 34664 9392 34670 9444
rect 36004 9376 36032 9540
rect 32088 9336 34100 9364
rect 32088 9324 32094 9336
rect 34790 9324 34796 9376
rect 34848 9364 34854 9376
rect 35345 9367 35403 9373
rect 35345 9364 35357 9367
rect 34848 9336 35357 9364
rect 34848 9324 34854 9336
rect 35345 9333 35357 9336
rect 35391 9333 35403 9367
rect 35345 9327 35403 9333
rect 35986 9324 35992 9376
rect 36044 9324 36050 9376
rect 1104 9274 41400 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 41400 9274
rect 1104 9200 41400 9222
rect 4420 9163 4478 9169
rect 4420 9129 4432 9163
rect 4466 9160 4478 9163
rect 6178 9160 6184 9172
rect 4466 9132 6184 9160
rect 4466 9129 4478 9132
rect 4420 9123 4478 9129
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 6546 9120 6552 9172
rect 6604 9120 6610 9172
rect 6825 9163 6883 9169
rect 6825 9129 6837 9163
rect 6871 9160 6883 9163
rect 6914 9160 6920 9172
rect 6871 9132 6920 9160
rect 6871 9129 6883 9132
rect 6825 9123 6883 9129
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 7377 9163 7435 9169
rect 7377 9129 7389 9163
rect 7423 9160 7435 9163
rect 7650 9160 7656 9172
rect 7423 9132 7656 9160
rect 7423 9129 7435 9132
rect 7377 9123 7435 9129
rect 7650 9120 7656 9132
rect 7708 9120 7714 9172
rect 8018 9120 8024 9172
rect 8076 9120 8082 9172
rect 9493 9163 9551 9169
rect 9493 9160 9505 9163
rect 8128 9132 9505 9160
rect 5442 9052 5448 9104
rect 5500 9092 5506 9104
rect 5905 9095 5963 9101
rect 5905 9092 5917 9095
rect 5500 9064 5917 9092
rect 5500 9052 5506 9064
rect 5905 9061 5917 9064
rect 5951 9061 5963 9095
rect 5905 9055 5963 9061
rect 7190 9052 7196 9104
rect 7248 9092 7254 9104
rect 8128 9092 8156 9132
rect 9493 9129 9505 9132
rect 9539 9129 9551 9163
rect 9493 9123 9551 9129
rect 9582 9120 9588 9172
rect 9640 9120 9646 9172
rect 11606 9120 11612 9172
rect 11664 9160 11670 9172
rect 11701 9163 11759 9169
rect 11701 9160 11713 9163
rect 11664 9132 11713 9160
rect 11664 9120 11670 9132
rect 11701 9129 11713 9132
rect 11747 9129 11759 9163
rect 11701 9123 11759 9129
rect 12250 9120 12256 9172
rect 12308 9120 12314 9172
rect 13170 9120 13176 9172
rect 13228 9120 13234 9172
rect 13814 9120 13820 9172
rect 13872 9160 13878 9172
rect 16482 9160 16488 9172
rect 13872 9132 16488 9160
rect 13872 9120 13878 9132
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 16574 9120 16580 9172
rect 16632 9120 16638 9172
rect 16850 9120 16856 9172
rect 16908 9120 16914 9172
rect 19150 9120 19156 9172
rect 19208 9120 19214 9172
rect 20806 9120 20812 9172
rect 20864 9120 20870 9172
rect 21818 9120 21824 9172
rect 21876 9120 21882 9172
rect 24486 9120 24492 9172
rect 24544 9160 24550 9172
rect 24857 9163 24915 9169
rect 24857 9160 24869 9163
rect 24544 9132 24869 9160
rect 24544 9120 24550 9132
rect 24857 9129 24869 9132
rect 24903 9129 24915 9163
rect 26418 9160 26424 9172
rect 24857 9123 24915 9129
rect 25056 9132 26424 9160
rect 9600 9092 9628 9120
rect 7248 9064 8156 9092
rect 8956 9064 9628 9092
rect 7248 9052 7254 9064
rect 6638 9024 6644 9036
rect 4172 8996 6644 9024
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 4172 8965 4200 8996
rect 6638 8984 6644 8996
rect 6696 8984 6702 9036
rect 7024 8996 8248 9024
rect 7024 8965 7052 8996
rect 4157 8959 4215 8965
rect 4157 8956 4169 8959
rect 4120 8928 4169 8956
rect 4120 8916 4126 8928
rect 4157 8925 4169 8928
rect 4203 8925 4215 8959
rect 6733 8959 6791 8965
rect 5566 8928 6592 8956
rect 4157 8919 4215 8925
rect 6564 8900 6592 8928
rect 6733 8925 6745 8959
rect 6779 8956 6791 8959
rect 7009 8959 7067 8965
rect 7009 8956 7021 8959
rect 6779 8928 7021 8956
rect 6779 8925 6791 8928
rect 6733 8919 6791 8925
rect 7009 8925 7021 8928
rect 7055 8925 7067 8959
rect 7009 8919 7067 8925
rect 7098 8916 7104 8968
rect 7156 8956 7162 8968
rect 7576 8965 7604 8996
rect 8220 8968 8248 8996
rect 7285 8959 7343 8965
rect 7285 8956 7297 8959
rect 7156 8928 7297 8956
rect 7156 8916 7162 8928
rect 7285 8925 7297 8928
rect 7331 8925 7343 8959
rect 7285 8919 7343 8925
rect 7561 8959 7619 8965
rect 7561 8925 7573 8959
rect 7607 8925 7619 8959
rect 7561 8919 7619 8925
rect 7837 8959 7895 8965
rect 7837 8925 7849 8959
rect 7883 8956 7895 8959
rect 7883 8928 7972 8956
rect 7883 8925 7895 8928
rect 7837 8919 7895 8925
rect 6457 8891 6515 8897
rect 6457 8857 6469 8891
rect 6503 8857 6515 8891
rect 6457 8851 6515 8857
rect 6472 8820 6500 8851
rect 6546 8848 6552 8900
rect 6604 8848 6610 8900
rect 7944 8897 7972 8928
rect 8202 8916 8208 8968
rect 8260 8916 8266 8968
rect 8956 8965 8984 9064
rect 11514 9052 11520 9104
rect 11572 9052 11578 9104
rect 9953 9027 10011 9033
rect 9953 9024 9965 9027
rect 9140 8996 9965 9024
rect 9140 8965 9168 8996
rect 9953 8993 9965 8996
rect 9999 8993 10011 9027
rect 9953 8987 10011 8993
rect 11238 8984 11244 9036
rect 11296 8984 11302 9036
rect 11885 9027 11943 9033
rect 11885 8993 11897 9027
rect 11931 9024 11943 9027
rect 12268 9024 12296 9120
rect 11931 8996 12296 9024
rect 13188 9024 13216 9120
rect 13538 9052 13544 9104
rect 13596 9092 13602 9104
rect 14921 9095 14979 9101
rect 14921 9092 14933 9095
rect 13596 9064 14933 9092
rect 13596 9052 13602 9064
rect 14921 9061 14933 9064
rect 14967 9061 14979 9095
rect 14921 9055 14979 9061
rect 15194 9052 15200 9104
rect 15252 9092 15258 9104
rect 16114 9092 16120 9104
rect 15252 9064 16120 9092
rect 15252 9052 15258 9064
rect 16114 9052 16120 9064
rect 16172 9052 16178 9104
rect 15841 9027 15899 9033
rect 13188 8996 14596 9024
rect 11931 8993 11943 8996
rect 11885 8987 11943 8993
rect 8941 8959 8999 8965
rect 8941 8925 8953 8959
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 6641 8891 6699 8897
rect 6641 8857 6653 8891
rect 6687 8888 6699 8891
rect 7193 8891 7251 8897
rect 7193 8888 7205 8891
rect 6687 8860 7205 8888
rect 6687 8857 6699 8860
rect 6641 8851 6699 8857
rect 7193 8857 7205 8860
rect 7239 8888 7251 8891
rect 7929 8891 7987 8897
rect 7239 8860 7788 8888
rect 7239 8857 7251 8860
rect 7193 8851 7251 8857
rect 7098 8820 7104 8832
rect 6472 8792 7104 8820
rect 7098 8780 7104 8792
rect 7156 8820 7162 8832
rect 7650 8820 7656 8832
rect 7156 8792 7656 8820
rect 7156 8780 7162 8792
rect 7650 8780 7656 8792
rect 7708 8780 7714 8832
rect 7760 8829 7788 8860
rect 7929 8857 7941 8891
rect 7975 8888 7987 8891
rect 8018 8888 8024 8900
rect 7975 8860 8024 8888
rect 7975 8857 7987 8860
rect 7929 8851 7987 8857
rect 8018 8848 8024 8860
rect 8076 8848 8082 8900
rect 8113 8891 8171 8897
rect 8113 8857 8125 8891
rect 8159 8888 8171 8891
rect 9232 8888 9260 8919
rect 9306 8916 9312 8968
rect 9364 8916 9370 8968
rect 9766 8916 9772 8968
rect 9824 8916 9830 8968
rect 9858 8916 9864 8968
rect 9916 8916 9922 8968
rect 11054 8916 11060 8968
rect 11112 8956 11118 8968
rect 11149 8959 11207 8965
rect 11149 8956 11161 8959
rect 11112 8928 11161 8956
rect 11112 8916 11118 8928
rect 11149 8925 11161 8928
rect 11195 8956 11207 8959
rect 11422 8956 11428 8968
rect 11195 8928 11428 8956
rect 11195 8925 11207 8928
rect 11149 8919 11207 8925
rect 11422 8916 11428 8928
rect 11480 8916 11486 8968
rect 11514 8916 11520 8968
rect 11572 8956 11578 8968
rect 11609 8959 11667 8965
rect 11609 8956 11621 8959
rect 11572 8928 11621 8956
rect 11572 8916 11578 8928
rect 11609 8925 11621 8928
rect 11655 8925 11667 8959
rect 11609 8919 11667 8925
rect 11790 8916 11796 8968
rect 11848 8956 11854 8968
rect 11848 8928 11928 8956
rect 11848 8916 11854 8928
rect 8159 8860 9352 8888
rect 8159 8857 8171 8860
rect 8113 8851 8171 8857
rect 7745 8823 7803 8829
rect 7745 8789 7757 8823
rect 7791 8820 7803 8823
rect 8128 8820 8156 8851
rect 8956 8832 8984 8860
rect 7791 8792 8156 8820
rect 7791 8789 7803 8792
rect 7745 8783 7803 8789
rect 8938 8780 8944 8832
rect 8996 8780 9002 8832
rect 9324 8820 9352 8860
rect 9490 8848 9496 8900
rect 9548 8888 9554 8900
rect 9585 8891 9643 8897
rect 9585 8888 9597 8891
rect 9548 8860 9597 8888
rect 9548 8848 9554 8860
rect 9585 8857 9597 8860
rect 9631 8857 9643 8891
rect 9585 8851 9643 8857
rect 9876 8820 9904 8916
rect 11330 8848 11336 8900
rect 11388 8848 11394 8900
rect 11900 8897 11928 8928
rect 11974 8916 11980 8968
rect 12032 8916 12038 8968
rect 12066 8916 12072 8968
rect 12124 8916 12130 8968
rect 12158 8916 12164 8968
rect 12216 8916 12222 8968
rect 13998 8916 14004 8968
rect 14056 8956 14062 8968
rect 14568 8965 14596 8996
rect 14660 8996 15516 9024
rect 14369 8959 14427 8965
rect 14369 8956 14381 8959
rect 14056 8928 14381 8956
rect 14056 8916 14062 8928
rect 14369 8925 14381 8928
rect 14415 8925 14427 8959
rect 14369 8919 14427 8925
rect 14461 8959 14519 8965
rect 14461 8925 14473 8959
rect 14507 8925 14519 8959
rect 14461 8919 14519 8925
rect 14553 8959 14611 8965
rect 14553 8925 14565 8959
rect 14599 8925 14611 8959
rect 14553 8919 14611 8925
rect 11885 8891 11943 8897
rect 11885 8857 11897 8891
rect 11931 8857 11943 8891
rect 14476 8888 14504 8919
rect 14660 8888 14688 8996
rect 14737 8959 14795 8965
rect 14737 8925 14749 8959
rect 14783 8925 14795 8959
rect 14737 8919 14795 8925
rect 15013 8959 15071 8965
rect 15013 8925 15025 8959
rect 15059 8925 15071 8959
rect 15013 8919 15071 8925
rect 11885 8851 11943 8857
rect 12406 8860 14688 8888
rect 9324 8792 9904 8820
rect 11348 8820 11376 8848
rect 12406 8820 12434 8860
rect 11348 8792 12434 8820
rect 14090 8780 14096 8832
rect 14148 8780 14154 8832
rect 14752 8820 14780 8919
rect 15028 8888 15056 8919
rect 15286 8916 15292 8968
rect 15344 8956 15350 8968
rect 15381 8959 15439 8965
rect 15381 8956 15393 8959
rect 15344 8928 15393 8956
rect 15344 8916 15350 8928
rect 15381 8925 15393 8928
rect 15427 8925 15439 8959
rect 15488 8956 15516 8996
rect 15841 8993 15853 9027
rect 15887 9024 15899 9027
rect 16022 9024 16028 9036
rect 15887 8996 16028 9024
rect 15887 8993 15899 8996
rect 15841 8987 15899 8993
rect 16022 8984 16028 8996
rect 16080 8984 16086 9036
rect 16592 9024 16620 9120
rect 16132 8996 16620 9024
rect 16132 8965 16160 8996
rect 16117 8959 16175 8965
rect 16117 8956 16129 8959
rect 15488 8928 16129 8956
rect 15381 8919 15439 8925
rect 16117 8925 16129 8928
rect 16163 8925 16175 8959
rect 16117 8919 16175 8925
rect 16206 8916 16212 8968
rect 16264 8916 16270 8968
rect 16301 8959 16359 8965
rect 16301 8925 16313 8959
rect 16347 8956 16359 8959
rect 16868 8956 16896 9120
rect 19168 9092 19196 9120
rect 21177 9095 21235 9101
rect 21177 9092 21189 9095
rect 19168 9064 21189 9092
rect 21177 9061 21189 9064
rect 21223 9092 21235 9095
rect 21266 9092 21272 9104
rect 21223 9064 21272 9092
rect 21223 9061 21235 9064
rect 21177 9055 21235 9061
rect 21266 9052 21272 9064
rect 21324 9052 21330 9104
rect 17313 9027 17371 9033
rect 17313 8993 17325 9027
rect 17359 9024 17371 9027
rect 19334 9024 19340 9036
rect 17359 8996 19340 9024
rect 17359 8993 17371 8996
rect 17313 8987 17371 8993
rect 19334 8984 19340 8996
rect 19392 9024 19398 9036
rect 19702 9024 19708 9036
rect 19392 8996 19708 9024
rect 19392 8984 19398 8996
rect 19702 8984 19708 8996
rect 19760 8984 19766 9036
rect 20901 9027 20959 9033
rect 20901 8993 20913 9027
rect 20947 9024 20959 9027
rect 20990 9024 20996 9036
rect 20947 8996 20996 9024
rect 20947 8993 20959 8996
rect 20901 8987 20959 8993
rect 20990 8984 20996 8996
rect 21048 8984 21054 9036
rect 21729 9027 21787 9033
rect 21729 8993 21741 9027
rect 21775 9024 21787 9027
rect 21836 9024 21864 9120
rect 21775 8996 21864 9024
rect 22005 9027 22063 9033
rect 21775 8993 21787 8996
rect 21729 8987 21787 8993
rect 22005 8993 22017 9027
rect 22051 9024 22063 9027
rect 22094 9024 22100 9036
rect 22051 8996 22100 9024
rect 22051 8993 22063 8996
rect 22005 8987 22063 8993
rect 22094 8984 22100 8996
rect 22152 8984 22158 9036
rect 23750 8984 23756 9036
rect 23808 8984 23814 9036
rect 18966 8956 18972 8968
rect 16347 8928 16896 8956
rect 18722 8928 18972 8956
rect 16347 8925 16359 8928
rect 16301 8919 16359 8925
rect 16316 8888 16344 8919
rect 18966 8916 18972 8928
rect 19024 8916 19030 8968
rect 19058 8916 19064 8968
rect 19116 8956 19122 8968
rect 25056 8965 25084 9132
rect 26418 9120 26424 9132
rect 26476 9120 26482 9172
rect 27614 9120 27620 9172
rect 27672 9120 27678 9172
rect 27801 9163 27859 9169
rect 27801 9129 27813 9163
rect 27847 9160 27859 9163
rect 27890 9160 27896 9172
rect 27847 9132 27896 9160
rect 27847 9129 27859 9132
rect 27801 9123 27859 9129
rect 27890 9120 27896 9132
rect 27948 9120 27954 9172
rect 30282 9120 30288 9172
rect 30340 9160 30346 9172
rect 30558 9160 30564 9172
rect 30340 9132 30564 9160
rect 30340 9120 30346 9132
rect 30558 9120 30564 9132
rect 30616 9120 30622 9172
rect 30653 9163 30711 9169
rect 30653 9129 30665 9163
rect 30699 9160 30711 9163
rect 32674 9160 32680 9172
rect 30699 9132 32680 9160
rect 30699 9129 30711 9132
rect 30653 9123 30711 9129
rect 32674 9120 32680 9132
rect 32732 9120 32738 9172
rect 33410 9120 33416 9172
rect 33468 9120 33474 9172
rect 33502 9120 33508 9172
rect 33560 9120 33566 9172
rect 33965 9163 34023 9169
rect 33965 9129 33977 9163
rect 34011 9160 34023 9163
rect 34422 9160 34428 9172
rect 34011 9132 34428 9160
rect 34011 9129 34023 9132
rect 33965 9123 34023 9129
rect 34422 9120 34428 9132
rect 34480 9120 34486 9172
rect 35986 9120 35992 9172
rect 36044 9120 36050 9172
rect 37458 9120 37464 9172
rect 37516 9120 37522 9172
rect 25222 8984 25228 9036
rect 25280 9024 25286 9036
rect 26053 9027 26111 9033
rect 26053 9024 26065 9027
rect 25280 8996 26065 9024
rect 25280 8984 25286 8996
rect 26053 8993 26065 8996
rect 26099 8993 26111 9027
rect 26053 8987 26111 8993
rect 26329 9027 26387 9033
rect 26329 8993 26341 9027
rect 26375 9024 26387 9027
rect 27632 9024 27660 9120
rect 28074 9052 28080 9104
rect 28132 9052 28138 9104
rect 28184 9064 28994 9092
rect 28184 9024 28212 9064
rect 26375 8996 27660 9024
rect 28092 8996 28212 9024
rect 26375 8993 26387 8996
rect 26329 8987 26387 8993
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 19116 8928 19441 8956
rect 19116 8916 19122 8928
rect 19429 8925 19441 8928
rect 19475 8925 19487 8959
rect 19429 8919 19487 8925
rect 20809 8959 20867 8965
rect 20809 8925 20821 8959
rect 20855 8925 20867 8959
rect 20809 8919 20867 8925
rect 25041 8959 25099 8965
rect 25041 8925 25053 8959
rect 25087 8925 25099 8959
rect 25041 8919 25099 8925
rect 15028 8860 16344 8888
rect 17586 8848 17592 8900
rect 17644 8848 17650 8900
rect 20824 8888 20852 8919
rect 21910 8888 21916 8900
rect 18892 8860 20208 8888
rect 20824 8860 21916 8888
rect 14826 8820 14832 8832
rect 14752 8792 14832 8820
rect 14826 8780 14832 8792
rect 14884 8820 14890 8832
rect 18892 8820 18920 8860
rect 14884 8792 18920 8820
rect 14884 8780 14890 8792
rect 18966 8780 18972 8832
rect 19024 8820 19030 8832
rect 19061 8823 19119 8829
rect 19061 8820 19073 8823
rect 19024 8792 19073 8820
rect 19024 8780 19030 8792
rect 19061 8789 19073 8792
rect 19107 8789 19119 8823
rect 19061 8783 19119 8789
rect 19242 8780 19248 8832
rect 19300 8820 19306 8832
rect 20073 8823 20131 8829
rect 20073 8820 20085 8823
rect 19300 8792 20085 8820
rect 19300 8780 19306 8792
rect 20073 8789 20085 8792
rect 20119 8789 20131 8823
rect 20180 8820 20208 8860
rect 21910 8848 21916 8860
rect 21968 8888 21974 8900
rect 22094 8888 22100 8900
rect 21968 8860 22100 8888
rect 21968 8848 21974 8860
rect 22094 8848 22100 8860
rect 22152 8848 22158 8900
rect 22554 8848 22560 8900
rect 22612 8848 22618 8900
rect 27338 8848 27344 8900
rect 27396 8848 27402 8900
rect 28092 8897 28120 8996
rect 28258 8984 28264 9036
rect 28316 9024 28322 9036
rect 28629 9027 28687 9033
rect 28629 9024 28641 9027
rect 28316 8996 28641 9024
rect 28316 8984 28322 8996
rect 28629 8993 28641 8996
rect 28675 8993 28687 9027
rect 28966 9024 28994 9064
rect 29546 9052 29552 9104
rect 29604 9092 29610 9104
rect 31662 9092 31668 9104
rect 29604 9064 30236 9092
rect 29604 9052 29610 9064
rect 28966 8996 29684 9024
rect 28629 8987 28687 8993
rect 29656 8965 29684 8996
rect 28813 8959 28871 8965
rect 28813 8956 28825 8959
rect 28184 8928 28825 8956
rect 28077 8891 28135 8897
rect 28077 8857 28089 8891
rect 28123 8857 28135 8891
rect 28077 8851 28135 8857
rect 21082 8820 21088 8832
rect 20180 8792 21088 8820
rect 20073 8783 20131 8789
rect 21082 8780 21088 8792
rect 21140 8780 21146 8832
rect 27246 8780 27252 8832
rect 27304 8820 27310 8832
rect 28184 8820 28212 8928
rect 28813 8925 28825 8928
rect 28859 8925 28871 8959
rect 28813 8919 28871 8925
rect 29549 8959 29607 8965
rect 29549 8925 29561 8959
rect 29595 8925 29607 8959
rect 29549 8919 29607 8925
rect 29641 8959 29699 8965
rect 29641 8925 29653 8959
rect 29687 8956 29699 8959
rect 29730 8956 29736 8968
rect 29687 8928 29736 8956
rect 29687 8925 29699 8928
rect 29641 8919 29699 8925
rect 28534 8848 28540 8900
rect 28592 8848 28598 8900
rect 29564 8888 29592 8919
rect 29730 8916 29736 8928
rect 29788 8916 29794 8968
rect 29914 8916 29920 8968
rect 29972 8916 29978 8968
rect 30024 8965 30052 9064
rect 30208 9036 30236 9064
rect 31496 9064 31668 9092
rect 30098 8984 30104 9036
rect 30156 8984 30162 9036
rect 30190 8984 30196 9036
rect 30248 8984 30254 9036
rect 30466 8984 30472 9036
rect 30524 9024 30530 9036
rect 31496 9033 31524 9064
rect 31662 9052 31668 9064
rect 31720 9052 31726 9104
rect 31849 9095 31907 9101
rect 31849 9061 31861 9095
rect 31895 9092 31907 9095
rect 33428 9092 33456 9120
rect 33873 9095 33931 9101
rect 33873 9092 33885 9095
rect 31895 9064 32260 9092
rect 33428 9064 33885 9092
rect 31895 9061 31907 9064
rect 31849 9055 31907 9061
rect 31481 9027 31539 9033
rect 30524 8996 30880 9024
rect 30524 8984 30530 8996
rect 30852 8965 30880 8996
rect 31481 8993 31493 9027
rect 31527 8993 31539 9027
rect 31481 8987 31539 8993
rect 30009 8959 30067 8965
rect 30009 8925 30021 8959
rect 30055 8925 30067 8959
rect 30653 8959 30711 8965
rect 30653 8956 30665 8959
rect 30009 8919 30067 8925
rect 30208 8928 30665 8956
rect 30208 8900 30236 8928
rect 30653 8925 30665 8928
rect 30699 8925 30711 8959
rect 30653 8919 30711 8925
rect 30837 8959 30895 8965
rect 30837 8925 30849 8959
rect 30883 8925 30895 8959
rect 30837 8919 30895 8925
rect 31846 8916 31852 8968
rect 31904 8916 31910 8968
rect 32030 8916 32036 8968
rect 32088 8956 32094 8968
rect 32125 8959 32183 8965
rect 32125 8956 32137 8959
rect 32088 8928 32137 8956
rect 32088 8916 32094 8928
rect 32125 8925 32137 8928
rect 32171 8925 32183 8959
rect 32125 8919 32183 8925
rect 28644 8860 29592 8888
rect 29825 8891 29883 8897
rect 28644 8832 28672 8860
rect 29825 8857 29837 8891
rect 29871 8857 29883 8891
rect 29825 8851 29883 8857
rect 27304 8792 28212 8820
rect 27304 8780 27310 8792
rect 28626 8780 28632 8832
rect 28684 8780 28690 8832
rect 29840 8820 29868 8851
rect 30190 8848 30196 8900
rect 30248 8848 30254 8900
rect 30282 8848 30288 8900
rect 30340 8848 30346 8900
rect 30377 8891 30435 8897
rect 30377 8857 30389 8891
rect 30423 8888 30435 8891
rect 30466 8888 30472 8900
rect 30423 8860 30472 8888
rect 30423 8857 30435 8860
rect 30377 8851 30435 8857
rect 30466 8848 30472 8860
rect 30524 8848 30530 8900
rect 30300 8820 30328 8848
rect 29840 8792 30328 8820
rect 31864 8820 31892 8916
rect 32232 8832 32260 9064
rect 33873 9061 33885 9064
rect 33919 9092 33931 9095
rect 34054 9092 34060 9104
rect 33919 9064 34060 9092
rect 33919 9061 33931 9064
rect 33873 9055 33931 9061
rect 34054 9052 34060 9064
rect 34112 9052 34118 9104
rect 34330 9052 34336 9104
rect 34388 9052 34394 9104
rect 34238 9024 34244 9036
rect 33520 8996 34244 9024
rect 32306 8916 32312 8968
rect 32364 8916 32370 8968
rect 33042 8916 33048 8968
rect 33100 8916 33106 8968
rect 33520 8965 33548 8996
rect 34238 8984 34244 8996
rect 34296 8984 34302 9036
rect 34348 9024 34376 9052
rect 34348 8996 35848 9024
rect 33505 8959 33563 8965
rect 33505 8925 33517 8959
rect 33551 8925 33563 8959
rect 33505 8919 33563 8925
rect 33597 8959 33655 8965
rect 33597 8925 33609 8959
rect 33643 8925 33655 8959
rect 33597 8919 33655 8925
rect 33060 8888 33088 8916
rect 33612 8888 33640 8919
rect 33686 8916 33692 8968
rect 33744 8956 33750 8968
rect 34149 8959 34207 8965
rect 34149 8956 34161 8959
rect 33744 8928 34161 8956
rect 33744 8916 33750 8928
rect 34149 8925 34161 8928
rect 34195 8925 34207 8959
rect 34149 8919 34207 8925
rect 33778 8888 33784 8900
rect 33060 8860 33784 8888
rect 33778 8848 33784 8860
rect 33836 8848 33842 8900
rect 34348 8888 34376 8996
rect 35820 8968 35848 8996
rect 37366 8984 37372 9036
rect 37424 9024 37430 9036
rect 37424 8996 37780 9024
rect 37424 8984 37430 8996
rect 34425 8959 34483 8965
rect 34425 8925 34437 8959
rect 34471 8956 34483 8959
rect 34606 8956 34612 8968
rect 34471 8928 34612 8956
rect 34471 8925 34483 8928
rect 34425 8919 34483 8925
rect 34606 8916 34612 8928
rect 34664 8916 34670 8968
rect 35802 8916 35808 8968
rect 35860 8916 35866 8968
rect 37752 8965 37780 8996
rect 37645 8959 37703 8965
rect 37645 8925 37657 8959
rect 37691 8925 37703 8959
rect 37645 8919 37703 8925
rect 37737 8959 37795 8965
rect 37737 8925 37749 8959
rect 37783 8925 37795 8959
rect 37737 8919 37795 8925
rect 35621 8891 35679 8897
rect 35621 8888 35633 8891
rect 33888 8860 34376 8888
rect 34440 8860 35633 8888
rect 31941 8823 31999 8829
rect 31941 8820 31953 8823
rect 31864 8792 31953 8820
rect 31941 8789 31953 8792
rect 31987 8789 31999 8823
rect 31941 8783 31999 8789
rect 32214 8780 32220 8832
rect 32272 8780 32278 8832
rect 33686 8780 33692 8832
rect 33744 8820 33750 8832
rect 33888 8820 33916 8860
rect 34440 8832 34468 8860
rect 35621 8857 35633 8860
rect 35667 8888 35679 8891
rect 35986 8888 35992 8900
rect 35667 8860 35992 8888
rect 35667 8857 35679 8860
rect 35621 8851 35679 8857
rect 35986 8848 35992 8860
rect 36044 8848 36050 8900
rect 37660 8888 37688 8919
rect 37826 8916 37832 8968
rect 37884 8916 37890 8968
rect 37918 8916 37924 8968
rect 37976 8916 37982 8968
rect 38013 8959 38071 8965
rect 38013 8925 38025 8959
rect 38059 8925 38071 8959
rect 38013 8919 38071 8925
rect 37844 8888 37872 8916
rect 38028 8888 38056 8919
rect 38930 8916 38936 8968
rect 38988 8916 38994 8968
rect 37660 8860 37780 8888
rect 37844 8860 38056 8888
rect 33744 8792 33916 8820
rect 33744 8780 33750 8792
rect 34330 8780 34336 8832
rect 34388 8780 34394 8832
rect 34422 8780 34428 8832
rect 34480 8780 34486 8832
rect 37752 8820 37780 8860
rect 38948 8820 38976 8916
rect 37752 8792 38976 8820
rect 1104 8730 41400 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 41400 8730
rect 1104 8656 41400 8678
rect 8938 8576 8944 8628
rect 8996 8576 9002 8628
rect 9030 8576 9036 8628
rect 9088 8576 9094 8628
rect 11330 8576 11336 8628
rect 11388 8576 11394 8628
rect 11974 8576 11980 8628
rect 12032 8576 12038 8628
rect 12710 8576 12716 8628
rect 12768 8616 12774 8628
rect 13722 8616 13728 8628
rect 12768 8588 13728 8616
rect 12768 8576 12774 8588
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 17586 8576 17592 8628
rect 17644 8576 17650 8628
rect 19242 8576 19248 8628
rect 19300 8576 19306 8628
rect 19426 8576 19432 8628
rect 19484 8576 19490 8628
rect 27154 8576 27160 8628
rect 27212 8616 27218 8628
rect 28537 8619 28595 8625
rect 28537 8616 28549 8619
rect 27212 8588 28549 8616
rect 27212 8576 27218 8588
rect 28537 8585 28549 8588
rect 28583 8616 28595 8619
rect 28626 8616 28632 8628
rect 28583 8588 28632 8616
rect 28583 8585 28595 8588
rect 28537 8579 28595 8585
rect 28626 8576 28632 8588
rect 28684 8576 28690 8628
rect 28718 8576 28724 8628
rect 28776 8616 28782 8628
rect 28905 8619 28963 8625
rect 28905 8616 28917 8619
rect 28776 8588 28917 8616
rect 28776 8576 28782 8588
rect 28905 8585 28917 8588
rect 28951 8616 28963 8619
rect 30466 8616 30472 8628
rect 28951 8588 30472 8616
rect 28951 8585 28963 8588
rect 28905 8579 28963 8585
rect 30466 8576 30472 8588
rect 30524 8576 30530 8628
rect 33413 8619 33471 8625
rect 30576 8588 32444 8616
rect 8849 8483 8907 8489
rect 8849 8449 8861 8483
rect 8895 8449 8907 8483
rect 8956 8480 8984 8576
rect 9048 8548 9076 8576
rect 11348 8548 11376 8576
rect 11992 8548 12020 8576
rect 14366 8548 14372 8560
rect 9048 8520 11928 8548
rect 11992 8520 12296 8548
rect 14214 8520 14372 8548
rect 9033 8483 9091 8489
rect 9033 8480 9045 8483
rect 8956 8452 9045 8480
rect 8849 8443 8907 8449
rect 9033 8449 9045 8452
rect 9079 8449 9091 8483
rect 9033 8443 9091 8449
rect 8864 8412 8892 8443
rect 9122 8440 9128 8492
rect 9180 8440 9186 8492
rect 11514 8480 11520 8492
rect 9646 8452 11520 8480
rect 9217 8415 9275 8421
rect 9217 8412 9229 8415
rect 8864 8384 9229 8412
rect 9217 8381 9229 8384
rect 9263 8381 9275 8415
rect 9646 8412 9674 8452
rect 11514 8440 11520 8452
rect 11572 8440 11578 8492
rect 11606 8440 11612 8492
rect 11664 8480 11670 8492
rect 11900 8489 11928 8520
rect 11793 8483 11851 8489
rect 11793 8480 11805 8483
rect 11664 8452 11805 8480
rect 11664 8440 11670 8452
rect 11793 8449 11805 8452
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8449 11943 8483
rect 11885 8443 11943 8449
rect 11974 8440 11980 8492
rect 12032 8440 12038 8492
rect 12158 8440 12164 8492
rect 12216 8440 12222 8492
rect 12268 8489 12296 8520
rect 14366 8508 14372 8520
rect 14424 8508 14430 8560
rect 16758 8508 16764 8560
rect 16816 8548 16822 8560
rect 17310 8548 17316 8560
rect 16816 8520 17316 8548
rect 16816 8508 16822 8520
rect 17310 8508 17316 8520
rect 17368 8508 17374 8560
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8449 12311 8483
rect 12253 8443 12311 8449
rect 13538 8440 13544 8492
rect 13596 8440 13602 8492
rect 13722 8440 13728 8492
rect 13780 8480 13786 8492
rect 13817 8483 13875 8489
rect 13817 8480 13829 8483
rect 13780 8452 13829 8480
rect 13780 8440 13786 8452
rect 13817 8449 13829 8452
rect 13863 8449 13875 8483
rect 13817 8443 13875 8449
rect 15102 8440 15108 8492
rect 15160 8440 15166 8492
rect 15286 8440 15292 8492
rect 15344 8480 15350 8492
rect 15565 8483 15623 8489
rect 15565 8480 15577 8483
rect 15344 8452 15577 8480
rect 15344 8440 15350 8452
rect 15565 8449 15577 8452
rect 15611 8449 15623 8483
rect 15565 8443 15623 8449
rect 16022 8440 16028 8492
rect 16080 8440 16086 8492
rect 16206 8440 16212 8492
rect 16264 8480 16270 8492
rect 16945 8483 17003 8489
rect 16945 8480 16957 8483
rect 16264 8452 16957 8480
rect 16264 8440 16270 8452
rect 16945 8449 16957 8452
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 9217 8375 9275 8381
rect 9324 8384 9674 8412
rect 7558 8304 7564 8356
rect 7616 8344 7622 8356
rect 9324 8344 9352 8384
rect 9766 8344 9772 8356
rect 7616 8316 9352 8344
rect 9416 8316 9772 8344
rect 7616 8304 7622 8316
rect 6086 8236 6092 8288
rect 6144 8276 6150 8288
rect 8294 8276 8300 8288
rect 6144 8248 8300 8276
rect 6144 8236 6150 8248
rect 8294 8236 8300 8248
rect 8352 8236 8358 8288
rect 8941 8279 8999 8285
rect 8941 8245 8953 8279
rect 8987 8276 8999 8279
rect 9122 8276 9128 8288
rect 8987 8248 9128 8276
rect 8987 8245 8999 8248
rect 8941 8239 8999 8245
rect 9122 8236 9128 8248
rect 9180 8276 9186 8288
rect 9416 8276 9444 8316
rect 9766 8304 9772 8316
rect 9824 8304 9830 8356
rect 11330 8304 11336 8356
rect 11388 8344 11394 8356
rect 11517 8347 11575 8353
rect 11517 8344 11529 8347
rect 11388 8316 11529 8344
rect 11388 8304 11394 8316
rect 11517 8313 11529 8316
rect 11563 8313 11575 8347
rect 12158 8344 12164 8356
rect 11517 8307 11575 8313
rect 11624 8316 12164 8344
rect 9180 8248 9444 8276
rect 9180 8236 9186 8248
rect 11146 8236 11152 8288
rect 11204 8276 11210 8288
rect 11624 8276 11652 8316
rect 12158 8304 12164 8316
rect 12216 8304 12222 8356
rect 15120 8344 15148 8440
rect 16298 8372 16304 8424
rect 16356 8372 16362 8424
rect 16390 8372 16396 8424
rect 16448 8412 16454 8424
rect 16853 8415 16911 8421
rect 16853 8412 16865 8415
rect 16448 8384 16865 8412
rect 16448 8372 16454 8384
rect 16853 8381 16865 8384
rect 16899 8381 16911 8415
rect 16853 8375 16911 8381
rect 17221 8415 17279 8421
rect 17221 8381 17233 8415
rect 17267 8381 17279 8415
rect 17221 8375 17279 8381
rect 17236 8344 17264 8375
rect 15120 8316 17264 8344
rect 17604 8344 17632 8576
rect 19260 8489 19288 8576
rect 19444 8489 19472 8576
rect 19978 8548 19984 8560
rect 19536 8520 19984 8548
rect 19536 8492 19564 8520
rect 19978 8508 19984 8520
rect 20036 8508 20042 8560
rect 27246 8508 27252 8560
rect 27304 8548 27310 8560
rect 27986 8551 28044 8557
rect 27986 8548 27998 8551
rect 27304 8520 27998 8548
rect 27304 8508 27310 8520
rect 27986 8517 27998 8520
rect 28032 8517 28044 8551
rect 27986 8511 28044 8517
rect 28215 8551 28273 8557
rect 28215 8517 28227 8551
rect 28261 8548 28273 8551
rect 28350 8548 28356 8560
rect 28261 8520 28356 8548
rect 28261 8517 28273 8520
rect 28215 8511 28273 8517
rect 28350 8508 28356 8520
rect 28408 8508 28414 8560
rect 30576 8548 30604 8588
rect 32030 8548 32036 8560
rect 28966 8520 30604 8548
rect 31772 8520 32036 8548
rect 19245 8483 19303 8489
rect 19245 8449 19257 8483
rect 19291 8449 19303 8483
rect 19245 8443 19303 8449
rect 19429 8483 19487 8489
rect 19429 8449 19441 8483
rect 19475 8449 19487 8483
rect 19429 8443 19487 8449
rect 19518 8440 19524 8492
rect 19576 8440 19582 8492
rect 19613 8483 19671 8489
rect 19613 8449 19625 8483
rect 19659 8480 19671 8483
rect 20070 8480 20076 8492
rect 19659 8452 20076 8480
rect 19659 8449 19671 8452
rect 19613 8443 19671 8449
rect 20070 8440 20076 8452
rect 20128 8440 20134 8492
rect 27893 8483 27951 8489
rect 27893 8449 27905 8483
rect 27939 8480 27951 8483
rect 27939 8452 28029 8480
rect 27939 8449 27951 8452
rect 27893 8443 27951 8449
rect 18322 8372 18328 8424
rect 18380 8412 18386 8424
rect 18380 8384 26924 8412
rect 18380 8372 18386 8384
rect 19797 8347 19855 8353
rect 19797 8344 19809 8347
rect 17604 8316 19809 8344
rect 19797 8313 19809 8316
rect 19843 8313 19855 8347
rect 26896 8344 26924 8384
rect 26970 8372 26976 8424
rect 27028 8372 27034 8424
rect 28001 8412 28029 8452
rect 28074 8440 28080 8492
rect 28132 8440 28138 8492
rect 28445 8483 28503 8489
rect 28445 8480 28457 8483
rect 28276 8452 28457 8480
rect 28276 8412 28304 8452
rect 28445 8449 28457 8452
rect 28491 8449 28503 8483
rect 28445 8443 28503 8449
rect 28001 8384 28304 8412
rect 28350 8372 28356 8424
rect 28408 8372 28414 8424
rect 28460 8412 28488 8443
rect 28626 8440 28632 8492
rect 28684 8440 28690 8492
rect 28721 8483 28779 8489
rect 28966 8486 28994 8520
rect 28721 8449 28733 8483
rect 28767 8478 28779 8483
rect 28849 8478 28994 8486
rect 28767 8458 28994 8478
rect 28767 8450 28877 8458
rect 28767 8449 28779 8450
rect 28721 8443 28779 8449
rect 29454 8440 29460 8492
rect 29512 8480 29518 8492
rect 29638 8480 29644 8492
rect 29512 8452 29644 8480
rect 29512 8440 29518 8452
rect 29638 8440 29644 8452
rect 29696 8480 29702 8492
rect 30116 8489 30144 8520
rect 29825 8483 29883 8489
rect 29825 8480 29837 8483
rect 29696 8452 29837 8480
rect 29696 8440 29702 8452
rect 29825 8449 29837 8452
rect 29871 8449 29883 8483
rect 29825 8443 29883 8449
rect 30101 8483 30159 8489
rect 30101 8449 30113 8483
rect 30147 8449 30159 8483
rect 30101 8443 30159 8449
rect 31386 8440 31392 8492
rect 31444 8440 31450 8492
rect 31662 8440 31668 8492
rect 31720 8440 31726 8492
rect 31772 8489 31800 8520
rect 32030 8508 32036 8520
rect 32088 8508 32094 8560
rect 31757 8483 31815 8489
rect 31757 8449 31769 8483
rect 31803 8449 31815 8483
rect 32214 8480 32220 8492
rect 31757 8443 31815 8449
rect 31864 8452 32220 8480
rect 31202 8412 31208 8424
rect 28460 8384 31208 8412
rect 31202 8372 31208 8384
rect 31260 8412 31266 8424
rect 31864 8412 31892 8452
rect 32214 8440 32220 8452
rect 32272 8480 32278 8492
rect 32309 8483 32367 8489
rect 32309 8480 32321 8483
rect 32272 8452 32321 8480
rect 32272 8440 32278 8452
rect 32309 8449 32321 8452
rect 32355 8449 32367 8483
rect 32416 8480 32444 8588
rect 33413 8585 33425 8619
rect 33459 8616 33471 8619
rect 33502 8616 33508 8628
rect 33459 8588 33508 8616
rect 33459 8585 33471 8588
rect 33413 8579 33471 8585
rect 33502 8576 33508 8588
rect 33560 8576 33566 8628
rect 33686 8576 33692 8628
rect 33744 8576 33750 8628
rect 35802 8576 35808 8628
rect 35860 8616 35866 8628
rect 37645 8619 37703 8625
rect 37645 8616 37657 8619
rect 35860 8588 37657 8616
rect 35860 8576 35866 8588
rect 37645 8585 37657 8588
rect 37691 8585 37703 8619
rect 37645 8579 37703 8585
rect 37829 8619 37887 8625
rect 37829 8585 37841 8619
rect 37875 8616 37887 8619
rect 37918 8616 37924 8628
rect 37875 8588 37924 8616
rect 37875 8585 37887 8588
rect 37829 8579 37887 8585
rect 37918 8576 37924 8588
rect 37976 8576 37982 8628
rect 32493 8551 32551 8557
rect 32493 8517 32505 8551
rect 32539 8548 32551 8551
rect 34422 8548 34428 8560
rect 32539 8520 34428 8548
rect 32539 8517 32551 8520
rect 32493 8511 32551 8517
rect 34422 8508 34428 8520
rect 34480 8508 34486 8560
rect 34514 8508 34520 8560
rect 34572 8548 34578 8560
rect 35894 8548 35900 8560
rect 34572 8520 35900 8548
rect 34572 8508 34578 8520
rect 35894 8508 35900 8520
rect 35952 8548 35958 8560
rect 37277 8551 37335 8557
rect 37277 8548 37289 8551
rect 35952 8520 37289 8548
rect 35952 8508 35958 8520
rect 37277 8517 37289 8520
rect 37323 8548 37335 8551
rect 38289 8551 38347 8557
rect 38289 8548 38301 8551
rect 37323 8520 38301 8548
rect 37323 8517 37335 8520
rect 37277 8511 37335 8517
rect 38289 8517 38301 8520
rect 38335 8517 38347 8551
rect 38289 8511 38347 8517
rect 32416 8452 33456 8480
rect 32309 8443 32367 8449
rect 31260 8384 31892 8412
rect 31260 8372 31266 8384
rect 32030 8372 32036 8424
rect 32088 8412 32094 8424
rect 32125 8415 32183 8421
rect 32125 8412 32137 8415
rect 32088 8384 32137 8412
rect 32088 8372 32094 8384
rect 32125 8381 32137 8384
rect 32171 8412 32183 8415
rect 33042 8412 33048 8424
rect 32171 8384 33048 8412
rect 32171 8381 32183 8384
rect 32125 8375 32183 8381
rect 33042 8372 33048 8384
rect 33100 8372 33106 8424
rect 33321 8415 33379 8421
rect 33321 8381 33333 8415
rect 33367 8381 33379 8415
rect 33321 8375 33379 8381
rect 30006 8344 30012 8356
rect 26896 8316 27953 8344
rect 19797 8307 19855 8313
rect 11204 8248 11652 8276
rect 11204 8236 11210 8248
rect 11790 8236 11796 8288
rect 11848 8276 11854 8288
rect 12345 8279 12403 8285
rect 12345 8276 12357 8279
rect 11848 8248 12357 8276
rect 11848 8236 11854 8248
rect 12345 8245 12357 8248
rect 12391 8245 12403 8279
rect 12345 8239 12403 8245
rect 16666 8236 16672 8288
rect 16724 8236 16730 8288
rect 18598 8236 18604 8288
rect 18656 8276 18662 8288
rect 20622 8276 20628 8288
rect 18656 8248 20628 8276
rect 18656 8236 18662 8248
rect 20622 8236 20628 8248
rect 20680 8236 20686 8288
rect 27430 8236 27436 8288
rect 27488 8276 27494 8288
rect 27617 8279 27675 8285
rect 27617 8276 27629 8279
rect 27488 8248 27629 8276
rect 27488 8236 27494 8248
rect 27617 8245 27629 8248
rect 27663 8245 27675 8279
rect 27617 8239 27675 8245
rect 27706 8236 27712 8288
rect 27764 8236 27770 8288
rect 27925 8276 27953 8316
rect 28736 8316 30012 8344
rect 28074 8276 28080 8288
rect 27925 8248 28080 8276
rect 28074 8236 28080 8248
rect 28132 8276 28138 8288
rect 28626 8276 28632 8288
rect 28132 8248 28632 8276
rect 28132 8236 28138 8248
rect 28626 8236 28632 8248
rect 28684 8276 28690 8288
rect 28736 8276 28764 8316
rect 30006 8304 30012 8316
rect 30064 8344 30070 8356
rect 30064 8316 31616 8344
rect 30064 8304 30070 8316
rect 28684 8248 28764 8276
rect 29917 8279 29975 8285
rect 28684 8236 28690 8248
rect 29917 8245 29929 8279
rect 29963 8276 29975 8279
rect 30282 8276 30288 8288
rect 29963 8248 30288 8276
rect 29963 8245 29975 8248
rect 29917 8239 29975 8245
rect 30282 8236 30288 8248
rect 30340 8236 30346 8288
rect 31588 8276 31616 8316
rect 31662 8304 31668 8356
rect 31720 8344 31726 8356
rect 33226 8344 33232 8356
rect 31720 8316 33232 8344
rect 31720 8304 31726 8316
rect 33226 8304 33232 8316
rect 33284 8344 33290 8356
rect 33336 8344 33364 8375
rect 33284 8316 33364 8344
rect 33428 8344 33456 8452
rect 34238 8440 34244 8492
rect 34296 8480 34302 8492
rect 35342 8480 35348 8492
rect 34296 8452 35348 8480
rect 34296 8440 34302 8452
rect 35342 8440 35348 8452
rect 35400 8440 35406 8492
rect 37458 8440 37464 8492
rect 37516 8440 37522 8492
rect 37550 8440 37556 8492
rect 37608 8440 37614 8492
rect 38102 8440 38108 8492
rect 38160 8440 38166 8492
rect 38378 8440 38384 8492
rect 38436 8440 38442 8492
rect 33505 8415 33563 8421
rect 33505 8381 33517 8415
rect 33551 8412 33563 8415
rect 33962 8412 33968 8424
rect 33551 8384 33968 8412
rect 33551 8381 33563 8384
rect 33505 8375 33563 8381
rect 33962 8372 33968 8384
rect 34020 8412 34026 8424
rect 34790 8412 34796 8424
rect 34020 8384 34796 8412
rect 34020 8372 34026 8384
rect 34790 8372 34796 8384
rect 34848 8372 34854 8424
rect 37921 8415 37979 8421
rect 37921 8381 37933 8415
rect 37967 8412 37979 8415
rect 38194 8412 38200 8424
rect 37967 8384 38200 8412
rect 37967 8381 37979 8384
rect 37921 8375 37979 8381
rect 38194 8372 38200 8384
rect 38252 8372 38258 8424
rect 41138 8344 41144 8356
rect 33428 8316 41144 8344
rect 33284 8304 33290 8316
rect 41138 8304 41144 8316
rect 41196 8304 41202 8356
rect 32766 8276 32772 8288
rect 31588 8248 32772 8276
rect 32766 8236 32772 8248
rect 32824 8236 32830 8288
rect 33870 8236 33876 8288
rect 33928 8276 33934 8288
rect 34330 8276 34336 8288
rect 33928 8248 34336 8276
rect 33928 8236 33934 8248
rect 34330 8236 34336 8248
rect 34388 8236 34394 8288
rect 35710 8236 35716 8288
rect 35768 8276 35774 8288
rect 41046 8276 41052 8288
rect 35768 8248 41052 8276
rect 35768 8236 35774 8248
rect 41046 8236 41052 8248
rect 41104 8236 41110 8288
rect 1104 8186 41400 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 41400 8186
rect 1104 8112 41400 8134
rect 1765 8075 1823 8081
rect 1765 8041 1777 8075
rect 1811 8072 1823 8075
rect 7558 8072 7564 8084
rect 1811 8044 7564 8072
rect 1811 8041 1823 8044
rect 1765 8035 1823 8041
rect 7558 8032 7564 8044
rect 7616 8032 7622 8084
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 8110 8072 8116 8084
rect 7800 8044 8116 8072
rect 7800 8032 7806 8044
rect 8110 8032 8116 8044
rect 8168 8072 8174 8084
rect 18693 8075 18751 8081
rect 8168 8044 12388 8072
rect 8168 8032 8174 8044
rect 7466 7964 7472 8016
rect 7524 8004 7530 8016
rect 8202 8004 8208 8016
rect 7524 7976 8208 8004
rect 7524 7964 7530 7976
rect 8202 7964 8208 7976
rect 8260 7964 8266 8016
rect 11054 7964 11060 8016
rect 11112 7964 11118 8016
rect 8018 7896 8024 7948
rect 8076 7936 8082 7948
rect 8573 7939 8631 7945
rect 8573 7936 8585 7939
rect 8076 7908 8585 7936
rect 8076 7896 8082 7908
rect 8573 7905 8585 7908
rect 8619 7905 8631 7939
rect 8573 7899 8631 7905
rect 11256 7908 11744 7936
rect 7935 7871 7993 7877
rect 7935 7837 7947 7871
rect 7981 7868 7993 7871
rect 8036 7868 8064 7896
rect 7981 7840 8064 7868
rect 7981 7837 7993 7840
rect 7935 7831 7993 7837
rect 8110 7828 8116 7880
rect 8168 7828 8174 7880
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7868 8263 7871
rect 11057 7871 11115 7877
rect 8251 7840 8708 7868
rect 8251 7837 8263 7840
rect 8205 7831 8263 7837
rect 8680 7812 8708 7840
rect 11057 7837 11069 7871
rect 11103 7868 11115 7871
rect 11146 7868 11152 7880
rect 11103 7840 11152 7868
rect 11103 7837 11115 7840
rect 11057 7831 11115 7837
rect 11146 7828 11152 7840
rect 11204 7828 11210 7880
rect 11256 7877 11284 7908
rect 11716 7877 11744 7908
rect 11241 7871 11299 7877
rect 11241 7837 11253 7871
rect 11287 7837 11299 7871
rect 11241 7831 11299 7837
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7868 11391 7871
rect 11609 7871 11667 7877
rect 11609 7868 11621 7871
rect 11379 7840 11621 7868
rect 11379 7837 11391 7840
rect 11333 7831 11391 7837
rect 934 7760 940 7812
rect 992 7800 998 7812
rect 1489 7803 1547 7809
rect 1489 7800 1501 7803
rect 992 7772 1501 7800
rect 992 7760 998 7772
rect 1489 7769 1501 7772
rect 1535 7769 1547 7803
rect 1489 7763 1547 7769
rect 8386 7760 8392 7812
rect 8444 7760 8450 7812
rect 8662 7760 8668 7812
rect 8720 7760 8726 7812
rect 11532 7744 11560 7840
rect 11609 7837 11621 7840
rect 11655 7837 11667 7871
rect 11609 7831 11667 7837
rect 11701 7871 11759 7877
rect 11701 7837 11713 7871
rect 11747 7868 11759 7871
rect 11790 7868 11796 7880
rect 11747 7840 11796 7868
rect 11747 7837 11759 7840
rect 11701 7831 11759 7837
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 11882 7828 11888 7880
rect 11940 7828 11946 7880
rect 11977 7871 12035 7877
rect 11977 7837 11989 7871
rect 12023 7868 12035 7871
rect 12066 7868 12072 7880
rect 12023 7840 12072 7868
rect 12023 7837 12035 7840
rect 11977 7831 12035 7837
rect 11992 7800 12020 7831
rect 12066 7828 12072 7840
rect 12124 7828 12130 7880
rect 12360 7868 12388 8044
rect 18693 8041 18705 8075
rect 18739 8072 18751 8075
rect 18966 8072 18972 8084
rect 18739 8044 18972 8072
rect 18739 8041 18751 8044
rect 18693 8035 18751 8041
rect 18966 8032 18972 8044
rect 19024 8032 19030 8084
rect 20254 8072 20260 8084
rect 19720 8044 20260 8072
rect 12710 7964 12716 8016
rect 12768 7964 12774 8016
rect 13538 8004 13544 8016
rect 12820 7976 13544 8004
rect 12437 7939 12495 7945
rect 12437 7905 12449 7939
rect 12483 7936 12495 7939
rect 12728 7936 12756 7964
rect 12483 7908 12756 7936
rect 12483 7905 12495 7908
rect 12437 7899 12495 7905
rect 12710 7868 12716 7880
rect 12360 7840 12716 7868
rect 12710 7828 12716 7840
rect 12768 7828 12774 7880
rect 12820 7877 12848 7976
rect 13538 7964 13544 7976
rect 13596 7964 13602 8016
rect 13173 7939 13231 7945
rect 13173 7936 13185 7939
rect 12912 7908 13185 7936
rect 12805 7871 12863 7877
rect 12805 7837 12817 7871
rect 12851 7837 12863 7871
rect 12805 7831 12863 7837
rect 11716 7772 12020 7800
rect 11716 7744 11744 7772
rect 12250 7760 12256 7812
rect 12308 7800 12314 7812
rect 12912 7800 12940 7908
rect 13173 7905 13185 7908
rect 13219 7905 13231 7939
rect 13173 7899 13231 7905
rect 18601 7939 18659 7945
rect 18601 7905 18613 7939
rect 18647 7936 18659 7939
rect 19426 7936 19432 7948
rect 18647 7908 19432 7936
rect 18647 7905 18659 7908
rect 18601 7899 18659 7905
rect 19426 7896 19432 7908
rect 19484 7936 19490 7948
rect 19720 7945 19748 8044
rect 20254 8032 20260 8044
rect 20312 8032 20318 8084
rect 20806 8032 20812 8084
rect 20864 8072 20870 8084
rect 21729 8075 21787 8081
rect 21729 8072 21741 8075
rect 20864 8044 21741 8072
rect 20864 8032 20870 8044
rect 21729 8041 21741 8044
rect 21775 8041 21787 8075
rect 26145 8075 26203 8081
rect 21729 8035 21787 8041
rect 23584 8044 26096 8072
rect 23584 8016 23612 8044
rect 23566 7964 23572 8016
rect 23624 7964 23630 8016
rect 26068 8004 26096 8044
rect 26145 8041 26157 8075
rect 26191 8072 26203 8075
rect 26970 8072 26976 8084
rect 26191 8044 26976 8072
rect 26191 8041 26203 8044
rect 26145 8035 26203 8041
rect 26970 8032 26976 8044
rect 27028 8032 27034 8084
rect 29546 8072 29552 8084
rect 27632 8044 29552 8072
rect 27632 8004 27660 8044
rect 29546 8032 29552 8044
rect 29604 8032 29610 8084
rect 29822 8032 29828 8084
rect 29880 8072 29886 8084
rect 30926 8072 30932 8084
rect 29880 8044 30932 8072
rect 29880 8032 29886 8044
rect 30926 8032 30932 8044
rect 30984 8032 30990 8084
rect 32398 8072 32404 8084
rect 31726 8044 32404 8072
rect 26068 7976 27660 8004
rect 27706 7964 27712 8016
rect 27764 7964 27770 8016
rect 31726 8004 31754 8044
rect 32398 8032 32404 8044
rect 32456 8032 32462 8084
rect 34054 8032 34060 8084
rect 34112 8072 34118 8084
rect 35345 8075 35403 8081
rect 35345 8072 35357 8075
rect 34112 8044 35357 8072
rect 34112 8032 34118 8044
rect 35345 8041 35357 8044
rect 35391 8041 35403 8075
rect 35345 8035 35403 8041
rect 36633 8075 36691 8081
rect 36633 8041 36645 8075
rect 36679 8072 36691 8075
rect 38378 8072 38384 8084
rect 36679 8044 38384 8072
rect 36679 8041 36691 8044
rect 36633 8035 36691 8041
rect 38378 8032 38384 8044
rect 38436 8032 38442 8084
rect 28966 7976 31754 8004
rect 19613 7939 19671 7945
rect 19613 7936 19625 7939
rect 19484 7908 19625 7936
rect 19484 7896 19490 7908
rect 19613 7905 19625 7908
rect 19659 7905 19671 7939
rect 19613 7899 19671 7905
rect 19705 7939 19763 7945
rect 19705 7905 19717 7939
rect 19751 7905 19763 7939
rect 19705 7899 19763 7905
rect 19981 7939 20039 7945
rect 19981 7905 19993 7939
rect 20027 7936 20039 7939
rect 21818 7936 21824 7948
rect 20027 7908 21824 7936
rect 20027 7905 20039 7908
rect 19981 7899 20039 7905
rect 21818 7896 21824 7908
rect 21876 7936 21882 7948
rect 22741 7939 22799 7945
rect 22741 7936 22753 7939
rect 21876 7908 22753 7936
rect 21876 7896 21882 7908
rect 22741 7905 22753 7908
rect 22787 7936 22799 7939
rect 24210 7936 24216 7948
rect 22787 7908 24216 7936
rect 22787 7905 22799 7908
rect 22741 7899 22799 7905
rect 24210 7896 24216 7908
rect 24268 7936 24274 7948
rect 24397 7939 24455 7945
rect 24397 7936 24409 7939
rect 24268 7908 24409 7936
rect 24268 7896 24274 7908
rect 24397 7905 24409 7908
rect 24443 7905 24455 7939
rect 24397 7899 24455 7905
rect 24673 7939 24731 7945
rect 24673 7905 24685 7939
rect 24719 7936 24731 7939
rect 27724 7936 27752 7964
rect 24719 7908 27752 7936
rect 24719 7905 24731 7908
rect 24673 7899 24731 7905
rect 13081 7871 13139 7877
rect 13081 7837 13093 7871
rect 13127 7868 13139 7871
rect 13998 7868 14004 7880
rect 13127 7840 14004 7868
rect 13127 7837 13139 7840
rect 13081 7831 13139 7837
rect 13998 7828 14004 7840
rect 14056 7828 14062 7880
rect 17770 7828 17776 7880
rect 17828 7868 17834 7880
rect 18325 7871 18383 7877
rect 18325 7868 18337 7871
rect 17828 7840 18337 7868
rect 17828 7828 17834 7840
rect 18325 7837 18337 7840
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 18874 7828 18880 7880
rect 18932 7868 18938 7880
rect 18932 7840 20024 7868
rect 18932 7828 18938 7840
rect 12308 7772 12940 7800
rect 12308 7760 12314 7772
rect 18690 7760 18696 7812
rect 18748 7800 18754 7812
rect 19889 7803 19947 7809
rect 19889 7800 19901 7803
rect 18748 7772 19901 7800
rect 18748 7760 18754 7772
rect 19889 7769 19901 7772
rect 19935 7769 19947 7803
rect 19889 7763 19947 7769
rect 8110 7692 8116 7744
rect 8168 7692 8174 7744
rect 11422 7692 11428 7744
rect 11480 7692 11486 7744
rect 11514 7692 11520 7744
rect 11572 7692 11578 7744
rect 11698 7692 11704 7744
rect 11756 7692 11762 7744
rect 15470 7692 15476 7744
rect 15528 7732 15534 7744
rect 16206 7732 16212 7744
rect 15528 7704 16212 7732
rect 15528 7692 15534 7704
rect 16206 7692 16212 7704
rect 16264 7692 16270 7744
rect 18877 7735 18935 7741
rect 18877 7701 18889 7735
rect 18923 7732 18935 7735
rect 19245 7735 19303 7741
rect 19245 7732 19257 7735
rect 18923 7704 19257 7732
rect 18923 7701 18935 7704
rect 18877 7695 18935 7701
rect 19245 7701 19257 7704
rect 19291 7701 19303 7735
rect 19996 7732 20024 7840
rect 23382 7828 23388 7880
rect 23440 7868 23446 7880
rect 23477 7871 23535 7877
rect 23477 7868 23489 7871
rect 23440 7840 23489 7868
rect 23440 7828 23446 7840
rect 23477 7837 23489 7840
rect 23523 7837 23535 7871
rect 28966 7868 28994 7976
rect 32030 7964 32036 8016
rect 32088 8004 32094 8016
rect 32088 7976 37228 8004
rect 32088 7964 32094 7976
rect 29730 7896 29736 7948
rect 29788 7936 29794 7948
rect 34701 7939 34759 7945
rect 29788 7908 30512 7936
rect 29788 7896 29794 7908
rect 23477 7831 23535 7837
rect 27172 7840 28994 7868
rect 20254 7760 20260 7812
rect 20312 7760 20318 7812
rect 20714 7800 20720 7812
rect 20364 7772 20720 7800
rect 20364 7732 20392 7772
rect 20714 7760 20720 7772
rect 20772 7760 20778 7812
rect 21910 7800 21916 7812
rect 21560 7772 21916 7800
rect 19996 7704 20392 7732
rect 19245 7695 19303 7701
rect 20898 7692 20904 7744
rect 20956 7732 20962 7744
rect 21560 7732 21588 7772
rect 21910 7760 21916 7772
rect 21968 7760 21974 7812
rect 23492 7800 23520 7831
rect 27172 7812 27200 7840
rect 29270 7828 29276 7880
rect 29328 7868 29334 7880
rect 29825 7871 29883 7877
rect 29825 7868 29837 7871
rect 29328 7840 29837 7868
rect 29328 7828 29334 7840
rect 29825 7837 29837 7840
rect 29871 7868 29883 7871
rect 30098 7868 30104 7880
rect 29871 7840 30104 7868
rect 29871 7837 29883 7840
rect 29825 7831 29883 7837
rect 30098 7828 30104 7840
rect 30156 7828 30162 7880
rect 30484 7812 30512 7908
rect 34701 7905 34713 7939
rect 34747 7936 34759 7939
rect 37093 7939 37151 7945
rect 37093 7936 37105 7939
rect 34747 7908 37105 7936
rect 34747 7905 34759 7908
rect 34701 7899 34759 7905
rect 37093 7905 37105 7908
rect 37139 7905 37151 7939
rect 37093 7899 37151 7905
rect 31570 7828 31576 7880
rect 31628 7868 31634 7880
rect 34882 7868 34888 7880
rect 31628 7840 34888 7868
rect 31628 7828 31634 7840
rect 34882 7828 34888 7840
rect 34940 7828 34946 7880
rect 34974 7828 34980 7880
rect 35032 7878 35038 7880
rect 35032 7877 35204 7878
rect 35032 7871 35219 7877
rect 35032 7850 35173 7871
rect 35032 7828 35038 7850
rect 35161 7837 35173 7850
rect 35207 7837 35219 7871
rect 35161 7831 35219 7837
rect 35437 7871 35495 7877
rect 35437 7837 35449 7871
rect 35483 7868 35495 7871
rect 35483 7840 35664 7868
rect 35483 7837 35495 7840
rect 35437 7831 35495 7837
rect 23492 7772 24900 7800
rect 20956 7704 21588 7732
rect 20956 7692 20962 7704
rect 23566 7692 23572 7744
rect 23624 7692 23630 7744
rect 24872 7732 24900 7772
rect 24946 7760 24952 7812
rect 25004 7800 25010 7812
rect 25004 7772 25162 7800
rect 25004 7760 25010 7772
rect 26050 7760 26056 7812
rect 26108 7800 26114 7812
rect 27154 7800 27160 7812
rect 26108 7772 27160 7800
rect 26108 7760 26114 7772
rect 27154 7760 27160 7772
rect 27212 7760 27218 7812
rect 29454 7800 29460 7812
rect 28368 7772 29460 7800
rect 28368 7744 28396 7772
rect 29454 7760 29460 7772
rect 29512 7760 29518 7812
rect 29546 7760 29552 7812
rect 29604 7760 29610 7812
rect 29730 7760 29736 7812
rect 29788 7760 29794 7812
rect 30466 7760 30472 7812
rect 30524 7800 30530 7812
rect 33778 7800 33784 7812
rect 30524 7772 33784 7800
rect 30524 7760 30530 7772
rect 33778 7760 33784 7772
rect 33836 7760 33842 7812
rect 35066 7760 35072 7812
rect 35124 7760 35130 7812
rect 35529 7803 35587 7809
rect 35529 7769 35541 7803
rect 35575 7769 35587 7803
rect 35529 7763 35587 7769
rect 28350 7732 28356 7744
rect 24872 7704 28356 7732
rect 28350 7692 28356 7704
rect 28408 7692 28414 7744
rect 29086 7692 29092 7744
rect 29144 7732 29150 7744
rect 29641 7735 29699 7741
rect 29641 7732 29653 7735
rect 29144 7704 29653 7732
rect 29144 7692 29150 7704
rect 29641 7701 29653 7704
rect 29687 7732 29699 7735
rect 30190 7732 30196 7744
rect 29687 7704 30196 7732
rect 29687 7701 29699 7704
rect 29641 7695 29699 7701
rect 30190 7692 30196 7704
rect 30248 7692 30254 7744
rect 30650 7692 30656 7744
rect 30708 7732 30714 7744
rect 32122 7732 32128 7744
rect 30708 7704 32128 7732
rect 30708 7692 30714 7704
rect 32122 7692 32128 7704
rect 32180 7732 32186 7744
rect 34698 7732 34704 7744
rect 32180 7704 34704 7732
rect 32180 7692 32186 7704
rect 34698 7692 34704 7704
rect 34756 7692 34762 7744
rect 34974 7692 34980 7744
rect 35032 7741 35038 7744
rect 35032 7732 35041 7741
rect 35032 7704 35077 7732
rect 35032 7695 35041 7704
rect 35032 7692 35038 7695
rect 35342 7692 35348 7744
rect 35400 7732 35406 7744
rect 35544 7732 35572 7763
rect 35400 7704 35572 7732
rect 35636 7732 35664 7840
rect 35986 7828 35992 7880
rect 36044 7868 36050 7880
rect 36817 7871 36875 7877
rect 36817 7868 36829 7871
rect 36044 7840 36829 7868
rect 36044 7828 36050 7840
rect 36817 7837 36829 7840
rect 36863 7837 36875 7871
rect 36817 7831 36875 7837
rect 36909 7871 36967 7877
rect 36909 7837 36921 7871
rect 36955 7837 36967 7871
rect 36909 7831 36967 7837
rect 37001 7871 37059 7877
rect 37001 7837 37013 7871
rect 37047 7868 37059 7871
rect 37200 7868 37228 7976
rect 37458 7896 37464 7948
rect 37516 7896 37522 7948
rect 37550 7896 37556 7948
rect 37608 7896 37614 7948
rect 37476 7868 37504 7896
rect 37047 7840 37504 7868
rect 37047 7837 37059 7840
rect 37001 7831 37059 7837
rect 35710 7760 35716 7812
rect 35768 7760 35774 7812
rect 35802 7760 35808 7812
rect 35860 7800 35866 7812
rect 35897 7803 35955 7809
rect 35897 7800 35909 7803
rect 35860 7772 35909 7800
rect 35860 7760 35866 7772
rect 35897 7769 35909 7772
rect 35943 7800 35955 7803
rect 36924 7800 36952 7831
rect 37568 7800 37596 7896
rect 35943 7772 37596 7800
rect 35943 7769 35955 7772
rect 35897 7763 35955 7769
rect 36078 7732 36084 7744
rect 35636 7704 36084 7732
rect 35400 7692 35406 7704
rect 36078 7692 36084 7704
rect 36136 7732 36142 7744
rect 40770 7732 40776 7744
rect 36136 7704 40776 7732
rect 36136 7692 36142 7704
rect 40770 7692 40776 7704
rect 40828 7692 40834 7744
rect 1104 7642 41400 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 41400 7642
rect 1104 7568 41400 7590
rect 7834 7528 7840 7540
rect 7116 7500 7840 7528
rect 7116 7469 7144 7500
rect 7834 7488 7840 7500
rect 7892 7488 7898 7540
rect 8110 7488 8116 7540
rect 8168 7488 8174 7540
rect 8573 7531 8631 7537
rect 8573 7497 8585 7531
rect 8619 7528 8631 7531
rect 8662 7528 8668 7540
rect 8619 7500 8668 7528
rect 8619 7497 8631 7500
rect 8573 7491 8631 7497
rect 8662 7488 8668 7500
rect 8720 7528 8726 7540
rect 10873 7531 10931 7537
rect 8720 7500 9260 7528
rect 8720 7488 8726 7500
rect 7101 7463 7159 7469
rect 7101 7429 7113 7463
rect 7147 7429 7159 7463
rect 7101 7423 7159 7429
rect 7190 7420 7196 7472
rect 7248 7460 7254 7472
rect 8128 7460 8156 7488
rect 7248 7432 7420 7460
rect 8128 7432 8984 7460
rect 7248 7420 7254 7432
rect 7392 7401 7420 7432
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7361 7343 7395
rect 7285 7355 7343 7361
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7361 7435 7395
rect 7653 7395 7711 7401
rect 7653 7392 7665 7395
rect 7377 7355 7435 7361
rect 7576 7364 7665 7392
rect 7300 7256 7328 7355
rect 7576 7336 7604 7364
rect 7653 7361 7665 7364
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 7742 7352 7748 7404
rect 7800 7352 7806 7404
rect 7834 7352 7840 7404
rect 7892 7352 7898 7404
rect 7975 7395 8033 7401
rect 7975 7361 7987 7395
rect 8021 7392 8033 7395
rect 8294 7392 8300 7404
rect 8021 7364 8300 7392
rect 8021 7361 8033 7364
rect 7975 7355 8033 7361
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 8386 7352 8392 7404
rect 8444 7352 8450 7404
rect 8478 7352 8484 7404
rect 8536 7392 8542 7404
rect 8956 7401 8984 7432
rect 9122 7420 9128 7472
rect 9180 7420 9186 7472
rect 9232 7460 9260 7500
rect 10873 7497 10885 7531
rect 10919 7497 10931 7531
rect 11790 7528 11796 7540
rect 10873 7491 10931 7497
rect 10980 7500 11796 7528
rect 10888 7460 10916 7491
rect 9232 7432 10916 7460
rect 8665 7395 8723 7401
rect 8665 7392 8677 7395
rect 8536 7364 8677 7392
rect 8536 7352 8542 7364
rect 8665 7361 8677 7364
rect 8711 7361 8723 7395
rect 8665 7355 8723 7361
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7361 8999 7395
rect 8941 7355 8999 7361
rect 7558 7284 7564 7336
rect 7616 7284 7622 7336
rect 8113 7327 8171 7333
rect 8113 7293 8125 7327
rect 8159 7324 8171 7327
rect 8202 7324 8208 7336
rect 8159 7296 8208 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 8404 7324 8432 7352
rect 8846 7324 8852 7336
rect 8404 7296 8852 7324
rect 8846 7284 8852 7296
rect 8904 7324 8910 7336
rect 9140 7324 9168 7420
rect 9232 7401 9260 7432
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7361 9275 7395
rect 9217 7355 9275 7361
rect 10873 7395 10931 7401
rect 10873 7361 10885 7395
rect 10919 7392 10931 7395
rect 10980 7392 11008 7500
rect 11790 7488 11796 7500
rect 11848 7528 11854 7540
rect 11848 7500 12480 7528
rect 11848 7488 11854 7500
rect 11514 7460 11520 7472
rect 10919 7364 11008 7392
rect 11164 7432 11520 7460
rect 10919 7361 10931 7364
rect 10873 7355 10931 7361
rect 8904 7296 9168 7324
rect 10689 7327 10747 7333
rect 8904 7284 8910 7296
rect 10689 7293 10701 7327
rect 10735 7324 10747 7327
rect 11164 7324 11192 7432
rect 11514 7420 11520 7432
rect 11572 7460 11578 7472
rect 11572 7432 12296 7460
rect 11572 7420 11578 7432
rect 12268 7404 12296 7432
rect 11241 7395 11299 7401
rect 11241 7361 11253 7395
rect 11287 7392 11299 7395
rect 11698 7392 11704 7404
rect 11287 7364 11704 7392
rect 11287 7361 11299 7364
rect 11241 7355 11299 7361
rect 11698 7352 11704 7364
rect 11756 7352 11762 7404
rect 11793 7395 11851 7401
rect 11793 7361 11805 7395
rect 11839 7361 11851 7395
rect 11793 7355 11851 7361
rect 11977 7395 12035 7401
rect 11977 7361 11989 7395
rect 12023 7392 12035 7395
rect 12023 7364 12204 7392
rect 12023 7361 12035 7364
rect 11977 7355 12035 7361
rect 10735 7296 11192 7324
rect 10735 7293 10747 7296
rect 10689 7287 10747 7293
rect 8757 7259 8815 7265
rect 8757 7256 8769 7259
rect 7300 7228 8769 7256
rect 8757 7225 8769 7228
rect 8803 7225 8815 7259
rect 8757 7219 8815 7225
rect 11606 7216 11612 7268
rect 11664 7256 11670 7268
rect 11808 7256 11836 7355
rect 11882 7284 11888 7336
rect 11940 7324 11946 7336
rect 12069 7327 12127 7333
rect 12069 7324 12081 7327
rect 11940 7296 12081 7324
rect 11940 7284 11946 7296
rect 12069 7293 12081 7296
rect 12115 7293 12127 7327
rect 12176 7324 12204 7364
rect 12250 7352 12256 7404
rect 12308 7352 12314 7404
rect 12452 7401 12480 7500
rect 14090 7488 14096 7540
rect 14148 7488 14154 7540
rect 16022 7528 16028 7540
rect 15028 7500 16028 7528
rect 12710 7420 12716 7472
rect 12768 7420 12774 7472
rect 13998 7420 14004 7472
rect 14056 7420 14062 7472
rect 12437 7395 12495 7401
rect 12437 7361 12449 7395
rect 12483 7361 12495 7395
rect 12437 7355 12495 7361
rect 12526 7352 12532 7404
rect 12584 7392 12590 7404
rect 12621 7395 12679 7401
rect 12621 7392 12633 7395
rect 12584 7364 12633 7392
rect 12584 7352 12590 7364
rect 12621 7361 12633 7364
rect 12667 7392 12679 7395
rect 14108 7392 14136 7488
rect 14660 7432 14872 7460
rect 14185 7395 14243 7401
rect 14185 7392 14197 7395
rect 12667 7364 13676 7392
rect 14108 7364 14197 7392
rect 12667 7361 12679 7364
rect 12621 7355 12679 7361
rect 12802 7324 12808 7336
rect 12176 7296 12808 7324
rect 12069 7287 12127 7293
rect 11664 7228 11836 7256
rect 11664 7216 11670 7228
rect 7101 7191 7159 7197
rect 7101 7157 7113 7191
rect 7147 7188 7159 7191
rect 7374 7188 7380 7200
rect 7147 7160 7380 7188
rect 7147 7157 7159 7160
rect 7101 7151 7159 7157
rect 7374 7148 7380 7160
rect 7432 7148 7438 7200
rect 7466 7148 7472 7200
rect 7524 7148 7530 7200
rect 7742 7148 7748 7200
rect 7800 7188 7806 7200
rect 8205 7191 8263 7197
rect 8205 7188 8217 7191
rect 7800 7160 8217 7188
rect 7800 7148 7806 7160
rect 8205 7157 8217 7160
rect 8251 7157 8263 7191
rect 8205 7151 8263 7157
rect 8478 7148 8484 7200
rect 8536 7188 8542 7200
rect 12084 7188 12112 7287
rect 12802 7284 12808 7296
rect 12860 7284 12866 7336
rect 13648 7324 13676 7364
rect 14185 7361 14197 7364
rect 14231 7361 14243 7395
rect 14185 7355 14243 7361
rect 14366 7352 14372 7404
rect 14424 7392 14430 7404
rect 14660 7401 14688 7432
rect 14844 7404 14872 7432
rect 14461 7395 14519 7401
rect 14461 7392 14473 7395
rect 14424 7364 14473 7392
rect 14424 7352 14430 7364
rect 14461 7361 14473 7364
rect 14507 7361 14519 7395
rect 14461 7355 14519 7361
rect 14645 7395 14703 7401
rect 14645 7361 14657 7395
rect 14691 7361 14703 7395
rect 14645 7355 14703 7361
rect 14660 7324 14688 7355
rect 14826 7352 14832 7404
rect 14884 7352 14890 7404
rect 15028 7336 15056 7500
rect 16022 7488 16028 7500
rect 16080 7488 16086 7540
rect 16485 7531 16543 7537
rect 16485 7497 16497 7531
rect 16531 7497 16543 7531
rect 19334 7528 19340 7540
rect 16485 7491 16543 7497
rect 18156 7500 19340 7528
rect 15381 7463 15439 7469
rect 15381 7429 15393 7463
rect 15427 7460 15439 7463
rect 16500 7460 16528 7491
rect 15427 7432 15700 7460
rect 15427 7429 15439 7432
rect 15381 7423 15439 7429
rect 15105 7395 15163 7401
rect 15105 7361 15117 7395
rect 15151 7392 15163 7395
rect 15470 7392 15476 7404
rect 15151 7390 15240 7392
rect 15304 7390 15476 7392
rect 15151 7364 15476 7390
rect 15151 7361 15163 7364
rect 15212 7362 15332 7364
rect 15105 7355 15163 7361
rect 13648 7296 14688 7324
rect 15010 7284 15016 7336
rect 15068 7324 15074 7336
rect 15197 7327 15255 7333
rect 15197 7324 15209 7327
rect 15068 7296 15209 7324
rect 15068 7284 15074 7296
rect 15197 7293 15209 7296
rect 15243 7293 15255 7327
rect 15197 7287 15255 7293
rect 13814 7216 13820 7268
rect 13872 7256 13878 7268
rect 15304 7256 15332 7362
rect 15470 7352 15476 7364
rect 15528 7352 15534 7404
rect 15672 7401 15700 7432
rect 15856 7432 16528 7460
rect 15657 7395 15715 7401
rect 15657 7361 15669 7395
rect 15703 7361 15715 7395
rect 15657 7355 15715 7361
rect 15750 7395 15808 7401
rect 15750 7361 15762 7395
rect 15796 7392 15808 7395
rect 15856 7392 15884 7432
rect 15796 7364 15884 7392
rect 15933 7395 15991 7401
rect 15796 7361 15808 7364
rect 15750 7355 15808 7361
rect 15933 7361 15945 7395
rect 15979 7361 15991 7395
rect 15933 7355 15991 7361
rect 15378 7284 15384 7336
rect 15436 7284 15442 7336
rect 15838 7284 15844 7336
rect 15896 7284 15902 7336
rect 15948 7324 15976 7355
rect 16022 7352 16028 7404
rect 16080 7392 16086 7404
rect 16117 7395 16175 7401
rect 16117 7392 16129 7395
rect 16080 7364 16129 7392
rect 16080 7352 16086 7364
rect 16117 7361 16129 7364
rect 16163 7361 16175 7395
rect 16117 7355 16175 7361
rect 16206 7352 16212 7404
rect 16264 7352 16270 7404
rect 16666 7352 16672 7404
rect 16724 7352 16730 7404
rect 18156 7401 18184 7500
rect 19334 7488 19340 7500
rect 19392 7488 19398 7540
rect 20254 7488 20260 7540
rect 20312 7528 20318 7540
rect 21085 7531 21143 7537
rect 21085 7528 21097 7531
rect 20312 7500 21097 7528
rect 20312 7488 20318 7500
rect 21085 7497 21097 7500
rect 21131 7497 21143 7531
rect 23566 7528 23572 7540
rect 21085 7491 21143 7497
rect 21928 7500 23572 7528
rect 18417 7463 18475 7469
rect 18417 7429 18429 7463
rect 18463 7460 18475 7463
rect 18690 7460 18696 7472
rect 18463 7432 18696 7460
rect 18463 7429 18475 7432
rect 18417 7423 18475 7429
rect 18690 7420 18696 7432
rect 18748 7420 18754 7472
rect 18874 7420 18880 7472
rect 18932 7420 18938 7472
rect 20346 7420 20352 7472
rect 20404 7460 20410 7472
rect 20404 7432 21312 7460
rect 20404 7420 20410 7432
rect 18141 7395 18199 7401
rect 18141 7361 18153 7395
rect 18187 7361 18199 7395
rect 18141 7355 18199 7361
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7392 20499 7395
rect 20806 7392 20812 7404
rect 20487 7364 20812 7392
rect 20487 7361 20499 7364
rect 20441 7355 20499 7361
rect 20806 7352 20812 7364
rect 20864 7352 20870 7404
rect 21284 7401 21312 7432
rect 21928 7401 21956 7500
rect 23566 7488 23572 7500
rect 23624 7488 23630 7540
rect 24118 7488 24124 7540
rect 24176 7488 24182 7540
rect 25774 7528 25780 7540
rect 25516 7500 25780 7528
rect 24136 7460 24164 7488
rect 25516 7469 25544 7500
rect 25774 7488 25780 7500
rect 25832 7528 25838 7540
rect 34330 7528 34336 7540
rect 25832 7500 26372 7528
rect 25832 7488 25838 7500
rect 23492 7432 24164 7460
rect 25501 7463 25559 7469
rect 21269 7395 21327 7401
rect 21269 7361 21281 7395
rect 21315 7361 21327 7395
rect 21269 7355 21327 7361
rect 21913 7395 21971 7401
rect 21913 7361 21925 7395
rect 21959 7361 21971 7395
rect 21913 7355 21971 7361
rect 22094 7352 22100 7404
rect 22152 7352 22158 7404
rect 23492 7401 23520 7432
rect 25501 7429 25513 7463
rect 25547 7429 25559 7463
rect 25501 7423 25559 7429
rect 26142 7420 26148 7472
rect 26200 7460 26206 7472
rect 26344 7469 26372 7500
rect 26988 7500 34336 7528
rect 26237 7463 26295 7469
rect 26237 7460 26249 7463
rect 26200 7432 26249 7460
rect 26200 7420 26206 7432
rect 26237 7429 26249 7432
rect 26283 7429 26295 7463
rect 26237 7423 26295 7429
rect 26329 7463 26387 7469
rect 26329 7429 26341 7463
rect 26375 7429 26387 7463
rect 26329 7423 26387 7429
rect 23477 7395 23535 7401
rect 23477 7361 23489 7395
rect 23523 7361 23535 7395
rect 23477 7355 23535 7361
rect 24854 7352 24860 7404
rect 24912 7392 24918 7404
rect 25222 7392 25228 7404
rect 24912 7364 25228 7392
rect 24912 7352 24918 7364
rect 25222 7352 25228 7364
rect 25280 7352 25286 7404
rect 26988 7401 27016 7500
rect 27154 7420 27160 7472
rect 27212 7420 27218 7472
rect 27249 7463 27307 7469
rect 27249 7429 27261 7463
rect 27295 7460 27307 7463
rect 28261 7463 28319 7469
rect 28261 7460 28273 7463
rect 27295 7432 28273 7460
rect 27295 7429 27307 7432
rect 27249 7423 27307 7429
rect 28261 7429 28273 7432
rect 28307 7429 28319 7463
rect 28261 7423 28319 7429
rect 28350 7420 28356 7472
rect 28408 7460 28414 7472
rect 29546 7460 29552 7472
rect 28408 7432 28580 7460
rect 28408 7420 28414 7432
rect 26053 7395 26111 7401
rect 26053 7361 26065 7395
rect 26099 7361 26111 7395
rect 26053 7355 26111 7361
rect 26467 7395 26525 7401
rect 26467 7361 26479 7395
rect 26513 7392 26525 7395
rect 26973 7395 27031 7401
rect 26513 7364 26924 7392
rect 26513 7361 26525 7364
rect 26467 7355 26525 7361
rect 16684 7324 16712 7352
rect 15948 7296 16712 7324
rect 19426 7284 19432 7336
rect 19484 7324 19490 7336
rect 20165 7327 20223 7333
rect 20165 7324 20177 7327
rect 19484 7296 20177 7324
rect 19484 7284 19490 7296
rect 20165 7293 20177 7296
rect 20211 7293 20223 7327
rect 20165 7287 20223 7293
rect 20993 7327 21051 7333
rect 20993 7293 21005 7327
rect 21039 7324 21051 7327
rect 21545 7327 21603 7333
rect 21545 7324 21557 7327
rect 21039 7296 21557 7324
rect 21039 7293 21051 7296
rect 20993 7287 21051 7293
rect 21545 7293 21557 7296
rect 21591 7293 21603 7327
rect 21545 7287 21603 7293
rect 13872 7228 15332 7256
rect 13872 7216 13878 7228
rect 8536 7160 12112 7188
rect 8536 7148 8542 7160
rect 15470 7148 15476 7200
rect 15528 7148 15534 7200
rect 15562 7148 15568 7200
rect 15620 7188 15626 7200
rect 16298 7188 16304 7200
rect 15620 7160 16304 7188
rect 15620 7148 15626 7160
rect 16298 7148 16304 7160
rect 16356 7148 16362 7200
rect 21453 7191 21511 7197
rect 21453 7157 21465 7191
rect 21499 7188 21511 7191
rect 21913 7191 21971 7197
rect 21913 7188 21925 7191
rect 21499 7160 21925 7188
rect 21499 7157 21511 7160
rect 21453 7151 21511 7157
rect 21913 7157 21925 7160
rect 21959 7157 21971 7191
rect 22112 7188 22140 7352
rect 23753 7327 23811 7333
rect 23753 7293 23765 7327
rect 23799 7324 23811 7327
rect 26068 7324 26096 7355
rect 26786 7324 26792 7336
rect 23799 7296 25176 7324
rect 26068 7296 26792 7324
rect 23799 7293 23811 7296
rect 23753 7287 23811 7293
rect 25148 7256 25176 7296
rect 26786 7284 26792 7296
rect 26844 7284 26850 7336
rect 26896 7324 26924 7364
rect 26973 7361 26985 7395
rect 27019 7361 27031 7395
rect 26973 7355 27031 7361
rect 27341 7395 27399 7401
rect 27341 7361 27353 7395
rect 27387 7392 27399 7395
rect 27430 7392 27436 7404
rect 27387 7364 27436 7392
rect 27387 7361 27399 7364
rect 27341 7355 27399 7361
rect 27356 7324 27384 7355
rect 27430 7352 27436 7364
rect 27488 7352 27494 7404
rect 27614 7352 27620 7404
rect 27672 7352 27678 7404
rect 28552 7401 28580 7432
rect 28920 7432 29552 7460
rect 28920 7401 28948 7432
rect 29546 7420 29552 7432
rect 29604 7460 29610 7472
rect 29604 7432 30880 7460
rect 29604 7420 29610 7432
rect 28537 7395 28595 7401
rect 28537 7361 28549 7395
rect 28583 7361 28595 7395
rect 28721 7395 28779 7401
rect 28721 7392 28733 7395
rect 28537 7355 28595 7361
rect 28644 7364 28733 7392
rect 28644 7336 28672 7364
rect 28721 7361 28733 7364
rect 28767 7361 28779 7395
rect 28721 7355 28779 7361
rect 28813 7395 28871 7401
rect 28813 7361 28825 7395
rect 28859 7361 28871 7395
rect 28813 7355 28871 7361
rect 28905 7395 28963 7401
rect 28905 7361 28917 7395
rect 28951 7361 28963 7395
rect 28905 7355 28963 7361
rect 26896 7296 27384 7324
rect 28626 7284 28632 7336
rect 28684 7284 28690 7336
rect 28828 7324 28856 7355
rect 29178 7352 29184 7404
rect 29236 7352 29242 7404
rect 29270 7352 29276 7404
rect 29328 7392 29334 7404
rect 29365 7395 29423 7401
rect 29365 7392 29377 7395
rect 29328 7364 29377 7392
rect 29328 7352 29334 7364
rect 29365 7361 29377 7364
rect 29411 7361 29423 7395
rect 29365 7355 29423 7361
rect 29454 7352 29460 7404
rect 29512 7392 29518 7404
rect 29641 7395 29699 7401
rect 29641 7392 29653 7395
rect 29512 7364 29653 7392
rect 29512 7352 29518 7364
rect 29641 7361 29653 7364
rect 29687 7361 29699 7395
rect 29641 7355 29699 7361
rect 29822 7352 29828 7404
rect 29880 7352 29886 7404
rect 29914 7352 29920 7404
rect 29972 7352 29978 7404
rect 30208 7401 30236 7432
rect 30193 7395 30251 7401
rect 30193 7361 30205 7395
rect 30239 7361 30251 7395
rect 30193 7355 30251 7361
rect 30282 7352 30288 7404
rect 30340 7392 30346 7404
rect 30377 7395 30435 7401
rect 30377 7392 30389 7395
rect 30340 7364 30389 7392
rect 30340 7352 30346 7364
rect 30377 7361 30389 7364
rect 30423 7361 30435 7395
rect 30377 7355 30435 7361
rect 28828 7296 28948 7324
rect 26605 7259 26663 7265
rect 26605 7256 26617 7259
rect 25148 7228 26617 7256
rect 26605 7225 26617 7228
rect 26651 7225 26663 7259
rect 28920 7256 28948 7296
rect 29086 7284 29092 7336
rect 29144 7284 29150 7336
rect 29840 7324 29868 7352
rect 30009 7327 30067 7333
rect 30009 7324 30021 7327
rect 29472 7296 30021 7324
rect 28920 7228 29132 7256
rect 26605 7219 26663 7225
rect 27246 7188 27252 7200
rect 22112 7160 27252 7188
rect 21913 7151 21971 7157
rect 27246 7148 27252 7160
rect 27304 7148 27310 7200
rect 27522 7148 27528 7200
rect 27580 7148 27586 7200
rect 28626 7148 28632 7200
rect 28684 7148 28690 7200
rect 28902 7148 28908 7200
rect 28960 7188 28966 7200
rect 28997 7191 29055 7197
rect 28997 7188 29009 7191
rect 28960 7160 29009 7188
rect 28960 7148 28966 7160
rect 28997 7157 29009 7160
rect 29043 7157 29055 7191
rect 29104 7188 29132 7228
rect 29472 7188 29500 7296
rect 30009 7293 30021 7296
rect 30055 7293 30067 7327
rect 30392 7324 30420 7355
rect 30466 7352 30472 7404
rect 30524 7392 30530 7404
rect 30561 7395 30619 7401
rect 30561 7392 30573 7395
rect 30524 7364 30573 7392
rect 30524 7352 30530 7364
rect 30561 7361 30573 7364
rect 30607 7361 30619 7395
rect 30561 7355 30619 7361
rect 30650 7352 30656 7404
rect 30708 7392 30714 7404
rect 30852 7401 30880 7432
rect 31036 7432 31524 7460
rect 30745 7395 30803 7401
rect 30745 7392 30757 7395
rect 30708 7364 30757 7392
rect 30708 7352 30714 7364
rect 30745 7361 30757 7364
rect 30791 7361 30803 7395
rect 30745 7355 30803 7361
rect 30837 7395 30895 7401
rect 30837 7361 30849 7395
rect 30883 7361 30895 7395
rect 30837 7355 30895 7361
rect 30926 7352 30932 7404
rect 30984 7392 30990 7404
rect 31036 7401 31064 7432
rect 31021 7395 31079 7401
rect 31021 7392 31033 7395
rect 30984 7364 31033 7392
rect 30984 7352 30990 7364
rect 31021 7361 31033 7364
rect 31067 7361 31079 7395
rect 31021 7355 31079 7361
rect 31202 7352 31208 7404
rect 31260 7392 31266 7404
rect 31496 7401 31524 7432
rect 31570 7420 31576 7472
rect 31628 7420 31634 7472
rect 31803 7429 31861 7435
rect 31803 7426 31815 7429
rect 31297 7395 31355 7401
rect 31297 7392 31309 7395
rect 31260 7364 31309 7392
rect 31260 7352 31266 7364
rect 31297 7361 31309 7364
rect 31343 7361 31355 7395
rect 31297 7355 31355 7361
rect 31481 7395 31539 7401
rect 31481 7361 31493 7395
rect 31527 7392 31539 7395
rect 31662 7392 31668 7404
rect 31527 7364 31668 7392
rect 31527 7361 31539 7364
rect 31481 7355 31539 7361
rect 31662 7352 31668 7364
rect 31720 7352 31726 7404
rect 31793 7395 31815 7426
rect 31849 7395 31861 7429
rect 32030 7420 32036 7472
rect 32088 7420 32094 7472
rect 32122 7420 32128 7472
rect 32180 7460 32186 7472
rect 32401 7463 32459 7469
rect 32401 7460 32413 7463
rect 32180 7432 32413 7460
rect 32180 7420 32186 7432
rect 32401 7429 32413 7432
rect 32447 7429 32459 7463
rect 32401 7423 32459 7429
rect 32490 7420 32496 7472
rect 32548 7420 32554 7472
rect 32600 7469 32628 7500
rect 34330 7488 34336 7500
rect 34388 7488 34394 7540
rect 35066 7488 35072 7540
rect 35124 7488 35130 7540
rect 35710 7528 35716 7540
rect 35504 7500 35716 7528
rect 32600 7463 32669 7469
rect 32600 7432 32623 7463
rect 32611 7429 32623 7432
rect 32657 7429 32669 7463
rect 33505 7463 33563 7469
rect 33505 7460 33517 7463
rect 32611 7423 32669 7429
rect 32876 7432 33517 7460
rect 31793 7392 31861 7395
rect 32048 7392 32076 7420
rect 31793 7364 32076 7392
rect 32309 7395 32367 7401
rect 31793 7324 31821 7364
rect 32309 7361 32321 7395
rect 32355 7392 32367 7395
rect 32355 7364 32674 7392
rect 32355 7361 32367 7364
rect 32309 7355 32367 7361
rect 30392 7316 30512 7324
rect 30576 7316 31821 7324
rect 30392 7296 31821 7316
rect 30009 7287 30067 7293
rect 30484 7288 30604 7296
rect 32030 7284 32036 7336
rect 32088 7324 32094 7336
rect 32646 7324 32674 7364
rect 32766 7352 32772 7404
rect 32824 7352 32830 7404
rect 32876 7324 32904 7432
rect 33505 7429 33517 7432
rect 33551 7429 33563 7463
rect 33505 7423 33563 7429
rect 33686 7420 33692 7472
rect 33744 7460 33750 7472
rect 34974 7460 34980 7472
rect 33744 7432 34980 7460
rect 33744 7420 33750 7432
rect 33045 7395 33103 7401
rect 33045 7361 33057 7395
rect 33091 7392 33103 7395
rect 33134 7392 33140 7404
rect 33091 7364 33140 7392
rect 33091 7361 33103 7364
rect 33045 7355 33103 7361
rect 33134 7352 33140 7364
rect 33192 7352 33198 7404
rect 33226 7352 33232 7404
rect 33284 7352 33290 7404
rect 33410 7352 33416 7404
rect 33468 7352 33474 7404
rect 33597 7395 33655 7401
rect 33597 7361 33609 7395
rect 33643 7392 33655 7395
rect 33870 7392 33876 7404
rect 33643 7364 33876 7392
rect 33643 7361 33655 7364
rect 33597 7355 33655 7361
rect 33870 7352 33876 7364
rect 33928 7352 33934 7404
rect 34716 7401 34744 7432
rect 34974 7420 34980 7432
rect 35032 7420 35038 7472
rect 35084 7460 35112 7488
rect 35342 7460 35348 7472
rect 35084 7432 35348 7460
rect 35342 7420 35348 7432
rect 35400 7420 35406 7472
rect 34517 7395 34575 7401
rect 34517 7361 34529 7395
rect 34563 7361 34575 7395
rect 34517 7355 34575 7361
rect 34701 7395 34759 7401
rect 34701 7361 34713 7395
rect 34747 7361 34759 7395
rect 34701 7355 34759 7361
rect 34793 7395 34851 7401
rect 34793 7361 34805 7395
rect 34839 7392 34851 7395
rect 34882 7392 34888 7404
rect 34839 7364 34888 7392
rect 34839 7361 34851 7364
rect 34793 7355 34851 7361
rect 32088 7296 32444 7324
rect 32646 7296 32904 7324
rect 33244 7324 33272 7352
rect 33321 7327 33379 7333
rect 33321 7324 33333 7327
rect 33244 7296 33333 7324
rect 32088 7284 32094 7296
rect 29549 7259 29607 7265
rect 29549 7225 29561 7259
rect 29595 7256 29607 7259
rect 29638 7256 29644 7268
rect 29595 7228 29644 7256
rect 29595 7225 29607 7228
rect 29549 7219 29607 7225
rect 29638 7216 29644 7228
rect 29696 7216 29702 7268
rect 30374 7216 30380 7268
rect 30432 7216 30438 7268
rect 30837 7259 30895 7265
rect 30837 7225 30849 7259
rect 30883 7256 30895 7259
rect 31941 7259 31999 7265
rect 30883 7228 31800 7256
rect 30883 7225 30895 7228
rect 30837 7219 30895 7225
rect 29104 7160 29500 7188
rect 30561 7191 30619 7197
rect 28997 7151 29055 7157
rect 30561 7157 30573 7191
rect 30607 7188 30619 7191
rect 30742 7188 30748 7200
rect 30607 7160 30748 7188
rect 30607 7157 30619 7160
rect 30561 7151 30619 7157
rect 30742 7148 30748 7160
rect 30800 7188 30806 7200
rect 31202 7188 31208 7200
rect 30800 7160 31208 7188
rect 30800 7148 30806 7160
rect 31202 7148 31208 7160
rect 31260 7148 31266 7200
rect 31294 7148 31300 7200
rect 31352 7148 31358 7200
rect 31772 7197 31800 7228
rect 31941 7225 31953 7259
rect 31987 7256 31999 7259
rect 32416 7256 32444 7296
rect 33321 7293 33333 7296
rect 33367 7293 33379 7327
rect 33321 7287 33379 7293
rect 34532 7324 34560 7355
rect 34882 7352 34888 7364
rect 34940 7352 34946 7404
rect 35069 7395 35127 7401
rect 35069 7361 35081 7395
rect 35115 7392 35127 7395
rect 35158 7392 35164 7404
rect 35115 7364 35164 7392
rect 35115 7361 35127 7364
rect 35069 7355 35127 7361
rect 35158 7352 35164 7364
rect 35216 7352 35222 7404
rect 35250 7352 35256 7404
rect 35308 7352 35314 7404
rect 35268 7324 35296 7352
rect 34532 7296 35296 7324
rect 34532 7256 34560 7296
rect 31987 7228 32352 7256
rect 32416 7228 34560 7256
rect 31987 7225 31999 7228
rect 31941 7219 31999 7225
rect 32324 7200 32352 7228
rect 34882 7216 34888 7268
rect 34940 7216 34946 7268
rect 34974 7216 34980 7268
rect 35032 7256 35038 7268
rect 35504 7256 35532 7500
rect 35710 7488 35716 7500
rect 35768 7488 35774 7540
rect 36170 7488 36176 7540
rect 36228 7528 36234 7540
rect 36446 7528 36452 7540
rect 36228 7500 36452 7528
rect 36228 7488 36234 7500
rect 36446 7488 36452 7500
rect 36504 7488 36510 7540
rect 36906 7488 36912 7540
rect 36964 7488 36970 7540
rect 35805 7463 35863 7469
rect 35805 7460 35817 7463
rect 35575 7429 35633 7435
rect 35575 7426 35587 7429
rect 35560 7395 35587 7426
rect 35621 7395 35633 7429
rect 35728 7432 35817 7460
rect 35728 7404 35756 7432
rect 35805 7429 35817 7432
rect 35851 7429 35863 7463
rect 35805 7423 35863 7429
rect 35986 7420 35992 7472
rect 36044 7460 36050 7472
rect 36924 7460 36952 7488
rect 36044 7432 36952 7460
rect 36044 7420 36050 7432
rect 35560 7389 35633 7395
rect 35560 7324 35588 7389
rect 35710 7352 35716 7404
rect 35768 7352 35774 7404
rect 36446 7352 36452 7404
rect 36504 7352 36510 7404
rect 35560 7296 35664 7324
rect 35032 7228 35532 7256
rect 35032 7216 35038 7228
rect 31757 7191 31815 7197
rect 31757 7157 31769 7191
rect 31803 7157 31815 7191
rect 31757 7151 31815 7157
rect 32122 7148 32128 7200
rect 32180 7148 32186 7200
rect 32306 7148 32312 7200
rect 32364 7148 32370 7200
rect 32398 7148 32404 7200
rect 32456 7188 32462 7200
rect 32861 7191 32919 7197
rect 32861 7188 32873 7191
rect 32456 7160 32873 7188
rect 32456 7148 32462 7160
rect 32861 7157 32873 7160
rect 32907 7157 32919 7191
rect 32861 7151 32919 7157
rect 33229 7191 33287 7197
rect 33229 7157 33241 7191
rect 33275 7188 33287 7191
rect 33778 7188 33784 7200
rect 33275 7160 33784 7188
rect 33275 7157 33287 7160
rect 33229 7151 33287 7157
rect 33778 7148 33784 7160
rect 33836 7148 33842 7200
rect 34517 7191 34575 7197
rect 34517 7157 34529 7191
rect 34563 7188 34575 7191
rect 34790 7188 34796 7200
rect 34563 7160 34796 7188
rect 34563 7157 34575 7160
rect 34517 7151 34575 7157
rect 34790 7148 34796 7160
rect 34848 7148 34854 7200
rect 34900 7188 34928 7216
rect 35636 7200 35664 7296
rect 35710 7216 35716 7268
rect 35768 7216 35774 7268
rect 35489 7191 35547 7197
rect 35489 7188 35501 7191
rect 34900 7160 35501 7188
rect 35489 7157 35501 7160
rect 35535 7157 35547 7191
rect 35489 7151 35547 7157
rect 35618 7148 35624 7200
rect 35676 7148 35682 7200
rect 35894 7148 35900 7200
rect 35952 7188 35958 7200
rect 35989 7191 36047 7197
rect 35989 7188 36001 7191
rect 35952 7160 36001 7188
rect 35952 7148 35958 7160
rect 35989 7157 36001 7160
rect 36035 7157 36047 7191
rect 35989 7151 36047 7157
rect 36538 7148 36544 7200
rect 36596 7148 36602 7200
rect 1104 7098 41400 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 41400 7098
rect 1104 7024 41400 7046
rect 7558 6944 7564 6996
rect 7616 6984 7622 6996
rect 8573 6987 8631 6993
rect 8573 6984 8585 6987
rect 7616 6956 8585 6984
rect 7616 6944 7622 6956
rect 8573 6953 8585 6956
rect 8619 6953 8631 6987
rect 8573 6947 8631 6953
rect 11422 6944 11428 6996
rect 11480 6984 11486 6996
rect 12161 6987 12219 6993
rect 12161 6984 12173 6987
rect 11480 6956 12173 6984
rect 11480 6944 11486 6956
rect 12161 6953 12173 6956
rect 12207 6984 12219 6987
rect 12618 6984 12624 6996
rect 12207 6956 12624 6984
rect 12207 6953 12219 6956
rect 12161 6947 12219 6953
rect 12618 6944 12624 6956
rect 12676 6944 12682 6996
rect 12802 6944 12808 6996
rect 12860 6984 12866 6996
rect 12989 6987 13047 6993
rect 12989 6984 13001 6987
rect 12860 6956 13001 6984
rect 12860 6944 12866 6956
rect 12989 6953 13001 6956
rect 13035 6953 13047 6987
rect 14921 6987 14979 6993
rect 14921 6984 14933 6987
rect 12989 6947 13047 6953
rect 13832 6956 14933 6984
rect 6840 6888 7236 6916
rect 1854 6740 1860 6792
rect 1912 6780 1918 6792
rect 4062 6780 4068 6792
rect 1912 6752 4068 6780
rect 1912 6740 1918 6752
rect 4062 6740 4068 6752
rect 4120 6780 4126 6792
rect 5166 6780 5172 6792
rect 4120 6752 5172 6780
rect 4120 6740 4126 6752
rect 5166 6740 5172 6752
rect 5224 6740 5230 6792
rect 6546 6740 6552 6792
rect 6604 6780 6610 6792
rect 6840 6780 6868 6888
rect 6917 6851 6975 6857
rect 6917 6817 6929 6851
rect 6963 6848 6975 6851
rect 7208 6848 7236 6888
rect 8202 6876 8208 6928
rect 8260 6916 8266 6928
rect 10318 6916 10324 6928
rect 8260 6888 10324 6916
rect 8260 6876 8266 6888
rect 10318 6876 10324 6888
rect 10376 6876 10382 6928
rect 12713 6919 12771 6925
rect 12713 6916 12725 6919
rect 12360 6888 12725 6916
rect 12360 6848 12388 6888
rect 12713 6885 12725 6888
rect 12759 6885 12771 6919
rect 12713 6879 12771 6885
rect 13173 6919 13231 6925
rect 13173 6885 13185 6919
rect 13219 6885 13231 6919
rect 13173 6879 13231 6885
rect 6963 6820 7144 6848
rect 7208 6820 9720 6848
rect 6963 6817 6975 6820
rect 6917 6811 6975 6817
rect 7116 6789 7144 6820
rect 9692 6792 9720 6820
rect 11624 6820 12388 6848
rect 12437 6851 12495 6857
rect 6604 6752 6868 6780
rect 7101 6783 7159 6789
rect 6604 6740 6610 6752
rect 7101 6749 7113 6783
rect 7147 6780 7159 6783
rect 7282 6780 7288 6792
rect 7147 6752 7288 6780
rect 7147 6749 7159 6752
rect 7101 6743 7159 6749
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 8021 6783 8079 6789
rect 8021 6780 8033 6783
rect 7524 6752 8033 6780
rect 7524 6740 7530 6752
rect 8021 6749 8033 6752
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 8478 6740 8484 6792
rect 8536 6740 8542 6792
rect 8662 6740 8668 6792
rect 8720 6740 8726 6792
rect 8757 6783 8815 6789
rect 8757 6749 8769 6783
rect 8803 6780 8815 6783
rect 8846 6780 8852 6792
rect 8803 6752 8852 6780
rect 8803 6749 8815 6752
rect 8757 6743 8815 6749
rect 8846 6740 8852 6752
rect 8904 6740 8910 6792
rect 9674 6740 9680 6792
rect 9732 6740 9738 6792
rect 11238 6740 11244 6792
rect 11296 6740 11302 6792
rect 11330 6740 11336 6792
rect 11388 6740 11394 6792
rect 11514 6789 11520 6792
rect 11481 6783 11520 6789
rect 11481 6749 11493 6783
rect 11481 6743 11520 6749
rect 11514 6740 11520 6743
rect 11572 6740 11578 6792
rect 11624 6789 11652 6820
rect 12437 6817 12449 6851
rect 12483 6848 12495 6851
rect 13188 6848 13216 6879
rect 12483 6820 13216 6848
rect 13357 6851 13415 6857
rect 12483 6817 12495 6820
rect 12437 6811 12495 6817
rect 13357 6817 13369 6851
rect 13403 6848 13415 6851
rect 13832 6848 13860 6956
rect 14921 6953 14933 6956
rect 14967 6953 14979 6987
rect 14921 6947 14979 6953
rect 15470 6944 15476 6996
rect 15528 6984 15534 6996
rect 15914 6987 15972 6993
rect 15914 6984 15926 6987
rect 15528 6956 15926 6984
rect 15528 6944 15534 6956
rect 15914 6953 15926 6956
rect 15960 6953 15972 6987
rect 15914 6947 15972 6953
rect 26316 6987 26374 6993
rect 26316 6953 26328 6987
rect 26362 6984 26374 6987
rect 27522 6984 27528 6996
rect 26362 6956 27528 6984
rect 26362 6953 26374 6956
rect 26316 6947 26374 6953
rect 27522 6944 27528 6956
rect 27580 6944 27586 6996
rect 27614 6944 27620 6996
rect 27672 6984 27678 6996
rect 27801 6987 27859 6993
rect 27801 6984 27813 6987
rect 27672 6956 27813 6984
rect 27672 6944 27678 6956
rect 27801 6953 27813 6956
rect 27847 6953 27859 6987
rect 27801 6947 27859 6953
rect 28166 6944 28172 6996
rect 28224 6984 28230 6996
rect 28813 6987 28871 6993
rect 28813 6984 28825 6987
rect 28224 6956 28825 6984
rect 28224 6944 28230 6956
rect 28813 6953 28825 6956
rect 28859 6953 28871 6987
rect 29178 6984 29184 6996
rect 28813 6947 28871 6953
rect 28966 6956 29184 6984
rect 27706 6876 27712 6928
rect 27764 6916 27770 6928
rect 28184 6916 28212 6944
rect 27764 6888 28212 6916
rect 27764 6876 27770 6888
rect 28626 6876 28632 6928
rect 28684 6916 28690 6928
rect 28966 6916 28994 6956
rect 29178 6944 29184 6956
rect 29236 6984 29242 6996
rect 29733 6987 29791 6993
rect 29733 6984 29745 6987
rect 29236 6956 29745 6984
rect 29236 6944 29242 6956
rect 29733 6953 29745 6956
rect 29779 6953 29791 6987
rect 32030 6984 32036 6996
rect 29733 6947 29791 6953
rect 29837 6956 32036 6984
rect 28684 6888 28994 6916
rect 29273 6919 29331 6925
rect 28684 6876 28690 6888
rect 29273 6885 29285 6919
rect 29319 6916 29331 6919
rect 29638 6916 29644 6928
rect 29319 6888 29644 6916
rect 29319 6885 29331 6888
rect 29273 6879 29331 6885
rect 29638 6876 29644 6888
rect 29696 6916 29702 6928
rect 29837 6916 29865 6956
rect 32030 6944 32036 6956
rect 32088 6944 32094 6996
rect 32214 6944 32220 6996
rect 32272 6944 32278 6996
rect 32306 6944 32312 6996
rect 32364 6984 32370 6996
rect 34146 6984 34152 6996
rect 32364 6956 34152 6984
rect 32364 6944 32370 6956
rect 29696 6888 29865 6916
rect 29696 6876 29702 6888
rect 31662 6876 31668 6928
rect 31720 6916 31726 6928
rect 31720 6888 32352 6916
rect 31720 6876 31726 6888
rect 13403 6820 13860 6848
rect 13403 6817 13415 6820
rect 13357 6811 13415 6817
rect 14274 6808 14280 6860
rect 14332 6848 14338 6860
rect 14645 6851 14703 6857
rect 14645 6848 14657 6851
rect 14332 6820 14657 6848
rect 14332 6808 14338 6820
rect 14645 6817 14657 6820
rect 14691 6817 14703 6851
rect 14645 6811 14703 6817
rect 15010 6808 15016 6860
rect 15068 6808 15074 6860
rect 15657 6851 15715 6857
rect 15657 6817 15669 6851
rect 15703 6848 15715 6851
rect 16298 6848 16304 6860
rect 15703 6820 16304 6848
rect 15703 6817 15715 6820
rect 15657 6811 15715 6817
rect 16298 6808 16304 6820
rect 16356 6808 16362 6860
rect 17310 6808 17316 6860
rect 17368 6848 17374 6860
rect 17405 6851 17463 6857
rect 17405 6848 17417 6851
rect 17368 6820 17417 6848
rect 17368 6808 17374 6820
rect 17405 6817 17417 6820
rect 17451 6817 17463 6851
rect 17405 6811 17463 6817
rect 18414 6808 18420 6860
rect 18472 6808 18478 6860
rect 19058 6808 19064 6860
rect 19116 6848 19122 6860
rect 20898 6848 20904 6860
rect 19116 6820 20904 6848
rect 19116 6808 19122 6820
rect 20898 6808 20904 6820
rect 20956 6808 20962 6860
rect 21192 6820 21772 6848
rect 11609 6783 11667 6789
rect 11609 6749 11621 6783
rect 11655 6749 11667 6783
rect 11609 6743 11667 6749
rect 11798 6783 11856 6789
rect 11798 6749 11810 6783
rect 11844 6749 11856 6783
rect 11798 6743 11856 6749
rect 12529 6783 12587 6789
rect 12529 6749 12541 6783
rect 12575 6780 12587 6783
rect 13265 6783 13323 6789
rect 12575 6752 12940 6780
rect 12575 6749 12587 6752
rect 12529 6743 12587 6749
rect 5445 6715 5503 6721
rect 5445 6681 5457 6715
rect 5491 6712 5503 6715
rect 5534 6712 5540 6724
rect 5491 6684 5540 6712
rect 5491 6681 5503 6684
rect 5445 6675 5503 6681
rect 5534 6672 5540 6684
rect 5592 6672 5598 6724
rect 7374 6672 7380 6724
rect 7432 6712 7438 6724
rect 8205 6715 8263 6721
rect 8205 6712 8217 6715
rect 7432 6684 8217 6712
rect 7432 6672 7438 6684
rect 8205 6681 8217 6684
rect 8251 6681 8263 6715
rect 10962 6712 10968 6724
rect 8205 6675 8263 6681
rect 8312 6684 10968 6712
rect 7650 6604 7656 6656
rect 7708 6604 7714 6656
rect 7926 6604 7932 6656
rect 7984 6644 7990 6656
rect 8312 6644 8340 6684
rect 10962 6672 10968 6684
rect 11020 6672 11026 6724
rect 11256 6712 11284 6740
rect 11698 6712 11704 6724
rect 11256 6684 11704 6712
rect 11698 6672 11704 6684
rect 11756 6672 11762 6724
rect 7984 6616 8340 6644
rect 7984 6604 7990 6616
rect 8386 6604 8392 6656
rect 8444 6604 8450 6656
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 11808 6644 11836 6743
rect 12066 6672 12072 6724
rect 12124 6672 12130 6724
rect 12250 6672 12256 6724
rect 12308 6712 12314 6724
rect 12805 6715 12863 6721
rect 12805 6712 12817 6715
rect 12308 6684 12817 6712
rect 12308 6672 12314 6684
rect 12805 6681 12817 6684
rect 12851 6681 12863 6715
rect 12805 6675 12863 6681
rect 11204 6616 11836 6644
rect 11204 6604 11210 6616
rect 11974 6604 11980 6656
rect 12032 6604 12038 6656
rect 12912 6644 12940 6752
rect 13265 6749 13277 6783
rect 13311 6749 13323 6783
rect 13265 6743 13323 6749
rect 13449 6783 13507 6789
rect 13449 6749 13461 6783
rect 13495 6780 13507 6783
rect 13630 6780 13636 6792
rect 13495 6752 13636 6780
rect 13495 6749 13507 6752
rect 13449 6743 13507 6749
rect 12986 6672 12992 6724
rect 13044 6721 13050 6724
rect 13044 6715 13068 6721
rect 13056 6712 13068 6715
rect 13280 6712 13308 6743
rect 13630 6740 13636 6752
rect 13688 6740 13694 6792
rect 13722 6740 13728 6792
rect 13780 6740 13786 6792
rect 13998 6740 14004 6792
rect 14056 6780 14062 6792
rect 14461 6783 14519 6789
rect 14461 6780 14473 6783
rect 14056 6752 14473 6780
rect 14056 6740 14062 6752
rect 14461 6749 14473 6752
rect 14507 6749 14519 6783
rect 14461 6743 14519 6749
rect 14921 6783 14979 6789
rect 14921 6749 14933 6783
rect 14967 6749 14979 6783
rect 14921 6743 14979 6749
rect 13538 6712 13544 6724
rect 13056 6684 13544 6712
rect 13056 6681 13068 6684
rect 13044 6675 13068 6681
rect 13044 6672 13050 6675
rect 13538 6672 13544 6684
rect 13596 6672 13602 6724
rect 13909 6715 13967 6721
rect 13909 6681 13921 6715
rect 13955 6712 13967 6715
rect 14936 6712 14964 6743
rect 17494 6740 17500 6792
rect 17552 6780 17558 6792
rect 17552 6752 18000 6780
rect 17552 6740 17558 6752
rect 17862 6712 17868 6724
rect 13955 6684 14964 6712
rect 17158 6684 17868 6712
rect 13955 6681 13967 6684
rect 13909 6675 13967 6681
rect 17862 6672 17868 6684
rect 17920 6672 17926 6724
rect 17972 6712 18000 6752
rect 18046 6740 18052 6792
rect 18104 6780 18110 6792
rect 18233 6783 18291 6789
rect 18233 6780 18245 6783
rect 18104 6752 18245 6780
rect 18104 6740 18110 6752
rect 18233 6749 18245 6752
rect 18279 6749 18291 6783
rect 18233 6743 18291 6749
rect 19426 6740 19432 6792
rect 19484 6740 19490 6792
rect 20073 6783 20131 6789
rect 20073 6749 20085 6783
rect 20119 6780 20131 6783
rect 21082 6780 21088 6792
rect 20119 6752 21088 6780
rect 20119 6749 20131 6752
rect 20073 6743 20131 6749
rect 21082 6740 21088 6752
rect 21140 6740 21146 6792
rect 21192 6712 21220 6820
rect 21744 6789 21772 6820
rect 21818 6808 21824 6860
rect 21876 6808 21882 6860
rect 26050 6848 26056 6860
rect 24504 6820 26056 6848
rect 24504 6792 24532 6820
rect 26050 6808 26056 6820
rect 26108 6808 26114 6860
rect 26786 6808 26792 6860
rect 26844 6848 26850 6860
rect 30374 6848 30380 6860
rect 26844 6820 30380 6848
rect 26844 6808 26850 6820
rect 30374 6808 30380 6820
rect 30432 6808 30438 6860
rect 31478 6808 31484 6860
rect 31536 6848 31542 6860
rect 31849 6851 31907 6857
rect 31849 6848 31861 6851
rect 31536 6820 31861 6848
rect 31536 6808 31542 6820
rect 31849 6817 31861 6820
rect 31895 6817 31907 6851
rect 31849 6811 31907 6817
rect 32033 6851 32091 6857
rect 32033 6817 32045 6851
rect 32079 6848 32091 6851
rect 32122 6848 32128 6860
rect 32079 6820 32128 6848
rect 32079 6817 32091 6820
rect 32033 6811 32091 6817
rect 32122 6808 32128 6820
rect 32180 6808 32186 6860
rect 32324 6857 32352 6888
rect 32490 6876 32496 6928
rect 32548 6876 32554 6928
rect 33137 6919 33195 6925
rect 33137 6885 33149 6919
rect 33183 6916 33195 6919
rect 33502 6916 33508 6928
rect 33183 6888 33508 6916
rect 33183 6885 33195 6888
rect 33137 6879 33195 6885
rect 33502 6876 33508 6888
rect 33560 6876 33566 6928
rect 32309 6851 32367 6857
rect 32309 6817 32321 6851
rect 32355 6817 32367 6851
rect 32508 6848 32536 6876
rect 32508 6820 33456 6848
rect 32309 6811 32367 6817
rect 21729 6783 21787 6789
rect 21545 6773 21603 6779
rect 21545 6739 21557 6773
rect 21591 6739 21603 6773
rect 21729 6749 21741 6783
rect 21775 6749 21787 6783
rect 21729 6743 21787 6749
rect 24486 6740 24492 6792
rect 24544 6740 24550 6792
rect 25409 6783 25467 6789
rect 25409 6749 25421 6783
rect 25455 6780 25467 6783
rect 25455 6752 26004 6780
rect 25455 6749 25467 6752
rect 25409 6743 25467 6749
rect 21545 6733 21603 6739
rect 17972 6684 21220 6712
rect 13814 6644 13820 6656
rect 12912 6616 13820 6644
rect 13814 6604 13820 6616
rect 13872 6604 13878 6656
rect 14090 6604 14096 6656
rect 14148 6604 14154 6656
rect 14550 6604 14556 6656
rect 14608 6604 14614 6656
rect 15286 6604 15292 6656
rect 15344 6604 15350 6656
rect 18690 6604 18696 6656
rect 18748 6644 18754 6656
rect 19245 6647 19303 6653
rect 19245 6644 19257 6647
rect 18748 6616 19257 6644
rect 18748 6604 18754 6616
rect 19245 6613 19257 6616
rect 19291 6613 19303 6647
rect 19245 6607 19303 6613
rect 20438 6604 20444 6656
rect 20496 6644 20502 6656
rect 20625 6647 20683 6653
rect 20625 6644 20637 6647
rect 20496 6616 20637 6644
rect 20496 6604 20502 6616
rect 20625 6613 20637 6616
rect 20671 6613 20683 6647
rect 21560 6644 21588 6733
rect 21637 6715 21695 6721
rect 21637 6681 21649 6715
rect 21683 6712 21695 6715
rect 22097 6715 22155 6721
rect 22097 6712 22109 6715
rect 21683 6684 22109 6712
rect 21683 6681 21695 6684
rect 21637 6675 21695 6681
rect 22097 6681 22109 6684
rect 22143 6681 22155 6715
rect 22097 6675 22155 6681
rect 22554 6672 22560 6724
rect 22612 6672 22618 6724
rect 23842 6672 23848 6724
rect 23900 6712 23906 6724
rect 25774 6712 25780 6724
rect 23900 6684 25780 6712
rect 23900 6672 23906 6684
rect 25774 6672 25780 6684
rect 25832 6672 25838 6724
rect 25976 6712 26004 6752
rect 27430 6740 27436 6792
rect 27488 6740 27494 6792
rect 28718 6740 28724 6792
rect 28776 6740 28782 6792
rect 28902 6740 28908 6792
rect 28960 6740 28966 6792
rect 29181 6783 29239 6789
rect 29181 6749 29193 6783
rect 29227 6749 29239 6783
rect 29181 6743 29239 6749
rect 26234 6712 26240 6724
rect 25976 6684 26240 6712
rect 26234 6672 26240 6684
rect 26292 6672 26298 6724
rect 28629 6715 28687 6721
rect 28629 6681 28641 6715
rect 28675 6712 28687 6715
rect 28736 6712 28764 6740
rect 28675 6684 28764 6712
rect 28675 6681 28687 6684
rect 28629 6675 28687 6681
rect 22370 6644 22376 6656
rect 21560 6616 22376 6644
rect 20625 6607 20683 6613
rect 22370 6604 22376 6616
rect 22428 6604 22434 6656
rect 25961 6647 26019 6653
rect 25961 6613 25973 6647
rect 26007 6644 26019 6647
rect 26694 6644 26700 6656
rect 26007 6616 26700 6644
rect 26007 6613 26019 6616
rect 25961 6607 26019 6613
rect 26694 6604 26700 6616
rect 26752 6604 26758 6656
rect 28834 6647 28892 6653
rect 28834 6613 28846 6647
rect 28880 6644 28892 6647
rect 28920 6644 28948 6740
rect 29196 6712 29224 6743
rect 29270 6740 29276 6792
rect 29328 6780 29334 6792
rect 29365 6783 29423 6789
rect 29365 6780 29377 6783
rect 29328 6752 29377 6780
rect 29328 6740 29334 6752
rect 29365 6749 29377 6752
rect 29411 6749 29423 6783
rect 29365 6743 29423 6749
rect 29454 6740 29460 6792
rect 29512 6740 29518 6792
rect 30282 6780 30288 6792
rect 29794 6755 30288 6780
rect 29779 6752 30288 6755
rect 29779 6749 29837 6752
rect 29472 6712 29500 6740
rect 29196 6684 29500 6712
rect 29549 6715 29607 6721
rect 29549 6681 29561 6715
rect 29595 6712 29607 6715
rect 29638 6712 29644 6724
rect 29595 6684 29644 6712
rect 29595 6681 29607 6684
rect 29549 6675 29607 6681
rect 29638 6672 29644 6684
rect 29696 6672 29702 6724
rect 29779 6715 29791 6749
rect 29825 6715 29837 6749
rect 30282 6740 30288 6752
rect 30340 6740 30346 6792
rect 30650 6740 30656 6792
rect 30708 6740 30714 6792
rect 31294 6740 31300 6792
rect 31352 6780 31358 6792
rect 31757 6783 31815 6789
rect 31757 6780 31769 6783
rect 31352 6752 31769 6780
rect 31352 6740 31358 6752
rect 31757 6749 31769 6752
rect 31803 6749 31815 6783
rect 31757 6743 31815 6749
rect 31941 6783 31999 6789
rect 31941 6749 31953 6783
rect 31987 6749 31999 6783
rect 31941 6743 31999 6749
rect 32217 6783 32275 6789
rect 32217 6749 32229 6783
rect 32263 6780 32275 6783
rect 32398 6780 32404 6792
rect 32263 6752 32404 6780
rect 32263 6749 32275 6752
rect 32217 6743 32275 6749
rect 29779 6709 29837 6715
rect 30101 6715 30159 6721
rect 30101 6712 30113 6715
rect 29932 6684 30113 6712
rect 28880 6616 28948 6644
rect 28880 6613 28892 6616
rect 28834 6607 28892 6613
rect 28994 6604 29000 6656
rect 29052 6604 29058 6656
rect 29932 6653 29960 6684
rect 30101 6681 30113 6684
rect 30147 6681 30159 6715
rect 30668 6712 30696 6740
rect 31956 6712 31984 6743
rect 32398 6740 32404 6752
rect 32456 6740 32462 6792
rect 32490 6740 32496 6792
rect 32548 6780 32554 6792
rect 32548 6752 33180 6780
rect 32548 6740 32554 6752
rect 33042 6712 33048 6724
rect 30668 6684 31892 6712
rect 31956 6684 33048 6712
rect 30101 6675 30159 6681
rect 29917 6647 29975 6653
rect 29917 6613 29929 6647
rect 29963 6613 29975 6647
rect 29917 6607 29975 6613
rect 31570 6604 31576 6656
rect 31628 6604 31634 6656
rect 31864 6644 31892 6684
rect 33042 6672 33048 6684
rect 33100 6672 33106 6724
rect 32490 6644 32496 6656
rect 31864 6616 32496 6644
rect 32490 6604 32496 6616
rect 32548 6604 32554 6656
rect 32674 6604 32680 6656
rect 32732 6604 32738 6656
rect 33152 6644 33180 6752
rect 33318 6740 33324 6792
rect 33376 6740 33382 6792
rect 33428 6789 33456 6820
rect 33612 6789 33640 6956
rect 34146 6944 34152 6956
rect 34204 6944 34210 6996
rect 34330 6944 34336 6996
rect 34388 6944 34394 6996
rect 34698 6944 34704 6996
rect 34756 6984 34762 6996
rect 35161 6987 35219 6993
rect 35161 6984 35173 6987
rect 34756 6956 35173 6984
rect 34756 6944 34762 6956
rect 35161 6953 35173 6956
rect 35207 6953 35219 6987
rect 35161 6947 35219 6953
rect 36265 6987 36323 6993
rect 36265 6953 36277 6987
rect 36311 6984 36323 6987
rect 36446 6984 36452 6996
rect 36311 6956 36452 6984
rect 36311 6953 36323 6956
rect 36265 6947 36323 6953
rect 36446 6944 36452 6956
rect 36504 6944 36510 6996
rect 34348 6916 34376 6944
rect 36538 6916 36544 6928
rect 34348 6888 36544 6916
rect 36538 6876 36544 6888
rect 36596 6876 36602 6928
rect 34606 6848 34612 6860
rect 33980 6820 34612 6848
rect 33980 6792 34008 6820
rect 34606 6808 34612 6820
rect 34664 6848 34670 6860
rect 35618 6848 35624 6860
rect 34664 6820 34928 6848
rect 34664 6808 34670 6820
rect 33413 6783 33471 6789
rect 33413 6749 33425 6783
rect 33459 6749 33471 6783
rect 33413 6743 33471 6749
rect 33597 6783 33655 6789
rect 33597 6749 33609 6783
rect 33643 6749 33655 6783
rect 33597 6743 33655 6749
rect 33689 6783 33747 6789
rect 33689 6749 33701 6783
rect 33735 6780 33747 6783
rect 33781 6783 33839 6789
rect 33781 6780 33793 6783
rect 33735 6752 33793 6780
rect 33735 6749 33747 6752
rect 33689 6743 33747 6749
rect 33781 6749 33793 6752
rect 33827 6749 33839 6783
rect 33781 6743 33839 6749
rect 33962 6740 33968 6792
rect 34020 6740 34026 6792
rect 34146 6740 34152 6792
rect 34204 6740 34210 6792
rect 34422 6740 34428 6792
rect 34480 6740 34486 6792
rect 33226 6672 33232 6724
rect 33284 6712 33290 6724
rect 33870 6712 33876 6724
rect 33284 6684 33876 6712
rect 33284 6672 33290 6684
rect 33870 6672 33876 6684
rect 33928 6712 33934 6724
rect 34330 6721 34336 6724
rect 34057 6715 34115 6721
rect 34057 6712 34069 6715
rect 33928 6684 34069 6712
rect 33928 6672 33934 6684
rect 34057 6681 34069 6684
rect 34103 6681 34115 6715
rect 34057 6675 34115 6681
rect 34287 6715 34336 6721
rect 34287 6681 34299 6715
rect 34333 6681 34336 6715
rect 34287 6675 34336 6681
rect 34330 6672 34336 6675
rect 34388 6672 34394 6724
rect 34900 6721 34928 6820
rect 35084 6820 35624 6848
rect 34974 6740 34980 6792
rect 35032 6780 35038 6792
rect 35084 6789 35112 6820
rect 35618 6808 35624 6820
rect 35676 6848 35682 6860
rect 35676 6820 36124 6848
rect 35676 6808 35682 6820
rect 35069 6783 35127 6789
rect 35069 6780 35081 6783
rect 35032 6752 35081 6780
rect 35032 6740 35038 6752
rect 35069 6749 35081 6752
rect 35115 6749 35127 6783
rect 35069 6743 35127 6749
rect 35342 6740 35348 6792
rect 35400 6780 35406 6792
rect 35437 6783 35495 6789
rect 35437 6780 35449 6783
rect 35400 6752 35449 6780
rect 35400 6740 35406 6752
rect 35437 6749 35449 6752
rect 35483 6749 35495 6783
rect 35437 6743 35495 6749
rect 35713 6783 35771 6789
rect 35713 6749 35725 6783
rect 35759 6780 35771 6783
rect 35802 6780 35808 6792
rect 35759 6752 35808 6780
rect 35759 6749 35771 6752
rect 35713 6743 35771 6749
rect 34885 6715 34943 6721
rect 34885 6681 34897 6715
rect 34931 6681 34943 6715
rect 34885 6675 34943 6681
rect 35452 6712 35480 6743
rect 35802 6740 35808 6752
rect 35860 6740 35866 6792
rect 36096 6789 36124 6820
rect 35897 6783 35955 6789
rect 35897 6749 35909 6783
rect 35943 6749 35955 6783
rect 35897 6743 35955 6749
rect 36081 6783 36139 6789
rect 36081 6749 36093 6783
rect 36127 6749 36139 6783
rect 36081 6743 36139 6749
rect 35912 6712 35940 6743
rect 35452 6684 35940 6712
rect 35452 6644 35480 6684
rect 33152 6616 35480 6644
rect 35526 6604 35532 6656
rect 35584 6604 35590 6656
rect 1104 6554 41400 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 41400 6554
rect 1104 6480 41400 6502
rect 5534 6400 5540 6452
rect 5592 6400 5598 6452
rect 6365 6443 6423 6449
rect 6365 6409 6377 6443
rect 6411 6409 6423 6443
rect 6365 6403 6423 6409
rect 6733 6443 6791 6449
rect 6733 6409 6745 6443
rect 6779 6440 6791 6443
rect 7650 6440 7656 6452
rect 6779 6412 7656 6440
rect 6779 6409 6791 6412
rect 6733 6403 6791 6409
rect 5166 6264 5172 6316
rect 5224 6264 5230 6316
rect 5721 6307 5779 6313
rect 5721 6273 5733 6307
rect 5767 6304 5779 6307
rect 6380 6304 6408 6403
rect 7650 6400 7656 6412
rect 7708 6400 7714 6452
rect 8386 6400 8392 6452
rect 8444 6400 8450 6452
rect 10042 6400 10048 6452
rect 10100 6440 10106 6452
rect 10870 6440 10876 6452
rect 10100 6412 10876 6440
rect 10100 6400 10106 6412
rect 10870 6400 10876 6412
rect 10928 6400 10934 6452
rect 11514 6400 11520 6452
rect 11572 6400 11578 6452
rect 11698 6400 11704 6452
rect 11756 6400 11762 6452
rect 12066 6400 12072 6452
rect 12124 6440 12130 6452
rect 12437 6443 12495 6449
rect 12437 6440 12449 6443
rect 12124 6412 12449 6440
rect 12124 6400 12130 6412
rect 12437 6409 12449 6412
rect 12483 6409 12495 6443
rect 12437 6403 12495 6409
rect 12802 6400 12808 6452
rect 12860 6440 12866 6452
rect 13265 6443 13323 6449
rect 13265 6440 13277 6443
rect 12860 6412 13277 6440
rect 12860 6400 12866 6412
rect 13265 6409 13277 6412
rect 13311 6409 13323 6443
rect 13265 6403 13323 6409
rect 13630 6400 13636 6452
rect 13688 6400 13694 6452
rect 14461 6443 14519 6449
rect 14461 6409 14473 6443
rect 14507 6440 14519 6443
rect 14550 6440 14556 6452
rect 14507 6412 14556 6440
rect 14507 6409 14519 6412
rect 14461 6403 14519 6409
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 15286 6400 15292 6452
rect 15344 6400 15350 6452
rect 18325 6443 18383 6449
rect 18325 6409 18337 6443
rect 18371 6440 18383 6443
rect 19426 6440 19432 6452
rect 18371 6412 19432 6440
rect 18371 6409 18383 6412
rect 18325 6403 18383 6409
rect 19426 6400 19432 6412
rect 19484 6400 19490 6452
rect 20438 6400 20444 6452
rect 20496 6440 20502 6452
rect 20533 6443 20591 6449
rect 20533 6440 20545 6443
rect 20496 6412 20545 6440
rect 20496 6400 20502 6412
rect 20533 6409 20545 6412
rect 20579 6409 20591 6443
rect 20533 6403 20591 6409
rect 20622 6400 20628 6452
rect 20680 6400 20686 6452
rect 20732 6412 26096 6440
rect 6825 6375 6883 6381
rect 6825 6341 6837 6375
rect 6871 6372 6883 6375
rect 7926 6372 7932 6384
rect 6871 6344 7932 6372
rect 6871 6341 6883 6344
rect 6825 6335 6883 6341
rect 7926 6332 7932 6344
rect 7984 6332 7990 6384
rect 8404 6372 8432 6400
rect 8036 6344 8432 6372
rect 8036 6313 8064 6344
rect 10318 6332 10324 6384
rect 10376 6332 10382 6384
rect 11146 6372 11152 6384
rect 10704 6344 11152 6372
rect 5767 6276 6408 6304
rect 8021 6307 8079 6313
rect 5767 6273 5779 6276
rect 5721 6267 5779 6273
rect 8021 6273 8033 6307
rect 8067 6273 8079 6307
rect 8297 6307 8355 6313
rect 8297 6304 8309 6307
rect 8021 6267 8079 6273
rect 8128 6276 8309 6304
rect 5184 6168 5212 6264
rect 8128 6248 8156 6276
rect 8297 6273 8309 6276
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 9674 6264 9680 6316
rect 9732 6264 9738 6316
rect 6270 6196 6276 6248
rect 6328 6236 6334 6248
rect 6822 6236 6828 6248
rect 6328 6208 6828 6236
rect 6328 6196 6334 6208
rect 6822 6196 6828 6208
rect 6880 6236 6886 6248
rect 6917 6239 6975 6245
rect 6917 6236 6929 6239
rect 6880 6208 6929 6236
rect 6880 6196 6886 6208
rect 6917 6205 6929 6208
rect 6963 6205 6975 6239
rect 8110 6236 8116 6248
rect 6917 6199 6975 6205
rect 7024 6208 8116 6236
rect 7024 6168 7052 6208
rect 8110 6196 8116 6208
rect 8168 6196 8174 6248
rect 8573 6239 8631 6245
rect 8573 6236 8585 6239
rect 8404 6208 8585 6236
rect 5184 6140 7052 6168
rect 7837 6103 7895 6109
rect 7837 6069 7849 6103
rect 7883 6100 7895 6103
rect 8404 6100 8432 6208
rect 8573 6205 8585 6208
rect 8619 6205 8631 6239
rect 8573 6199 8631 6205
rect 8662 6196 8668 6248
rect 8720 6236 8726 6248
rect 10704 6236 10732 6344
rect 10781 6307 10839 6313
rect 10781 6273 10793 6307
rect 10827 6273 10839 6307
rect 10781 6267 10839 6273
rect 8720 6208 10732 6236
rect 8720 6196 8726 6208
rect 10796 6168 10824 6267
rect 10980 6245 11008 6344
rect 11146 6332 11152 6344
rect 11204 6332 11210 6384
rect 11716 6372 11744 6400
rect 12342 6372 12348 6384
rect 11716 6344 12348 6372
rect 12342 6332 12348 6344
rect 12400 6332 12406 6384
rect 11054 6264 11060 6316
rect 11112 6304 11118 6316
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 11112 6276 11713 6304
rect 11112 6264 11118 6276
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 11790 6264 11796 6316
rect 11848 6304 11854 6316
rect 11977 6307 12035 6313
rect 11977 6304 11989 6307
rect 11848 6276 11989 6304
rect 11848 6264 11854 6276
rect 11977 6273 11989 6276
rect 12023 6273 12035 6307
rect 11977 6267 12035 6273
rect 12069 6307 12127 6313
rect 12069 6273 12081 6307
rect 12115 6304 12127 6307
rect 12986 6304 12992 6316
rect 12115 6276 12992 6304
rect 12115 6273 12127 6276
rect 12069 6267 12127 6273
rect 12986 6264 12992 6276
rect 13044 6264 13050 6316
rect 13173 6307 13231 6313
rect 13173 6273 13185 6307
rect 13219 6304 13231 6307
rect 13648 6304 13676 6400
rect 13219 6276 13676 6304
rect 14093 6307 14151 6313
rect 13219 6273 13231 6276
rect 13173 6267 13231 6273
rect 14093 6273 14105 6307
rect 14139 6304 14151 6307
rect 14366 6304 14372 6316
rect 14139 6276 14372 6304
rect 14139 6273 14151 6276
rect 14093 6267 14151 6273
rect 10965 6239 11023 6245
rect 10965 6205 10977 6239
rect 11011 6205 11023 6239
rect 10965 6199 11023 6205
rect 11606 6196 11612 6248
rect 11664 6236 11670 6248
rect 12161 6239 12219 6245
rect 12161 6236 12173 6239
rect 11664 6208 12173 6236
rect 11664 6196 11670 6208
rect 12161 6205 12173 6208
rect 12207 6236 12219 6239
rect 12250 6236 12256 6248
rect 12207 6208 12256 6236
rect 12207 6205 12219 6208
rect 12161 6199 12219 6205
rect 12250 6196 12256 6208
rect 12308 6236 12314 6248
rect 14108 6236 14136 6267
rect 14366 6264 14372 6276
rect 14424 6264 14430 6316
rect 12308 6208 14136 6236
rect 14185 6239 14243 6245
rect 12308 6196 12314 6208
rect 14185 6205 14197 6239
rect 14231 6236 14243 6239
rect 15304 6236 15332 6400
rect 17954 6332 17960 6384
rect 18012 6372 18018 6384
rect 18785 6375 18843 6381
rect 18785 6372 18797 6375
rect 18012 6344 18797 6372
rect 18012 6332 18018 6344
rect 18785 6341 18797 6344
rect 18831 6341 18843 6375
rect 18785 6335 18843 6341
rect 19058 6332 19064 6384
rect 19116 6372 19122 6384
rect 19153 6375 19211 6381
rect 19153 6372 19165 6375
rect 19116 6344 19165 6372
rect 19116 6332 19122 6344
rect 19153 6341 19165 6344
rect 19199 6341 19211 6375
rect 19153 6335 19211 6341
rect 19334 6332 19340 6384
rect 19392 6372 19398 6384
rect 19889 6375 19947 6381
rect 19889 6372 19901 6375
rect 19392 6344 19901 6372
rect 19392 6332 19398 6344
rect 19889 6341 19901 6344
rect 19935 6341 19947 6375
rect 20732 6372 20760 6412
rect 19889 6335 19947 6341
rect 20640 6344 20760 6372
rect 18693 6307 18751 6313
rect 18693 6273 18705 6307
rect 18739 6304 18751 6307
rect 20070 6304 20076 6316
rect 18739 6276 20076 6304
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 20070 6264 20076 6276
rect 20128 6264 20134 6316
rect 14231 6208 15332 6236
rect 14231 6205 14243 6208
rect 14185 6199 14243 6205
rect 18966 6196 18972 6248
rect 19024 6196 19030 6248
rect 20640 6236 20668 6344
rect 22370 6332 22376 6384
rect 22428 6332 22434 6384
rect 23842 6372 23848 6384
rect 22480 6344 23848 6372
rect 21177 6307 21235 6313
rect 21177 6304 21189 6307
rect 20916 6276 21189 6304
rect 19168 6208 20668 6236
rect 10796 6140 13308 6168
rect 7883 6072 8432 6100
rect 7883 6069 7895 6072
rect 7837 6063 7895 6069
rect 10410 6060 10416 6112
rect 10468 6060 10474 6112
rect 11885 6103 11943 6109
rect 11885 6069 11897 6103
rect 11931 6100 11943 6103
rect 12158 6100 12164 6112
rect 11931 6072 12164 6100
rect 11931 6069 11943 6072
rect 11885 6063 11943 6069
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 12253 6103 12311 6109
rect 12253 6069 12265 6103
rect 12299 6100 12311 6103
rect 12802 6100 12808 6112
rect 12299 6072 12808 6100
rect 12299 6069 12311 6072
rect 12253 6063 12311 6069
rect 12802 6060 12808 6072
rect 12860 6060 12866 6112
rect 13280 6100 13308 6140
rect 13446 6128 13452 6180
rect 13504 6168 13510 6180
rect 18046 6168 18052 6180
rect 13504 6140 18052 6168
rect 13504 6128 13510 6140
rect 18046 6128 18052 6140
rect 18104 6168 18110 6180
rect 19168 6168 19196 6208
rect 20806 6196 20812 6248
rect 20864 6196 20870 6248
rect 18104 6140 19196 6168
rect 20165 6171 20223 6177
rect 18104 6128 18110 6140
rect 20165 6137 20177 6171
rect 20211 6168 20223 6171
rect 20211 6140 20576 6168
rect 20211 6137 20223 6140
rect 20165 6131 20223 6137
rect 14090 6100 14096 6112
rect 13280 6072 14096 6100
rect 14090 6060 14096 6072
rect 14148 6060 14154 6112
rect 18966 6060 18972 6112
rect 19024 6100 19030 6112
rect 20254 6100 20260 6112
rect 19024 6072 20260 6100
rect 19024 6060 19030 6072
rect 20254 6060 20260 6072
rect 20312 6060 20318 6112
rect 20548 6100 20576 6140
rect 20916 6100 20944 6276
rect 21177 6273 21189 6276
rect 21223 6273 21235 6307
rect 21177 6267 21235 6273
rect 22278 6264 22284 6316
rect 22336 6264 22342 6316
rect 22480 6313 22508 6344
rect 23842 6332 23848 6344
rect 23900 6332 23906 6384
rect 25222 6332 25228 6384
rect 25280 6332 25286 6384
rect 26068 6372 26096 6412
rect 26234 6400 26240 6452
rect 26292 6400 26298 6452
rect 26694 6400 26700 6452
rect 26752 6400 26758 6452
rect 26804 6412 34376 6440
rect 26804 6372 26832 6412
rect 26068 6344 26832 6372
rect 28994 6332 29000 6384
rect 29052 6332 29058 6384
rect 29546 6332 29552 6384
rect 29604 6332 29610 6384
rect 33686 6332 33692 6384
rect 33744 6332 33750 6384
rect 34348 6372 34376 6412
rect 34422 6400 34428 6452
rect 34480 6440 34486 6452
rect 35437 6443 35495 6449
rect 35437 6440 35449 6443
rect 34480 6412 35449 6440
rect 34480 6400 34486 6412
rect 35437 6409 35449 6412
rect 35483 6409 35495 6443
rect 35437 6403 35495 6409
rect 40954 6372 40960 6384
rect 34348 6344 40960 6372
rect 40954 6332 40960 6344
rect 41012 6332 41018 6384
rect 22465 6307 22523 6313
rect 22465 6273 22477 6307
rect 22511 6273 22523 6307
rect 22465 6267 22523 6273
rect 24486 6264 24492 6316
rect 24544 6264 24550 6316
rect 26513 6307 26571 6313
rect 26513 6273 26525 6307
rect 26559 6273 26571 6307
rect 26513 6267 26571 6273
rect 26789 6307 26847 6313
rect 26789 6273 26801 6307
rect 26835 6304 26847 6307
rect 27522 6304 27528 6316
rect 26835 6276 27528 6304
rect 26835 6273 26847 6276
rect 26789 6267 26847 6273
rect 24765 6239 24823 6245
rect 24765 6205 24777 6239
rect 24811 6236 24823 6239
rect 26329 6239 26387 6245
rect 26329 6236 26341 6239
rect 24811 6208 26341 6236
rect 24811 6205 24823 6208
rect 24765 6199 24823 6205
rect 26329 6205 26341 6208
rect 26375 6205 26387 6239
rect 26528 6236 26556 6267
rect 27522 6264 27528 6276
rect 27580 6264 27586 6316
rect 29012 6236 29040 6332
rect 29178 6264 29184 6316
rect 29236 6304 29242 6316
rect 29457 6307 29515 6313
rect 29457 6304 29469 6307
rect 29236 6276 29469 6304
rect 29236 6264 29242 6276
rect 29457 6273 29469 6276
rect 29503 6273 29515 6307
rect 29457 6267 29515 6273
rect 29638 6264 29644 6316
rect 29696 6302 29702 6316
rect 31205 6307 31263 6313
rect 29696 6274 29739 6302
rect 29696 6264 29702 6274
rect 31205 6273 31217 6307
rect 31251 6304 31263 6307
rect 31294 6304 31300 6316
rect 31251 6276 31300 6304
rect 31251 6273 31263 6276
rect 31205 6267 31263 6273
rect 31294 6264 31300 6276
rect 31352 6264 31358 6316
rect 31389 6307 31447 6313
rect 31389 6273 31401 6307
rect 31435 6304 31447 6307
rect 32214 6304 32220 6316
rect 31435 6276 32220 6304
rect 31435 6273 31447 6276
rect 31389 6267 31447 6273
rect 32214 6264 32220 6276
rect 32272 6304 32278 6316
rect 35621 6307 35679 6313
rect 32272 6276 34205 6304
rect 32272 6264 32278 6276
rect 26528 6208 29040 6236
rect 34057 6239 34115 6245
rect 26329 6199 26387 6205
rect 34057 6205 34069 6239
rect 34103 6205 34115 6239
rect 34177 6236 34205 6276
rect 35621 6273 35633 6307
rect 35667 6273 35679 6307
rect 35621 6267 35679 6273
rect 34330 6236 34336 6248
rect 34177 6208 34336 6236
rect 34057 6199 34115 6205
rect 33689 6171 33747 6177
rect 33689 6168 33701 6171
rect 28736 6140 33701 6168
rect 28736 6112 28764 6140
rect 33689 6137 33701 6140
rect 33735 6137 33747 6171
rect 33965 6171 34023 6177
rect 33965 6168 33977 6171
rect 33689 6131 33747 6137
rect 33796 6140 33977 6168
rect 20548 6072 20944 6100
rect 20990 6060 20996 6112
rect 21048 6060 21054 6112
rect 21082 6060 21088 6112
rect 21140 6100 21146 6112
rect 22002 6100 22008 6112
rect 21140 6072 22008 6100
rect 21140 6060 21146 6072
rect 22002 6060 22008 6072
rect 22060 6060 22066 6112
rect 28718 6060 28724 6112
rect 28776 6060 28782 6112
rect 30834 6060 30840 6112
rect 30892 6100 30898 6112
rect 31205 6103 31263 6109
rect 31205 6100 31217 6103
rect 30892 6072 31217 6100
rect 30892 6060 30898 6072
rect 31205 6069 31217 6072
rect 31251 6069 31263 6103
rect 31205 6063 31263 6069
rect 33594 6060 33600 6112
rect 33652 6100 33658 6112
rect 33796 6100 33824 6140
rect 33965 6137 33977 6140
rect 34011 6137 34023 6171
rect 34072 6168 34100 6199
rect 34330 6196 34336 6208
rect 34388 6236 34394 6248
rect 34388 6208 34744 6236
rect 34388 6196 34394 6208
rect 34146 6168 34152 6180
rect 34072 6140 34152 6168
rect 33965 6131 34023 6137
rect 34146 6128 34152 6140
rect 34204 6128 34210 6180
rect 34716 6168 34744 6208
rect 34790 6196 34796 6248
rect 34848 6196 34854 6248
rect 35636 6168 35664 6267
rect 34716 6140 35664 6168
rect 33652 6072 33824 6100
rect 33873 6103 33931 6109
rect 33652 6060 33658 6072
rect 33873 6069 33885 6103
rect 33919 6100 33931 6103
rect 34606 6100 34612 6112
rect 33919 6072 34612 6100
rect 33919 6069 33931 6072
rect 33873 6063 33931 6069
rect 34606 6060 34612 6072
rect 34664 6060 34670 6112
rect 35710 6060 35716 6112
rect 35768 6060 35774 6112
rect 1104 6010 41400 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 41400 6010
rect 1104 5936 41400 5958
rect 6822 5856 6828 5908
rect 6880 5896 6886 5908
rect 6880 5868 10824 5896
rect 6880 5856 6886 5868
rect 10796 5828 10824 5868
rect 10870 5856 10876 5908
rect 10928 5856 10934 5908
rect 18966 5896 18972 5908
rect 10980 5868 18972 5896
rect 10980 5828 11008 5868
rect 18966 5856 18972 5868
rect 19024 5856 19030 5908
rect 20254 5856 20260 5908
rect 20312 5896 20318 5908
rect 20806 5896 20812 5908
rect 20312 5868 20812 5896
rect 20312 5856 20318 5868
rect 20806 5856 20812 5868
rect 20864 5856 20870 5908
rect 20990 5856 20996 5908
rect 21048 5856 21054 5908
rect 21082 5856 21088 5908
rect 21140 5856 21146 5908
rect 22002 5856 22008 5908
rect 22060 5896 22066 5908
rect 22094 5896 22100 5908
rect 22060 5868 22100 5896
rect 22060 5856 22066 5868
rect 22094 5856 22100 5868
rect 22152 5856 22158 5908
rect 27798 5856 27804 5908
rect 27856 5896 27862 5908
rect 28629 5899 28687 5905
rect 28629 5896 28641 5899
rect 27856 5868 28641 5896
rect 27856 5856 27862 5868
rect 28629 5865 28641 5868
rect 28675 5865 28687 5899
rect 28629 5859 28687 5865
rect 33594 5856 33600 5908
rect 33652 5896 33658 5908
rect 33873 5899 33931 5905
rect 33873 5896 33885 5899
rect 33652 5868 33885 5896
rect 33652 5856 33658 5868
rect 33873 5865 33885 5868
rect 33919 5865 33931 5899
rect 36170 5896 36176 5908
rect 33873 5859 33931 5865
rect 35360 5868 36176 5896
rect 10796 5800 11008 5828
rect 11146 5788 11152 5840
rect 11204 5828 11210 5840
rect 15102 5828 15108 5840
rect 11204 5800 15108 5828
rect 11204 5788 11210 5800
rect 15102 5788 15108 5800
rect 15160 5788 15166 5840
rect 8110 5720 8116 5772
rect 8168 5760 8174 5772
rect 9125 5763 9183 5769
rect 9125 5760 9137 5763
rect 8168 5732 9137 5760
rect 8168 5720 8174 5732
rect 9125 5729 9137 5732
rect 9171 5760 9183 5763
rect 9766 5760 9772 5772
rect 9171 5732 9772 5760
rect 9171 5729 9183 5732
rect 9125 5723 9183 5729
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 19334 5720 19340 5772
rect 19392 5720 19398 5772
rect 19613 5763 19671 5769
rect 19613 5729 19625 5763
rect 19659 5760 19671 5763
rect 21008 5760 21036 5856
rect 27522 5788 27528 5840
rect 27580 5828 27586 5840
rect 27580 5800 30972 5828
rect 27580 5788 27586 5800
rect 19659 5732 21036 5760
rect 21177 5763 21235 5769
rect 19659 5729 19671 5732
rect 19613 5723 19671 5729
rect 21177 5729 21189 5763
rect 21223 5760 21235 5763
rect 21818 5760 21824 5772
rect 21223 5732 21824 5760
rect 21223 5729 21235 5732
rect 21177 5723 21235 5729
rect 21818 5720 21824 5732
rect 21876 5720 21882 5772
rect 21910 5720 21916 5772
rect 21968 5760 21974 5772
rect 30834 5760 30840 5772
rect 21968 5732 29592 5760
rect 21968 5720 21974 5732
rect 16117 5695 16175 5701
rect 16117 5661 16129 5695
rect 16163 5661 16175 5695
rect 16117 5655 16175 5661
rect 9398 5584 9404 5636
rect 9456 5584 9462 5636
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 16132 5624 16160 5655
rect 20714 5652 20720 5704
rect 20772 5652 20778 5704
rect 22554 5652 22560 5704
rect 22612 5652 22618 5704
rect 27709 5695 27767 5701
rect 27709 5661 27721 5695
rect 27755 5661 27767 5695
rect 27709 5655 27767 5661
rect 27801 5695 27859 5701
rect 27801 5661 27813 5695
rect 27847 5692 27859 5695
rect 27982 5692 27988 5704
rect 27847 5664 27988 5692
rect 27847 5661 27859 5664
rect 27801 5655 27859 5661
rect 16298 5624 16304 5636
rect 9732 5596 9890 5624
rect 16132 5596 16304 5624
rect 9732 5584 9738 5596
rect 16298 5584 16304 5596
rect 16356 5584 16362 5636
rect 16393 5627 16451 5633
rect 16393 5593 16405 5627
rect 16439 5624 16451 5627
rect 16666 5624 16672 5636
rect 16439 5596 16672 5624
rect 16439 5593 16451 5596
rect 16393 5587 16451 5593
rect 16666 5584 16672 5596
rect 16724 5584 16730 5636
rect 17862 5624 17868 5636
rect 17618 5596 17868 5624
rect 17862 5584 17868 5596
rect 17920 5584 17926 5636
rect 18046 5584 18052 5636
rect 18104 5624 18110 5636
rect 18141 5627 18199 5633
rect 18141 5624 18153 5627
rect 18104 5596 18153 5624
rect 18104 5584 18110 5596
rect 18141 5593 18153 5596
rect 18187 5593 18199 5627
rect 18141 5587 18199 5593
rect 21453 5627 21511 5633
rect 21453 5593 21465 5627
rect 21499 5593 21511 5627
rect 21453 5587 21511 5593
rect 21468 5556 21496 5587
rect 23198 5584 23204 5636
rect 23256 5584 23262 5636
rect 27724 5624 27752 5655
rect 27982 5652 27988 5664
rect 28040 5652 28046 5704
rect 28166 5652 28172 5704
rect 28224 5692 28230 5704
rect 28261 5695 28319 5701
rect 28261 5692 28273 5695
rect 28224 5664 28273 5692
rect 28224 5652 28230 5664
rect 28261 5661 28273 5664
rect 28307 5661 28319 5695
rect 28261 5655 28319 5661
rect 28445 5695 28503 5701
rect 28445 5661 28457 5695
rect 28491 5661 28503 5695
rect 28445 5655 28503 5661
rect 28460 5624 28488 5655
rect 28718 5652 28724 5704
rect 28776 5652 28782 5704
rect 29362 5652 29368 5704
rect 29420 5652 29426 5704
rect 29564 5701 29592 5732
rect 30576 5732 30840 5760
rect 30576 5701 30604 5732
rect 30834 5720 30840 5732
rect 30892 5720 30898 5772
rect 29549 5695 29607 5701
rect 29549 5661 29561 5695
rect 29595 5661 29607 5695
rect 30561 5695 30619 5701
rect 29549 5655 29607 5661
rect 29656 5664 30420 5692
rect 29380 5624 29408 5652
rect 29656 5624 29684 5664
rect 27724 5596 28948 5624
rect 29380 5596 29684 5624
rect 22462 5556 22468 5568
rect 21468 5528 22468 5556
rect 22462 5516 22468 5528
rect 22520 5516 22526 5568
rect 26050 5516 26056 5568
rect 26108 5556 26114 5568
rect 28258 5556 28264 5568
rect 26108 5528 28264 5556
rect 26108 5516 26114 5528
rect 28258 5516 28264 5528
rect 28316 5516 28322 5568
rect 28920 5565 28948 5596
rect 30006 5584 30012 5636
rect 30064 5624 30070 5636
rect 30285 5627 30343 5633
rect 30285 5624 30297 5627
rect 30064 5596 30297 5624
rect 30064 5584 30070 5596
rect 30285 5593 30297 5596
rect 30331 5593 30343 5627
rect 30392 5624 30420 5664
rect 30561 5661 30573 5695
rect 30607 5661 30619 5695
rect 30561 5655 30619 5661
rect 30742 5652 30748 5704
rect 30800 5652 30806 5704
rect 30944 5701 30972 5800
rect 34057 5763 34115 5769
rect 34057 5729 34069 5763
rect 34103 5760 34115 5763
rect 34790 5760 34796 5772
rect 34103 5732 34796 5760
rect 34103 5729 34115 5732
rect 34057 5723 34115 5729
rect 34790 5720 34796 5732
rect 34848 5720 34854 5772
rect 30929 5695 30987 5701
rect 30929 5661 30941 5695
rect 30975 5692 30987 5695
rect 32582 5692 32588 5704
rect 30975 5664 32588 5692
rect 30975 5661 30987 5664
rect 30929 5655 30987 5661
rect 32582 5652 32588 5664
rect 32640 5652 32646 5704
rect 33229 5695 33287 5701
rect 33229 5661 33241 5695
rect 33275 5692 33287 5695
rect 33594 5692 33600 5704
rect 33275 5664 33600 5692
rect 33275 5661 33287 5664
rect 33229 5655 33287 5661
rect 33594 5652 33600 5664
rect 33652 5652 33658 5704
rect 33686 5652 33692 5704
rect 33744 5692 33750 5704
rect 33873 5695 33931 5701
rect 33873 5692 33885 5695
rect 33744 5664 33885 5692
rect 33744 5652 33750 5664
rect 33873 5661 33885 5664
rect 33919 5661 33931 5695
rect 33873 5655 33931 5661
rect 34146 5652 34152 5704
rect 34204 5692 34210 5704
rect 35360 5701 35388 5868
rect 36170 5856 36176 5868
rect 36228 5856 36234 5908
rect 40954 5856 40960 5908
rect 41012 5856 41018 5908
rect 35345 5695 35403 5701
rect 34204 5664 35296 5692
rect 34204 5652 34210 5664
rect 30837 5627 30895 5633
rect 30837 5624 30849 5627
rect 30392 5596 30849 5624
rect 30285 5587 30343 5593
rect 30837 5593 30849 5596
rect 30883 5593 30895 5627
rect 30837 5587 30895 5593
rect 32766 5584 32772 5636
rect 32824 5624 32830 5636
rect 33704 5624 33732 5652
rect 32824 5596 33732 5624
rect 35268 5624 35296 5664
rect 35345 5661 35357 5695
rect 35391 5661 35403 5695
rect 35345 5655 35403 5661
rect 35621 5695 35679 5701
rect 35621 5661 35633 5695
rect 35667 5692 35679 5695
rect 35710 5692 35716 5704
rect 35667 5664 35716 5692
rect 35667 5661 35679 5664
rect 35621 5655 35679 5661
rect 35710 5652 35716 5664
rect 35768 5652 35774 5704
rect 36265 5695 36323 5701
rect 36265 5661 36277 5695
rect 36311 5692 36323 5695
rect 36906 5692 36912 5704
rect 36311 5664 36912 5692
rect 36311 5661 36323 5664
rect 36265 5655 36323 5661
rect 36280 5624 36308 5655
rect 36906 5652 36912 5664
rect 36964 5652 36970 5704
rect 40773 5695 40831 5701
rect 40773 5661 40785 5695
rect 40819 5692 40831 5695
rect 40819 5664 41368 5692
rect 40819 5661 40831 5664
rect 40773 5655 40831 5661
rect 35268 5596 36308 5624
rect 32824 5584 32830 5596
rect 41340 5568 41368 5664
rect 28905 5559 28963 5565
rect 28905 5525 28917 5559
rect 28951 5525 28963 5559
rect 28905 5519 28963 5525
rect 29914 5516 29920 5568
rect 29972 5556 29978 5568
rect 31113 5559 31171 5565
rect 31113 5556 31125 5559
rect 29972 5528 31125 5556
rect 29972 5516 29978 5528
rect 31113 5525 31125 5528
rect 31159 5525 31171 5559
rect 31113 5519 31171 5525
rect 33226 5516 33232 5568
rect 33284 5556 33290 5568
rect 33781 5559 33839 5565
rect 33781 5556 33793 5559
rect 33284 5528 33793 5556
rect 33284 5516 33290 5528
rect 33781 5525 33793 5528
rect 33827 5525 33839 5559
rect 33781 5519 33839 5525
rect 34330 5516 34336 5568
rect 34388 5516 34394 5568
rect 35161 5559 35219 5565
rect 35161 5525 35173 5559
rect 35207 5556 35219 5559
rect 35342 5556 35348 5568
rect 35207 5528 35348 5556
rect 35207 5525 35219 5528
rect 35161 5519 35219 5525
rect 35342 5516 35348 5528
rect 35400 5516 35406 5568
rect 35529 5559 35587 5565
rect 35529 5525 35541 5559
rect 35575 5556 35587 5559
rect 36817 5559 36875 5565
rect 36817 5556 36829 5559
rect 35575 5528 36829 5556
rect 35575 5525 35587 5528
rect 35529 5519 35587 5525
rect 36817 5525 36829 5528
rect 36863 5525 36875 5559
rect 36817 5519 36875 5525
rect 41322 5516 41328 5568
rect 41380 5516 41386 5568
rect 1104 5466 41400 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 41400 5466
rect 1104 5392 41400 5414
rect 9398 5312 9404 5364
rect 9456 5352 9462 5364
rect 9585 5355 9643 5361
rect 9585 5352 9597 5355
rect 9456 5324 9597 5352
rect 9456 5312 9462 5324
rect 9585 5321 9597 5324
rect 9631 5321 9643 5355
rect 9585 5315 9643 5321
rect 10410 5312 10416 5364
rect 10468 5312 10474 5364
rect 11974 5352 11980 5364
rect 11808 5324 11980 5352
rect 9769 5219 9827 5225
rect 9769 5185 9781 5219
rect 9815 5216 9827 5219
rect 10428 5216 10456 5312
rect 11808 5293 11836 5324
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 13265 5355 13323 5361
rect 13265 5352 13277 5355
rect 12492 5324 13277 5352
rect 12492 5312 12498 5324
rect 13265 5321 13277 5324
rect 13311 5321 13323 5355
rect 13265 5315 13323 5321
rect 16298 5312 16304 5364
rect 16356 5352 16362 5364
rect 19334 5352 19340 5364
rect 16356 5324 19340 5352
rect 16356 5312 16362 5324
rect 11793 5287 11851 5293
rect 11793 5253 11805 5287
rect 11839 5253 11851 5287
rect 13078 5284 13084 5296
rect 13018 5256 13084 5284
rect 11793 5247 11851 5253
rect 13078 5244 13084 5256
rect 13136 5244 13142 5296
rect 16666 5244 16672 5296
rect 16724 5244 16730 5296
rect 17037 5287 17095 5293
rect 17037 5253 17049 5287
rect 17083 5284 17095 5287
rect 17083 5256 18092 5284
rect 17083 5253 17095 5256
rect 17037 5247 17095 5253
rect 18064 5228 18092 5256
rect 9815 5188 10456 5216
rect 16853 5219 16911 5225
rect 9815 5185 9827 5188
rect 9769 5179 9827 5185
rect 16853 5185 16865 5219
rect 16899 5216 16911 5219
rect 16942 5216 16948 5228
rect 16899 5188 16948 5216
rect 16899 5185 16911 5188
rect 16853 5179 16911 5185
rect 16942 5176 16948 5188
rect 17000 5176 17006 5228
rect 17126 5176 17132 5228
rect 17184 5176 17190 5228
rect 18046 5176 18052 5228
rect 18104 5176 18110 5228
rect 18156 5225 18184 5324
rect 19334 5312 19340 5324
rect 19392 5312 19398 5364
rect 20162 5312 20168 5364
rect 20220 5352 20226 5364
rect 21821 5355 21879 5361
rect 21821 5352 21833 5355
rect 20220 5324 21833 5352
rect 20220 5312 20226 5324
rect 21821 5321 21833 5324
rect 21867 5321 21879 5355
rect 21821 5315 21879 5321
rect 22462 5312 22468 5364
rect 22520 5312 22526 5364
rect 31389 5355 31447 5361
rect 27632 5324 31340 5352
rect 18417 5287 18475 5293
rect 18417 5253 18429 5287
rect 18463 5284 18475 5287
rect 18690 5284 18696 5296
rect 18463 5256 18696 5284
rect 18463 5253 18475 5256
rect 18417 5247 18475 5253
rect 18690 5244 18696 5256
rect 18748 5244 18754 5296
rect 20622 5284 20628 5296
rect 19642 5270 20628 5284
rect 19628 5256 20628 5270
rect 18141 5219 18199 5225
rect 18141 5185 18153 5219
rect 18187 5185 18199 5219
rect 18141 5179 18199 5185
rect 9950 5108 9956 5160
rect 10008 5108 10014 5160
rect 11517 5151 11575 5157
rect 11517 5117 11529 5151
rect 11563 5117 11575 5151
rect 11517 5111 11575 5117
rect 11624 5120 14412 5148
rect 9766 5040 9772 5092
rect 9824 5080 9830 5092
rect 11532 5080 11560 5111
rect 9824 5052 11560 5080
rect 9824 5040 9830 5052
rect 10597 5015 10655 5021
rect 10597 4981 10609 5015
rect 10643 5012 10655 5015
rect 11624 5012 11652 5120
rect 14384 5024 14412 5120
rect 10643 4984 11652 5012
rect 10643 4981 10655 4984
rect 10597 4975 10655 4981
rect 14366 4972 14372 5024
rect 14424 4972 14430 5024
rect 17144 5012 17172 5176
rect 17862 5108 17868 5160
rect 17920 5148 17926 5160
rect 19628 5148 19656 5256
rect 20622 5244 20628 5256
rect 20680 5244 20686 5296
rect 27632 5231 27660 5324
rect 29086 5244 29092 5296
rect 29144 5244 29150 5296
rect 31312 5284 31340 5324
rect 31389 5321 31401 5355
rect 31435 5352 31447 5355
rect 31570 5352 31576 5364
rect 31435 5324 31576 5352
rect 31435 5321 31447 5324
rect 31389 5315 31447 5321
rect 31570 5312 31576 5324
rect 31628 5312 31634 5364
rect 31662 5312 31668 5364
rect 31720 5312 31726 5364
rect 32309 5355 32367 5361
rect 32309 5321 32321 5355
rect 32355 5352 32367 5355
rect 32674 5352 32680 5364
rect 32355 5324 32680 5352
rect 32355 5321 32367 5324
rect 32309 5315 32367 5321
rect 32674 5312 32680 5324
rect 32732 5312 32738 5364
rect 32766 5312 32772 5364
rect 32824 5312 32830 5364
rect 33336 5324 35204 5352
rect 31680 5284 31708 5312
rect 32784 5284 32812 5312
rect 31312 5256 31708 5284
rect 32509 5256 32812 5284
rect 22278 5216 22284 5228
rect 17920 5120 19656 5148
rect 22066 5188 22284 5216
rect 17920 5108 17926 5120
rect 22066 5080 22094 5188
rect 22278 5176 22284 5188
rect 22336 5176 22342 5228
rect 27157 5219 27215 5225
rect 27157 5185 27169 5219
rect 27203 5185 27215 5219
rect 27157 5179 27215 5185
rect 22189 5151 22247 5157
rect 22189 5117 22201 5151
rect 22235 5148 22247 5151
rect 23198 5148 23204 5160
rect 22235 5120 23204 5148
rect 22235 5117 22247 5120
rect 22189 5111 22247 5117
rect 23198 5108 23204 5120
rect 23256 5108 23262 5160
rect 27172 5148 27200 5179
rect 27246 5176 27252 5228
rect 27304 5176 27310 5228
rect 27522 5176 27528 5228
rect 27580 5176 27586 5228
rect 27617 5225 27675 5231
rect 27617 5191 27629 5225
rect 27663 5191 27675 5225
rect 27617 5185 27675 5191
rect 28166 5176 28172 5228
rect 28224 5176 28230 5228
rect 28258 5176 28264 5228
rect 28316 5216 28322 5228
rect 28353 5219 28411 5225
rect 28353 5216 28365 5219
rect 28316 5188 28365 5216
rect 28316 5176 28322 5188
rect 28353 5185 28365 5188
rect 28399 5185 28411 5219
rect 28353 5179 28411 5185
rect 27893 5151 27951 5157
rect 27172 5120 27844 5148
rect 27614 5080 27620 5092
rect 19444 5052 22094 5080
rect 27448 5052 27620 5080
rect 19444 5012 19472 5052
rect 17144 4984 19472 5012
rect 19889 5015 19947 5021
rect 19889 4981 19901 5015
rect 19935 5012 19947 5015
rect 20070 5012 20076 5024
rect 19935 4984 20076 5012
rect 19935 4981 19947 4984
rect 19889 4975 19947 4981
rect 20070 4972 20076 4984
rect 20128 5012 20134 5024
rect 20622 5012 20628 5024
rect 20128 4984 20628 5012
rect 20128 4972 20134 4984
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 26970 4972 26976 5024
rect 27028 4972 27034 5024
rect 27448 5021 27476 5052
rect 27614 5040 27620 5052
rect 27672 5040 27678 5092
rect 27433 5015 27491 5021
rect 27433 4981 27445 5015
rect 27479 4981 27491 5015
rect 27433 4975 27491 4981
rect 27706 4972 27712 5024
rect 27764 4972 27770 5024
rect 27816 5021 27844 5120
rect 27893 5117 27905 5151
rect 27939 5148 27951 5151
rect 28184 5148 28212 5176
rect 27939 5120 28212 5148
rect 27939 5117 27951 5120
rect 27893 5111 27951 5117
rect 27801 5015 27859 5021
rect 27801 4981 27813 5015
rect 27847 4981 27859 5015
rect 28368 5012 28396 5179
rect 29914 5176 29920 5228
rect 29972 5176 29978 5228
rect 31018 5176 31024 5228
rect 31076 5176 31082 5228
rect 31297 5219 31355 5225
rect 31297 5185 31309 5219
rect 31343 5216 31355 5219
rect 31754 5216 31760 5228
rect 31343 5188 31760 5216
rect 31343 5185 31355 5188
rect 31297 5179 31355 5185
rect 31754 5176 31760 5188
rect 31812 5216 31818 5228
rect 32509 5216 32537 5256
rect 31812 5188 32537 5216
rect 31812 5176 31818 5188
rect 32582 5176 32588 5228
rect 32640 5176 32646 5228
rect 32677 5219 32735 5225
rect 32677 5185 32689 5219
rect 32723 5216 32735 5219
rect 33226 5216 33232 5228
rect 32723 5188 33232 5216
rect 32723 5185 32735 5188
rect 32677 5179 32735 5185
rect 33226 5176 33232 5188
rect 33284 5176 33290 5228
rect 33336 5225 33364 5324
rect 33502 5244 33508 5296
rect 33560 5284 33566 5296
rect 33597 5287 33655 5293
rect 33597 5284 33609 5287
rect 33560 5256 33609 5284
rect 33560 5244 33566 5256
rect 33597 5253 33609 5256
rect 33643 5253 33655 5287
rect 33597 5247 33655 5253
rect 34054 5244 34060 5296
rect 34112 5244 34118 5296
rect 35176 5225 35204 5324
rect 36906 5312 36912 5364
rect 36964 5312 36970 5364
rect 35342 5244 35348 5296
rect 35400 5284 35406 5296
rect 35437 5287 35495 5293
rect 35437 5284 35449 5287
rect 35400 5256 35449 5284
rect 35400 5244 35406 5256
rect 35437 5253 35449 5256
rect 35483 5253 35495 5287
rect 35437 5247 35495 5253
rect 33321 5219 33379 5225
rect 33321 5185 33333 5219
rect 33367 5185 33379 5219
rect 33321 5179 33379 5185
rect 35161 5219 35219 5225
rect 35161 5185 35173 5219
rect 35207 5185 35219 5219
rect 35161 5179 35219 5185
rect 28629 5151 28687 5157
rect 28629 5117 28641 5151
rect 28675 5148 28687 5151
rect 29932 5148 29960 5176
rect 30377 5151 30435 5157
rect 30377 5148 30389 5151
rect 28675 5120 29960 5148
rect 30024 5120 30389 5148
rect 28675 5117 28687 5120
rect 28629 5111 28687 5117
rect 28994 5012 29000 5024
rect 28368 4984 29000 5012
rect 27801 4975 27859 4981
rect 28994 4972 29000 4984
rect 29052 4972 29058 5024
rect 29362 4972 29368 5024
rect 29420 5012 29426 5024
rect 30024 5012 30052 5120
rect 30377 5117 30389 5120
rect 30423 5117 30435 5151
rect 31036 5148 31064 5176
rect 31481 5151 31539 5157
rect 31481 5148 31493 5151
rect 31036 5120 31493 5148
rect 30377 5111 30435 5117
rect 31481 5117 31493 5120
rect 31527 5117 31539 5151
rect 32600 5148 32628 5176
rect 32769 5151 32827 5157
rect 32769 5148 32781 5151
rect 32600 5120 32781 5148
rect 31481 5111 31539 5117
rect 32769 5117 32781 5120
rect 32815 5117 32827 5151
rect 32769 5111 32827 5117
rect 33336 5080 33364 5179
rect 34790 5108 34796 5160
rect 34848 5148 34854 5160
rect 35069 5151 35127 5157
rect 35069 5148 35081 5151
rect 34848 5120 35081 5148
rect 34848 5108 34854 5120
rect 35069 5117 35081 5120
rect 35115 5117 35127 5151
rect 35069 5111 35127 5117
rect 36170 5108 36176 5160
rect 36228 5148 36234 5160
rect 36556 5148 36584 5202
rect 36228 5120 36584 5148
rect 36228 5108 36234 5120
rect 31726 5052 33364 5080
rect 31726 5024 31754 5052
rect 29420 4984 30052 5012
rect 29420 4972 29426 4984
rect 30926 4972 30932 5024
rect 30984 4972 30990 5024
rect 31662 4972 31668 5024
rect 31720 4984 31754 5024
rect 31720 4972 31726 4984
rect 32950 4972 32956 5024
rect 33008 4972 33014 5024
rect 1104 4922 41400 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 41400 4922
rect 1104 4848 41400 4870
rect 3605 4811 3663 4817
rect 3605 4777 3617 4811
rect 3651 4808 3663 4811
rect 9950 4808 9956 4820
rect 3651 4780 9956 4808
rect 3651 4777 3663 4780
rect 3605 4771 3663 4777
rect 9950 4768 9956 4780
rect 10008 4768 10014 4820
rect 14366 4768 14372 4820
rect 14424 4808 14430 4820
rect 16282 4811 16340 4817
rect 16282 4808 16294 4811
rect 14424 4780 16294 4808
rect 14424 4768 14430 4780
rect 16282 4777 16294 4780
rect 16328 4777 16340 4811
rect 16282 4771 16340 4777
rect 17770 4768 17776 4820
rect 17828 4768 17834 4820
rect 27522 4768 27528 4820
rect 27580 4808 27586 4820
rect 27939 4811 27997 4817
rect 27939 4808 27951 4811
rect 27580 4780 27951 4808
rect 27580 4768 27586 4780
rect 27939 4777 27951 4780
rect 27985 4808 27997 4811
rect 28166 4808 28172 4820
rect 27985 4780 28172 4808
rect 27985 4777 27997 4780
rect 27939 4771 27997 4777
rect 28166 4768 28172 4780
rect 28224 4768 28230 4820
rect 29086 4768 29092 4820
rect 29144 4768 29150 4820
rect 31754 4768 31760 4820
rect 31812 4768 31818 4820
rect 33594 4768 33600 4820
rect 33652 4817 33658 4820
rect 33652 4811 33701 4817
rect 33652 4777 33655 4811
rect 33689 4777 33701 4811
rect 33652 4771 33701 4777
rect 33652 4768 33658 4771
rect 29104 4740 29132 4768
rect 28000 4712 29132 4740
rect 1854 4632 1860 4684
rect 1912 4632 1918 4684
rect 16025 4675 16083 4681
rect 16025 4641 16037 4675
rect 16071 4672 16083 4675
rect 16298 4672 16304 4684
rect 16071 4644 16304 4672
rect 16071 4641 16083 4644
rect 16025 4635 16083 4641
rect 16298 4632 16304 4644
rect 16356 4632 16362 4684
rect 26050 4632 26056 4684
rect 26108 4672 26114 4684
rect 26145 4675 26203 4681
rect 26145 4672 26157 4675
rect 26108 4644 26157 4672
rect 26108 4632 26114 4644
rect 26145 4641 26157 4644
rect 26191 4641 26203 4675
rect 26145 4635 26203 4641
rect 26513 4675 26571 4681
rect 26513 4641 26525 4675
rect 26559 4672 26571 4675
rect 26970 4672 26976 4684
rect 26559 4644 26976 4672
rect 26559 4641 26571 4644
rect 26513 4635 26571 4641
rect 26970 4632 26976 4644
rect 27028 4632 27034 4684
rect 6546 4604 6552 4616
rect 3266 4576 6552 4604
rect 6546 4564 6552 4576
rect 6604 4564 6610 4616
rect 17862 4604 17868 4616
rect 17434 4576 17868 4604
rect 17862 4564 17868 4576
rect 17920 4564 17926 4616
rect 27430 4564 27436 4616
rect 27488 4604 27494 4616
rect 27488 4576 27568 4604
rect 27488 4564 27494 4576
rect 2130 4496 2136 4548
rect 2188 4496 2194 4548
rect 27540 4536 27568 4576
rect 28000 4536 28028 4712
rect 28994 4632 29000 4684
rect 29052 4672 29058 4684
rect 30006 4672 30012 4684
rect 29052 4644 30012 4672
rect 29052 4632 29058 4644
rect 30006 4632 30012 4644
rect 30064 4672 30070 4684
rect 31662 4672 31668 4684
rect 30064 4644 31668 4672
rect 30064 4632 30070 4644
rect 31662 4632 31668 4644
rect 31720 4672 31726 4684
rect 31849 4675 31907 4681
rect 31849 4672 31861 4675
rect 31720 4644 31861 4672
rect 31720 4632 31726 4644
rect 31849 4641 31861 4644
rect 31895 4641 31907 4675
rect 31849 4635 31907 4641
rect 32217 4675 32275 4681
rect 32217 4641 32229 4675
rect 32263 4672 32275 4675
rect 32950 4672 32956 4684
rect 32263 4644 32956 4672
rect 32263 4641 32275 4644
rect 32217 4635 32275 4641
rect 32950 4632 32956 4644
rect 33008 4632 33014 4684
rect 29178 4564 29184 4616
rect 29236 4564 29242 4616
rect 35986 4564 35992 4616
rect 36044 4564 36050 4616
rect 27540 4522 28028 4536
rect 27554 4508 28028 4522
rect 29196 4468 29224 4564
rect 30285 4539 30343 4545
rect 30285 4505 30297 4539
rect 30331 4536 30343 4539
rect 30558 4536 30564 4548
rect 30331 4508 30564 4536
rect 30331 4505 30343 4508
rect 30285 4499 30343 4505
rect 30558 4496 30564 4508
rect 30616 4496 30622 4548
rect 30668 4508 30774 4536
rect 31726 4508 31984 4536
rect 30668 4468 30696 4508
rect 31726 4468 31754 4508
rect 29196 4440 31754 4468
rect 31956 4468 31984 4508
rect 32508 4508 32614 4536
rect 32508 4468 32536 4508
rect 34054 4468 34060 4480
rect 31956 4440 34060 4468
rect 34054 4428 34060 4440
rect 34112 4468 34118 4480
rect 36170 4468 36176 4480
rect 34112 4440 36176 4468
rect 34112 4428 34118 4440
rect 36170 4428 36176 4440
rect 36228 4428 36234 4480
rect 1104 4378 41400 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 41400 4378
rect 1104 4304 41400 4326
rect 1949 4267 2007 4273
rect 1949 4233 1961 4267
rect 1995 4264 2007 4267
rect 2130 4264 2136 4276
rect 1995 4236 2136 4264
rect 1995 4233 2007 4236
rect 1949 4227 2007 4233
rect 2130 4224 2136 4236
rect 2188 4224 2194 4276
rect 30558 4224 30564 4276
rect 30616 4224 30622 4276
rect 30926 4224 30932 4276
rect 30984 4224 30990 4276
rect 934 4088 940 4140
rect 992 4128 998 4140
rect 1857 4131 1915 4137
rect 1857 4128 1869 4131
rect 992 4100 1869 4128
rect 992 4088 998 4100
rect 1857 4097 1869 4100
rect 1903 4097 1915 4131
rect 1857 4091 1915 4097
rect 9766 4088 9772 4140
rect 9824 4128 9830 4140
rect 10781 4131 10839 4137
rect 10781 4128 10793 4131
rect 9824 4100 10793 4128
rect 9824 4088 9830 4100
rect 10781 4097 10793 4100
rect 10827 4097 10839 4131
rect 10781 4091 10839 4097
rect 30745 4131 30803 4137
rect 30745 4097 30757 4131
rect 30791 4128 30803 4131
rect 30944 4128 30972 4224
rect 30791 4100 30972 4128
rect 30791 4097 30803 4100
rect 30745 4091 30803 4097
rect 10962 3884 10968 3936
rect 11020 3884 11026 3936
rect 1104 3834 41400 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 41400 3834
rect 1104 3760 41400 3782
rect 15010 3544 15016 3596
rect 15068 3544 15074 3596
rect 14 3476 20 3528
rect 72 3516 78 3528
rect 3602 3516 3608 3528
rect 72 3488 3608 3516
rect 72 3476 78 3488
rect 3602 3476 3608 3488
rect 3660 3476 3666 3528
rect 14734 3476 14740 3528
rect 14792 3476 14798 3528
rect 14829 3519 14887 3525
rect 14829 3485 14841 3519
rect 14875 3485 14887 3519
rect 14829 3479 14887 3485
rect 14182 3408 14188 3460
rect 14240 3448 14246 3460
rect 14844 3448 14872 3479
rect 14240 3420 14872 3448
rect 14240 3408 14246 3420
rect 23198 3408 23204 3460
rect 23256 3448 23262 3460
rect 36722 3448 36728 3460
rect 23256 3420 36728 3448
rect 23256 3408 23262 3420
rect 36722 3408 36728 3420
rect 36780 3408 36786 3460
rect 1104 3290 41400 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 41400 3290
rect 1104 3216 41400 3238
rect 14734 3136 14740 3188
rect 14792 3136 14798 3188
rect 14093 3043 14151 3049
rect 14093 3009 14105 3043
rect 14139 3040 14151 3043
rect 14752 3040 14780 3136
rect 14139 3012 14780 3040
rect 14139 3009 14151 3012
rect 14093 3003 14151 3009
rect 3234 2796 3240 2848
rect 3292 2836 3298 2848
rect 14185 2839 14243 2845
rect 14185 2836 14197 2839
rect 3292 2808 14197 2836
rect 3292 2796 3298 2808
rect 14185 2805 14197 2808
rect 14231 2805 14243 2839
rect 14185 2799 14243 2805
rect 1104 2746 41400 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 41400 2746
rect 1104 2672 41400 2694
rect 40770 2592 40776 2644
rect 40828 2592 40834 2644
rect 20622 2456 20628 2508
rect 20680 2496 20686 2508
rect 20680 2468 29684 2496
rect 20680 2456 20686 2468
rect 7282 2388 7288 2440
rect 7340 2388 7346 2440
rect 22094 2388 22100 2440
rect 22152 2388 22158 2440
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29549 2431 29607 2437
rect 29549 2428 29561 2431
rect 29052 2400 29561 2428
rect 29052 2388 29058 2400
rect 29549 2397 29561 2400
rect 29595 2397 29607 2431
rect 29656 2428 29684 2468
rect 29822 2456 29828 2508
rect 29880 2456 29886 2508
rect 33045 2431 33103 2437
rect 33045 2428 33057 2431
rect 29656 2400 33057 2428
rect 29549 2391 29607 2397
rect 33045 2397 33057 2400
rect 33091 2397 33103 2431
rect 33045 2391 33103 2397
rect 40678 2320 40684 2372
rect 40736 2320 40742 2372
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7377 2295 7435 2301
rect 7377 2292 7389 2295
rect 7156 2264 7389 2292
rect 7156 2252 7162 2264
rect 7377 2261 7389 2264
rect 7423 2261 7435 2295
rect 7377 2255 7435 2261
rect 22002 2252 22008 2304
rect 22060 2292 22066 2304
rect 22189 2295 22247 2301
rect 22189 2292 22201 2295
rect 22060 2264 22201 2292
rect 22060 2252 22066 2264
rect 22189 2261 22201 2264
rect 22235 2261 22247 2295
rect 22189 2255 22247 2261
rect 33134 2252 33140 2304
rect 33192 2252 33198 2304
rect 1104 2202 41400 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 41400 2202
rect 1104 2128 41400 2150
<< via1 >>
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 1308 42304 1360 42356
rect 35072 42347 35124 42356
rect 35072 42313 35081 42347
rect 35081 42313 35115 42347
rect 35115 42313 35124 42347
rect 35072 42304 35124 42313
rect 9036 42236 9088 42288
rect 1492 42211 1544 42220
rect 1492 42177 1501 42211
rect 1501 42177 1535 42211
rect 1535 42177 1544 42211
rect 1492 42168 1544 42177
rect 17500 42211 17552 42220
rect 17500 42177 17509 42211
rect 17509 42177 17543 42211
rect 17543 42177 17552 42211
rect 17500 42168 17552 42177
rect 19432 42168 19484 42220
rect 30932 42168 30984 42220
rect 34520 42168 34572 42220
rect 38660 42168 38712 42220
rect 31300 42143 31352 42152
rect 31300 42109 31309 42143
rect 31309 42109 31343 42143
rect 31343 42109 31352 42143
rect 31300 42100 31352 42109
rect 37188 42100 37240 42152
rect 9312 42007 9364 42016
rect 9312 41973 9321 42007
rect 9321 41973 9355 42007
rect 9355 41973 9364 42007
rect 9312 41964 9364 41973
rect 17316 42007 17368 42016
rect 17316 41973 17325 42007
rect 17325 41973 17359 42007
rect 17359 41973 17368 42007
rect 17316 41964 17368 41973
rect 19616 41964 19668 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 17316 41760 17368 41812
rect 11152 41624 11204 41676
rect 19340 41667 19392 41676
rect 19340 41633 19349 41667
rect 19349 41633 19383 41667
rect 19383 41633 19392 41667
rect 19340 41624 19392 41633
rect 19616 41667 19668 41676
rect 19616 41633 19625 41667
rect 19625 41633 19659 41667
rect 19659 41633 19668 41667
rect 19616 41624 19668 41633
rect 19984 41624 20036 41676
rect 10600 41488 10652 41540
rect 10968 41420 11020 41472
rect 16120 41599 16172 41608
rect 16120 41565 16129 41599
rect 16129 41565 16163 41599
rect 16163 41565 16172 41599
rect 16120 41556 16172 41565
rect 18788 41556 18840 41608
rect 12072 41531 12124 41540
rect 12072 41497 12081 41531
rect 12081 41497 12115 41531
rect 12115 41497 12124 41531
rect 12072 41488 12124 41497
rect 11520 41420 11572 41472
rect 12900 41420 12952 41472
rect 14004 41488 14056 41540
rect 14372 41531 14424 41540
rect 14372 41497 14381 41531
rect 14381 41497 14415 41531
rect 14415 41497 14424 41531
rect 14372 41488 14424 41497
rect 17408 41488 17460 41540
rect 22100 41556 22152 41608
rect 20904 41488 20956 41540
rect 22468 41531 22520 41540
rect 22468 41497 22477 41531
rect 22477 41497 22511 41531
rect 22511 41497 22520 41531
rect 22468 41488 22520 41497
rect 23940 41488 23992 41540
rect 24216 41531 24268 41540
rect 24216 41497 24225 41531
rect 24225 41497 24259 41531
rect 24259 41497 24268 41531
rect 24216 41488 24268 41497
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 12072 41216 12124 41268
rect 14372 41216 14424 41268
rect 17500 41216 17552 41268
rect 19432 41259 19484 41268
rect 19432 41225 19441 41259
rect 19441 41225 19475 41259
rect 19475 41225 19484 41259
rect 19432 41216 19484 41225
rect 19984 41216 20036 41268
rect 23848 41216 23900 41268
rect 24216 41216 24268 41268
rect 41880 41216 41932 41268
rect 1676 41191 1728 41200
rect 1676 41157 1685 41191
rect 1685 41157 1719 41191
rect 1719 41157 1728 41191
rect 1676 41148 1728 41157
rect 3608 41080 3660 41132
rect 2688 41012 2740 41064
rect 2872 41012 2924 41064
rect 3424 41055 3476 41064
rect 3424 41021 3433 41055
rect 3433 41021 3467 41055
rect 3467 41021 3476 41055
rect 3424 41012 3476 41021
rect 4068 41055 4120 41064
rect 4068 41021 4077 41055
rect 4077 41021 4111 41055
rect 4111 41021 4120 41055
rect 4068 41012 4120 41021
rect 12532 41080 12584 41132
rect 5356 41012 5408 41064
rect 11520 41012 11572 41064
rect 12808 41123 12860 41132
rect 12808 41089 12817 41123
rect 12817 41089 12851 41123
rect 12851 41089 12860 41123
rect 12808 41080 12860 41089
rect 14280 41123 14332 41132
rect 14280 41089 14289 41123
rect 14289 41089 14323 41123
rect 14323 41089 14332 41123
rect 14280 41080 14332 41089
rect 16120 41080 16172 41132
rect 17224 41123 17276 41132
rect 17224 41089 17233 41123
rect 17233 41089 17267 41123
rect 17267 41089 17276 41123
rect 17224 41080 17276 41089
rect 17316 41055 17368 41064
rect 17316 41021 17325 41055
rect 17325 41021 17359 41055
rect 17359 41021 17368 41055
rect 17316 41012 17368 41021
rect 15384 40944 15436 40996
rect 17592 41012 17644 41064
rect 21364 41123 21416 41132
rect 21364 41089 21373 41123
rect 21373 41089 21407 41123
rect 21407 41089 21416 41123
rect 21364 41080 21416 41089
rect 21640 41123 21692 41132
rect 21640 41089 21649 41123
rect 21649 41089 21683 41123
rect 21683 41089 21692 41123
rect 21640 41080 21692 41089
rect 22100 41148 22152 41200
rect 23388 41080 23440 41132
rect 23940 41080 23992 41132
rect 40776 41123 40828 41132
rect 40776 41089 40785 41123
rect 40785 41089 40819 41123
rect 40819 41089 40828 41123
rect 40776 41080 40828 41089
rect 5264 40876 5316 40928
rect 11060 40919 11112 40928
rect 11060 40885 11069 40919
rect 11069 40885 11103 40919
rect 11103 40885 11112 40919
rect 11060 40876 11112 40885
rect 16028 40876 16080 40928
rect 21088 41012 21140 41064
rect 21824 41055 21876 41064
rect 21824 41021 21833 41055
rect 21833 41021 21867 41055
rect 21867 41021 21876 41055
rect 21824 41012 21876 41021
rect 23848 41055 23900 41064
rect 23848 41021 23857 41055
rect 23857 41021 23891 41055
rect 23891 41021 23900 41055
rect 23848 41012 23900 41021
rect 40960 40919 41012 40928
rect 40960 40885 40969 40919
rect 40969 40885 41003 40919
rect 41003 40885 41012 40919
rect 40960 40876 41012 40885
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 1676 40672 1728 40724
rect 4068 40672 4120 40724
rect 3424 40536 3476 40588
rect 2872 40511 2924 40520
rect 2872 40477 2881 40511
rect 2881 40477 2915 40511
rect 2915 40477 2924 40511
rect 2872 40468 2924 40477
rect 4620 40468 4672 40520
rect 5356 40468 5408 40520
rect 9772 40604 9824 40656
rect 11152 40672 11204 40724
rect 15384 40672 15436 40724
rect 15476 40672 15528 40724
rect 15660 40647 15712 40656
rect 8024 40443 8076 40452
rect 8024 40409 8033 40443
rect 8033 40409 8067 40443
rect 8067 40409 8076 40443
rect 8024 40400 8076 40409
rect 10416 40511 10468 40520
rect 10416 40477 10425 40511
rect 10425 40477 10459 40511
rect 10459 40477 10468 40511
rect 10416 40468 10468 40477
rect 13268 40536 13320 40588
rect 4620 40375 4672 40384
rect 4620 40341 4629 40375
rect 4629 40341 4663 40375
rect 4663 40341 4672 40375
rect 4620 40332 4672 40341
rect 4804 40332 4856 40384
rect 8852 40332 8904 40384
rect 9956 40332 10008 40384
rect 11060 40468 11112 40520
rect 10692 40443 10744 40452
rect 10692 40409 10701 40443
rect 10701 40409 10735 40443
rect 10735 40409 10744 40443
rect 10692 40400 10744 40409
rect 11520 40468 11572 40520
rect 14188 40468 14240 40520
rect 11244 40332 11296 40384
rect 11336 40375 11388 40384
rect 11336 40341 11345 40375
rect 11345 40341 11379 40375
rect 11379 40341 11388 40375
rect 11336 40332 11388 40341
rect 11428 40332 11480 40384
rect 12348 40332 12400 40384
rect 14280 40332 14332 40384
rect 14740 40511 14792 40520
rect 14740 40477 14749 40511
rect 14749 40477 14783 40511
rect 14783 40477 14792 40511
rect 14740 40468 14792 40477
rect 15660 40613 15669 40647
rect 15669 40613 15703 40647
rect 15703 40613 15712 40647
rect 15660 40604 15712 40613
rect 17224 40672 17276 40724
rect 21364 40672 21416 40724
rect 22468 40715 22520 40724
rect 22468 40681 22477 40715
rect 22477 40681 22511 40715
rect 22511 40681 22520 40715
rect 22468 40672 22520 40681
rect 15016 40511 15068 40520
rect 15016 40477 15025 40511
rect 15025 40477 15059 40511
rect 15059 40477 15068 40511
rect 15016 40468 15068 40477
rect 15384 40468 15436 40520
rect 16580 40536 16632 40588
rect 16948 40468 17000 40520
rect 19432 40579 19484 40588
rect 19432 40545 19441 40579
rect 19441 40545 19475 40579
rect 19475 40545 19484 40579
rect 19432 40536 19484 40545
rect 21640 40536 21692 40588
rect 22284 40536 22336 40588
rect 20720 40468 20772 40520
rect 14740 40332 14792 40384
rect 15292 40332 15344 40384
rect 19432 40400 19484 40452
rect 21180 40400 21232 40452
rect 22468 40468 22520 40520
rect 24216 40468 24268 40520
rect 15844 40332 15896 40384
rect 17500 40375 17552 40384
rect 17500 40341 17509 40375
rect 17509 40341 17543 40375
rect 17543 40341 17552 40375
rect 17500 40332 17552 40341
rect 18328 40375 18380 40384
rect 18328 40341 18337 40375
rect 18337 40341 18371 40375
rect 18371 40341 18380 40375
rect 18328 40332 18380 40341
rect 20076 40332 20128 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 9864 40128 9916 40180
rect 7472 40103 7524 40112
rect 7472 40069 7481 40103
rect 7481 40069 7515 40103
rect 7515 40069 7524 40103
rect 7472 40060 7524 40069
rect 8208 40060 8260 40112
rect 7288 39992 7340 40044
rect 10140 40103 10192 40112
rect 10140 40069 10175 40103
rect 10175 40069 10192 40103
rect 10508 40171 10560 40180
rect 10508 40137 10517 40171
rect 10517 40137 10551 40171
rect 10551 40137 10560 40171
rect 10508 40128 10560 40137
rect 10600 40128 10652 40180
rect 11152 40128 11204 40180
rect 11336 40128 11388 40180
rect 10140 40060 10192 40069
rect 8484 40035 8536 40044
rect 8484 40001 8493 40035
rect 8493 40001 8527 40035
rect 8527 40001 8536 40035
rect 8484 39992 8536 40001
rect 2688 39924 2740 39976
rect 8576 39924 8628 39976
rect 10048 40035 10100 40044
rect 10048 40001 10057 40035
rect 10057 40001 10091 40035
rect 10091 40001 10100 40035
rect 10048 39992 10100 40001
rect 11060 40060 11112 40112
rect 10784 40035 10836 40044
rect 10784 40001 10793 40035
rect 10793 40001 10827 40035
rect 10827 40001 10836 40035
rect 11428 40060 11480 40112
rect 10784 39992 10836 40001
rect 10140 39924 10192 39976
rect 10416 39924 10468 39976
rect 11520 39967 11572 39976
rect 11520 39933 11529 39967
rect 11529 39933 11563 39967
rect 11563 39933 11572 39967
rect 11520 39924 11572 39933
rect 14188 40128 14240 40180
rect 15844 40128 15896 40180
rect 19432 40128 19484 40180
rect 13912 40060 13964 40112
rect 15384 40103 15436 40112
rect 15384 40069 15393 40103
rect 15393 40069 15427 40103
rect 15427 40069 15436 40103
rect 15384 40060 15436 40069
rect 15568 40060 15620 40112
rect 15016 39992 15068 40044
rect 15292 40035 15344 40044
rect 15292 40001 15301 40035
rect 15301 40001 15335 40035
rect 15335 40001 15344 40035
rect 15292 39992 15344 40001
rect 15476 40035 15528 40044
rect 15476 40001 15485 40035
rect 15485 40001 15519 40035
rect 15519 40001 15528 40035
rect 15476 39992 15528 40001
rect 16212 40103 16264 40112
rect 16212 40069 16221 40103
rect 16221 40069 16255 40103
rect 16255 40069 16264 40103
rect 16212 40060 16264 40069
rect 19340 40060 19392 40112
rect 24952 40171 25004 40180
rect 24952 40137 24961 40171
rect 24961 40137 24995 40171
rect 24995 40137 25004 40171
rect 24952 40128 25004 40137
rect 40776 40128 40828 40180
rect 23572 40060 23624 40112
rect 11888 39967 11940 39976
rect 11888 39933 11897 39967
rect 11897 39933 11931 39967
rect 11931 39933 11940 39967
rect 11888 39924 11940 39933
rect 10876 39856 10928 39908
rect 13176 39967 13228 39976
rect 13176 39933 13185 39967
rect 13185 39933 13219 39967
rect 13219 39933 13228 39967
rect 13176 39924 13228 39933
rect 14740 39924 14792 39976
rect 15844 39992 15896 40044
rect 18880 40035 18932 40044
rect 18880 40001 18889 40035
rect 18889 40001 18923 40035
rect 18923 40001 18932 40035
rect 18880 39992 18932 40001
rect 22008 40035 22060 40044
rect 22008 40001 22017 40035
rect 22017 40001 22051 40035
rect 22051 40001 22060 40035
rect 22008 39992 22060 40001
rect 23112 40035 23164 40044
rect 23112 40001 23121 40035
rect 23121 40001 23155 40035
rect 23155 40001 23164 40035
rect 23112 39992 23164 40001
rect 16672 39967 16724 39976
rect 16672 39933 16681 39967
rect 16681 39933 16715 39967
rect 16715 39933 16724 39967
rect 16672 39924 16724 39933
rect 17408 39924 17460 39976
rect 18052 39924 18104 39976
rect 18328 39924 18380 39976
rect 20720 39967 20772 39976
rect 20720 39933 20729 39967
rect 20729 39933 20763 39967
rect 20763 39933 20772 39967
rect 20720 39924 20772 39933
rect 21824 39924 21876 39976
rect 15660 39856 15712 39908
rect 8116 39788 8168 39840
rect 12624 39788 12676 39840
rect 12716 39788 12768 39840
rect 15936 39788 15988 39840
rect 16396 39831 16448 39840
rect 16396 39797 16405 39831
rect 16405 39797 16439 39831
rect 16439 39797 16448 39831
rect 16396 39788 16448 39797
rect 21824 39831 21876 39840
rect 21824 39797 21833 39831
rect 21833 39797 21867 39831
rect 21867 39797 21876 39831
rect 21824 39788 21876 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 7380 39584 7432 39636
rect 8208 39627 8260 39636
rect 8208 39593 8217 39627
rect 8217 39593 8251 39627
rect 8251 39593 8260 39627
rect 8208 39584 8260 39593
rect 8576 39584 8628 39636
rect 8668 39584 8720 39636
rect 11244 39584 11296 39636
rect 12900 39584 12952 39636
rect 13176 39584 13228 39636
rect 15016 39584 15068 39636
rect 16212 39584 16264 39636
rect 1492 39448 1544 39500
rect 4068 39448 4120 39500
rect 7288 39448 7340 39500
rect 8484 39448 8536 39500
rect 11796 39559 11848 39568
rect 11796 39525 11805 39559
rect 11805 39525 11839 39559
rect 11839 39525 11848 39559
rect 11796 39516 11848 39525
rect 12716 39516 12768 39568
rect 15200 39516 15252 39568
rect 9220 39491 9272 39500
rect 9220 39457 9229 39491
rect 9229 39457 9263 39491
rect 9263 39457 9272 39491
rect 9220 39448 9272 39457
rect 9588 39448 9640 39500
rect 7840 39423 7892 39432
rect 7840 39389 7849 39423
rect 7849 39389 7883 39423
rect 7883 39389 7892 39423
rect 7840 39380 7892 39389
rect 5724 39312 5776 39364
rect 8116 39312 8168 39364
rect 9680 39312 9732 39364
rect 10784 39380 10836 39432
rect 11244 39423 11296 39432
rect 11244 39389 11253 39423
rect 11253 39389 11287 39423
rect 11287 39389 11296 39423
rect 11244 39380 11296 39389
rect 11888 39448 11940 39500
rect 11060 39312 11112 39364
rect 11612 39423 11664 39432
rect 11612 39389 11621 39423
rect 11621 39389 11655 39423
rect 11655 39389 11664 39423
rect 11612 39380 11664 39389
rect 16396 39448 16448 39500
rect 21824 39448 21876 39500
rect 23112 39584 23164 39636
rect 22836 39516 22888 39568
rect 26148 39448 26200 39500
rect 4620 39244 4672 39296
rect 7012 39244 7064 39296
rect 7840 39244 7892 39296
rect 8392 39287 8444 39296
rect 8392 39253 8401 39287
rect 8401 39253 8435 39287
rect 8435 39253 8444 39287
rect 8392 39244 8444 39253
rect 8484 39244 8536 39296
rect 9956 39244 10008 39296
rect 10140 39244 10192 39296
rect 12900 39423 12952 39432
rect 12900 39389 12910 39423
rect 12910 39389 12944 39423
rect 12944 39389 12952 39423
rect 12900 39380 12952 39389
rect 13268 39423 13320 39432
rect 13268 39389 13282 39423
rect 13282 39389 13316 39423
rect 13316 39389 13320 39423
rect 13268 39380 13320 39389
rect 14740 39423 14792 39432
rect 14740 39389 14749 39423
rect 14749 39389 14783 39423
rect 14783 39389 14792 39423
rect 14740 39380 14792 39389
rect 13084 39355 13136 39364
rect 13084 39321 13093 39355
rect 13093 39321 13127 39355
rect 13127 39321 13136 39355
rect 13084 39312 13136 39321
rect 12992 39244 13044 39296
rect 14188 39244 14240 39296
rect 15476 39380 15528 39432
rect 16672 39380 16724 39432
rect 17224 39380 17276 39432
rect 20168 39380 20220 39432
rect 20720 39380 20772 39432
rect 24952 39380 25004 39432
rect 15292 39312 15344 39364
rect 15568 39355 15620 39364
rect 15568 39321 15577 39355
rect 15577 39321 15611 39355
rect 15611 39321 15620 39355
rect 15568 39312 15620 39321
rect 15844 39355 15896 39364
rect 15844 39321 15853 39355
rect 15853 39321 15887 39355
rect 15887 39321 15896 39355
rect 15844 39312 15896 39321
rect 26056 39312 26108 39364
rect 27712 39312 27764 39364
rect 18236 39244 18288 39296
rect 18788 39244 18840 39296
rect 20628 39244 20680 39296
rect 22928 39287 22980 39296
rect 22928 39253 22937 39287
rect 22937 39253 22971 39287
rect 22971 39253 22980 39287
rect 22928 39244 22980 39253
rect 23388 39244 23440 39296
rect 27804 39244 27856 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 3608 39040 3660 39092
rect 4068 39083 4120 39092
rect 4068 39049 4077 39083
rect 4077 39049 4111 39083
rect 4111 39049 4120 39083
rect 4068 39040 4120 39049
rect 4712 38972 4764 39024
rect 7288 39040 7340 39092
rect 5724 38904 5776 38956
rect 7012 38947 7064 38956
rect 7012 38913 7021 38947
rect 7021 38913 7055 38947
rect 7055 38913 7064 38947
rect 7012 38904 7064 38913
rect 1768 38836 1820 38888
rect 3056 38836 3108 38888
rect 6460 38836 6512 38888
rect 2688 38700 2740 38752
rect 6736 38700 6788 38752
rect 8392 39040 8444 39092
rect 9220 39040 9272 39092
rect 11244 39083 11296 39092
rect 11244 39049 11253 39083
rect 11253 39049 11287 39083
rect 11287 39049 11296 39083
rect 11244 39040 11296 39049
rect 11796 39040 11848 39092
rect 12900 39040 12952 39092
rect 16580 39040 16632 39092
rect 17224 39083 17276 39092
rect 17224 39049 17233 39083
rect 17233 39049 17267 39083
rect 17267 39049 17276 39083
rect 17224 39040 17276 39049
rect 17960 39040 18012 39092
rect 8484 38947 8536 38956
rect 8484 38913 8494 38947
rect 8494 38913 8528 38947
rect 8528 38913 8536 38947
rect 8484 38904 8536 38913
rect 8668 38947 8720 38956
rect 8668 38913 8677 38947
rect 8677 38913 8711 38947
rect 8711 38913 8720 38947
rect 8668 38904 8720 38913
rect 8852 38947 8904 38956
rect 8852 38913 8866 38947
rect 8866 38913 8900 38947
rect 8900 38913 8904 38947
rect 8852 38904 8904 38913
rect 9588 38904 9640 38956
rect 10784 38904 10836 38956
rect 11428 38972 11480 39024
rect 11336 38904 11388 38956
rect 11704 38947 11756 38956
rect 11704 38913 11713 38947
rect 11713 38913 11747 38947
rect 11747 38913 11756 38947
rect 11704 38904 11756 38913
rect 12992 38972 13044 39024
rect 12624 38947 12676 38956
rect 12624 38913 12633 38947
rect 12633 38913 12667 38947
rect 12667 38913 12676 38947
rect 12624 38904 12676 38913
rect 13912 38904 13964 38956
rect 12900 38879 12952 38888
rect 12900 38845 12909 38879
rect 12909 38845 12943 38879
rect 12943 38845 12952 38879
rect 12900 38836 12952 38845
rect 14372 38836 14424 38888
rect 8208 38700 8260 38752
rect 8484 38700 8536 38752
rect 12256 38768 12308 38820
rect 11336 38700 11388 38752
rect 15476 38836 15528 38888
rect 17316 38836 17368 38888
rect 17592 38836 17644 38888
rect 20168 39040 20220 39092
rect 22008 39040 22060 39092
rect 22928 39040 22980 39092
rect 26056 39040 26108 39092
rect 18236 38972 18288 39024
rect 18788 38972 18840 39024
rect 22008 38904 22060 38956
rect 25596 38947 25648 38956
rect 25596 38913 25605 38947
rect 25605 38913 25639 38947
rect 25639 38913 25648 38947
rect 25596 38904 25648 38913
rect 25780 38947 25832 38956
rect 25780 38913 25789 38947
rect 25789 38913 25823 38947
rect 25823 38913 25832 38947
rect 25780 38904 25832 38913
rect 26056 38904 26108 38956
rect 27804 38904 27856 38956
rect 19432 38768 19484 38820
rect 15384 38743 15436 38752
rect 15384 38709 15393 38743
rect 15393 38709 15427 38743
rect 15427 38709 15436 38743
rect 15384 38700 15436 38709
rect 20904 38700 20956 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 3056 38496 3108 38548
rect 4712 38539 4764 38548
rect 4712 38505 4721 38539
rect 4721 38505 4755 38539
rect 4755 38505 4764 38539
rect 4712 38496 4764 38505
rect 6552 38539 6604 38548
rect 6552 38505 6561 38539
rect 6561 38505 6595 38539
rect 6595 38505 6604 38539
rect 6552 38496 6604 38505
rect 6736 38496 6788 38548
rect 11704 38496 11756 38548
rect 12900 38496 12952 38548
rect 17960 38496 18012 38548
rect 22008 38539 22060 38548
rect 22008 38505 22017 38539
rect 22017 38505 22051 38539
rect 22051 38505 22060 38539
rect 22008 38496 22060 38505
rect 23204 38496 23256 38548
rect 27620 38496 27672 38548
rect 4620 38292 4672 38344
rect 5356 38360 5408 38412
rect 6736 38360 6788 38412
rect 6828 38360 6880 38412
rect 8024 38428 8076 38480
rect 6644 38335 6696 38344
rect 6644 38301 6653 38335
rect 6653 38301 6687 38335
rect 6687 38301 6696 38335
rect 6644 38292 6696 38301
rect 4620 38156 4672 38208
rect 5540 38156 5592 38208
rect 6460 38156 6512 38208
rect 6828 38199 6880 38208
rect 6828 38165 6837 38199
rect 6837 38165 6871 38199
rect 6871 38165 6880 38199
rect 6828 38156 6880 38165
rect 7288 38335 7340 38344
rect 7288 38301 7297 38335
rect 7297 38301 7331 38335
rect 7331 38301 7340 38335
rect 7288 38292 7340 38301
rect 7748 38292 7800 38344
rect 9404 38360 9456 38412
rect 8208 38292 8260 38344
rect 11060 38335 11112 38344
rect 11060 38301 11069 38335
rect 11069 38301 11103 38335
rect 11103 38301 11112 38335
rect 11060 38292 11112 38301
rect 11152 38292 11204 38344
rect 11244 38292 11296 38344
rect 11612 38428 11664 38480
rect 14832 38428 14884 38480
rect 11520 38335 11572 38344
rect 11520 38301 11529 38335
rect 11529 38301 11563 38335
rect 11563 38301 11572 38335
rect 11520 38292 11572 38301
rect 11980 38335 12032 38344
rect 11980 38301 11989 38335
rect 11989 38301 12023 38335
rect 12023 38301 12032 38335
rect 11980 38292 12032 38301
rect 15936 38360 15988 38412
rect 16580 38360 16632 38412
rect 13268 38292 13320 38344
rect 14464 38292 14516 38344
rect 17040 38335 17092 38344
rect 17040 38301 17049 38335
rect 17049 38301 17083 38335
rect 17083 38301 17092 38335
rect 17040 38292 17092 38301
rect 22468 38360 22520 38412
rect 24952 38360 25004 38412
rect 26148 38360 26200 38412
rect 12256 38267 12308 38276
rect 12256 38233 12265 38267
rect 12265 38233 12299 38267
rect 12299 38233 12308 38267
rect 12256 38224 12308 38233
rect 15384 38224 15436 38276
rect 14280 38156 14332 38208
rect 17316 38199 17368 38208
rect 17316 38165 17325 38199
rect 17325 38165 17359 38199
rect 17359 38165 17368 38199
rect 17316 38156 17368 38165
rect 17592 38292 17644 38344
rect 18144 38292 18196 38344
rect 20168 38292 20220 38344
rect 17684 38267 17736 38276
rect 17684 38233 17693 38267
rect 17693 38233 17727 38267
rect 17727 38233 17736 38267
rect 17684 38224 17736 38233
rect 17776 38267 17828 38276
rect 17776 38233 17785 38267
rect 17785 38233 17819 38267
rect 17819 38233 17828 38267
rect 17776 38224 17828 38233
rect 18604 38156 18656 38208
rect 20352 38156 20404 38208
rect 20628 38224 20680 38276
rect 20996 38224 21048 38276
rect 25044 38224 25096 38276
rect 23388 38156 23440 38208
rect 25320 38156 25372 38208
rect 27896 38267 27948 38276
rect 27896 38233 27905 38267
rect 27905 38233 27939 38267
rect 27939 38233 27948 38267
rect 27896 38224 27948 38233
rect 31208 38224 31260 38276
rect 26424 38199 26476 38208
rect 26424 38165 26433 38199
rect 26433 38165 26467 38199
rect 26467 38165 26476 38199
rect 26424 38156 26476 38165
rect 27804 38156 27856 38208
rect 30012 38156 30064 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 6644 37952 6696 38004
rect 8116 37952 8168 38004
rect 6276 37816 6328 37868
rect 6460 37816 6512 37868
rect 6736 37816 6788 37868
rect 7012 37816 7064 37868
rect 8208 37884 8260 37936
rect 8944 37859 8996 37868
rect 8944 37825 8953 37859
rect 8953 37825 8987 37859
rect 8987 37825 8996 37859
rect 8944 37816 8996 37825
rect 9404 37952 9456 38004
rect 11060 37952 11112 38004
rect 11980 37952 12032 38004
rect 15844 37952 15896 38004
rect 17776 37952 17828 38004
rect 18144 37995 18196 38004
rect 18144 37961 18153 37995
rect 18153 37961 18187 37995
rect 18187 37961 18196 37995
rect 18144 37952 18196 37961
rect 11336 37884 11388 37936
rect 16028 37884 16080 37936
rect 17040 37884 17092 37936
rect 17868 37884 17920 37936
rect 9496 37816 9548 37868
rect 9680 37748 9732 37800
rect 10784 37859 10836 37868
rect 10784 37825 10793 37859
rect 10793 37825 10827 37859
rect 10827 37825 10836 37859
rect 10784 37816 10836 37825
rect 11060 37816 11112 37868
rect 13728 37816 13780 37868
rect 14556 37859 14608 37868
rect 14556 37825 14565 37859
rect 14565 37825 14599 37859
rect 14599 37825 14608 37859
rect 14556 37816 14608 37825
rect 14740 37859 14792 37868
rect 14740 37825 14749 37859
rect 14749 37825 14783 37859
rect 14783 37825 14792 37859
rect 14740 37816 14792 37825
rect 16488 37816 16540 37868
rect 18512 37816 18564 37868
rect 19064 37884 19116 37936
rect 19524 37816 19576 37868
rect 12992 37680 13044 37732
rect 18328 37680 18380 37732
rect 19432 37791 19484 37800
rect 19432 37757 19441 37791
rect 19441 37757 19475 37791
rect 19475 37757 19484 37791
rect 19432 37748 19484 37757
rect 20904 37748 20956 37800
rect 22008 37859 22060 37868
rect 22008 37825 22017 37859
rect 22017 37825 22051 37859
rect 22051 37825 22060 37859
rect 22008 37816 22060 37825
rect 22652 37859 22704 37868
rect 22652 37825 22661 37859
rect 22661 37825 22695 37859
rect 22695 37825 22704 37859
rect 22652 37816 22704 37825
rect 23112 37859 23164 37868
rect 23112 37825 23121 37859
rect 23121 37825 23155 37859
rect 23155 37825 23164 37859
rect 23112 37816 23164 37825
rect 23204 37816 23256 37868
rect 6736 37655 6788 37664
rect 6736 37621 6745 37655
rect 6745 37621 6779 37655
rect 6779 37621 6788 37655
rect 6736 37612 6788 37621
rect 7104 37612 7156 37664
rect 7748 37612 7800 37664
rect 8116 37655 8168 37664
rect 8116 37621 8125 37655
rect 8125 37621 8159 37655
rect 8159 37621 8168 37655
rect 8116 37612 8168 37621
rect 10416 37612 10468 37664
rect 14648 37655 14700 37664
rect 14648 37621 14657 37655
rect 14657 37621 14691 37655
rect 14691 37621 14700 37655
rect 14648 37612 14700 37621
rect 16580 37612 16632 37664
rect 17684 37612 17736 37664
rect 19248 37723 19300 37732
rect 19248 37689 19257 37723
rect 19257 37689 19291 37723
rect 19291 37689 19300 37723
rect 19248 37680 19300 37689
rect 22100 37723 22152 37732
rect 22100 37689 22109 37723
rect 22109 37689 22143 37723
rect 22143 37689 22152 37723
rect 22100 37680 22152 37689
rect 20352 37612 20404 37664
rect 22376 37612 22428 37664
rect 23480 37859 23532 37868
rect 23480 37825 23489 37859
rect 23489 37825 23523 37859
rect 23523 37825 23532 37859
rect 23480 37816 23532 37825
rect 23572 37816 23624 37868
rect 24952 37952 25004 38004
rect 25320 37952 25372 38004
rect 25688 37884 25740 37936
rect 26424 37884 26476 37936
rect 27712 37884 27764 37936
rect 25504 37748 25556 37800
rect 26148 37748 26200 37800
rect 24584 37612 24636 37664
rect 24768 37612 24820 37664
rect 25596 37612 25648 37664
rect 27252 37791 27304 37800
rect 27252 37757 27261 37791
rect 27261 37757 27295 37791
rect 27295 37757 27304 37791
rect 27252 37748 27304 37757
rect 27804 37612 27856 37664
rect 29368 37612 29420 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 6552 37408 6604 37460
rect 6736 37408 6788 37460
rect 7288 37408 7340 37460
rect 7656 37408 7708 37460
rect 9496 37408 9548 37460
rect 11060 37408 11112 37460
rect 11520 37408 11572 37460
rect 14556 37408 14608 37460
rect 8024 37340 8076 37392
rect 6920 37272 6972 37324
rect 10324 37315 10376 37324
rect 10324 37281 10333 37315
rect 10333 37281 10367 37315
rect 10367 37281 10376 37315
rect 10324 37272 10376 37281
rect 14280 37340 14332 37392
rect 15844 37408 15896 37460
rect 17684 37408 17736 37460
rect 19248 37408 19300 37460
rect 23480 37408 23532 37460
rect 27252 37408 27304 37460
rect 27896 37451 27948 37460
rect 27896 37417 27905 37451
rect 27905 37417 27939 37451
rect 27939 37417 27948 37451
rect 27896 37408 27948 37417
rect 15292 37383 15344 37392
rect 15292 37349 15301 37383
rect 15301 37349 15335 37383
rect 15335 37349 15344 37383
rect 15292 37340 15344 37349
rect 7104 37204 7156 37256
rect 9956 37204 10008 37256
rect 5540 37136 5592 37188
rect 7196 37068 7248 37120
rect 8300 37068 8352 37120
rect 9036 37068 9088 37120
rect 11060 37204 11112 37256
rect 11244 37204 11296 37256
rect 14096 37204 14148 37256
rect 14280 37179 14332 37188
rect 14280 37145 14289 37179
rect 14289 37145 14323 37179
rect 14323 37145 14332 37179
rect 14280 37136 14332 37145
rect 16212 37247 16264 37256
rect 16212 37213 16221 37247
rect 16221 37213 16255 37247
rect 16255 37213 16264 37247
rect 16212 37204 16264 37213
rect 16304 37204 16356 37256
rect 16488 37204 16540 37256
rect 18512 37272 18564 37324
rect 18236 37204 18288 37256
rect 19248 37272 19300 37324
rect 19064 37247 19116 37256
rect 19064 37213 19073 37247
rect 19073 37213 19107 37247
rect 19107 37213 19116 37247
rect 19064 37204 19116 37213
rect 12440 37111 12492 37120
rect 12440 37077 12449 37111
rect 12449 37077 12483 37111
rect 12483 37077 12492 37111
rect 12440 37068 12492 37077
rect 12808 37111 12860 37120
rect 12808 37077 12817 37111
rect 12817 37077 12851 37111
rect 12851 37077 12860 37111
rect 12808 37068 12860 37077
rect 14740 37068 14792 37120
rect 19432 37272 19484 37324
rect 20168 37272 20220 37324
rect 22376 37272 22428 37324
rect 24952 37383 25004 37392
rect 24952 37349 24961 37383
rect 24961 37349 24995 37383
rect 24995 37349 25004 37383
rect 24952 37340 25004 37349
rect 23388 37204 23440 37256
rect 23572 37204 23624 37256
rect 24492 37204 24544 37256
rect 24676 37247 24728 37256
rect 24676 37213 24685 37247
rect 24685 37213 24719 37247
rect 24719 37213 24728 37247
rect 24676 37204 24728 37213
rect 25228 37272 25280 37324
rect 27620 37340 27672 37392
rect 17316 37068 17368 37120
rect 18052 37068 18104 37120
rect 18972 37068 19024 37120
rect 19524 37136 19576 37188
rect 24584 37179 24636 37188
rect 24584 37145 24593 37179
rect 24593 37145 24627 37179
rect 24627 37145 24636 37179
rect 24584 37136 24636 37145
rect 23756 37111 23808 37120
rect 23756 37077 23765 37111
rect 23765 37077 23799 37111
rect 23799 37077 23808 37111
rect 23756 37068 23808 37077
rect 25504 37136 25556 37188
rect 25964 37247 26016 37256
rect 25964 37213 25973 37247
rect 25973 37213 26007 37247
rect 26007 37213 26016 37247
rect 25964 37204 26016 37213
rect 26056 37204 26108 37256
rect 27528 37272 27580 37324
rect 25780 37068 25832 37120
rect 26240 37179 26292 37188
rect 26240 37145 26249 37179
rect 26249 37145 26283 37179
rect 26283 37145 26292 37179
rect 26240 37136 26292 37145
rect 28448 37204 28500 37256
rect 31208 37272 31260 37324
rect 27436 37136 27488 37188
rect 27344 37068 27396 37120
rect 27620 37179 27672 37188
rect 27620 37145 27629 37179
rect 27629 37145 27663 37179
rect 27663 37145 27672 37179
rect 27620 37136 27672 37145
rect 40776 37247 40828 37256
rect 40776 37213 40785 37247
rect 40785 37213 40819 37247
rect 40819 37213 40828 37247
rect 40776 37204 40828 37213
rect 31852 37179 31904 37188
rect 31852 37145 31861 37179
rect 31861 37145 31895 37179
rect 31895 37145 31904 37179
rect 31852 37136 31904 37145
rect 35624 37136 35676 37188
rect 31484 37068 31536 37120
rect 40960 37111 41012 37120
rect 40960 37077 40969 37111
rect 40969 37077 41003 37111
rect 41003 37077 41012 37111
rect 40960 37068 41012 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 5264 36864 5316 36916
rect 3792 36839 3844 36848
rect 3792 36805 3801 36839
rect 3801 36805 3835 36839
rect 3835 36805 3844 36839
rect 3792 36796 3844 36805
rect 1768 36771 1820 36780
rect 1768 36737 1777 36771
rect 1777 36737 1811 36771
rect 1811 36737 1820 36771
rect 1768 36728 1820 36737
rect 5724 36728 5776 36780
rect 6368 36728 6420 36780
rect 6920 36864 6972 36916
rect 7288 36864 7340 36916
rect 10692 36864 10744 36916
rect 6736 36728 6788 36780
rect 7104 36728 7156 36780
rect 7288 36771 7340 36780
rect 7288 36737 7298 36771
rect 7298 36737 7332 36771
rect 7332 36737 7340 36771
rect 7288 36728 7340 36737
rect 8300 36796 8352 36848
rect 7748 36771 7800 36780
rect 7748 36737 7757 36771
rect 7757 36737 7791 36771
rect 7791 36737 7800 36771
rect 7748 36728 7800 36737
rect 10232 36728 10284 36780
rect 12440 36796 12492 36848
rect 14096 36839 14148 36848
rect 14096 36805 14105 36839
rect 14105 36805 14139 36839
rect 14139 36805 14148 36839
rect 14096 36796 14148 36805
rect 2044 36703 2096 36712
rect 2044 36669 2053 36703
rect 2053 36669 2087 36703
rect 2087 36669 2096 36703
rect 2044 36660 2096 36669
rect 4068 36524 4120 36576
rect 7196 36703 7248 36712
rect 7196 36669 7205 36703
rect 7205 36669 7239 36703
rect 7239 36669 7248 36703
rect 7196 36660 7248 36669
rect 7380 36703 7432 36712
rect 7380 36669 7389 36703
rect 7389 36669 7423 36703
rect 7423 36669 7432 36703
rect 7380 36660 7432 36669
rect 7564 36660 7616 36712
rect 10784 36660 10836 36712
rect 8668 36592 8720 36644
rect 6092 36567 6144 36576
rect 6092 36533 6101 36567
rect 6101 36533 6135 36567
rect 6135 36533 6144 36567
rect 6092 36524 6144 36533
rect 6460 36567 6512 36576
rect 6460 36533 6469 36567
rect 6469 36533 6503 36567
rect 6503 36533 6512 36567
rect 6460 36524 6512 36533
rect 6920 36524 6972 36576
rect 13912 36660 13964 36712
rect 15016 36728 15068 36780
rect 14648 36703 14700 36712
rect 14648 36669 14657 36703
rect 14657 36669 14691 36703
rect 14691 36669 14700 36703
rect 14648 36660 14700 36669
rect 15752 36728 15804 36780
rect 16212 36728 16264 36780
rect 16856 36771 16908 36780
rect 16856 36737 16865 36771
rect 16865 36737 16899 36771
rect 16899 36737 16908 36771
rect 16856 36728 16908 36737
rect 17684 36796 17736 36848
rect 14280 36592 14332 36644
rect 16488 36660 16540 36712
rect 18052 36771 18104 36780
rect 18052 36737 18061 36771
rect 18061 36737 18095 36771
rect 18095 36737 18104 36771
rect 18052 36728 18104 36737
rect 18328 36771 18380 36780
rect 18328 36737 18337 36771
rect 18337 36737 18371 36771
rect 18371 36737 18380 36771
rect 18328 36728 18380 36737
rect 18420 36771 18472 36780
rect 18420 36737 18429 36771
rect 18429 36737 18463 36771
rect 18463 36737 18472 36771
rect 18420 36728 18472 36737
rect 14832 36567 14884 36576
rect 14832 36533 14841 36567
rect 14841 36533 14875 36567
rect 14875 36533 14884 36567
rect 14832 36524 14884 36533
rect 14924 36524 14976 36576
rect 15200 36567 15252 36576
rect 15200 36533 15209 36567
rect 15209 36533 15243 36567
rect 15243 36533 15252 36567
rect 15200 36524 15252 36533
rect 15384 36524 15436 36576
rect 17040 36524 17092 36576
rect 17316 36567 17368 36576
rect 17316 36533 17325 36567
rect 17325 36533 17359 36567
rect 17359 36533 17368 36567
rect 17316 36524 17368 36533
rect 18236 36592 18288 36644
rect 18604 36703 18656 36712
rect 18604 36669 18613 36703
rect 18613 36669 18647 36703
rect 18647 36669 18656 36703
rect 18604 36660 18656 36669
rect 18972 36592 19024 36644
rect 19156 36771 19208 36780
rect 19156 36737 19165 36771
rect 19165 36737 19199 36771
rect 19199 36737 19208 36771
rect 19156 36728 19208 36737
rect 20168 36796 20220 36848
rect 22652 36864 22704 36916
rect 24768 36864 24820 36916
rect 25228 36864 25280 36916
rect 27436 36864 27488 36916
rect 28172 36864 28224 36916
rect 20996 36728 21048 36780
rect 23756 36728 23808 36780
rect 23940 36728 23992 36780
rect 27252 36771 27304 36780
rect 27252 36737 27261 36771
rect 27261 36737 27295 36771
rect 27295 36737 27304 36771
rect 27252 36728 27304 36737
rect 27344 36728 27396 36780
rect 19432 36660 19484 36712
rect 19892 36703 19944 36712
rect 19892 36669 19901 36703
rect 19901 36669 19935 36703
rect 19935 36669 19944 36703
rect 19892 36660 19944 36669
rect 19616 36592 19668 36644
rect 17592 36524 17644 36576
rect 18880 36567 18932 36576
rect 18880 36533 18889 36567
rect 18889 36533 18923 36567
rect 18923 36533 18932 36567
rect 18880 36524 18932 36533
rect 20536 36524 20588 36576
rect 22836 36703 22888 36712
rect 22836 36669 22845 36703
rect 22845 36669 22879 36703
rect 22879 36669 22888 36703
rect 22836 36660 22888 36669
rect 27528 36771 27580 36780
rect 27528 36737 27537 36771
rect 27537 36737 27571 36771
rect 27571 36737 27580 36771
rect 27528 36728 27580 36737
rect 27712 36796 27764 36848
rect 31852 36864 31904 36916
rect 40040 36864 40092 36916
rect 30012 36771 30064 36780
rect 30012 36737 30021 36771
rect 30021 36737 30055 36771
rect 30055 36737 30064 36771
rect 30012 36728 30064 36737
rect 27804 36660 27856 36712
rect 28172 36703 28224 36712
rect 28172 36669 28181 36703
rect 28181 36669 28215 36703
rect 28215 36669 28224 36703
rect 28172 36660 28224 36669
rect 29828 36660 29880 36712
rect 30196 36592 30248 36644
rect 28724 36524 28776 36576
rect 29368 36524 29420 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2044 36320 2096 36372
rect 3424 36227 3476 36236
rect 3424 36193 3433 36227
rect 3433 36193 3467 36227
rect 3467 36193 3476 36227
rect 3424 36184 3476 36193
rect 4068 36320 4120 36372
rect 6920 36363 6972 36372
rect 6920 36329 6929 36363
rect 6929 36329 6963 36363
rect 6963 36329 6972 36363
rect 6920 36320 6972 36329
rect 7564 36320 7616 36372
rect 10324 36320 10376 36372
rect 10784 36363 10836 36372
rect 10784 36329 10793 36363
rect 10793 36329 10827 36363
rect 10827 36329 10836 36363
rect 10784 36320 10836 36329
rect 12808 36320 12860 36372
rect 14832 36320 14884 36372
rect 15016 36320 15068 36372
rect 16304 36320 16356 36372
rect 16856 36320 16908 36372
rect 17316 36320 17368 36372
rect 18420 36320 18472 36372
rect 19892 36320 19944 36372
rect 23756 36320 23808 36372
rect 5724 36252 5776 36304
rect 7932 36252 7984 36304
rect 7012 36184 7064 36236
rect 6092 36116 6144 36168
rect 3792 36048 3844 36100
rect 4160 36048 4212 36100
rect 3976 35980 4028 36032
rect 5540 36023 5592 36032
rect 5540 35989 5549 36023
rect 5549 35989 5583 36023
rect 5583 35989 5592 36023
rect 5540 35980 5592 35989
rect 8208 36116 8260 36168
rect 8300 36116 8352 36168
rect 10232 36252 10284 36304
rect 12716 36227 12768 36236
rect 12716 36193 12725 36227
rect 12725 36193 12759 36227
rect 12759 36193 12768 36227
rect 12716 36184 12768 36193
rect 15844 36252 15896 36304
rect 13728 36227 13780 36236
rect 13728 36193 13737 36227
rect 13737 36193 13771 36227
rect 13771 36193 13780 36227
rect 13728 36184 13780 36193
rect 7748 36091 7800 36100
rect 7748 36057 7757 36091
rect 7757 36057 7791 36091
rect 7791 36057 7800 36091
rect 7748 36048 7800 36057
rect 8116 36048 8168 36100
rect 8852 36048 8904 36100
rect 10048 36048 10100 36100
rect 10508 36159 10560 36168
rect 10508 36125 10517 36159
rect 10517 36125 10551 36159
rect 10551 36125 10560 36159
rect 10508 36116 10560 36125
rect 10968 36116 11020 36168
rect 12532 36116 12584 36168
rect 11060 36048 11112 36100
rect 10692 35980 10744 36032
rect 18512 36295 18564 36304
rect 18512 36261 18521 36295
rect 18521 36261 18555 36295
rect 18555 36261 18564 36295
rect 18512 36252 18564 36261
rect 15936 36116 15988 36168
rect 16488 36116 16540 36168
rect 18052 36116 18104 36168
rect 19432 36252 19484 36304
rect 19616 36252 19668 36304
rect 20168 36252 20220 36304
rect 22836 36252 22888 36304
rect 24216 36252 24268 36304
rect 25964 36252 26016 36304
rect 28356 36320 28408 36372
rect 28448 36363 28500 36372
rect 28448 36329 28457 36363
rect 28457 36329 28491 36363
rect 28491 36329 28500 36363
rect 28448 36320 28500 36329
rect 28724 36363 28776 36372
rect 28724 36329 28733 36363
rect 28733 36329 28767 36363
rect 28767 36329 28776 36363
rect 28724 36320 28776 36329
rect 29736 36363 29788 36372
rect 29736 36329 29745 36363
rect 29745 36329 29779 36363
rect 29779 36329 29788 36363
rect 29736 36320 29788 36329
rect 40776 36320 40828 36372
rect 18880 36184 18932 36236
rect 16212 36048 16264 36100
rect 17868 36048 17920 36100
rect 18236 36048 18288 36100
rect 18972 36159 19024 36168
rect 18972 36125 18981 36159
rect 18981 36125 19015 36159
rect 19015 36125 19024 36159
rect 18972 36116 19024 36125
rect 19248 36159 19300 36168
rect 19248 36125 19257 36159
rect 19257 36125 19291 36159
rect 19291 36125 19300 36159
rect 19248 36116 19300 36125
rect 22376 36184 22428 36236
rect 27988 36184 28040 36236
rect 19984 36116 20036 36168
rect 25596 36116 25648 36168
rect 27528 36116 27580 36168
rect 29368 36184 29420 36236
rect 25872 36048 25924 36100
rect 25964 36048 26016 36100
rect 26516 36048 26568 36100
rect 28264 36159 28316 36168
rect 28264 36125 28273 36159
rect 28273 36125 28307 36159
rect 28307 36125 28316 36159
rect 28264 36116 28316 36125
rect 29000 36116 29052 36168
rect 28632 36091 28684 36100
rect 28632 36057 28641 36091
rect 28641 36057 28675 36091
rect 28675 36057 28684 36091
rect 28632 36048 28684 36057
rect 29828 36159 29880 36168
rect 29828 36125 29837 36159
rect 29837 36125 29871 36159
rect 29871 36125 29880 36159
rect 29828 36116 29880 36125
rect 30012 36184 30064 36236
rect 31852 36159 31904 36168
rect 31852 36125 31861 36159
rect 31861 36125 31895 36159
rect 31895 36125 31904 36159
rect 31852 36116 31904 36125
rect 31944 36159 31996 36168
rect 31944 36125 31953 36159
rect 31953 36125 31987 36159
rect 31987 36125 31996 36159
rect 31944 36116 31996 36125
rect 24124 35980 24176 36032
rect 26240 35980 26292 36032
rect 27252 35980 27304 36032
rect 28080 35980 28132 36032
rect 28908 35980 28960 36032
rect 31116 36048 31168 36100
rect 34152 36116 34204 36168
rect 32128 36023 32180 36032
rect 32128 35989 32137 36023
rect 32137 35989 32171 36023
rect 32171 35989 32180 36023
rect 32128 35980 32180 35989
rect 33140 35980 33192 36032
rect 33876 35980 33928 36032
rect 33968 36023 34020 36032
rect 33968 35989 33977 36023
rect 33977 35989 34011 36023
rect 34011 35989 34020 36023
rect 33968 35980 34020 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4160 35776 4212 35828
rect 8116 35776 8168 35828
rect 5080 35683 5132 35692
rect 5080 35649 5089 35683
rect 5089 35649 5123 35683
rect 5123 35649 5132 35683
rect 5080 35640 5132 35649
rect 5540 35640 5592 35692
rect 5356 35615 5408 35624
rect 5356 35581 5365 35615
rect 5365 35581 5399 35615
rect 5399 35581 5408 35615
rect 5356 35572 5408 35581
rect 6460 35640 6512 35692
rect 7012 35640 7064 35692
rect 10968 35776 11020 35828
rect 14464 35776 14516 35828
rect 16212 35776 16264 35828
rect 10416 35708 10468 35760
rect 19432 35776 19484 35828
rect 6552 35572 6604 35624
rect 9956 35572 10008 35624
rect 10232 35615 10284 35624
rect 10232 35581 10241 35615
rect 10241 35581 10275 35615
rect 10275 35581 10284 35615
rect 10232 35572 10284 35581
rect 10968 35640 11020 35692
rect 17316 35708 17368 35760
rect 14924 35640 14976 35692
rect 13636 35572 13688 35624
rect 15936 35640 15988 35692
rect 18052 35640 18104 35692
rect 19156 35640 19208 35692
rect 20628 35640 20680 35692
rect 21916 35640 21968 35692
rect 22376 35640 22428 35692
rect 23480 35776 23532 35828
rect 24676 35776 24728 35828
rect 24952 35776 25004 35828
rect 25320 35776 25372 35828
rect 23940 35708 23992 35760
rect 24124 35683 24176 35692
rect 24124 35649 24133 35683
rect 24133 35649 24167 35683
rect 24167 35649 24176 35683
rect 24124 35640 24176 35649
rect 14280 35504 14332 35556
rect 15384 35504 15436 35556
rect 17408 35572 17460 35624
rect 19248 35572 19300 35624
rect 22560 35615 22612 35624
rect 22560 35581 22569 35615
rect 22569 35581 22603 35615
rect 22603 35581 22612 35615
rect 22560 35572 22612 35581
rect 15568 35504 15620 35556
rect 23112 35572 23164 35624
rect 24584 35640 24636 35692
rect 24676 35683 24728 35692
rect 24676 35649 24685 35683
rect 24685 35649 24719 35683
rect 24719 35649 24728 35683
rect 24676 35640 24728 35649
rect 24768 35615 24820 35624
rect 24768 35581 24777 35615
rect 24777 35581 24811 35615
rect 24811 35581 24820 35615
rect 24768 35572 24820 35581
rect 24860 35615 24912 35624
rect 24860 35581 24869 35615
rect 24869 35581 24903 35615
rect 24903 35581 24912 35615
rect 24860 35572 24912 35581
rect 25228 35751 25280 35760
rect 25228 35717 25237 35751
rect 25237 35717 25271 35751
rect 25271 35717 25280 35751
rect 26240 35776 26292 35828
rect 25228 35708 25280 35717
rect 27528 35708 27580 35760
rect 28172 35708 28224 35760
rect 29736 35708 29788 35760
rect 23296 35504 23348 35556
rect 25596 35640 25648 35692
rect 25688 35683 25740 35692
rect 25688 35649 25697 35683
rect 25697 35649 25731 35683
rect 25731 35649 25740 35683
rect 25688 35640 25740 35649
rect 26424 35640 26476 35692
rect 29920 35683 29972 35692
rect 29920 35649 29929 35683
rect 29929 35649 29963 35683
rect 29963 35649 29972 35683
rect 29920 35640 29972 35649
rect 30104 35683 30156 35692
rect 30104 35649 30134 35683
rect 30134 35649 30156 35683
rect 30104 35640 30156 35649
rect 25872 35572 25924 35624
rect 26056 35572 26108 35624
rect 27528 35572 27580 35624
rect 29276 35572 29328 35624
rect 29828 35572 29880 35624
rect 30288 35683 30340 35692
rect 30288 35649 30297 35683
rect 30297 35649 30331 35683
rect 30331 35649 30340 35683
rect 30288 35640 30340 35649
rect 31852 35708 31904 35760
rect 31116 35683 31168 35692
rect 31116 35649 31150 35683
rect 31150 35649 31168 35683
rect 31116 35640 31168 35649
rect 31760 35640 31812 35692
rect 32128 35708 32180 35760
rect 33140 35751 33192 35760
rect 33140 35717 33149 35751
rect 33149 35717 33183 35751
rect 33183 35717 33192 35751
rect 33140 35708 33192 35717
rect 6828 35436 6880 35488
rect 9864 35479 9916 35488
rect 9864 35445 9873 35479
rect 9873 35445 9907 35479
rect 9907 35445 9916 35479
rect 9864 35436 9916 35445
rect 10140 35436 10192 35488
rect 15108 35479 15160 35488
rect 15108 35445 15117 35479
rect 15117 35445 15151 35479
rect 15151 35445 15160 35479
rect 15108 35436 15160 35445
rect 16488 35436 16540 35488
rect 17224 35436 17276 35488
rect 17960 35436 18012 35488
rect 21824 35479 21876 35488
rect 21824 35445 21833 35479
rect 21833 35445 21867 35479
rect 21867 35445 21876 35479
rect 21824 35436 21876 35445
rect 22652 35436 22704 35488
rect 24400 35436 24452 35488
rect 24584 35436 24636 35488
rect 25136 35436 25188 35488
rect 25688 35479 25740 35488
rect 25688 35445 25697 35479
rect 25697 35445 25731 35479
rect 25731 35445 25740 35479
rect 25688 35436 25740 35445
rect 31116 35504 31168 35556
rect 32128 35572 32180 35624
rect 34520 35640 34572 35692
rect 34244 35572 34296 35624
rect 31944 35504 31996 35556
rect 33784 35547 33836 35556
rect 33784 35513 33793 35547
rect 33793 35513 33827 35547
rect 33827 35513 33836 35547
rect 33784 35504 33836 35513
rect 30472 35436 30524 35488
rect 31024 35479 31076 35488
rect 31024 35445 31033 35479
rect 31033 35445 31067 35479
rect 31067 35445 31076 35479
rect 31024 35436 31076 35445
rect 31392 35436 31444 35488
rect 34152 35436 34204 35488
rect 34336 35479 34388 35488
rect 34336 35445 34345 35479
rect 34345 35445 34379 35479
rect 34379 35445 34388 35479
rect 34336 35436 34388 35445
rect 34704 35436 34756 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 7748 35232 7800 35284
rect 8760 35232 8812 35284
rect 9864 35232 9916 35284
rect 4712 35096 4764 35148
rect 7564 35096 7616 35148
rect 11520 35096 11572 35148
rect 12256 35096 12308 35148
rect 4068 35028 4120 35080
rect 7288 35028 7340 35080
rect 10048 35071 10100 35080
rect 10048 35037 10057 35071
rect 10057 35037 10091 35071
rect 10091 35037 10100 35071
rect 10048 35028 10100 35037
rect 10140 35071 10192 35080
rect 10140 35037 10149 35071
rect 10149 35037 10183 35071
rect 10183 35037 10192 35071
rect 10140 35028 10192 35037
rect 10600 35028 10652 35080
rect 10508 34960 10560 35012
rect 11244 35028 11296 35080
rect 11704 35071 11756 35080
rect 11704 35037 11713 35071
rect 11713 35037 11747 35071
rect 11747 35037 11756 35071
rect 11704 35028 11756 35037
rect 13544 35232 13596 35284
rect 15568 35232 15620 35284
rect 17500 35232 17552 35284
rect 21088 35232 21140 35284
rect 23020 35232 23072 35284
rect 15844 35164 15896 35216
rect 16304 35096 16356 35148
rect 15752 35028 15804 35080
rect 16212 35028 16264 35080
rect 14556 34960 14608 35012
rect 16488 35071 16540 35080
rect 16488 35037 16497 35071
rect 16497 35037 16531 35071
rect 16531 35037 16540 35071
rect 16488 35028 16540 35037
rect 19432 35028 19484 35080
rect 21824 35096 21876 35148
rect 23388 35164 23440 35216
rect 23572 35164 23624 35216
rect 24584 35164 24636 35216
rect 25136 35232 25188 35284
rect 26424 35275 26476 35284
rect 26424 35241 26433 35275
rect 26433 35241 26467 35275
rect 26467 35241 26476 35275
rect 26424 35232 26476 35241
rect 26792 35275 26844 35284
rect 26792 35241 26801 35275
rect 26801 35241 26835 35275
rect 26835 35241 26844 35275
rect 26792 35232 26844 35241
rect 27068 35275 27120 35284
rect 27068 35241 27077 35275
rect 27077 35241 27111 35275
rect 27111 35241 27120 35275
rect 27068 35232 27120 35241
rect 27160 35275 27212 35284
rect 27160 35241 27169 35275
rect 27169 35241 27203 35275
rect 27203 35241 27212 35275
rect 27160 35232 27212 35241
rect 29184 35275 29236 35284
rect 29184 35241 29193 35275
rect 29193 35241 29227 35275
rect 29227 35241 29236 35275
rect 29184 35232 29236 35241
rect 31024 35232 31076 35284
rect 31116 35232 31168 35284
rect 9772 34935 9824 34944
rect 9772 34901 9797 34935
rect 9797 34901 9824 34935
rect 9772 34892 9824 34901
rect 9956 34892 10008 34944
rect 10324 34935 10376 34944
rect 10324 34901 10333 34935
rect 10333 34901 10367 34935
rect 10367 34901 10376 34935
rect 10324 34892 10376 34901
rect 11612 34892 11664 34944
rect 11888 34935 11940 34944
rect 11888 34901 11897 34935
rect 11897 34901 11931 34935
rect 11931 34901 11940 34935
rect 11888 34892 11940 34901
rect 14096 34892 14148 34944
rect 20352 34960 20404 35012
rect 20260 34935 20312 34944
rect 20260 34901 20269 34935
rect 20269 34901 20303 34935
rect 20303 34901 20312 34935
rect 20260 34892 20312 34901
rect 21732 34892 21784 34944
rect 24216 35096 24268 35148
rect 23112 35071 23164 35080
rect 23112 35037 23121 35071
rect 23121 35037 23155 35071
rect 23155 35037 23164 35071
rect 23112 35028 23164 35037
rect 23204 35071 23256 35080
rect 23204 35037 23213 35071
rect 23213 35037 23247 35071
rect 23247 35037 23256 35071
rect 23204 35028 23256 35037
rect 22928 35003 22980 35012
rect 22928 34969 22937 35003
rect 22937 34969 22971 35003
rect 22971 34969 22980 35003
rect 22928 34960 22980 34969
rect 24124 35028 24176 35080
rect 24400 35071 24452 35080
rect 24400 35037 24409 35071
rect 24409 35037 24443 35071
rect 24443 35037 24452 35071
rect 24400 35028 24452 35037
rect 24584 35071 24636 35080
rect 24584 35037 24591 35071
rect 24591 35037 24636 35071
rect 24584 35028 24636 35037
rect 27344 35164 27396 35216
rect 25964 35096 26016 35148
rect 25044 35028 25096 35080
rect 25136 35071 25188 35080
rect 25136 35037 25145 35071
rect 25145 35037 25179 35071
rect 25179 35037 25188 35071
rect 25136 35028 25188 35037
rect 25320 35071 25372 35080
rect 25320 35037 25327 35071
rect 25327 35037 25372 35071
rect 25320 35028 25372 35037
rect 25412 35071 25464 35080
rect 25412 35037 25421 35071
rect 25421 35037 25455 35071
rect 25455 35037 25464 35071
rect 25412 35028 25464 35037
rect 25504 35071 25556 35080
rect 25504 35037 25513 35071
rect 25513 35037 25547 35071
rect 25547 35037 25556 35071
rect 25504 35028 25556 35037
rect 26148 35028 26200 35080
rect 26240 35071 26292 35080
rect 26240 35037 26249 35071
rect 26249 35037 26283 35071
rect 26283 35037 26292 35071
rect 26240 35028 26292 35037
rect 29552 35096 29604 35148
rect 25780 34960 25832 35012
rect 26608 35003 26660 35012
rect 26608 34969 26617 35003
rect 26617 34969 26651 35003
rect 26651 34969 26660 35003
rect 26608 34960 26660 34969
rect 22560 34935 22612 34944
rect 22560 34901 22569 34935
rect 22569 34901 22603 34935
rect 22603 34901 22612 34935
rect 22560 34892 22612 34901
rect 23664 34892 23716 34944
rect 24308 34892 24360 34944
rect 25044 34935 25096 34944
rect 25044 34901 25053 34935
rect 25053 34901 25087 34935
rect 25087 34901 25096 34935
rect 25044 34892 25096 34901
rect 25412 34892 25464 34944
rect 26240 34892 26292 34944
rect 26332 34892 26384 34944
rect 26976 35028 27028 35080
rect 27528 35028 27580 35080
rect 28908 35071 28960 35080
rect 28908 35037 28917 35071
rect 28917 35037 28951 35071
rect 28951 35037 28960 35071
rect 28908 35028 28960 35037
rect 29000 35028 29052 35080
rect 31024 35139 31076 35148
rect 31024 35105 31033 35139
rect 31033 35105 31067 35139
rect 31067 35105 31076 35139
rect 31024 35096 31076 35105
rect 33508 35275 33560 35284
rect 33508 35241 33517 35275
rect 33517 35241 33551 35275
rect 33551 35241 33560 35275
rect 33508 35232 33560 35241
rect 34704 35232 34756 35284
rect 36084 35275 36136 35284
rect 36084 35241 36093 35275
rect 36093 35241 36127 35275
rect 36127 35241 36136 35275
rect 36084 35232 36136 35241
rect 34244 35207 34296 35216
rect 34244 35173 34253 35207
rect 34253 35173 34287 35207
rect 34287 35173 34296 35207
rect 34244 35164 34296 35173
rect 28816 34960 28868 35012
rect 29736 34960 29788 35012
rect 31392 35071 31444 35080
rect 31392 35037 31401 35071
rect 31401 35037 31435 35071
rect 31435 35037 31444 35071
rect 31392 35028 31444 35037
rect 32588 35096 32640 35148
rect 33784 35096 33836 35148
rect 32864 35028 32916 35080
rect 33968 35028 34020 35080
rect 34336 35028 34388 35080
rect 27252 34892 27304 34944
rect 29460 34892 29512 34944
rect 30012 34892 30064 34944
rect 31116 34935 31168 34944
rect 31116 34901 31125 34935
rect 31125 34901 31159 34935
rect 31159 34901 31168 34935
rect 31116 34892 31168 34901
rect 31576 34960 31628 35012
rect 31668 35003 31720 35012
rect 31668 34969 31677 35003
rect 31677 34969 31711 35003
rect 31711 34969 31720 35003
rect 31668 34960 31720 34969
rect 31760 34960 31812 35012
rect 32588 34960 32640 35012
rect 34060 34892 34112 34944
rect 36360 34892 36412 34944
rect 36820 34892 36872 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 1032 34688 1084 34740
rect 7564 34688 7616 34740
rect 9680 34731 9732 34740
rect 9680 34697 9689 34731
rect 9689 34697 9723 34731
rect 9723 34697 9732 34731
rect 9680 34688 9732 34697
rect 10324 34688 10376 34740
rect 10968 34731 11020 34740
rect 10968 34697 10977 34731
rect 10977 34697 11011 34731
rect 11011 34697 11020 34731
rect 10968 34688 11020 34697
rect 11244 34688 11296 34740
rect 6552 34620 6604 34672
rect 1860 34595 1912 34604
rect 1860 34561 1869 34595
rect 1869 34561 1903 34595
rect 1903 34561 1912 34595
rect 1860 34552 1912 34561
rect 6920 34552 6972 34604
rect 11520 34663 11572 34672
rect 11520 34629 11529 34663
rect 11529 34629 11563 34663
rect 11563 34629 11572 34663
rect 11520 34620 11572 34629
rect 12072 34620 12124 34672
rect 13084 34688 13136 34740
rect 7564 34484 7616 34536
rect 10416 34552 10468 34604
rect 11612 34552 11664 34604
rect 11888 34552 11940 34604
rect 12348 34595 12400 34604
rect 12348 34561 12357 34595
rect 12357 34561 12391 34595
rect 12391 34561 12400 34595
rect 12348 34552 12400 34561
rect 12624 34552 12676 34604
rect 12808 34552 12860 34604
rect 13544 34552 13596 34604
rect 14280 34688 14332 34740
rect 14464 34663 14516 34672
rect 14464 34629 14473 34663
rect 14473 34629 14507 34663
rect 14507 34629 14516 34663
rect 14464 34620 14516 34629
rect 15108 34620 15160 34672
rect 17684 34688 17736 34740
rect 19984 34688 20036 34740
rect 20076 34731 20128 34740
rect 20076 34697 20085 34731
rect 20085 34697 20119 34731
rect 20119 34697 20128 34731
rect 20076 34688 20128 34697
rect 20628 34731 20680 34740
rect 20628 34697 20637 34731
rect 20637 34697 20671 34731
rect 20671 34697 20680 34731
rect 20628 34688 20680 34697
rect 22928 34688 22980 34740
rect 23112 34688 23164 34740
rect 23480 34688 23532 34740
rect 4988 34416 5040 34468
rect 6184 34416 6236 34468
rect 7656 34416 7708 34468
rect 8944 34416 8996 34468
rect 11704 34484 11756 34536
rect 11336 34416 11388 34468
rect 14096 34484 14148 34536
rect 6920 34348 6972 34400
rect 7380 34391 7432 34400
rect 7380 34357 7389 34391
rect 7389 34357 7423 34391
rect 7423 34357 7432 34391
rect 7380 34348 7432 34357
rect 11152 34348 11204 34400
rect 12348 34348 12400 34400
rect 14648 34595 14700 34604
rect 14648 34561 14662 34595
rect 14662 34561 14696 34595
rect 14696 34561 14700 34595
rect 14648 34552 14700 34561
rect 14556 34484 14608 34536
rect 17224 34595 17276 34604
rect 17224 34561 17233 34595
rect 17233 34561 17267 34595
rect 17267 34561 17276 34595
rect 17224 34552 17276 34561
rect 16120 34348 16172 34400
rect 16764 34348 16816 34400
rect 17316 34416 17368 34468
rect 17592 34527 17644 34536
rect 17592 34493 17601 34527
rect 17601 34493 17635 34527
rect 17635 34493 17644 34527
rect 17592 34484 17644 34493
rect 17868 34595 17920 34604
rect 17868 34561 17877 34595
rect 17877 34561 17911 34595
rect 17911 34561 17920 34595
rect 20444 34663 20496 34672
rect 20444 34629 20453 34663
rect 20453 34629 20487 34663
rect 20487 34629 20496 34663
rect 20444 34620 20496 34629
rect 17868 34552 17920 34561
rect 19892 34595 19944 34604
rect 19892 34561 19901 34595
rect 19901 34561 19935 34595
rect 19935 34561 19944 34595
rect 19892 34552 19944 34561
rect 17776 34484 17828 34536
rect 19064 34416 19116 34468
rect 19432 34416 19484 34468
rect 21548 34552 21600 34604
rect 22836 34595 22888 34604
rect 22836 34561 22845 34595
rect 22845 34561 22879 34595
rect 22879 34561 22888 34595
rect 22836 34552 22888 34561
rect 24768 34688 24820 34740
rect 23940 34620 23992 34672
rect 26148 34688 26200 34740
rect 26424 34688 26476 34740
rect 26792 34731 26844 34740
rect 26792 34697 26801 34731
rect 26801 34697 26835 34731
rect 26835 34697 26844 34731
rect 26792 34688 26844 34697
rect 27620 34731 27672 34740
rect 27620 34697 27629 34731
rect 27629 34697 27663 34731
rect 27663 34697 27672 34731
rect 27620 34688 27672 34697
rect 18972 34348 19024 34400
rect 19984 34348 20036 34400
rect 20260 34416 20312 34468
rect 25504 34552 25556 34604
rect 24308 34484 24360 34536
rect 26424 34595 26476 34604
rect 26424 34561 26433 34595
rect 26433 34561 26467 34595
rect 26467 34561 26476 34595
rect 26424 34552 26476 34561
rect 26516 34595 26568 34604
rect 26516 34561 26525 34595
rect 26525 34561 26559 34595
rect 26559 34561 26568 34595
rect 26516 34552 26568 34561
rect 26700 34552 26752 34604
rect 26884 34552 26936 34604
rect 28264 34620 28316 34672
rect 28908 34620 28960 34672
rect 29092 34688 29144 34740
rect 29552 34688 29604 34740
rect 30104 34688 30156 34740
rect 30472 34688 30524 34740
rect 32772 34688 32824 34740
rect 33968 34688 34020 34740
rect 35348 34731 35400 34740
rect 35348 34697 35357 34731
rect 35357 34697 35391 34731
rect 35391 34697 35400 34731
rect 35348 34688 35400 34697
rect 29276 34620 29328 34672
rect 27344 34595 27396 34604
rect 27344 34561 27350 34595
rect 27350 34561 27384 34595
rect 27384 34561 27396 34595
rect 27344 34552 27396 34561
rect 28816 34552 28868 34604
rect 29460 34552 29512 34604
rect 29552 34595 29604 34604
rect 29552 34561 29561 34595
rect 29561 34561 29595 34595
rect 29595 34561 29604 34595
rect 29552 34552 29604 34561
rect 24584 34416 24636 34468
rect 20536 34348 20588 34400
rect 22652 34348 22704 34400
rect 23848 34348 23900 34400
rect 24400 34348 24452 34400
rect 26608 34348 26660 34400
rect 28908 34484 28960 34536
rect 29736 34620 29788 34672
rect 30012 34620 30064 34672
rect 30196 34620 30248 34672
rect 31576 34620 31628 34672
rect 32312 34663 32364 34672
rect 32312 34629 32321 34663
rect 32321 34629 32355 34663
rect 32355 34629 32364 34663
rect 32312 34620 32364 34629
rect 31300 34552 31352 34604
rect 32680 34595 32732 34604
rect 32680 34561 32689 34595
rect 32689 34561 32723 34595
rect 32723 34561 32732 34595
rect 32680 34552 32732 34561
rect 28540 34416 28592 34468
rect 32220 34527 32272 34536
rect 32220 34493 32229 34527
rect 32229 34493 32263 34527
rect 32263 34493 32272 34527
rect 32220 34484 32272 34493
rect 27160 34348 27212 34400
rect 28724 34348 28776 34400
rect 29368 34416 29420 34468
rect 29736 34416 29788 34468
rect 30564 34416 30616 34468
rect 33692 34552 33744 34604
rect 34152 34552 34204 34604
rect 33416 34527 33468 34536
rect 33416 34493 33425 34527
rect 33425 34493 33459 34527
rect 33459 34493 33468 34527
rect 35716 34552 35768 34604
rect 36360 34552 36412 34604
rect 33416 34484 33468 34493
rect 34796 34416 34848 34468
rect 35532 34484 35584 34536
rect 36452 34527 36504 34536
rect 36452 34493 36461 34527
rect 36461 34493 36495 34527
rect 36495 34493 36504 34527
rect 36452 34484 36504 34493
rect 37740 34484 37792 34536
rect 35440 34416 35492 34468
rect 36360 34416 36412 34468
rect 30288 34348 30340 34400
rect 33876 34348 33928 34400
rect 37464 34348 37516 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 5080 34144 5132 34196
rect 8300 34187 8352 34196
rect 8300 34153 8309 34187
rect 8309 34153 8343 34187
rect 8343 34153 8352 34187
rect 8300 34144 8352 34153
rect 9772 34187 9824 34196
rect 9772 34153 9781 34187
rect 9781 34153 9815 34187
rect 9815 34153 9824 34187
rect 9772 34144 9824 34153
rect 11704 34144 11756 34196
rect 5264 34076 5316 34128
rect 4068 34051 4120 34060
rect 4068 34017 4077 34051
rect 4077 34017 4111 34051
rect 4111 34017 4120 34051
rect 4068 34008 4120 34017
rect 5816 34076 5868 34128
rect 6920 34076 6972 34128
rect 4436 33940 4488 33992
rect 4712 33983 4764 33992
rect 4712 33949 4721 33983
rect 4721 33949 4755 33983
rect 4755 33949 4764 33983
rect 4712 33940 4764 33949
rect 4988 33940 5040 33992
rect 7380 34008 7432 34060
rect 9680 34076 9732 34128
rect 5724 33983 5776 33992
rect 5724 33949 5733 33983
rect 5733 33949 5767 33983
rect 5767 33949 5776 33983
rect 5724 33940 5776 33949
rect 6828 33940 6880 33992
rect 7012 33983 7064 33992
rect 7012 33949 7021 33983
rect 7021 33949 7055 33983
rect 7055 33949 7064 33983
rect 7012 33940 7064 33949
rect 4896 33872 4948 33924
rect 5264 33872 5316 33924
rect 5908 33915 5960 33924
rect 5908 33881 5917 33915
rect 5917 33881 5951 33915
rect 5951 33881 5960 33915
rect 5908 33872 5960 33881
rect 9680 33983 9732 33992
rect 9680 33949 9689 33983
rect 9689 33949 9723 33983
rect 9723 33949 9732 33983
rect 9680 33940 9732 33949
rect 4528 33804 4580 33856
rect 6920 33804 6972 33856
rect 7196 33847 7248 33856
rect 7196 33813 7205 33847
rect 7205 33813 7239 33847
rect 7239 33813 7248 33847
rect 7196 33804 7248 33813
rect 10692 33940 10744 33992
rect 12716 34144 12768 34196
rect 14464 34144 14516 34196
rect 16212 34144 16264 34196
rect 19892 34187 19944 34196
rect 19892 34153 19901 34187
rect 19901 34153 19935 34187
rect 19935 34153 19944 34187
rect 19892 34144 19944 34153
rect 20444 34187 20496 34196
rect 20444 34153 20453 34187
rect 20453 34153 20487 34187
rect 20487 34153 20496 34187
rect 20444 34144 20496 34153
rect 20536 34144 20588 34196
rect 11152 34008 11204 34060
rect 11060 33940 11112 33992
rect 11888 33983 11940 33992
rect 11888 33949 11897 33983
rect 11897 33949 11931 33983
rect 11931 33949 11940 33983
rect 11888 33940 11940 33949
rect 12808 33940 12860 33992
rect 12624 33872 12676 33924
rect 13176 33940 13228 33992
rect 13544 33940 13596 33992
rect 13452 33872 13504 33924
rect 13912 33983 13964 33992
rect 13912 33949 13921 33983
rect 13921 33949 13955 33983
rect 13955 33949 13964 33983
rect 13912 33940 13964 33949
rect 18236 34076 18288 34128
rect 16304 34008 16356 34060
rect 18696 34008 18748 34060
rect 19064 34008 19116 34060
rect 20536 34008 20588 34060
rect 21456 34051 21508 34060
rect 21456 34017 21465 34051
rect 21465 34017 21499 34051
rect 21499 34017 21508 34051
rect 21456 34008 21508 34017
rect 22100 34008 22152 34060
rect 14464 33983 14516 33992
rect 14464 33949 14473 33983
rect 14473 33949 14507 33983
rect 14507 33949 14516 33983
rect 14464 33940 14516 33949
rect 14556 33983 14608 33992
rect 14556 33949 14565 33983
rect 14565 33949 14599 33983
rect 14599 33949 14608 33983
rect 14556 33940 14608 33949
rect 15752 33940 15804 33992
rect 16764 33940 16816 33992
rect 16856 33983 16908 33992
rect 16856 33949 16865 33983
rect 16865 33949 16899 33983
rect 16899 33949 16908 33983
rect 16856 33940 16908 33949
rect 15200 33872 15252 33924
rect 16120 33872 16172 33924
rect 16212 33804 16264 33856
rect 18236 33872 18288 33924
rect 17040 33804 17092 33856
rect 17132 33804 17184 33856
rect 19616 33940 19668 33992
rect 19984 33940 20036 33992
rect 20260 33983 20312 33992
rect 20260 33949 20269 33983
rect 20269 33949 20303 33983
rect 20303 33949 20312 33983
rect 20260 33940 20312 33949
rect 18972 33915 19024 33924
rect 18972 33881 18981 33915
rect 18981 33881 19015 33915
rect 19015 33881 19024 33915
rect 18972 33872 19024 33881
rect 19064 33872 19116 33924
rect 18604 33804 18656 33856
rect 20076 33804 20128 33856
rect 20536 33872 20588 33924
rect 21364 33983 21416 33992
rect 21364 33949 21373 33983
rect 21373 33949 21407 33983
rect 21407 33949 21416 33983
rect 21364 33940 21416 33949
rect 22284 33983 22336 33992
rect 22284 33949 22293 33983
rect 22293 33949 22327 33983
rect 22327 33949 22336 33983
rect 22284 33940 22336 33949
rect 22560 34144 22612 34196
rect 25044 34144 25096 34196
rect 22836 34076 22888 34128
rect 24860 34119 24912 34128
rect 24860 34085 24869 34119
rect 24869 34085 24903 34119
rect 24903 34085 24912 34119
rect 24860 34076 24912 34085
rect 25596 34076 25648 34128
rect 25228 34008 25280 34060
rect 27620 34144 27672 34196
rect 28540 34144 28592 34196
rect 22652 33983 22704 33992
rect 22652 33949 22661 33983
rect 22661 33949 22695 33983
rect 22695 33949 22704 33983
rect 22652 33940 22704 33949
rect 21640 33804 21692 33856
rect 23572 33940 23624 33992
rect 23204 33872 23256 33924
rect 24124 33940 24176 33992
rect 24860 33940 24912 33992
rect 25688 33940 25740 33992
rect 27436 34076 27488 34128
rect 27160 33983 27212 33992
rect 27160 33949 27169 33983
rect 27169 33949 27203 33983
rect 27203 33949 27212 33983
rect 27160 33940 27212 33949
rect 27528 33983 27580 33992
rect 27528 33949 27537 33983
rect 27537 33949 27571 33983
rect 27571 33949 27580 33983
rect 27528 33940 27580 33949
rect 27436 33915 27488 33924
rect 27436 33881 27445 33915
rect 27445 33881 27479 33915
rect 27479 33881 27488 33915
rect 27436 33872 27488 33881
rect 33784 34144 33836 34196
rect 37464 34187 37516 34196
rect 37464 34153 37473 34187
rect 37473 34153 37507 34187
rect 37507 34153 37516 34187
rect 37464 34144 37516 34153
rect 28724 34076 28776 34128
rect 29276 34076 29328 34128
rect 28540 33983 28592 33992
rect 28540 33949 28549 33983
rect 28549 33949 28583 33983
rect 28583 33949 28592 33983
rect 28540 33940 28592 33949
rect 28816 33983 28868 33992
rect 28816 33949 28825 33983
rect 28825 33949 28859 33983
rect 28859 33949 28868 33983
rect 28816 33940 28868 33949
rect 29000 33983 29052 33992
rect 29000 33949 29014 33983
rect 29014 33949 29048 33983
rect 29048 33949 29052 33983
rect 29000 33940 29052 33949
rect 29644 33983 29696 33992
rect 29644 33949 29654 33983
rect 29654 33949 29688 33983
rect 29688 33949 29696 33983
rect 29644 33940 29696 33949
rect 28908 33915 28960 33924
rect 28908 33881 28917 33915
rect 28917 33881 28951 33915
rect 28951 33881 28960 33915
rect 28908 33872 28960 33881
rect 29460 33872 29512 33924
rect 30012 33983 30064 33992
rect 30012 33949 30026 33983
rect 30026 33949 30060 33983
rect 30060 33949 30064 33983
rect 30288 34051 30340 34060
rect 30288 34017 30297 34051
rect 30297 34017 30331 34051
rect 30331 34017 30340 34051
rect 30288 34008 30340 34017
rect 32220 34076 32272 34128
rect 32956 34076 33008 34128
rect 32588 34008 32640 34060
rect 33048 34008 33100 34060
rect 30012 33940 30064 33949
rect 30564 33983 30616 33992
rect 30564 33949 30573 33983
rect 30573 33949 30607 33983
rect 30607 33949 30616 33983
rect 30564 33940 30616 33949
rect 30656 33983 30708 33992
rect 30656 33949 30665 33983
rect 30665 33949 30699 33983
rect 30699 33949 30708 33983
rect 30656 33940 30708 33949
rect 32772 33940 32824 33992
rect 33600 33940 33652 33992
rect 35440 34076 35492 34128
rect 34796 34008 34848 34060
rect 36176 34008 36228 34060
rect 22928 33847 22980 33856
rect 22928 33813 22937 33847
rect 22937 33813 22971 33847
rect 22971 33813 22980 33847
rect 22928 33804 22980 33813
rect 24216 33847 24268 33856
rect 24216 33813 24225 33847
rect 24225 33813 24259 33847
rect 24259 33813 24268 33847
rect 24216 33804 24268 33813
rect 24676 33804 24728 33856
rect 25688 33804 25740 33856
rect 26516 33847 26568 33856
rect 26516 33813 26525 33847
rect 26525 33813 26559 33847
rect 26559 33813 26568 33847
rect 26516 33804 26568 33813
rect 26700 33804 26752 33856
rect 26792 33804 26844 33856
rect 27344 33804 27396 33856
rect 27712 33804 27764 33856
rect 29184 33847 29236 33856
rect 29184 33813 29193 33847
rect 29193 33813 29227 33847
rect 29227 33813 29236 33847
rect 29184 33804 29236 33813
rect 29368 33804 29420 33856
rect 30472 33804 30524 33856
rect 32128 33915 32180 33924
rect 32128 33881 32162 33915
rect 32162 33881 32180 33915
rect 32128 33872 32180 33881
rect 32312 33847 32364 33856
rect 32312 33813 32321 33847
rect 32321 33813 32355 33847
rect 32355 33813 32364 33847
rect 32312 33804 32364 33813
rect 32680 33804 32732 33856
rect 33784 33804 33836 33856
rect 34520 33940 34572 33992
rect 34888 33983 34940 33992
rect 34888 33949 34897 33983
rect 34897 33949 34931 33983
rect 34931 33949 34940 33983
rect 34888 33940 34940 33949
rect 36360 33872 36412 33924
rect 34612 33804 34664 33856
rect 35348 33804 35400 33856
rect 35440 33804 35492 33856
rect 35716 33804 35768 33856
rect 37372 33915 37424 33924
rect 37372 33881 37381 33915
rect 37381 33881 37415 33915
rect 37415 33881 37424 33915
rect 37372 33872 37424 33881
rect 37832 33872 37884 33924
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 6828 33600 6880 33652
rect 6920 33600 6972 33652
rect 9680 33600 9732 33652
rect 4436 33507 4488 33516
rect 4436 33473 4445 33507
rect 4445 33473 4479 33507
rect 4479 33473 4488 33507
rect 4436 33464 4488 33473
rect 4896 33464 4948 33516
rect 5908 33532 5960 33584
rect 6736 33532 6788 33584
rect 5264 33507 5316 33516
rect 5264 33473 5273 33507
rect 5273 33473 5307 33507
rect 5307 33473 5316 33507
rect 5264 33464 5316 33473
rect 6276 33464 6328 33516
rect 7472 33532 7524 33584
rect 8668 33507 8720 33516
rect 8668 33473 8677 33507
rect 8677 33473 8711 33507
rect 8711 33473 8720 33507
rect 8668 33464 8720 33473
rect 9128 33464 9180 33516
rect 5816 33328 5868 33380
rect 4528 33303 4580 33312
rect 4528 33269 4537 33303
rect 4537 33269 4571 33303
rect 4571 33269 4580 33303
rect 4528 33260 4580 33269
rect 4988 33303 5040 33312
rect 4988 33269 4997 33303
rect 4997 33269 5031 33303
rect 5031 33269 5040 33303
rect 4988 33260 5040 33269
rect 9680 33507 9732 33516
rect 9680 33473 9689 33507
rect 9689 33473 9723 33507
rect 9723 33473 9732 33507
rect 9680 33464 9732 33473
rect 9864 33396 9916 33448
rect 11888 33600 11940 33652
rect 12072 33600 12124 33652
rect 12624 33643 12676 33652
rect 12624 33609 12633 33643
rect 12633 33609 12667 33643
rect 12667 33609 12676 33643
rect 12624 33600 12676 33609
rect 13452 33600 13504 33652
rect 14464 33600 14516 33652
rect 11520 33575 11572 33584
rect 11520 33541 11529 33575
rect 11529 33541 11563 33575
rect 11563 33541 11572 33575
rect 11520 33532 11572 33541
rect 11336 33464 11388 33516
rect 13176 33532 13228 33584
rect 14004 33532 14056 33584
rect 10324 33396 10376 33448
rect 10876 33396 10928 33448
rect 12624 33464 12676 33516
rect 13084 33507 13136 33516
rect 13084 33473 13093 33507
rect 13093 33473 13127 33507
rect 13127 33473 13136 33507
rect 13084 33464 13136 33473
rect 11152 33328 11204 33380
rect 14648 33464 14700 33516
rect 14832 33507 14884 33516
rect 14832 33473 14841 33507
rect 14841 33473 14875 33507
rect 14875 33473 14884 33507
rect 14832 33464 14884 33473
rect 14556 33328 14608 33380
rect 10048 33260 10100 33312
rect 10232 33303 10284 33312
rect 10232 33269 10241 33303
rect 10241 33269 10275 33303
rect 10275 33269 10284 33303
rect 10232 33260 10284 33269
rect 10416 33303 10468 33312
rect 10416 33269 10425 33303
rect 10425 33269 10459 33303
rect 10459 33269 10468 33303
rect 10416 33260 10468 33269
rect 12348 33303 12400 33312
rect 12348 33269 12357 33303
rect 12357 33269 12391 33303
rect 12391 33269 12400 33303
rect 12348 33260 12400 33269
rect 16856 33600 16908 33652
rect 17132 33600 17184 33652
rect 17684 33643 17736 33652
rect 17684 33609 17693 33643
rect 17693 33609 17727 33643
rect 17727 33609 17736 33643
rect 17684 33600 17736 33609
rect 17776 33600 17828 33652
rect 17868 33600 17920 33652
rect 16120 33507 16172 33516
rect 16120 33473 16129 33507
rect 16129 33473 16163 33507
rect 16163 33473 16172 33507
rect 16120 33464 16172 33473
rect 16212 33464 16264 33516
rect 16764 33507 16816 33516
rect 16764 33473 16773 33507
rect 16773 33473 16807 33507
rect 16807 33473 16816 33507
rect 16764 33464 16816 33473
rect 17316 33507 17368 33516
rect 17316 33473 17325 33507
rect 17325 33473 17359 33507
rect 17359 33473 17368 33507
rect 17316 33464 17368 33473
rect 16028 33439 16080 33448
rect 16028 33405 16037 33439
rect 16037 33405 16071 33439
rect 16071 33405 16080 33439
rect 16028 33396 16080 33405
rect 17224 33439 17276 33448
rect 17224 33405 17233 33439
rect 17233 33405 17267 33439
rect 17267 33405 17276 33439
rect 17224 33396 17276 33405
rect 18236 33532 18288 33584
rect 19432 33464 19484 33516
rect 19524 33507 19576 33516
rect 19524 33473 19533 33507
rect 19533 33473 19567 33507
rect 19567 33473 19576 33507
rect 19524 33464 19576 33473
rect 22284 33600 22336 33652
rect 25136 33600 25188 33652
rect 26700 33600 26752 33652
rect 27528 33600 27580 33652
rect 27988 33600 28040 33652
rect 30012 33600 30064 33652
rect 33232 33643 33284 33652
rect 33232 33609 33241 33643
rect 33241 33609 33275 33643
rect 33275 33609 33284 33643
rect 33232 33600 33284 33609
rect 34888 33600 34940 33652
rect 35348 33600 35400 33652
rect 21180 33464 21232 33516
rect 22008 33464 22060 33516
rect 23020 33532 23072 33584
rect 29000 33532 29052 33584
rect 24860 33464 24912 33516
rect 18604 33396 18656 33448
rect 17868 33328 17920 33380
rect 20260 33396 20312 33448
rect 24032 33396 24084 33448
rect 25596 33464 25648 33516
rect 26976 33396 27028 33448
rect 27344 33464 27396 33516
rect 30472 33464 30524 33516
rect 32220 33464 32272 33516
rect 33600 33532 33652 33584
rect 33784 33532 33836 33584
rect 32956 33464 33008 33516
rect 33968 33507 34020 33516
rect 33968 33473 33977 33507
rect 33977 33473 34011 33507
rect 34011 33473 34020 33507
rect 33968 33464 34020 33473
rect 28908 33396 28960 33448
rect 29460 33396 29512 33448
rect 30288 33396 30340 33448
rect 32680 33396 32732 33448
rect 33600 33396 33652 33448
rect 35716 33507 35768 33516
rect 35716 33473 35725 33507
rect 35725 33473 35759 33507
rect 35759 33473 35768 33507
rect 35716 33464 35768 33473
rect 36176 33532 36228 33584
rect 22100 33328 22152 33380
rect 22376 33328 22428 33380
rect 15660 33260 15712 33312
rect 16948 33260 17000 33312
rect 20260 33260 20312 33312
rect 20904 33260 20956 33312
rect 21364 33303 21416 33312
rect 21364 33269 21373 33303
rect 21373 33269 21407 33303
rect 21407 33269 21416 33303
rect 21364 33260 21416 33269
rect 25228 33260 25280 33312
rect 25320 33303 25372 33312
rect 25320 33269 25329 33303
rect 25329 33269 25363 33303
rect 25363 33269 25372 33303
rect 25320 33260 25372 33269
rect 25504 33328 25556 33380
rect 25688 33371 25740 33380
rect 25688 33337 25697 33371
rect 25697 33337 25731 33371
rect 25731 33337 25740 33371
rect 25688 33328 25740 33337
rect 28816 33328 28868 33380
rect 35992 33396 36044 33448
rect 37280 33507 37332 33516
rect 37280 33473 37289 33507
rect 37289 33473 37323 33507
rect 37323 33473 37332 33507
rect 37280 33464 37332 33473
rect 37832 33464 37884 33516
rect 36636 33396 36688 33448
rect 38016 33464 38068 33516
rect 40592 33464 40644 33516
rect 25780 33260 25832 33312
rect 26332 33260 26384 33312
rect 26792 33260 26844 33312
rect 27436 33303 27488 33312
rect 27436 33269 27445 33303
rect 27445 33269 27479 33303
rect 27479 33269 27488 33303
rect 27436 33260 27488 33269
rect 27620 33260 27672 33312
rect 30564 33260 30616 33312
rect 32128 33303 32180 33312
rect 32128 33269 32137 33303
rect 32137 33269 32171 33303
rect 32171 33269 32180 33303
rect 32128 33260 32180 33269
rect 32772 33260 32824 33312
rect 34336 33328 34388 33380
rect 36360 33328 36412 33380
rect 39212 33439 39264 33448
rect 39212 33405 39221 33439
rect 39221 33405 39255 33439
rect 39255 33405 39264 33439
rect 39212 33396 39264 33405
rect 41052 33396 41104 33448
rect 38384 33328 38436 33380
rect 35716 33260 35768 33312
rect 40960 33303 41012 33312
rect 40960 33269 40969 33303
rect 40969 33269 41003 33303
rect 41003 33269 41012 33303
rect 40960 33260 41012 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 7288 33099 7340 33108
rect 7288 33065 7297 33099
rect 7297 33065 7331 33099
rect 7331 33065 7340 33099
rect 7288 33056 7340 33065
rect 11152 33056 11204 33108
rect 14556 33056 14608 33108
rect 15844 33099 15896 33108
rect 15844 33065 15853 33099
rect 15853 33065 15887 33099
rect 15887 33065 15896 33099
rect 15844 33056 15896 33065
rect 16120 33056 16172 33108
rect 16764 33056 16816 33108
rect 19524 33099 19576 33108
rect 19524 33065 19533 33099
rect 19533 33065 19567 33099
rect 19567 33065 19576 33099
rect 19524 33056 19576 33065
rect 20444 33056 20496 33108
rect 24768 33056 24820 33108
rect 26516 33056 26568 33108
rect 7104 32988 7156 33040
rect 8024 32988 8076 33040
rect 10784 32920 10836 32972
rect 15936 32920 15988 32972
rect 23388 32988 23440 33040
rect 20168 32963 20220 32972
rect 20168 32929 20177 32963
rect 20177 32929 20211 32963
rect 20211 32929 20220 32963
rect 20168 32920 20220 32929
rect 7196 32895 7248 32904
rect 7196 32861 7205 32895
rect 7205 32861 7239 32895
rect 7239 32861 7248 32895
rect 7196 32852 7248 32861
rect 11612 32895 11664 32904
rect 11612 32861 11621 32895
rect 11621 32861 11655 32895
rect 11655 32861 11664 32895
rect 11612 32852 11664 32861
rect 12072 32895 12124 32904
rect 12072 32861 12081 32895
rect 12081 32861 12115 32895
rect 12115 32861 12124 32895
rect 12072 32852 12124 32861
rect 15660 32852 15712 32904
rect 11980 32784 12032 32836
rect 14004 32784 14056 32836
rect 17316 32852 17368 32904
rect 15936 32784 15988 32836
rect 7656 32759 7708 32768
rect 7656 32725 7665 32759
rect 7665 32725 7699 32759
rect 7699 32725 7708 32759
rect 7656 32716 7708 32725
rect 9864 32716 9916 32768
rect 15660 32716 15712 32768
rect 15844 32716 15896 32768
rect 21364 32920 21416 32972
rect 20996 32852 21048 32904
rect 21180 32852 21232 32904
rect 24676 32963 24728 32972
rect 24676 32929 24685 32963
rect 24685 32929 24719 32963
rect 24719 32929 24728 32963
rect 24676 32920 24728 32929
rect 25872 32920 25924 32972
rect 27252 32920 27304 32972
rect 35992 33056 36044 33108
rect 30288 32988 30340 33040
rect 36360 32988 36412 33040
rect 18052 32716 18104 32768
rect 19984 32759 20036 32768
rect 19984 32725 19993 32759
rect 19993 32725 20027 32759
rect 20027 32725 20036 32759
rect 19984 32716 20036 32725
rect 20076 32716 20128 32768
rect 21824 32716 21876 32768
rect 22284 32716 22336 32768
rect 22744 32827 22796 32836
rect 22744 32793 22753 32827
rect 22753 32793 22787 32827
rect 22787 32793 22796 32827
rect 22744 32784 22796 32793
rect 25320 32852 25372 32904
rect 24860 32827 24912 32836
rect 24860 32793 24869 32827
rect 24869 32793 24903 32827
rect 24903 32793 24912 32827
rect 24860 32784 24912 32793
rect 26056 32895 26108 32904
rect 26056 32861 26065 32895
rect 26065 32861 26099 32895
rect 26099 32861 26108 32895
rect 26056 32852 26108 32861
rect 26700 32852 26752 32904
rect 27160 32852 27212 32904
rect 27528 32852 27580 32904
rect 28080 32852 28132 32904
rect 30380 32852 30432 32904
rect 30656 32852 30708 32904
rect 26608 32784 26660 32836
rect 27436 32784 27488 32836
rect 28264 32784 28316 32836
rect 23480 32716 23532 32768
rect 24676 32716 24728 32768
rect 26240 32759 26292 32768
rect 26240 32725 26249 32759
rect 26249 32725 26283 32759
rect 26283 32725 26292 32759
rect 26240 32716 26292 32725
rect 26332 32716 26384 32768
rect 26884 32716 26936 32768
rect 29276 32716 29328 32768
rect 30840 32716 30892 32768
rect 34152 32852 34204 32904
rect 34796 32852 34848 32904
rect 37372 33056 37424 33108
rect 38016 33056 38068 33108
rect 38384 33056 38436 33108
rect 41052 33099 41104 33108
rect 41052 33065 41061 33099
rect 41061 33065 41095 33099
rect 41095 33065 41104 33099
rect 41052 33056 41104 33065
rect 37096 32963 37148 32972
rect 37096 32929 37105 32963
rect 37105 32929 37139 32963
rect 37139 32929 37148 32963
rect 37096 32920 37148 32929
rect 37280 32920 37332 32972
rect 38476 32920 38528 32972
rect 37832 32784 37884 32836
rect 38108 32852 38160 32904
rect 38660 32852 38712 32904
rect 39856 32895 39908 32904
rect 39856 32861 39865 32895
rect 39865 32861 39899 32895
rect 39899 32861 39908 32895
rect 39856 32852 39908 32861
rect 40500 32895 40552 32904
rect 40500 32861 40509 32895
rect 40509 32861 40543 32895
rect 40543 32861 40552 32895
rect 40500 32852 40552 32861
rect 34060 32716 34112 32768
rect 35348 32716 35400 32768
rect 37004 32759 37056 32768
rect 37004 32725 37013 32759
rect 37013 32725 37047 32759
rect 37047 32725 37056 32759
rect 37004 32716 37056 32725
rect 37280 32716 37332 32768
rect 37556 32716 37608 32768
rect 37648 32716 37700 32768
rect 38568 32759 38620 32768
rect 38568 32725 38577 32759
rect 38577 32725 38611 32759
rect 38611 32725 38620 32759
rect 38568 32716 38620 32725
rect 39580 32716 39632 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 5724 32512 5776 32564
rect 6828 32512 6880 32564
rect 6920 32555 6972 32564
rect 6920 32521 6929 32555
rect 6929 32521 6963 32555
rect 6963 32521 6972 32555
rect 6920 32512 6972 32521
rect 7288 32512 7340 32564
rect 7656 32512 7708 32564
rect 8024 32512 8076 32564
rect 4988 32444 5040 32496
rect 6092 32444 6144 32496
rect 6000 32419 6052 32428
rect 6000 32385 6009 32419
rect 6009 32385 6043 32419
rect 6043 32385 6052 32419
rect 6000 32376 6052 32385
rect 6184 32419 6236 32428
rect 6184 32385 6193 32419
rect 6193 32385 6227 32419
rect 6227 32385 6236 32419
rect 6184 32376 6236 32385
rect 8300 32444 8352 32496
rect 5080 32351 5132 32360
rect 5080 32317 5089 32351
rect 5089 32317 5123 32351
rect 5123 32317 5132 32351
rect 5080 32308 5132 32317
rect 6276 32308 6328 32360
rect 8300 32351 8352 32360
rect 8300 32317 8309 32351
rect 8309 32317 8343 32351
rect 8343 32317 8352 32351
rect 8300 32308 8352 32317
rect 9772 32512 9824 32564
rect 11336 32512 11388 32564
rect 12072 32512 12124 32564
rect 13912 32512 13964 32564
rect 14556 32512 14608 32564
rect 14832 32512 14884 32564
rect 16028 32555 16080 32564
rect 16028 32521 16037 32555
rect 16037 32521 16071 32555
rect 16071 32521 16080 32555
rect 16028 32512 16080 32521
rect 17960 32512 18012 32564
rect 22744 32512 22796 32564
rect 24768 32512 24820 32564
rect 27068 32512 27120 32564
rect 31208 32512 31260 32564
rect 9404 32419 9456 32428
rect 9404 32385 9413 32419
rect 9413 32385 9447 32419
rect 9447 32385 9456 32419
rect 9404 32376 9456 32385
rect 10600 32376 10652 32428
rect 9864 32351 9916 32360
rect 9864 32317 9873 32351
rect 9873 32317 9907 32351
rect 9907 32317 9916 32351
rect 9864 32308 9916 32317
rect 11888 32376 11940 32428
rect 12348 32308 12400 32360
rect 14004 32419 14056 32428
rect 14004 32385 14013 32419
rect 14013 32385 14047 32419
rect 14047 32385 14056 32419
rect 14004 32376 14056 32385
rect 15568 32444 15620 32496
rect 18052 32487 18104 32496
rect 18052 32453 18061 32487
rect 18061 32453 18095 32487
rect 18095 32453 18104 32487
rect 18052 32444 18104 32453
rect 21824 32444 21876 32496
rect 22284 32444 22336 32496
rect 22468 32444 22520 32496
rect 22836 32444 22888 32496
rect 24216 32487 24268 32496
rect 24216 32453 24225 32487
rect 24225 32453 24259 32487
rect 24259 32453 24268 32487
rect 24216 32444 24268 32453
rect 14280 32351 14332 32360
rect 14280 32317 14289 32351
rect 14289 32317 14323 32351
rect 14323 32317 14332 32351
rect 14280 32308 14332 32317
rect 4896 32215 4948 32224
rect 4896 32181 4905 32215
rect 4905 32181 4939 32215
rect 4939 32181 4948 32215
rect 4896 32172 4948 32181
rect 5908 32172 5960 32224
rect 6644 32172 6696 32224
rect 6828 32172 6880 32224
rect 7748 32215 7800 32224
rect 7748 32181 7757 32215
rect 7757 32181 7791 32215
rect 7791 32181 7800 32215
rect 7748 32172 7800 32181
rect 8208 32172 8260 32224
rect 12532 32240 12584 32292
rect 16212 32308 16264 32360
rect 21180 32376 21232 32428
rect 21640 32376 21692 32428
rect 24860 32444 24912 32496
rect 28264 32444 28316 32496
rect 28632 32444 28684 32496
rect 30656 32444 30708 32496
rect 19156 32308 19208 32360
rect 25412 32376 25464 32428
rect 16304 32240 16356 32292
rect 21364 32240 21416 32292
rect 22652 32308 22704 32360
rect 24400 32351 24452 32360
rect 24400 32317 24409 32351
rect 24409 32317 24443 32351
rect 24443 32317 24452 32351
rect 24400 32308 24452 32317
rect 26700 32419 26752 32428
rect 26700 32385 26709 32419
rect 26709 32385 26743 32419
rect 26743 32385 26752 32419
rect 26700 32376 26752 32385
rect 26608 32308 26660 32360
rect 27528 32419 27580 32428
rect 27528 32385 27537 32419
rect 27537 32385 27571 32419
rect 27571 32385 27580 32419
rect 27528 32376 27580 32385
rect 27620 32376 27672 32428
rect 27988 32308 28040 32360
rect 28816 32376 28868 32428
rect 29000 32419 29052 32428
rect 29000 32385 29029 32419
rect 29029 32385 29052 32419
rect 29000 32376 29052 32385
rect 29276 32419 29328 32428
rect 29276 32385 29285 32419
rect 29285 32385 29319 32419
rect 29319 32385 29328 32419
rect 29276 32376 29328 32385
rect 29460 32376 29512 32428
rect 29644 32376 29696 32428
rect 30288 32376 30340 32428
rect 30380 32419 30432 32428
rect 30380 32385 30389 32419
rect 30389 32385 30423 32419
rect 30423 32385 30432 32419
rect 30380 32376 30432 32385
rect 29920 32308 29972 32360
rect 32588 32555 32640 32564
rect 32588 32521 32597 32555
rect 32597 32521 32631 32555
rect 32631 32521 32640 32555
rect 32588 32512 32640 32521
rect 32864 32555 32916 32564
rect 32864 32521 32873 32555
rect 32873 32521 32907 32555
rect 32907 32521 32916 32555
rect 32864 32512 32916 32521
rect 33876 32512 33928 32564
rect 34796 32512 34848 32564
rect 35992 32512 36044 32564
rect 37096 32512 37148 32564
rect 38016 32512 38068 32564
rect 38660 32512 38712 32564
rect 40500 32512 40552 32564
rect 40960 32555 41012 32564
rect 40960 32521 40969 32555
rect 40969 32521 41003 32555
rect 41003 32521 41012 32555
rect 40960 32512 41012 32521
rect 32220 32351 32272 32360
rect 32220 32317 32229 32351
rect 32229 32317 32263 32351
rect 32263 32317 32272 32351
rect 32220 32308 32272 32317
rect 23756 32240 23808 32292
rect 24216 32240 24268 32292
rect 24768 32240 24820 32292
rect 8576 32215 8628 32224
rect 8576 32181 8585 32215
rect 8585 32181 8619 32215
rect 8619 32181 8628 32215
rect 8576 32172 8628 32181
rect 9680 32215 9732 32224
rect 9680 32181 9689 32215
rect 9689 32181 9723 32215
rect 9723 32181 9732 32215
rect 9680 32172 9732 32181
rect 12440 32172 12492 32224
rect 14188 32215 14240 32224
rect 14188 32181 14197 32215
rect 14197 32181 14231 32215
rect 14231 32181 14240 32215
rect 14188 32172 14240 32181
rect 15200 32172 15252 32224
rect 15936 32172 15988 32224
rect 16488 32172 16540 32224
rect 21456 32172 21508 32224
rect 24308 32172 24360 32224
rect 24676 32172 24728 32224
rect 25320 32172 25372 32224
rect 26332 32283 26384 32292
rect 26332 32249 26341 32283
rect 26341 32249 26375 32283
rect 26375 32249 26384 32283
rect 26332 32240 26384 32249
rect 27896 32240 27948 32292
rect 32680 32419 32732 32428
rect 32680 32385 32689 32419
rect 32689 32385 32723 32419
rect 32723 32385 32732 32419
rect 32680 32376 32732 32385
rect 33048 32376 33100 32428
rect 34244 32308 34296 32360
rect 34428 32444 34480 32496
rect 36268 32376 36320 32428
rect 36452 32376 36504 32428
rect 37832 32444 37884 32496
rect 37464 32376 37516 32428
rect 37280 32308 37332 32360
rect 38016 32376 38068 32428
rect 38384 32376 38436 32428
rect 38476 32376 38528 32428
rect 39212 32444 39264 32496
rect 40592 32376 40644 32428
rect 40776 32419 40828 32428
rect 40776 32385 40785 32419
rect 40785 32385 40819 32419
rect 40819 32385 40828 32419
rect 40776 32376 40828 32385
rect 27068 32172 27120 32224
rect 27160 32172 27212 32224
rect 27344 32215 27396 32224
rect 27344 32181 27353 32215
rect 27353 32181 27387 32215
rect 27387 32181 27396 32215
rect 27344 32172 27396 32181
rect 27528 32172 27580 32224
rect 29000 32172 29052 32224
rect 29644 32172 29696 32224
rect 30196 32215 30248 32224
rect 30196 32181 30205 32215
rect 30205 32181 30239 32215
rect 30239 32181 30248 32215
rect 30196 32172 30248 32181
rect 30748 32172 30800 32224
rect 32036 32172 32088 32224
rect 39580 32308 39632 32360
rect 38108 32240 38160 32292
rect 33140 32172 33192 32224
rect 33324 32172 33376 32224
rect 34612 32172 34664 32224
rect 37556 32172 37608 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 4804 31968 4856 32020
rect 4896 31968 4948 32020
rect 6000 31968 6052 32020
rect 6092 31968 6144 32020
rect 5908 31943 5960 31952
rect 5908 31909 5917 31943
rect 5917 31909 5951 31943
rect 5951 31909 5960 31943
rect 5908 31900 5960 31909
rect 5356 31875 5408 31884
rect 5356 31841 5365 31875
rect 5365 31841 5399 31875
rect 5399 31841 5408 31875
rect 5356 31832 5408 31841
rect 2964 31807 3016 31816
rect 2964 31773 2973 31807
rect 2973 31773 3007 31807
rect 3007 31773 3016 31807
rect 2964 31764 3016 31773
rect 4988 31764 5040 31816
rect 5724 31764 5776 31816
rect 6000 31764 6052 31816
rect 7196 31968 7248 32020
rect 7932 31968 7984 32020
rect 6644 31832 6696 31884
rect 6184 31807 6236 31816
rect 6184 31773 6193 31807
rect 6193 31773 6227 31807
rect 6227 31773 6236 31807
rect 6184 31764 6236 31773
rect 6920 31764 6972 31816
rect 7104 31807 7156 31816
rect 7104 31773 7114 31807
rect 7114 31773 7148 31807
rect 7148 31773 7156 31807
rect 7748 31832 7800 31884
rect 9680 31832 9732 31884
rect 12624 32011 12676 32020
rect 12624 31977 12633 32011
rect 12633 31977 12667 32011
rect 12667 31977 12676 32011
rect 12624 31968 12676 31977
rect 13084 31968 13136 32020
rect 14924 31968 14976 32020
rect 15200 32011 15252 32020
rect 15200 31977 15209 32011
rect 15209 31977 15243 32011
rect 15243 31977 15252 32011
rect 15200 31968 15252 31977
rect 15660 31968 15712 32020
rect 7104 31764 7156 31773
rect 2780 31671 2832 31680
rect 2780 31637 2789 31671
rect 2789 31637 2823 31671
rect 2823 31637 2832 31671
rect 2780 31628 2832 31637
rect 8208 31764 8260 31816
rect 11612 31832 11664 31884
rect 14556 31832 14608 31884
rect 14924 31875 14976 31884
rect 14924 31841 14932 31875
rect 14932 31841 14966 31875
rect 14966 31841 14976 31875
rect 14924 31832 14976 31841
rect 17408 31900 17460 31952
rect 12440 31807 12492 31816
rect 12440 31773 12449 31807
rect 12449 31773 12483 31807
rect 12483 31773 12492 31807
rect 12440 31764 12492 31773
rect 12532 31807 12584 31816
rect 12532 31773 12541 31807
rect 12541 31773 12575 31807
rect 12575 31773 12584 31807
rect 12532 31764 12584 31773
rect 14188 31764 14240 31816
rect 14648 31807 14700 31816
rect 14648 31773 14657 31807
rect 14657 31773 14691 31807
rect 14691 31773 14700 31807
rect 14648 31764 14700 31773
rect 7656 31671 7708 31680
rect 7656 31637 7665 31671
rect 7665 31637 7699 31671
rect 7699 31637 7708 31671
rect 7656 31628 7708 31637
rect 8944 31628 8996 31680
rect 9404 31628 9456 31680
rect 12440 31628 12492 31680
rect 14464 31671 14516 31680
rect 14464 31637 14473 31671
rect 14473 31637 14507 31671
rect 14507 31637 14516 31671
rect 14464 31628 14516 31637
rect 14648 31628 14700 31680
rect 15568 31764 15620 31816
rect 15752 31807 15804 31816
rect 15752 31773 15761 31807
rect 15761 31773 15795 31807
rect 15795 31773 15804 31807
rect 15752 31764 15804 31773
rect 16304 31764 16356 31816
rect 22192 31968 22244 32020
rect 23664 32011 23716 32020
rect 23664 31977 23673 32011
rect 23673 31977 23707 32011
rect 23707 31977 23716 32011
rect 23664 31968 23716 31977
rect 24124 31968 24176 32020
rect 24216 31968 24268 32020
rect 25320 32011 25372 32020
rect 25320 31977 25329 32011
rect 25329 31977 25363 32011
rect 25363 31977 25372 32011
rect 25320 31968 25372 31977
rect 25872 31968 25924 32020
rect 26608 31968 26660 32020
rect 27252 32011 27304 32020
rect 27252 31977 27261 32011
rect 27261 31977 27295 32011
rect 27295 31977 27304 32011
rect 27252 31968 27304 31977
rect 27344 31968 27396 32020
rect 27896 32011 27948 32020
rect 27896 31977 27905 32011
rect 27905 31977 27939 32011
rect 27939 31977 27948 32011
rect 27896 31968 27948 31977
rect 27988 31968 28040 32020
rect 33324 31968 33376 32020
rect 34612 31968 34664 32020
rect 35348 31968 35400 32020
rect 19340 31900 19392 31952
rect 25964 31900 26016 31952
rect 26332 31900 26384 31952
rect 18696 31875 18748 31884
rect 18696 31841 18705 31875
rect 18705 31841 18739 31875
rect 18739 31841 18748 31875
rect 18696 31832 18748 31841
rect 15660 31739 15712 31748
rect 15660 31705 15669 31739
rect 15669 31705 15703 31739
rect 15703 31705 15712 31739
rect 15660 31696 15712 31705
rect 16212 31696 16264 31748
rect 16120 31628 16172 31680
rect 19340 31764 19392 31816
rect 20904 31764 20956 31816
rect 21456 31807 21508 31816
rect 21456 31773 21465 31807
rect 21465 31773 21499 31807
rect 21499 31773 21508 31807
rect 21456 31764 21508 31773
rect 21548 31807 21600 31816
rect 21548 31773 21558 31807
rect 21558 31773 21592 31807
rect 21592 31773 21600 31807
rect 21548 31764 21600 31773
rect 20168 31696 20220 31748
rect 20352 31696 20404 31748
rect 22376 31696 22428 31748
rect 22836 31764 22888 31816
rect 23480 31764 23532 31816
rect 24492 31875 24544 31884
rect 24492 31841 24501 31875
rect 24501 31841 24535 31875
rect 24535 31841 24544 31875
rect 24492 31832 24544 31841
rect 23296 31696 23348 31748
rect 24860 31832 24912 31884
rect 25320 31832 25372 31884
rect 25872 31832 25924 31884
rect 26884 31900 26936 31952
rect 26976 31900 27028 31952
rect 24768 31764 24820 31816
rect 26424 31764 26476 31816
rect 26700 31764 26752 31816
rect 24952 31739 25004 31748
rect 24952 31705 24961 31739
rect 24961 31705 24995 31739
rect 24995 31705 25004 31739
rect 24952 31696 25004 31705
rect 16856 31628 16908 31680
rect 21088 31628 21140 31680
rect 21732 31628 21784 31680
rect 22100 31671 22152 31680
rect 22100 31637 22109 31671
rect 22109 31637 22143 31671
rect 22143 31637 22152 31671
rect 22100 31628 22152 31637
rect 23572 31628 23624 31680
rect 24860 31671 24912 31680
rect 24860 31637 24869 31671
rect 24869 31637 24903 31671
rect 24903 31637 24912 31671
rect 24860 31628 24912 31637
rect 26332 31739 26384 31748
rect 26332 31705 26341 31739
rect 26341 31705 26375 31739
rect 26375 31705 26384 31739
rect 26332 31696 26384 31705
rect 26424 31628 26476 31680
rect 27252 31807 27304 31816
rect 27252 31773 27261 31807
rect 27261 31773 27295 31807
rect 27295 31773 27304 31807
rect 27252 31764 27304 31773
rect 27528 31764 27580 31816
rect 27160 31696 27212 31748
rect 28080 31764 28132 31816
rect 28908 31900 28960 31952
rect 29092 31900 29144 31952
rect 30012 31900 30064 31952
rect 28172 31696 28224 31748
rect 29000 31807 29052 31816
rect 29000 31773 29009 31807
rect 29009 31773 29043 31807
rect 29043 31773 29052 31807
rect 29000 31764 29052 31773
rect 29644 31832 29696 31884
rect 30288 31832 30340 31884
rect 30380 31764 30432 31816
rect 29092 31696 29144 31748
rect 29552 31739 29604 31748
rect 29552 31705 29561 31739
rect 29561 31705 29595 31739
rect 29595 31705 29604 31739
rect 29552 31696 29604 31705
rect 30564 31696 30616 31748
rect 31760 31832 31812 31884
rect 34428 31900 34480 31952
rect 33600 31832 33652 31884
rect 36636 32011 36688 32020
rect 36636 31977 36645 32011
rect 36645 31977 36679 32011
rect 36679 31977 36688 32011
rect 36636 31968 36688 31977
rect 36728 31968 36780 32020
rect 37096 31968 37148 32020
rect 37464 31968 37516 32020
rect 31208 31764 31260 31816
rect 31484 31764 31536 31816
rect 32128 31764 32180 31816
rect 32404 31764 32456 31816
rect 33232 31764 33284 31816
rect 33968 31807 34020 31816
rect 33968 31773 33977 31807
rect 33977 31773 34011 31807
rect 34011 31773 34020 31807
rect 33968 31764 34020 31773
rect 34244 31764 34296 31816
rect 32680 31696 32732 31748
rect 34612 31764 34664 31816
rect 35716 31832 35768 31884
rect 34888 31807 34940 31816
rect 34888 31773 34897 31807
rect 34897 31773 34931 31807
rect 34931 31773 34940 31807
rect 34888 31764 34940 31773
rect 35348 31764 35400 31816
rect 36820 31832 36872 31884
rect 37004 31832 37056 31884
rect 26976 31628 27028 31680
rect 27896 31628 27948 31680
rect 29460 31628 29512 31680
rect 31484 31628 31536 31680
rect 32496 31628 32548 31680
rect 33508 31628 33560 31680
rect 33784 31671 33836 31680
rect 33784 31637 33793 31671
rect 33793 31637 33827 31671
rect 33827 31637 33836 31671
rect 33784 31628 33836 31637
rect 33876 31628 33928 31680
rect 34980 31696 35032 31748
rect 37280 31696 37332 31748
rect 37556 31807 37608 31816
rect 37556 31773 37565 31807
rect 37565 31773 37599 31807
rect 37599 31773 37608 31807
rect 37556 31764 37608 31773
rect 37648 31807 37700 31816
rect 37648 31773 37657 31807
rect 37657 31773 37691 31807
rect 37691 31773 37700 31807
rect 37648 31764 37700 31773
rect 38568 31900 38620 31952
rect 38200 31739 38252 31748
rect 38200 31705 38209 31739
rect 38209 31705 38243 31739
rect 38243 31705 38252 31739
rect 38200 31696 38252 31705
rect 41604 31764 41656 31816
rect 34520 31628 34572 31680
rect 35348 31628 35400 31680
rect 35716 31628 35768 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 2044 31331 2096 31340
rect 2044 31297 2053 31331
rect 2053 31297 2087 31331
rect 2087 31297 2096 31331
rect 2044 31288 2096 31297
rect 2780 31356 2832 31408
rect 3056 31356 3108 31408
rect 4896 31331 4948 31340
rect 4896 31297 4905 31331
rect 4905 31297 4939 31331
rect 4939 31297 4948 31331
rect 4896 31288 4948 31297
rect 4988 31331 5040 31340
rect 4988 31297 4997 31331
rect 4997 31297 5031 31331
rect 5031 31297 5040 31331
rect 4988 31288 5040 31297
rect 8944 31424 8996 31476
rect 10048 31424 10100 31476
rect 14372 31424 14424 31476
rect 7196 31356 7248 31408
rect 9496 31288 9548 31340
rect 15108 31356 15160 31408
rect 15476 31424 15528 31476
rect 16212 31467 16264 31476
rect 16212 31433 16221 31467
rect 16221 31433 16255 31467
rect 16255 31433 16264 31467
rect 16212 31424 16264 31433
rect 16304 31424 16356 31476
rect 14280 31288 14332 31340
rect 15200 31288 15252 31340
rect 15936 31356 15988 31408
rect 16948 31356 17000 31408
rect 17500 31356 17552 31408
rect 20996 31424 21048 31476
rect 21088 31424 21140 31476
rect 22192 31424 22244 31476
rect 16120 31288 16172 31340
rect 16488 31288 16540 31340
rect 22560 31424 22612 31476
rect 22928 31424 22980 31476
rect 23756 31424 23808 31476
rect 24032 31424 24084 31476
rect 24124 31424 24176 31476
rect 24952 31424 25004 31476
rect 27252 31424 27304 31476
rect 27344 31424 27396 31476
rect 24676 31356 24728 31408
rect 27804 31356 27856 31408
rect 29000 31424 29052 31476
rect 29368 31424 29420 31476
rect 29736 31467 29788 31476
rect 29736 31433 29745 31467
rect 29745 31433 29779 31467
rect 29779 31433 29788 31467
rect 29736 31424 29788 31433
rect 30932 31424 30984 31476
rect 31024 31424 31076 31476
rect 3700 31220 3752 31272
rect 7656 31220 7708 31272
rect 8576 31220 8628 31272
rect 9864 31220 9916 31272
rect 11796 31263 11848 31272
rect 11796 31229 11805 31263
rect 11805 31229 11839 31263
rect 11839 31229 11848 31263
rect 11796 31220 11848 31229
rect 13544 31263 13596 31272
rect 13544 31229 13553 31263
rect 13553 31229 13587 31263
rect 13587 31229 13596 31263
rect 13544 31220 13596 31229
rect 14188 31220 14240 31272
rect 14464 31263 14516 31272
rect 14464 31229 14473 31263
rect 14473 31229 14507 31263
rect 14507 31229 14516 31263
rect 14464 31220 14516 31229
rect 14740 31220 14792 31272
rect 6184 31152 6236 31204
rect 1768 31084 1820 31136
rect 5080 31127 5132 31136
rect 5080 31093 5089 31127
rect 5089 31093 5123 31127
rect 5123 31093 5132 31127
rect 5080 31084 5132 31093
rect 6736 31084 6788 31136
rect 7288 31084 7340 31136
rect 7932 31084 7984 31136
rect 8392 31127 8444 31136
rect 8392 31093 8401 31127
rect 8401 31093 8435 31127
rect 8435 31093 8444 31127
rect 8392 31084 8444 31093
rect 16580 31152 16632 31204
rect 16396 31127 16448 31136
rect 16396 31093 16405 31127
rect 16405 31093 16439 31127
rect 16439 31093 16448 31127
rect 16396 31084 16448 31093
rect 17224 31263 17276 31272
rect 17224 31229 17233 31263
rect 17233 31229 17267 31263
rect 17267 31229 17276 31263
rect 17224 31220 17276 31229
rect 18696 31220 18748 31272
rect 19064 31263 19116 31272
rect 19064 31229 19073 31263
rect 19073 31229 19107 31263
rect 19107 31229 19116 31263
rect 19064 31220 19116 31229
rect 19248 31084 19300 31136
rect 20444 31084 20496 31136
rect 22008 31220 22060 31272
rect 22192 31220 22244 31272
rect 20628 31084 20680 31136
rect 21272 31127 21324 31136
rect 21272 31093 21281 31127
rect 21281 31093 21315 31127
rect 21315 31093 21324 31127
rect 21272 31084 21324 31093
rect 21732 31084 21784 31136
rect 22100 31084 22152 31136
rect 22192 31127 22244 31136
rect 22192 31093 22201 31127
rect 22201 31093 22235 31127
rect 22235 31093 22244 31127
rect 22192 31084 22244 31093
rect 22284 31127 22336 31136
rect 22284 31093 22293 31127
rect 22293 31093 22327 31127
rect 22327 31093 22336 31127
rect 22284 31084 22336 31093
rect 22928 31288 22980 31340
rect 23572 31288 23624 31340
rect 23848 31331 23900 31340
rect 23848 31297 23855 31331
rect 23855 31297 23900 31331
rect 23848 31288 23900 31297
rect 24129 31331 24181 31340
rect 24129 31297 24138 31331
rect 24138 31297 24172 31331
rect 24172 31297 24181 31331
rect 24129 31288 24181 31297
rect 23940 31220 23992 31272
rect 24308 31220 24360 31272
rect 24584 31331 24636 31340
rect 24584 31297 24593 31331
rect 24593 31297 24627 31331
rect 24627 31297 24636 31331
rect 24584 31288 24636 31297
rect 25228 31288 25280 31340
rect 24768 31220 24820 31272
rect 25412 31152 25464 31204
rect 25780 31331 25832 31340
rect 25780 31297 25789 31331
rect 25789 31297 25823 31331
rect 25823 31297 25832 31331
rect 25780 31288 25832 31297
rect 25872 31331 25924 31340
rect 25872 31297 25881 31331
rect 25881 31297 25915 31331
rect 25915 31297 25924 31331
rect 25872 31288 25924 31297
rect 26516 31288 26568 31340
rect 27896 31288 27948 31340
rect 29092 31288 29144 31340
rect 28540 31220 28592 31272
rect 29552 31263 29604 31272
rect 29552 31229 29561 31263
rect 29561 31229 29595 31263
rect 29595 31229 29604 31263
rect 29552 31220 29604 31229
rect 31392 31288 31444 31340
rect 31484 31331 31536 31340
rect 31484 31297 31493 31331
rect 31493 31297 31527 31331
rect 31527 31297 31536 31331
rect 31484 31288 31536 31297
rect 31760 31288 31812 31340
rect 32404 31288 32456 31340
rect 32496 31288 32548 31340
rect 33508 31424 33560 31476
rect 33876 31424 33928 31476
rect 34888 31424 34940 31476
rect 35808 31424 35860 31476
rect 36912 31424 36964 31476
rect 41052 31424 41104 31476
rect 33784 31356 33836 31408
rect 34704 31356 34756 31408
rect 35532 31356 35584 31408
rect 25964 31152 26016 31204
rect 26332 31152 26384 31204
rect 26424 31152 26476 31204
rect 27528 31152 27580 31204
rect 30932 31220 30984 31272
rect 33416 31331 33468 31340
rect 33416 31297 33425 31331
rect 33425 31297 33459 31331
rect 33459 31297 33468 31331
rect 33416 31288 33468 31297
rect 34060 31288 34112 31340
rect 34980 31288 35032 31340
rect 38016 31331 38068 31340
rect 38016 31297 38025 31331
rect 38025 31297 38059 31331
rect 38059 31297 38068 31331
rect 38016 31288 38068 31297
rect 40040 31356 40092 31408
rect 38568 31288 38620 31340
rect 38936 31288 38988 31340
rect 33600 31220 33652 31272
rect 33968 31220 34020 31272
rect 34244 31263 34296 31272
rect 34244 31229 34253 31263
rect 34253 31229 34287 31263
rect 34287 31229 34296 31263
rect 34244 31220 34296 31229
rect 34336 31263 34388 31272
rect 34336 31229 34345 31263
rect 34345 31229 34379 31263
rect 34379 31229 34388 31263
rect 34336 31220 34388 31229
rect 34428 31263 34480 31272
rect 34428 31229 34437 31263
rect 34437 31229 34471 31263
rect 34471 31229 34480 31263
rect 34428 31220 34480 31229
rect 25688 31084 25740 31136
rect 25780 31084 25832 31136
rect 26792 31084 26844 31136
rect 27252 31127 27304 31136
rect 27252 31093 27261 31127
rect 27261 31093 27295 31127
rect 27295 31093 27304 31127
rect 27252 31084 27304 31093
rect 28264 31084 28316 31136
rect 28540 31084 28592 31136
rect 29276 31084 29328 31136
rect 29460 31127 29512 31136
rect 29460 31093 29469 31127
rect 29469 31093 29503 31127
rect 29503 31093 29512 31127
rect 29460 31084 29512 31093
rect 30104 31127 30156 31136
rect 30104 31093 30113 31127
rect 30113 31093 30147 31127
rect 30147 31093 30156 31127
rect 30104 31084 30156 31093
rect 31484 31084 31536 31136
rect 32128 31127 32180 31136
rect 32128 31093 32137 31127
rect 32137 31093 32171 31127
rect 32171 31093 32180 31127
rect 32128 31084 32180 31093
rect 32680 31127 32732 31136
rect 32680 31093 32689 31127
rect 32689 31093 32723 31127
rect 32723 31093 32732 31127
rect 32680 31084 32732 31093
rect 34796 31220 34848 31272
rect 38200 31220 38252 31272
rect 39028 31220 39080 31272
rect 39580 31263 39632 31272
rect 39580 31229 39589 31263
rect 39589 31229 39623 31263
rect 39623 31229 39632 31263
rect 39580 31220 39632 31229
rect 33600 31084 33652 31136
rect 37280 31084 37332 31136
rect 38384 31084 38436 31136
rect 38660 31127 38712 31136
rect 38660 31093 38669 31127
rect 38669 31093 38703 31127
rect 38703 31093 38712 31127
rect 38660 31084 38712 31093
rect 38752 31084 38804 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 2964 30880 3016 30932
rect 11796 30880 11848 30932
rect 13544 30880 13596 30932
rect 15108 30880 15160 30932
rect 17224 30880 17276 30932
rect 19064 30880 19116 30932
rect 21272 30880 21324 30932
rect 21824 30880 21876 30932
rect 22284 30880 22336 30932
rect 22836 30880 22888 30932
rect 23112 30880 23164 30932
rect 24216 30880 24268 30932
rect 24400 30923 24452 30932
rect 24400 30889 24409 30923
rect 24409 30889 24443 30923
rect 24443 30889 24452 30923
rect 24400 30880 24452 30889
rect 11612 30812 11664 30864
rect 12348 30855 12400 30864
rect 12348 30821 12357 30855
rect 12357 30821 12391 30855
rect 12391 30821 12400 30855
rect 12348 30812 12400 30821
rect 1768 30744 1820 30796
rect 3424 30744 3476 30796
rect 5080 30744 5132 30796
rect 1400 30719 1452 30728
rect 1400 30685 1409 30719
rect 1409 30685 1443 30719
rect 1443 30685 1452 30719
rect 1400 30676 1452 30685
rect 3056 30676 3108 30728
rect 2964 30608 3016 30660
rect 4068 30608 4120 30660
rect 3700 30540 3752 30592
rect 10232 30608 10284 30660
rect 10876 30676 10928 30728
rect 12072 30676 12124 30728
rect 12440 30676 12492 30728
rect 12532 30719 12584 30728
rect 12532 30685 12541 30719
rect 12541 30685 12575 30719
rect 12575 30685 12584 30719
rect 12532 30676 12584 30685
rect 11152 30608 11204 30660
rect 11428 30651 11480 30660
rect 11428 30617 11437 30651
rect 11437 30617 11471 30651
rect 11471 30617 11480 30651
rect 11428 30608 11480 30617
rect 11520 30651 11572 30660
rect 11520 30617 11529 30651
rect 11529 30617 11563 30651
rect 11563 30617 11572 30651
rect 11520 30608 11572 30617
rect 17132 30812 17184 30864
rect 17500 30812 17552 30864
rect 14648 30744 14700 30796
rect 16396 30744 16448 30796
rect 16580 30744 16632 30796
rect 17592 30744 17644 30796
rect 19156 30812 19208 30864
rect 17960 30676 18012 30728
rect 19340 30676 19392 30728
rect 18052 30608 18104 30660
rect 18144 30608 18196 30660
rect 18236 30651 18288 30660
rect 18236 30617 18245 30651
rect 18245 30617 18279 30651
rect 18279 30617 18288 30651
rect 18236 30608 18288 30617
rect 11980 30540 12032 30592
rect 12716 30540 12768 30592
rect 16856 30540 16908 30592
rect 18604 30583 18656 30592
rect 18604 30549 18613 30583
rect 18613 30549 18647 30583
rect 18647 30549 18656 30583
rect 18604 30540 18656 30549
rect 18696 30583 18748 30592
rect 18696 30549 18705 30583
rect 18705 30549 18739 30583
rect 18739 30549 18748 30583
rect 18696 30540 18748 30549
rect 19064 30540 19116 30592
rect 20444 30676 20496 30728
rect 21180 30719 21232 30728
rect 21180 30685 21189 30719
rect 21189 30685 21223 30719
rect 21223 30685 21232 30719
rect 22008 30812 22060 30864
rect 24492 30812 24544 30864
rect 24952 30855 25004 30864
rect 24952 30821 24961 30855
rect 24961 30821 24995 30855
rect 24995 30821 25004 30855
rect 24952 30812 25004 30821
rect 21180 30676 21232 30685
rect 20536 30608 20588 30660
rect 21640 30719 21692 30728
rect 21640 30685 21650 30719
rect 21650 30685 21684 30719
rect 21684 30685 21692 30719
rect 26424 30880 26476 30932
rect 26700 30880 26752 30932
rect 21640 30676 21692 30685
rect 22008 30676 22060 30728
rect 22836 30676 22888 30728
rect 23756 30676 23808 30728
rect 24676 30719 24728 30728
rect 24676 30685 24685 30719
rect 24685 30685 24719 30719
rect 24719 30685 24728 30719
rect 24676 30676 24728 30685
rect 25044 30676 25096 30728
rect 26608 30744 26660 30796
rect 29736 30880 29788 30932
rect 32588 30880 32640 30932
rect 32680 30880 32732 30932
rect 31024 30812 31076 30864
rect 31208 30812 31260 30864
rect 31668 30812 31720 30864
rect 28448 30744 28500 30796
rect 28816 30744 28868 30796
rect 30472 30744 30524 30796
rect 33140 30812 33192 30864
rect 23020 30608 23072 30660
rect 25780 30651 25832 30660
rect 25780 30617 25789 30651
rect 25789 30617 25823 30651
rect 25823 30617 25832 30651
rect 25780 30608 25832 30617
rect 25964 30651 26016 30660
rect 25964 30617 25973 30651
rect 25973 30617 26007 30651
rect 26007 30617 26016 30651
rect 25964 30608 26016 30617
rect 26332 30608 26384 30660
rect 26792 30676 26844 30728
rect 27068 30676 27120 30728
rect 27528 30676 27580 30728
rect 28908 30719 28960 30728
rect 28908 30685 28917 30719
rect 28917 30685 28951 30719
rect 28951 30685 28960 30719
rect 28908 30676 28960 30685
rect 29828 30676 29880 30728
rect 31208 30719 31260 30728
rect 31208 30685 31217 30719
rect 31217 30685 31251 30719
rect 31251 30685 31260 30719
rect 31208 30676 31260 30685
rect 31484 30719 31536 30728
rect 31484 30685 31493 30719
rect 31493 30685 31527 30719
rect 31527 30685 31536 30719
rect 31484 30676 31536 30685
rect 32128 30719 32180 30728
rect 32128 30685 32137 30719
rect 32137 30685 32171 30719
rect 32171 30685 32180 30719
rect 32128 30676 32180 30685
rect 32680 30744 32732 30796
rect 34796 30744 34848 30796
rect 36728 30787 36780 30796
rect 36728 30753 36737 30787
rect 36737 30753 36771 30787
rect 36771 30753 36780 30787
rect 36728 30744 36780 30753
rect 34060 30676 34112 30728
rect 35532 30676 35584 30728
rect 35716 30719 35768 30728
rect 35716 30685 35725 30719
rect 35725 30685 35759 30719
rect 35759 30685 35768 30719
rect 35716 30676 35768 30685
rect 37556 30880 37608 30932
rect 38200 30923 38252 30932
rect 38200 30889 38209 30923
rect 38209 30889 38243 30923
rect 38243 30889 38252 30923
rect 38200 30880 38252 30889
rect 38752 30923 38804 30932
rect 37648 30812 37700 30864
rect 37280 30787 37332 30796
rect 37280 30753 37289 30787
rect 37289 30753 37323 30787
rect 37323 30753 37332 30787
rect 37280 30744 37332 30753
rect 38752 30889 38761 30923
rect 38761 30889 38795 30923
rect 38795 30889 38804 30923
rect 38752 30880 38804 30889
rect 39580 30880 39632 30932
rect 20904 30540 20956 30592
rect 34704 30608 34756 30660
rect 38016 30676 38068 30728
rect 38384 30676 38436 30728
rect 38568 30744 38620 30796
rect 38844 30719 38896 30728
rect 38844 30685 38853 30719
rect 38853 30685 38887 30719
rect 38887 30685 38896 30719
rect 38844 30676 38896 30685
rect 38936 30608 38988 30660
rect 23296 30540 23348 30592
rect 25596 30583 25648 30592
rect 25596 30549 25605 30583
rect 25605 30549 25639 30583
rect 25639 30549 25648 30583
rect 25596 30540 25648 30549
rect 25688 30540 25740 30592
rect 27436 30540 27488 30592
rect 32404 30583 32456 30592
rect 32404 30549 32413 30583
rect 32413 30549 32447 30583
rect 32447 30549 32456 30583
rect 32404 30540 32456 30549
rect 33416 30540 33468 30592
rect 33876 30583 33928 30592
rect 33876 30549 33885 30583
rect 33885 30549 33919 30583
rect 33919 30549 33928 30583
rect 33876 30540 33928 30549
rect 34520 30540 34572 30592
rect 36912 30540 36964 30592
rect 38476 30583 38528 30592
rect 38476 30549 38485 30583
rect 38485 30549 38519 30583
rect 38519 30549 38528 30583
rect 38476 30540 38528 30549
rect 38844 30540 38896 30592
rect 41328 30676 41380 30728
rect 39212 30583 39264 30592
rect 39212 30549 39221 30583
rect 39221 30549 39255 30583
rect 39255 30549 39264 30583
rect 39212 30540 39264 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 2044 30336 2096 30388
rect 2780 30379 2832 30388
rect 2780 30345 2789 30379
rect 2789 30345 2823 30379
rect 2823 30345 2832 30379
rect 2780 30336 2832 30345
rect 4804 30200 4856 30252
rect 7932 30200 7984 30252
rect 2872 30175 2924 30184
rect 2872 30141 2881 30175
rect 2881 30141 2915 30175
rect 2915 30141 2924 30175
rect 2872 30132 2924 30141
rect 3332 30132 3384 30184
rect 7840 30132 7892 30184
rect 8208 30200 8260 30252
rect 8944 30336 8996 30388
rect 18052 30336 18104 30388
rect 8576 30200 8628 30252
rect 9312 30243 9364 30252
rect 9312 30209 9321 30243
rect 9321 30209 9355 30243
rect 9355 30209 9364 30243
rect 9312 30200 9364 30209
rect 9496 30243 9548 30252
rect 9496 30209 9503 30243
rect 9503 30209 9548 30243
rect 9496 30200 9548 30209
rect 10876 30268 10928 30320
rect 19064 30336 19116 30388
rect 8852 30132 8904 30184
rect 9956 30200 10008 30252
rect 17960 30243 18012 30252
rect 17960 30209 17969 30243
rect 17969 30209 18003 30243
rect 18003 30209 18012 30243
rect 17960 30200 18012 30209
rect 18236 30200 18288 30252
rect 18972 30268 19024 30320
rect 19248 30336 19300 30388
rect 18788 30200 18840 30252
rect 18604 30132 18656 30184
rect 20444 30268 20496 30320
rect 22192 30336 22244 30388
rect 22744 30336 22796 30388
rect 23756 30336 23808 30388
rect 24676 30336 24728 30388
rect 26332 30336 26384 30388
rect 21180 30268 21232 30320
rect 27252 30336 27304 30388
rect 27896 30336 27948 30388
rect 30104 30379 30156 30388
rect 30104 30345 30113 30379
rect 30113 30345 30147 30379
rect 30147 30345 30156 30379
rect 30104 30336 30156 30345
rect 31852 30336 31904 30388
rect 38568 30336 38620 30388
rect 19340 30200 19392 30252
rect 4896 30064 4948 30116
rect 6552 30064 6604 30116
rect 9772 30064 9824 30116
rect 19248 30132 19300 30184
rect 20628 30132 20680 30184
rect 20444 30064 20496 30116
rect 21180 30132 21232 30184
rect 21548 30200 21600 30252
rect 25964 30200 26016 30252
rect 27528 30200 27580 30252
rect 29368 30200 29420 30252
rect 29460 30243 29512 30252
rect 29460 30209 29469 30243
rect 29469 30209 29503 30243
rect 29503 30209 29512 30243
rect 29460 30200 29512 30209
rect 29644 30243 29696 30252
rect 29644 30209 29651 30243
rect 29651 30209 29696 30243
rect 29644 30200 29696 30209
rect 21916 30132 21968 30184
rect 24308 30132 24360 30184
rect 28264 30132 28316 30184
rect 5080 29996 5132 30048
rect 6184 29996 6236 30048
rect 6460 29996 6512 30048
rect 11244 29996 11296 30048
rect 13820 29996 13872 30048
rect 13912 29996 13964 30048
rect 14832 29996 14884 30048
rect 18052 30039 18104 30048
rect 18052 30005 18061 30039
rect 18061 30005 18095 30039
rect 18095 30005 18104 30039
rect 18052 29996 18104 30005
rect 21456 30064 21508 30116
rect 20812 29996 20864 30048
rect 21824 30064 21876 30116
rect 26516 30064 26568 30116
rect 28448 30064 28500 30116
rect 31760 30200 31812 30252
rect 32496 30200 32548 30252
rect 32864 30243 32916 30252
rect 32864 30209 32873 30243
rect 32873 30209 32907 30243
rect 32907 30209 32916 30243
rect 32864 30200 32916 30209
rect 30288 30132 30340 30184
rect 31576 30132 31628 30184
rect 32588 30132 32640 30184
rect 34796 30132 34848 30184
rect 33416 30064 33468 30116
rect 34612 30064 34664 30116
rect 35900 30175 35952 30184
rect 35900 30141 35909 30175
rect 35909 30141 35943 30175
rect 35943 30141 35952 30175
rect 35900 30132 35952 30141
rect 36268 30200 36320 30252
rect 36360 30243 36412 30252
rect 36360 30209 36369 30243
rect 36369 30209 36403 30243
rect 36403 30209 36412 30243
rect 36360 30200 36412 30209
rect 36176 30064 36228 30116
rect 38476 30268 38528 30320
rect 40040 30268 40092 30320
rect 37556 30107 37608 30116
rect 37556 30073 37565 30107
rect 37565 30073 37599 30107
rect 37599 30073 37608 30107
rect 37556 30064 37608 30073
rect 38752 30200 38804 30252
rect 39028 30132 39080 30184
rect 39580 30175 39632 30184
rect 39580 30141 39589 30175
rect 39589 30141 39623 30175
rect 39623 30141 39632 30175
rect 39580 30132 39632 30141
rect 38660 30064 38712 30116
rect 38936 30064 38988 30116
rect 21640 29996 21692 30048
rect 24768 29996 24820 30048
rect 30012 29996 30064 30048
rect 32220 30039 32272 30048
rect 32220 30005 32229 30039
rect 32229 30005 32263 30039
rect 32263 30005 32272 30039
rect 32220 29996 32272 30005
rect 32772 29996 32824 30048
rect 33876 29996 33928 30048
rect 34704 29996 34756 30048
rect 35808 29996 35860 30048
rect 35992 29996 36044 30048
rect 36636 29996 36688 30048
rect 38016 30039 38068 30048
rect 38016 30005 38025 30039
rect 38025 30005 38059 30039
rect 38059 30005 38068 30039
rect 38016 29996 38068 30005
rect 38844 30039 38896 30048
rect 38844 30005 38853 30039
rect 38853 30005 38887 30039
rect 38887 30005 38896 30039
rect 38844 29996 38896 30005
rect 39120 30039 39172 30048
rect 39120 30005 39129 30039
rect 39129 30005 39163 30039
rect 39163 30005 39172 30039
rect 39120 29996 39172 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2872 29792 2924 29844
rect 5264 29792 5316 29844
rect 6736 29835 6788 29844
rect 6736 29801 6745 29835
rect 6745 29801 6779 29835
rect 6779 29801 6788 29835
rect 6736 29792 6788 29801
rect 7380 29792 7432 29844
rect 7932 29792 7984 29844
rect 8668 29792 8720 29844
rect 4988 29724 5040 29776
rect 2688 29631 2740 29640
rect 2688 29597 2697 29631
rect 2697 29597 2731 29631
rect 2731 29597 2740 29631
rect 2688 29588 2740 29597
rect 4160 29520 4212 29572
rect 4804 29563 4856 29572
rect 4804 29529 4813 29563
rect 4813 29529 4847 29563
rect 4847 29529 4856 29563
rect 4804 29520 4856 29529
rect 7012 29724 7064 29776
rect 9680 29724 9732 29776
rect 5356 29631 5408 29640
rect 5356 29597 5365 29631
rect 5365 29597 5399 29631
rect 5399 29597 5408 29631
rect 5356 29588 5408 29597
rect 2504 29495 2556 29504
rect 2504 29461 2513 29495
rect 2513 29461 2547 29495
rect 2547 29461 2556 29495
rect 2504 29452 2556 29461
rect 5448 29452 5500 29504
rect 5816 29631 5868 29640
rect 6736 29656 6788 29708
rect 5816 29597 5830 29631
rect 5830 29597 5864 29631
rect 5864 29597 5868 29631
rect 5816 29588 5868 29597
rect 6184 29631 6236 29640
rect 6184 29597 6194 29631
rect 6194 29597 6228 29631
rect 6228 29597 6236 29631
rect 6184 29588 6236 29597
rect 6460 29631 6512 29640
rect 6460 29597 6469 29631
rect 6469 29597 6503 29631
rect 6503 29597 6512 29631
rect 6460 29588 6512 29597
rect 7104 29588 7156 29640
rect 7196 29631 7248 29640
rect 7196 29597 7205 29631
rect 7205 29597 7239 29631
rect 7239 29597 7248 29631
rect 7196 29588 7248 29597
rect 7380 29631 7432 29640
rect 7380 29597 7387 29631
rect 7387 29597 7432 29631
rect 7380 29588 7432 29597
rect 7748 29588 7800 29640
rect 7932 29588 7984 29640
rect 8208 29656 8260 29708
rect 9312 29656 9364 29708
rect 13820 29835 13872 29844
rect 13820 29801 13829 29835
rect 13829 29801 13863 29835
rect 13863 29801 13872 29835
rect 13820 29792 13872 29801
rect 14372 29792 14424 29844
rect 15016 29792 15068 29844
rect 18512 29792 18564 29844
rect 22192 29792 22244 29844
rect 22468 29835 22520 29844
rect 22468 29801 22477 29835
rect 22477 29801 22511 29835
rect 22511 29801 22520 29835
rect 22468 29792 22520 29801
rect 24400 29792 24452 29844
rect 24584 29792 24636 29844
rect 26056 29792 26108 29844
rect 26516 29835 26568 29844
rect 26516 29801 26525 29835
rect 26525 29801 26559 29835
rect 26559 29801 26568 29835
rect 26516 29792 26568 29801
rect 27620 29792 27672 29844
rect 8116 29631 8168 29640
rect 8116 29597 8126 29631
rect 8126 29597 8160 29631
rect 8160 29597 8168 29631
rect 8116 29588 8168 29597
rect 8576 29588 8628 29640
rect 5632 29563 5684 29572
rect 5632 29529 5641 29563
rect 5641 29529 5675 29563
rect 5675 29529 5684 29563
rect 5632 29520 5684 29529
rect 7012 29520 7064 29572
rect 8208 29520 8260 29572
rect 9220 29520 9272 29572
rect 6552 29452 6604 29504
rect 7840 29452 7892 29504
rect 9404 29588 9456 29640
rect 11520 29656 11572 29708
rect 12808 29724 12860 29776
rect 16396 29724 16448 29776
rect 21640 29724 21692 29776
rect 9588 29631 9640 29640
rect 9588 29597 9598 29631
rect 9598 29597 9632 29631
rect 9632 29597 9640 29631
rect 9588 29588 9640 29597
rect 9956 29588 10008 29640
rect 11980 29588 12032 29640
rect 12256 29631 12308 29640
rect 12256 29597 12265 29631
rect 12265 29597 12299 29631
rect 12299 29597 12308 29631
rect 12256 29588 12308 29597
rect 13176 29631 13228 29640
rect 13176 29597 13185 29631
rect 13185 29597 13219 29631
rect 13219 29597 13228 29631
rect 13176 29588 13228 29597
rect 13268 29631 13320 29640
rect 13268 29597 13278 29631
rect 13278 29597 13312 29631
rect 13312 29597 13320 29631
rect 13268 29588 13320 29597
rect 9772 29563 9824 29572
rect 9772 29529 9781 29563
rect 9781 29529 9815 29563
rect 9815 29529 9824 29563
rect 9772 29520 9824 29529
rect 9864 29563 9916 29572
rect 9864 29529 9873 29563
rect 9873 29529 9907 29563
rect 9907 29529 9916 29563
rect 9864 29520 9916 29529
rect 11704 29520 11756 29572
rect 11888 29520 11940 29572
rect 13360 29520 13412 29572
rect 13912 29588 13964 29640
rect 14096 29631 14148 29640
rect 14096 29597 14105 29631
rect 14105 29597 14139 29631
rect 14139 29597 14148 29631
rect 14096 29588 14148 29597
rect 14372 29656 14424 29708
rect 14832 29588 14884 29640
rect 15016 29588 15068 29640
rect 20812 29656 20864 29708
rect 21088 29656 21140 29708
rect 21732 29656 21784 29708
rect 22376 29656 22428 29708
rect 23020 29656 23072 29708
rect 10048 29452 10100 29504
rect 12348 29452 12400 29504
rect 12716 29452 12768 29504
rect 15108 29563 15160 29572
rect 15108 29529 15117 29563
rect 15117 29529 15151 29563
rect 15151 29529 15160 29563
rect 15108 29520 15160 29529
rect 14648 29452 14700 29504
rect 18144 29588 18196 29640
rect 23204 29631 23256 29640
rect 23204 29597 23213 29631
rect 23213 29597 23247 29631
rect 23247 29597 23256 29631
rect 23204 29588 23256 29597
rect 23388 29588 23440 29640
rect 23848 29656 23900 29708
rect 24676 29588 24728 29640
rect 26332 29724 26384 29776
rect 30564 29792 30616 29844
rect 31576 29792 31628 29844
rect 33140 29792 33192 29844
rect 34980 29792 35032 29844
rect 35808 29792 35860 29844
rect 36636 29792 36688 29844
rect 37464 29792 37516 29844
rect 38200 29792 38252 29844
rect 38936 29792 38988 29844
rect 39580 29792 39632 29844
rect 15568 29520 15620 29572
rect 16948 29563 17000 29572
rect 16948 29529 16957 29563
rect 16957 29529 16991 29563
rect 16991 29529 17000 29563
rect 16948 29520 17000 29529
rect 18236 29520 18288 29572
rect 22192 29520 22244 29572
rect 22744 29520 22796 29572
rect 15476 29495 15528 29504
rect 15476 29461 15485 29495
rect 15485 29461 15519 29495
rect 15519 29461 15528 29495
rect 15476 29452 15528 29461
rect 17684 29452 17736 29504
rect 21088 29452 21140 29504
rect 21824 29452 21876 29504
rect 22468 29495 22520 29504
rect 22468 29461 22477 29495
rect 22477 29461 22511 29495
rect 22511 29461 22520 29495
rect 22468 29452 22520 29461
rect 22652 29495 22704 29504
rect 22652 29461 22661 29495
rect 22661 29461 22695 29495
rect 22695 29461 22704 29495
rect 22652 29452 22704 29461
rect 23204 29452 23256 29504
rect 23664 29452 23716 29504
rect 24308 29520 24360 29572
rect 26516 29656 26568 29708
rect 26424 29588 26476 29640
rect 28632 29656 28684 29708
rect 26792 29588 26844 29640
rect 29736 29724 29788 29776
rect 30288 29724 30340 29776
rect 29368 29631 29420 29640
rect 29368 29597 29377 29631
rect 29377 29597 29411 29631
rect 29411 29597 29420 29631
rect 29368 29588 29420 29597
rect 29460 29588 29512 29640
rect 30012 29656 30064 29708
rect 30288 29588 30340 29640
rect 30380 29588 30432 29640
rect 30932 29588 30984 29640
rect 31024 29631 31076 29640
rect 31024 29597 31033 29631
rect 31033 29597 31067 29631
rect 31067 29597 31076 29631
rect 31024 29588 31076 29597
rect 31852 29724 31904 29776
rect 32312 29724 32364 29776
rect 33508 29724 33560 29776
rect 34336 29724 34388 29776
rect 38568 29724 38620 29776
rect 32772 29656 32824 29708
rect 31668 29631 31720 29640
rect 31668 29597 31677 29631
rect 31677 29597 31711 29631
rect 31711 29597 31720 29631
rect 31668 29588 31720 29597
rect 32864 29588 32916 29640
rect 27528 29452 27580 29504
rect 27804 29452 27856 29504
rect 29828 29452 29880 29504
rect 33232 29520 33284 29572
rect 33508 29588 33560 29640
rect 35992 29656 36044 29708
rect 34336 29631 34388 29640
rect 34336 29597 34345 29631
rect 34345 29597 34379 29631
rect 34379 29597 34388 29631
rect 34336 29588 34388 29597
rect 34704 29631 34756 29640
rect 34704 29597 34713 29631
rect 34713 29597 34747 29631
rect 34747 29597 34756 29631
rect 34704 29588 34756 29597
rect 34888 29588 34940 29640
rect 34980 29631 35032 29640
rect 34980 29597 34989 29631
rect 34989 29597 35023 29631
rect 35023 29597 35032 29631
rect 34980 29588 35032 29597
rect 30380 29452 30432 29504
rect 30472 29495 30524 29504
rect 30472 29461 30481 29495
rect 30481 29461 30515 29495
rect 30515 29461 30524 29495
rect 30472 29452 30524 29461
rect 31116 29452 31168 29504
rect 32772 29452 32824 29504
rect 34060 29495 34112 29504
rect 34060 29461 34069 29495
rect 34069 29461 34103 29495
rect 34103 29461 34112 29495
rect 34060 29452 34112 29461
rect 34980 29452 35032 29504
rect 35532 29588 35584 29640
rect 36912 29631 36964 29640
rect 36912 29597 36921 29631
rect 36921 29597 36955 29631
rect 36955 29597 36964 29631
rect 36912 29588 36964 29597
rect 39212 29656 39264 29708
rect 36268 29520 36320 29572
rect 37648 29520 37700 29572
rect 38476 29631 38528 29640
rect 38476 29597 38485 29631
rect 38485 29597 38519 29631
rect 38519 29597 38528 29631
rect 38476 29588 38528 29597
rect 38752 29588 38804 29640
rect 35808 29452 35860 29504
rect 36636 29452 36688 29504
rect 37004 29495 37056 29504
rect 37004 29461 37013 29495
rect 37013 29461 37047 29495
rect 37047 29461 37056 29495
rect 37004 29452 37056 29461
rect 38752 29452 38804 29504
rect 38844 29452 38896 29504
rect 41512 29588 41564 29640
rect 40684 29520 40736 29572
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 2688 29248 2740 29300
rect 4528 29248 4580 29300
rect 5356 29248 5408 29300
rect 5540 29248 5592 29300
rect 3608 29180 3660 29232
rect 4160 29223 4212 29232
rect 4160 29189 4169 29223
rect 4169 29189 4203 29223
rect 4203 29189 4212 29223
rect 4160 29180 4212 29189
rect 4896 29223 4948 29232
rect 4896 29189 4905 29223
rect 4905 29189 4939 29223
rect 4939 29189 4948 29223
rect 4896 29180 4948 29189
rect 3240 29112 3292 29164
rect 3424 29155 3476 29164
rect 3424 29121 3433 29155
rect 3433 29121 3467 29155
rect 3467 29121 3476 29155
rect 3424 29112 3476 29121
rect 5080 29155 5132 29164
rect 5080 29121 5089 29155
rect 5089 29121 5123 29155
rect 5123 29121 5132 29155
rect 5080 29112 5132 29121
rect 5172 29112 5224 29164
rect 5264 29112 5316 29164
rect 5356 29155 5408 29164
rect 5356 29121 5365 29155
rect 5365 29121 5399 29155
rect 5399 29121 5408 29155
rect 5356 29112 5408 29121
rect 5908 29180 5960 29232
rect 5632 29155 5684 29164
rect 5632 29121 5641 29155
rect 5641 29121 5675 29155
rect 5675 29121 5684 29155
rect 5632 29112 5684 29121
rect 5816 29155 5868 29164
rect 5816 29121 5830 29155
rect 5830 29121 5864 29155
rect 5864 29121 5868 29155
rect 7104 29248 7156 29300
rect 7840 29248 7892 29300
rect 5816 29112 5868 29121
rect 6276 29112 6328 29164
rect 6552 29155 6604 29164
rect 6552 29121 6561 29155
rect 6561 29121 6595 29155
rect 6595 29121 6604 29155
rect 6552 29112 6604 29121
rect 6644 29155 6696 29164
rect 6644 29121 6653 29155
rect 6653 29121 6687 29155
rect 6687 29121 6696 29155
rect 6644 29112 6696 29121
rect 6736 29155 6788 29164
rect 6736 29121 6745 29155
rect 6745 29121 6779 29155
rect 6779 29121 6788 29155
rect 6736 29112 6788 29121
rect 7380 29112 7432 29164
rect 7564 29155 7616 29164
rect 7564 29121 7573 29155
rect 7573 29121 7607 29155
rect 7607 29121 7616 29155
rect 7564 29112 7616 29121
rect 7656 29155 7708 29164
rect 7656 29121 7665 29155
rect 7665 29121 7699 29155
rect 7699 29121 7708 29155
rect 7656 29112 7708 29121
rect 7932 29155 7984 29164
rect 7932 29121 7941 29155
rect 7941 29121 7975 29155
rect 7975 29121 7984 29155
rect 7932 29112 7984 29121
rect 8392 29248 8444 29300
rect 9680 29248 9732 29300
rect 8208 29223 8260 29232
rect 8208 29189 8217 29223
rect 8217 29189 8251 29223
rect 8251 29189 8260 29223
rect 8208 29180 8260 29189
rect 8576 29180 8628 29232
rect 8668 29223 8720 29232
rect 8668 29189 8677 29223
rect 8677 29189 8711 29223
rect 8711 29189 8720 29223
rect 8668 29180 8720 29189
rect 9128 29180 9180 29232
rect 8300 29155 8352 29164
rect 8300 29121 8309 29155
rect 8309 29121 8343 29155
rect 8343 29121 8352 29155
rect 8300 29112 8352 29121
rect 9312 29112 9364 29164
rect 10048 29223 10100 29232
rect 10048 29189 10057 29223
rect 10057 29189 10091 29223
rect 10091 29189 10100 29223
rect 10048 29180 10100 29189
rect 11704 29248 11756 29300
rect 11520 29180 11572 29232
rect 9864 29155 9916 29164
rect 9864 29121 9871 29155
rect 9871 29121 9916 29155
rect 3332 28976 3384 29028
rect 1860 28951 1912 28960
rect 1860 28917 1869 28951
rect 1869 28917 1903 28951
rect 1903 28917 1912 28951
rect 1860 28908 1912 28917
rect 5724 28976 5776 29028
rect 5816 28976 5868 29028
rect 6828 28976 6880 29028
rect 7380 28976 7432 29028
rect 8300 28976 8352 29028
rect 8392 28976 8444 29028
rect 9036 29044 9088 29096
rect 9864 29112 9916 29121
rect 10140 29112 10192 29164
rect 11060 29112 11112 29164
rect 12348 29223 12400 29232
rect 12348 29189 12357 29223
rect 12357 29189 12391 29223
rect 12391 29189 12400 29223
rect 12348 29180 12400 29189
rect 12532 29248 12584 29300
rect 13360 29248 13412 29300
rect 13544 29248 13596 29300
rect 14096 29248 14148 29300
rect 14372 29248 14424 29300
rect 15108 29248 15160 29300
rect 16948 29248 17000 29300
rect 17684 29248 17736 29300
rect 10416 29044 10468 29096
rect 7012 28908 7064 28960
rect 7840 28951 7892 28960
rect 7840 28917 7849 28951
rect 7849 28917 7883 28951
rect 7883 28917 7892 28951
rect 7840 28908 7892 28917
rect 8208 28908 8260 28960
rect 8852 28908 8904 28960
rect 10324 28951 10376 28960
rect 10324 28917 10333 28951
rect 10333 28917 10367 28951
rect 10367 28917 10376 28951
rect 10324 28908 10376 28917
rect 11612 28908 11664 28960
rect 12716 29112 12768 29164
rect 12808 29155 12860 29164
rect 12808 29121 12817 29155
rect 12817 29121 12851 29155
rect 12851 29121 12860 29155
rect 12808 29112 12860 29121
rect 12992 29155 13044 29164
rect 12992 29121 12999 29155
rect 12999 29121 13044 29155
rect 12992 29112 13044 29121
rect 13176 29155 13228 29164
rect 13176 29121 13185 29155
rect 13185 29121 13219 29155
rect 13219 29121 13228 29155
rect 13176 29112 13228 29121
rect 13452 29112 13504 29164
rect 12808 28976 12860 29028
rect 13728 29155 13780 29164
rect 13728 29121 13737 29155
rect 13737 29121 13771 29155
rect 13771 29121 13780 29155
rect 13728 29112 13780 29121
rect 14280 29155 14332 29164
rect 14280 29121 14289 29155
rect 14289 29121 14323 29155
rect 14323 29121 14332 29155
rect 14280 29112 14332 29121
rect 14832 29155 14884 29164
rect 14832 29121 14841 29155
rect 14841 29121 14875 29155
rect 14875 29121 14884 29155
rect 14832 29112 14884 29121
rect 15108 29112 15160 29164
rect 13360 28976 13412 29028
rect 15016 29087 15068 29096
rect 15016 29053 15025 29087
rect 15025 29053 15059 29087
rect 15059 29053 15068 29087
rect 15016 29044 15068 29053
rect 15108 28976 15160 29028
rect 15384 29155 15436 29164
rect 15384 29121 15394 29155
rect 15394 29121 15428 29155
rect 15428 29121 15436 29155
rect 15844 29180 15896 29232
rect 15384 29112 15436 29121
rect 15660 29155 15712 29164
rect 15660 29121 15669 29155
rect 15669 29121 15703 29155
rect 15703 29121 15712 29155
rect 15660 29112 15712 29121
rect 16212 29155 16264 29164
rect 16212 29121 16221 29155
rect 16221 29121 16255 29155
rect 16255 29121 16264 29155
rect 16212 29112 16264 29121
rect 16488 29112 16540 29164
rect 17500 29180 17552 29232
rect 21640 29248 21692 29300
rect 15936 29044 15988 29096
rect 16948 29112 17000 29164
rect 17224 29155 17276 29164
rect 17224 29121 17233 29155
rect 17233 29121 17267 29155
rect 17267 29121 17276 29155
rect 17224 29112 17276 29121
rect 17408 29155 17460 29164
rect 17408 29121 17417 29155
rect 17417 29121 17451 29155
rect 17451 29121 17460 29155
rect 17408 29112 17460 29121
rect 15568 28976 15620 29028
rect 15752 28976 15804 29028
rect 16948 28976 17000 29028
rect 17040 29019 17092 29028
rect 17040 28985 17049 29019
rect 17049 28985 17083 29019
rect 17083 28985 17092 29019
rect 17040 28976 17092 28985
rect 17592 28976 17644 29028
rect 12532 28908 12584 28960
rect 13544 28908 13596 28960
rect 14188 28908 14240 28960
rect 18328 29112 18380 29164
rect 18512 29155 18564 29164
rect 18512 29121 18521 29155
rect 18521 29121 18555 29155
rect 18555 29121 18564 29155
rect 18512 29112 18564 29121
rect 18880 29112 18932 29164
rect 18420 28976 18472 29028
rect 18696 29019 18748 29028
rect 18696 28985 18705 29019
rect 18705 28985 18739 29019
rect 18739 28985 18748 29019
rect 18696 28976 18748 28985
rect 19432 29112 19484 29164
rect 20628 29180 20680 29232
rect 20536 29155 20588 29164
rect 20536 29121 20545 29155
rect 20545 29121 20579 29155
rect 20579 29121 20588 29155
rect 20536 29112 20588 29121
rect 21456 29112 21508 29164
rect 19524 29044 19576 29096
rect 19892 28976 19944 29028
rect 21272 29087 21324 29096
rect 21272 29053 21281 29087
rect 21281 29053 21315 29087
rect 21315 29053 21324 29087
rect 21272 29044 21324 29053
rect 22008 29180 22060 29232
rect 21916 29112 21968 29164
rect 22744 29180 22796 29232
rect 23480 29248 23532 29300
rect 26516 29248 26568 29300
rect 30472 29248 30524 29300
rect 30932 29248 30984 29300
rect 32956 29248 33008 29300
rect 22468 29155 22520 29164
rect 22468 29121 22477 29155
rect 22477 29121 22511 29155
rect 22511 29121 22520 29155
rect 22468 29112 22520 29121
rect 23480 29155 23532 29164
rect 23480 29121 23489 29155
rect 23489 29121 23523 29155
rect 23523 29121 23532 29155
rect 23480 29112 23532 29121
rect 24216 29155 24268 29164
rect 24216 29121 24225 29155
rect 24225 29121 24259 29155
rect 24259 29121 24268 29155
rect 24216 29112 24268 29121
rect 22560 29044 22612 29096
rect 24952 29180 25004 29232
rect 24860 29155 24912 29164
rect 24860 29121 24869 29155
rect 24869 29121 24903 29155
rect 24903 29121 24912 29155
rect 24860 29112 24912 29121
rect 25228 29155 25280 29164
rect 25228 29121 25237 29155
rect 25237 29121 25271 29155
rect 25271 29121 25280 29155
rect 25228 29112 25280 29121
rect 24492 29044 24544 29096
rect 22192 28976 22244 29028
rect 23388 28976 23440 29028
rect 25504 29112 25556 29164
rect 26976 29112 27028 29164
rect 29736 29155 29788 29164
rect 29736 29121 29745 29155
rect 29745 29121 29779 29155
rect 29779 29121 29788 29155
rect 29736 29112 29788 29121
rect 29828 29155 29880 29164
rect 29828 29121 29837 29155
rect 29837 29121 29871 29155
rect 29871 29121 29880 29155
rect 29828 29112 29880 29121
rect 31392 29180 31444 29232
rect 31116 29155 31168 29164
rect 31116 29121 31125 29155
rect 31125 29121 31159 29155
rect 31159 29121 31168 29155
rect 31116 29112 31168 29121
rect 31208 29155 31260 29164
rect 31208 29121 31217 29155
rect 31217 29121 31251 29155
rect 31251 29121 31260 29155
rect 31208 29112 31260 29121
rect 31668 29112 31720 29164
rect 31852 29155 31904 29164
rect 31852 29121 31861 29155
rect 31861 29121 31895 29155
rect 31895 29121 31904 29155
rect 31852 29112 31904 29121
rect 33140 29180 33192 29232
rect 32496 29155 32548 29164
rect 18512 28908 18564 28960
rect 19248 28908 19300 28960
rect 20720 28908 20772 28960
rect 25780 28976 25832 29028
rect 27344 28976 27396 29028
rect 24308 28908 24360 28960
rect 25964 28908 26016 28960
rect 26424 28908 26476 28960
rect 26608 28908 26660 28960
rect 27252 28908 27304 28960
rect 28264 28908 28316 28960
rect 29368 28908 29420 28960
rect 29460 28908 29512 28960
rect 29736 28976 29788 29028
rect 30472 28976 30524 29028
rect 30564 28976 30616 29028
rect 31116 28976 31168 29028
rect 32496 29121 32543 29155
rect 32543 29121 32548 29155
rect 32496 29112 32548 29121
rect 32864 29087 32916 29096
rect 32864 29053 32873 29087
rect 32873 29053 32907 29087
rect 32907 29053 32916 29087
rect 32864 29044 32916 29053
rect 33048 29112 33100 29164
rect 33416 29248 33468 29300
rect 35164 29248 35216 29300
rect 39120 29248 39172 29300
rect 33692 29223 33744 29232
rect 33692 29189 33701 29223
rect 33701 29189 33735 29223
rect 33735 29189 33744 29223
rect 33692 29180 33744 29189
rect 34428 29155 34480 29164
rect 34428 29121 34437 29155
rect 34437 29121 34471 29155
rect 34471 29121 34480 29155
rect 34428 29112 34480 29121
rect 35900 29180 35952 29232
rect 35992 29112 36044 29164
rect 37464 29112 37516 29164
rect 37648 29112 37700 29164
rect 34888 29087 34940 29096
rect 34888 29053 34897 29087
rect 34897 29053 34931 29087
rect 34931 29053 34940 29087
rect 34888 29044 34940 29053
rect 35164 29087 35216 29096
rect 35164 29053 35173 29087
rect 35173 29053 35207 29087
rect 35207 29053 35216 29087
rect 35164 29044 35216 29053
rect 35900 29044 35952 29096
rect 34980 28976 35032 29028
rect 29828 28908 29880 28960
rect 32036 28908 32088 28960
rect 32312 28908 32364 28960
rect 32588 28908 32640 28960
rect 32956 28908 33008 28960
rect 33600 28908 33652 28960
rect 35256 28908 35308 28960
rect 37372 28976 37424 29028
rect 38844 28976 38896 29028
rect 39488 28976 39540 29028
rect 37648 28908 37700 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 5356 28704 5408 28756
rect 5816 28704 5868 28756
rect 11060 28747 11112 28756
rect 11060 28713 11069 28747
rect 11069 28713 11103 28747
rect 11103 28713 11112 28747
rect 11060 28704 11112 28713
rect 12256 28704 12308 28756
rect 5540 28636 5592 28688
rect 2504 28568 2556 28620
rect 1400 28500 1452 28552
rect 3056 28568 3108 28620
rect 4804 28568 4856 28620
rect 5172 28500 5224 28552
rect 8300 28636 8352 28688
rect 7840 28568 7892 28620
rect 5908 28543 5960 28552
rect 5908 28509 5917 28543
rect 5917 28509 5951 28543
rect 5951 28509 5960 28543
rect 5908 28500 5960 28509
rect 6644 28500 6696 28552
rect 7564 28500 7616 28552
rect 10968 28636 11020 28688
rect 12716 28704 12768 28756
rect 14280 28704 14332 28756
rect 3608 28475 3660 28484
rect 3608 28441 3617 28475
rect 3617 28441 3651 28475
rect 3651 28441 3660 28475
rect 3608 28432 3660 28441
rect 5264 28432 5316 28484
rect 7380 28432 7432 28484
rect 10048 28543 10100 28552
rect 10048 28509 10057 28543
rect 10057 28509 10091 28543
rect 10091 28509 10100 28543
rect 10048 28500 10100 28509
rect 10232 28543 10284 28552
rect 10232 28509 10241 28543
rect 10241 28509 10275 28543
rect 10275 28509 10284 28543
rect 10232 28500 10284 28509
rect 11336 28500 11388 28552
rect 11704 28543 11756 28552
rect 11704 28509 11713 28543
rect 11713 28509 11747 28543
rect 11747 28509 11756 28543
rect 11704 28500 11756 28509
rect 11980 28500 12032 28552
rect 11612 28432 11664 28484
rect 12164 28500 12216 28552
rect 12716 28500 12768 28552
rect 13452 28636 13504 28688
rect 15016 28704 15068 28756
rect 15568 28747 15620 28756
rect 15568 28713 15577 28747
rect 15577 28713 15611 28747
rect 15611 28713 15620 28747
rect 15568 28704 15620 28713
rect 15752 28704 15804 28756
rect 16212 28704 16264 28756
rect 17040 28704 17092 28756
rect 17684 28704 17736 28756
rect 13084 28543 13136 28552
rect 13084 28509 13093 28543
rect 13093 28509 13127 28543
rect 13127 28509 13136 28543
rect 13084 28500 13136 28509
rect 14096 28500 14148 28552
rect 14372 28500 14424 28552
rect 14832 28636 14884 28688
rect 19432 28747 19484 28756
rect 19432 28713 19441 28747
rect 19441 28713 19475 28747
rect 19475 28713 19484 28747
rect 19432 28704 19484 28713
rect 19800 28704 19852 28756
rect 21272 28704 21324 28756
rect 21548 28704 21600 28756
rect 21732 28704 21784 28756
rect 21824 28747 21876 28756
rect 21824 28713 21833 28747
rect 21833 28713 21867 28747
rect 21867 28713 21876 28747
rect 21824 28704 21876 28713
rect 22100 28704 22152 28756
rect 23020 28704 23072 28756
rect 24032 28704 24084 28756
rect 24400 28704 24452 28756
rect 24952 28747 25004 28756
rect 24952 28713 24961 28747
rect 24961 28713 24995 28747
rect 24995 28713 25004 28747
rect 24952 28704 25004 28713
rect 25320 28704 25372 28756
rect 25964 28704 26016 28756
rect 26792 28704 26844 28756
rect 27712 28704 27764 28756
rect 28172 28704 28224 28756
rect 15016 28543 15068 28552
rect 15016 28509 15025 28543
rect 15025 28509 15059 28543
rect 15059 28509 15068 28543
rect 15016 28500 15068 28509
rect 15108 28543 15160 28552
rect 15108 28509 15117 28543
rect 15117 28509 15151 28543
rect 15151 28509 15160 28543
rect 15108 28500 15160 28509
rect 15384 28500 15436 28552
rect 15476 28500 15528 28552
rect 15936 28543 15988 28552
rect 15936 28509 15945 28543
rect 15945 28509 15979 28543
rect 15979 28509 15988 28543
rect 15936 28500 15988 28509
rect 5908 28364 5960 28416
rect 6184 28364 6236 28416
rect 7748 28407 7800 28416
rect 7748 28373 7757 28407
rect 7757 28373 7791 28407
rect 7791 28373 7800 28407
rect 7748 28364 7800 28373
rect 8852 28364 8904 28416
rect 9864 28364 9916 28416
rect 10232 28364 10284 28416
rect 10508 28364 10560 28416
rect 10968 28364 11020 28416
rect 11152 28364 11204 28416
rect 11244 28407 11296 28416
rect 11244 28373 11253 28407
rect 11253 28373 11287 28407
rect 11287 28373 11296 28407
rect 11244 28364 11296 28373
rect 11520 28364 11572 28416
rect 15568 28475 15620 28484
rect 15568 28441 15577 28475
rect 15577 28441 15611 28475
rect 15611 28441 15620 28475
rect 15568 28432 15620 28441
rect 15844 28432 15896 28484
rect 11980 28364 12032 28416
rect 12624 28364 12676 28416
rect 13268 28364 13320 28416
rect 14832 28364 14884 28416
rect 14924 28364 14976 28416
rect 17408 28500 17460 28552
rect 18144 28543 18196 28552
rect 18144 28509 18153 28543
rect 18153 28509 18187 28543
rect 18187 28509 18196 28543
rect 18144 28500 18196 28509
rect 18236 28500 18288 28552
rect 17500 28475 17552 28484
rect 17500 28441 17509 28475
rect 17509 28441 17543 28475
rect 17543 28441 17552 28475
rect 17500 28432 17552 28441
rect 17684 28475 17736 28484
rect 17684 28441 17693 28475
rect 17693 28441 17727 28475
rect 17727 28441 17736 28475
rect 17684 28432 17736 28441
rect 18512 28500 18564 28552
rect 19892 28636 19944 28688
rect 21180 28611 21232 28620
rect 21180 28577 21195 28611
rect 21195 28577 21229 28611
rect 21229 28577 21232 28611
rect 22560 28636 22612 28688
rect 21180 28568 21232 28577
rect 20352 28500 20404 28552
rect 19156 28432 19208 28484
rect 19248 28475 19300 28484
rect 19248 28441 19257 28475
rect 19257 28441 19291 28475
rect 19291 28441 19300 28475
rect 19248 28432 19300 28441
rect 19524 28432 19576 28484
rect 19800 28432 19852 28484
rect 20996 28500 21048 28552
rect 21088 28543 21140 28552
rect 21088 28509 21097 28543
rect 21097 28509 21131 28543
rect 21131 28509 21140 28543
rect 21088 28500 21140 28509
rect 21456 28543 21508 28552
rect 21456 28509 21465 28543
rect 21465 28509 21499 28543
rect 21499 28509 21508 28543
rect 21456 28500 21508 28509
rect 21548 28500 21600 28552
rect 22100 28568 22152 28620
rect 22468 28568 22520 28620
rect 21272 28475 21324 28484
rect 21272 28441 21281 28475
rect 21281 28441 21315 28475
rect 21315 28441 21324 28475
rect 21272 28432 21324 28441
rect 22192 28432 22244 28484
rect 22560 28500 22612 28552
rect 23020 28543 23072 28552
rect 23020 28509 23029 28543
rect 23029 28509 23063 28543
rect 23063 28509 23072 28543
rect 23020 28500 23072 28509
rect 23572 28679 23624 28688
rect 23572 28645 23581 28679
rect 23581 28645 23615 28679
rect 23615 28645 23624 28679
rect 23572 28636 23624 28645
rect 23388 28543 23440 28552
rect 23388 28509 23397 28543
rect 23397 28509 23431 28543
rect 23431 28509 23440 28543
rect 23388 28500 23440 28509
rect 23480 28543 23532 28552
rect 23480 28509 23489 28543
rect 23489 28509 23523 28543
rect 23523 28509 23532 28543
rect 23480 28500 23532 28509
rect 23664 28543 23716 28552
rect 23664 28509 23673 28543
rect 23673 28509 23707 28543
rect 23707 28509 23716 28543
rect 23664 28500 23716 28509
rect 23756 28543 23808 28552
rect 23756 28509 23765 28543
rect 23765 28509 23799 28543
rect 23799 28509 23808 28543
rect 23756 28500 23808 28509
rect 24492 28636 24544 28688
rect 28724 28704 28776 28756
rect 29184 28704 29236 28756
rect 29460 28704 29512 28756
rect 30012 28704 30064 28756
rect 31024 28704 31076 28756
rect 36268 28704 36320 28756
rect 36728 28704 36780 28756
rect 17408 28407 17460 28416
rect 17408 28373 17417 28407
rect 17417 28373 17451 28407
rect 17451 28373 17460 28407
rect 17408 28364 17460 28373
rect 18512 28364 18564 28416
rect 20720 28364 20772 28416
rect 22744 28364 22796 28416
rect 24032 28364 24084 28416
rect 24860 28500 24912 28552
rect 25044 28500 25096 28552
rect 25320 28500 25372 28552
rect 25504 28543 25556 28552
rect 25504 28509 25513 28543
rect 25513 28509 25547 28543
rect 25547 28509 25556 28543
rect 25504 28500 25556 28509
rect 24492 28432 24544 28484
rect 24952 28432 25004 28484
rect 26424 28543 26476 28552
rect 26424 28509 26433 28543
rect 26433 28509 26467 28543
rect 26467 28509 26476 28543
rect 26424 28500 26476 28509
rect 26608 28500 26660 28552
rect 26700 28500 26752 28552
rect 26884 28568 26936 28620
rect 24768 28364 24820 28416
rect 25228 28364 25280 28416
rect 25872 28407 25924 28416
rect 25872 28373 25897 28407
rect 25897 28373 25924 28407
rect 26240 28432 26292 28484
rect 26884 28466 26936 28518
rect 27160 28543 27212 28552
rect 27160 28509 27169 28543
rect 27169 28509 27203 28543
rect 27203 28509 27212 28543
rect 27160 28500 27212 28509
rect 27252 28500 27304 28552
rect 27436 28500 27488 28552
rect 27528 28543 27580 28552
rect 27528 28509 27537 28543
rect 27537 28509 27571 28543
rect 27571 28509 27580 28543
rect 27528 28500 27580 28509
rect 25872 28364 25924 28373
rect 26884 28364 26936 28416
rect 27252 28364 27304 28416
rect 27528 28364 27580 28416
rect 27712 28364 27764 28416
rect 28356 28500 28408 28552
rect 28172 28432 28224 28484
rect 28264 28407 28316 28416
rect 28264 28373 28273 28407
rect 28273 28373 28307 28407
rect 28307 28373 28316 28407
rect 28264 28364 28316 28373
rect 28356 28364 28408 28416
rect 28908 28500 28960 28552
rect 29092 28636 29144 28688
rect 29368 28568 29420 28620
rect 33692 28568 33744 28620
rect 29184 28543 29236 28552
rect 29184 28509 29198 28543
rect 29198 28509 29232 28543
rect 29232 28509 29236 28543
rect 29184 28500 29236 28509
rect 29828 28500 29880 28552
rect 31208 28500 31260 28552
rect 31392 28500 31444 28552
rect 32036 28500 32088 28552
rect 32772 28500 32824 28552
rect 34336 28636 34388 28688
rect 34704 28679 34756 28688
rect 34704 28645 34713 28679
rect 34713 28645 34747 28679
rect 34747 28645 34756 28679
rect 34704 28636 34756 28645
rect 34520 28568 34572 28620
rect 29000 28475 29052 28484
rect 29000 28441 29009 28475
rect 29009 28441 29043 28475
rect 29043 28441 29052 28475
rect 29000 28432 29052 28441
rect 29644 28432 29696 28484
rect 29184 28364 29236 28416
rect 31024 28364 31076 28416
rect 31392 28364 31444 28416
rect 32128 28432 32180 28484
rect 34152 28500 34204 28552
rect 34796 28500 34848 28552
rect 34980 28543 35032 28552
rect 34980 28509 34989 28543
rect 34989 28509 35023 28543
rect 35023 28509 35032 28543
rect 34980 28500 35032 28509
rect 35348 28568 35400 28620
rect 35532 28500 35584 28552
rect 37832 28636 37884 28688
rect 35808 28500 35860 28552
rect 32588 28364 32640 28416
rect 33968 28364 34020 28416
rect 34980 28364 35032 28416
rect 35624 28364 35676 28416
rect 37556 28500 37608 28552
rect 37832 28500 37884 28552
rect 36820 28432 36872 28484
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 1860 28160 1912 28212
rect 5448 28160 5500 28212
rect 6184 28160 6236 28212
rect 9312 28160 9364 28212
rect 3056 28092 3108 28144
rect 5724 28135 5776 28144
rect 5724 28101 5733 28135
rect 5733 28101 5767 28135
rect 5767 28101 5776 28135
rect 5724 28092 5776 28101
rect 1400 28067 1452 28076
rect 1400 28033 1409 28067
rect 1409 28033 1443 28067
rect 1443 28033 1452 28067
rect 1400 28024 1452 28033
rect 4988 28024 5040 28076
rect 5356 28024 5408 28076
rect 3332 27956 3384 28008
rect 6092 27956 6144 28008
rect 11244 28160 11296 28212
rect 12532 28160 12584 28212
rect 12716 28160 12768 28212
rect 13452 28160 13504 28212
rect 14188 28160 14240 28212
rect 20996 28160 21048 28212
rect 21180 28160 21232 28212
rect 22284 28160 22336 28212
rect 11888 28092 11940 28144
rect 12164 28067 12216 28076
rect 12164 28033 12173 28067
rect 12173 28033 12207 28067
rect 12207 28033 12216 28067
rect 12164 28024 12216 28033
rect 12256 28024 12308 28076
rect 14464 28092 14516 28144
rect 15568 28092 15620 28144
rect 19064 28092 19116 28144
rect 19248 28092 19300 28144
rect 12624 28024 12676 28076
rect 14188 28024 14240 28076
rect 15384 28024 15436 28076
rect 15844 28024 15896 28076
rect 18052 28024 18104 28076
rect 20812 28067 20864 28076
rect 20812 28033 20821 28067
rect 20821 28033 20855 28067
rect 20855 28033 20864 28067
rect 20812 28024 20864 28033
rect 21272 28092 21324 28144
rect 22836 28092 22888 28144
rect 23020 28092 23072 28144
rect 23388 28160 23440 28212
rect 23848 28160 23900 28212
rect 24952 28160 25004 28212
rect 25872 28160 25924 28212
rect 26424 28160 26476 28212
rect 27252 28160 27304 28212
rect 23756 28092 23808 28144
rect 25320 28092 25372 28144
rect 13544 27956 13596 28008
rect 17684 27956 17736 28008
rect 19340 27956 19392 28008
rect 20352 27956 20404 28008
rect 21824 28024 21876 28076
rect 22560 28024 22612 28076
rect 24032 28024 24084 28076
rect 26424 28067 26476 28076
rect 26424 28033 26433 28067
rect 26433 28033 26467 28067
rect 26467 28033 26476 28067
rect 26424 28024 26476 28033
rect 22744 27956 22796 28008
rect 23480 27956 23532 28008
rect 23664 27956 23716 28008
rect 24860 27956 24912 28008
rect 26700 27956 26752 28008
rect 27252 28024 27304 28076
rect 27528 28092 27580 28144
rect 27620 27956 27672 28008
rect 8668 27888 8720 27940
rect 13636 27888 13688 27940
rect 14280 27888 14332 27940
rect 15016 27888 15068 27940
rect 17224 27888 17276 27940
rect 4712 27820 4764 27872
rect 8300 27820 8352 27872
rect 10048 27820 10100 27872
rect 10324 27820 10376 27872
rect 12164 27820 12216 27872
rect 19524 27820 19576 27872
rect 25044 27888 25096 27940
rect 25136 27888 25188 27940
rect 27528 27888 27580 27940
rect 27988 28067 28040 28076
rect 27988 28033 27997 28067
rect 27997 28033 28031 28067
rect 28031 28033 28040 28067
rect 27988 28024 28040 28033
rect 28172 28067 28224 28076
rect 28172 28033 28181 28067
rect 28181 28033 28215 28067
rect 28215 28033 28224 28067
rect 28172 28024 28224 28033
rect 28356 28203 28408 28212
rect 28356 28169 28365 28203
rect 28365 28169 28399 28203
rect 28399 28169 28408 28203
rect 28356 28160 28408 28169
rect 28540 28160 28592 28212
rect 29092 28160 29144 28212
rect 32312 28160 32364 28212
rect 32588 28160 32640 28212
rect 31760 28092 31812 28144
rect 32772 28092 32824 28144
rect 34336 28160 34388 28212
rect 34704 28160 34756 28212
rect 37464 28160 37516 28212
rect 38384 28160 38436 28212
rect 28080 27956 28132 28008
rect 28540 27956 28592 28008
rect 28908 28067 28960 28076
rect 28908 28033 28917 28067
rect 28917 28033 28951 28067
rect 28951 28033 28960 28067
rect 28908 28024 28960 28033
rect 29276 28024 29328 28076
rect 31576 28024 31628 28076
rect 35716 28135 35768 28144
rect 35716 28101 35725 28135
rect 35725 28101 35759 28135
rect 35759 28101 35768 28135
rect 35716 28092 35768 28101
rect 21272 27820 21324 27872
rect 22284 27820 22336 27872
rect 25964 27820 26016 27872
rect 26148 27820 26200 27872
rect 26884 27820 26936 27872
rect 27712 27820 27764 27872
rect 28356 27888 28408 27940
rect 28264 27820 28316 27872
rect 28724 27863 28776 27872
rect 28724 27829 28733 27863
rect 28733 27829 28767 27863
rect 28767 27829 28776 27863
rect 28724 27820 28776 27829
rect 29092 27931 29144 27940
rect 29092 27897 29101 27931
rect 29101 27897 29135 27931
rect 29135 27897 29144 27931
rect 29092 27888 29144 27897
rect 34520 28024 34572 28076
rect 35900 28024 35952 28076
rect 36912 28024 36964 28076
rect 38016 28024 38068 28076
rect 38292 28067 38344 28076
rect 38292 28033 38301 28067
rect 38301 28033 38335 28067
rect 38335 28033 38344 28067
rect 38292 28024 38344 28033
rect 40040 28092 40092 28144
rect 40684 28092 40736 28144
rect 39028 28067 39080 28076
rect 33968 27999 34020 28008
rect 33968 27965 33977 27999
rect 33977 27965 34011 27999
rect 34011 27965 34020 27999
rect 33968 27956 34020 27965
rect 35532 27956 35584 28008
rect 36452 27956 36504 28008
rect 36544 27999 36596 28008
rect 36544 27965 36553 27999
rect 36553 27965 36587 27999
rect 36587 27965 36596 27999
rect 36544 27956 36596 27965
rect 31024 27820 31076 27872
rect 31300 27820 31352 27872
rect 31852 27820 31904 27872
rect 32588 27820 32640 27872
rect 33784 27863 33836 27872
rect 33784 27829 33793 27863
rect 33793 27829 33827 27863
rect 33827 27829 33836 27863
rect 33784 27820 33836 27829
rect 34704 27820 34756 27872
rect 35992 27888 36044 27940
rect 37372 27956 37424 28008
rect 39028 28033 39044 28067
rect 39044 28033 39078 28067
rect 39078 28033 39080 28067
rect 39028 28024 39080 28033
rect 36360 27820 36412 27872
rect 37280 27863 37332 27872
rect 37280 27829 37289 27863
rect 37289 27829 37323 27863
rect 37323 27829 37332 27863
rect 37280 27820 37332 27829
rect 37556 27820 37608 27872
rect 39304 27999 39356 28008
rect 39304 27965 39313 27999
rect 39313 27965 39347 27999
rect 39347 27965 39356 27999
rect 39304 27956 39356 27965
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 8300 27616 8352 27668
rect 10416 27616 10468 27668
rect 10968 27616 11020 27668
rect 12348 27616 12400 27668
rect 12624 27616 12676 27668
rect 13820 27616 13872 27668
rect 4620 27548 4672 27600
rect 4896 27344 4948 27396
rect 5080 27344 5132 27396
rect 6000 27548 6052 27600
rect 8852 27548 8904 27600
rect 15844 27616 15896 27668
rect 15936 27616 15988 27668
rect 19524 27659 19576 27668
rect 5632 27412 5684 27464
rect 5816 27412 5868 27464
rect 6000 27455 6052 27464
rect 6000 27421 6035 27455
rect 6035 27421 6052 27455
rect 6000 27412 6052 27421
rect 7748 27455 7800 27464
rect 7748 27421 7757 27455
rect 7757 27421 7791 27455
rect 7791 27421 7800 27455
rect 7748 27412 7800 27421
rect 5356 27387 5408 27396
rect 5356 27353 5365 27387
rect 5365 27353 5399 27387
rect 5399 27353 5408 27387
rect 5356 27344 5408 27353
rect 6368 27344 6420 27396
rect 7012 27344 7064 27396
rect 6276 27276 6328 27328
rect 7932 27344 7984 27396
rect 8300 27412 8352 27464
rect 8484 27455 8536 27464
rect 8484 27421 8493 27455
rect 8493 27421 8527 27455
rect 8527 27421 8536 27455
rect 8484 27412 8536 27421
rect 8576 27412 8628 27464
rect 8760 27455 8812 27464
rect 8760 27421 8769 27455
rect 8769 27421 8803 27455
rect 8803 27421 8812 27455
rect 8760 27412 8812 27421
rect 15108 27548 15160 27600
rect 9772 27455 9824 27464
rect 9772 27421 9781 27455
rect 9781 27421 9815 27455
rect 9815 27421 9824 27455
rect 9772 27412 9824 27421
rect 8392 27276 8444 27328
rect 10324 27480 10376 27532
rect 13544 27480 13596 27532
rect 12440 27412 12492 27464
rect 10324 27344 10376 27396
rect 15752 27412 15804 27464
rect 16212 27455 16264 27464
rect 16212 27421 16221 27455
rect 16221 27421 16255 27455
rect 16255 27421 16264 27455
rect 16212 27412 16264 27421
rect 13728 27344 13780 27396
rect 13912 27344 13964 27396
rect 15568 27344 15620 27396
rect 15936 27344 15988 27396
rect 16580 27412 16632 27464
rect 16764 27455 16816 27464
rect 16764 27421 16773 27455
rect 16773 27421 16807 27455
rect 16807 27421 16816 27455
rect 16764 27412 16816 27421
rect 17592 27455 17644 27464
rect 17592 27421 17601 27455
rect 17601 27421 17635 27455
rect 17635 27421 17644 27455
rect 17592 27412 17644 27421
rect 17960 27412 18012 27464
rect 19524 27625 19533 27659
rect 19533 27625 19567 27659
rect 19567 27625 19576 27659
rect 19524 27616 19576 27625
rect 19616 27548 19668 27600
rect 25964 27616 26016 27668
rect 26424 27616 26476 27668
rect 27252 27659 27304 27668
rect 27252 27625 27261 27659
rect 27261 27625 27295 27659
rect 27295 27625 27304 27659
rect 27252 27616 27304 27625
rect 27344 27616 27396 27668
rect 23112 27548 23164 27600
rect 23204 27548 23256 27600
rect 23388 27548 23440 27600
rect 26332 27548 26384 27600
rect 26608 27591 26660 27600
rect 26608 27557 26617 27591
rect 26617 27557 26651 27591
rect 26651 27557 26660 27591
rect 26608 27548 26660 27557
rect 10048 27276 10100 27328
rect 10416 27276 10468 27328
rect 10784 27276 10836 27328
rect 12808 27276 12860 27328
rect 14372 27276 14424 27328
rect 18144 27344 18196 27396
rect 18328 27344 18380 27396
rect 19984 27412 20036 27464
rect 20536 27412 20588 27464
rect 22376 27480 22428 27532
rect 27804 27548 27856 27600
rect 23848 27480 23900 27532
rect 24400 27480 24452 27532
rect 25044 27523 25096 27532
rect 25044 27489 25053 27523
rect 25053 27489 25087 27523
rect 25087 27489 25096 27523
rect 25044 27480 25096 27489
rect 25596 27480 25648 27532
rect 19248 27387 19300 27396
rect 19248 27353 19257 27387
rect 19257 27353 19291 27387
rect 19291 27353 19300 27387
rect 19248 27344 19300 27353
rect 22560 27344 22612 27396
rect 24768 27455 24820 27464
rect 24768 27421 24777 27455
rect 24777 27421 24811 27455
rect 24811 27421 24820 27455
rect 24768 27412 24820 27421
rect 25228 27412 25280 27464
rect 25872 27480 25924 27532
rect 26056 27412 26108 27464
rect 18880 27276 18932 27328
rect 19616 27276 19668 27328
rect 22100 27319 22152 27328
rect 22100 27285 22109 27319
rect 22109 27285 22143 27319
rect 22143 27285 22152 27319
rect 22100 27276 22152 27285
rect 22744 27276 22796 27328
rect 23020 27276 23072 27328
rect 26516 27455 26568 27464
rect 26516 27421 26525 27455
rect 26525 27421 26559 27455
rect 26559 27421 26568 27455
rect 26516 27412 26568 27421
rect 27252 27480 27304 27532
rect 28172 27480 28224 27532
rect 29184 27616 29236 27668
rect 30104 27616 30156 27668
rect 30288 27616 30340 27668
rect 31024 27616 31076 27668
rect 36084 27616 36136 27668
rect 30932 27591 30984 27600
rect 30932 27557 30941 27591
rect 30941 27557 30975 27591
rect 30975 27557 30984 27591
rect 30932 27548 30984 27557
rect 31668 27548 31720 27600
rect 32404 27548 32456 27600
rect 32772 27548 32824 27600
rect 37648 27659 37700 27668
rect 37648 27625 37657 27659
rect 37657 27625 37691 27659
rect 37691 27625 37700 27659
rect 37648 27616 37700 27625
rect 39304 27616 39356 27668
rect 29644 27480 29696 27532
rect 30288 27480 30340 27532
rect 31484 27480 31536 27532
rect 27436 27412 27488 27464
rect 28540 27412 28592 27464
rect 30840 27412 30892 27464
rect 31024 27455 31076 27464
rect 31024 27421 31033 27455
rect 31033 27421 31067 27455
rect 31067 27421 31076 27455
rect 31024 27412 31076 27421
rect 31208 27455 31260 27464
rect 31208 27421 31217 27455
rect 31217 27421 31251 27455
rect 31251 27421 31260 27455
rect 31208 27412 31260 27421
rect 31576 27412 31628 27464
rect 31852 27455 31904 27464
rect 31852 27421 31861 27455
rect 31861 27421 31895 27455
rect 31895 27421 31904 27455
rect 31852 27412 31904 27421
rect 26332 27344 26384 27396
rect 31116 27344 31168 27396
rect 32496 27412 32548 27464
rect 33324 27455 33376 27464
rect 33324 27421 33333 27455
rect 33333 27421 33367 27455
rect 33367 27421 33376 27455
rect 33324 27412 33376 27421
rect 33416 27412 33468 27464
rect 32588 27344 32640 27396
rect 34060 27412 34112 27464
rect 37372 27480 37424 27532
rect 34704 27455 34756 27464
rect 34704 27421 34713 27455
rect 34713 27421 34747 27455
rect 34747 27421 34756 27455
rect 34704 27412 34756 27421
rect 34980 27412 35032 27464
rect 34428 27387 34480 27396
rect 34428 27353 34437 27387
rect 34437 27353 34471 27387
rect 34471 27353 34480 27387
rect 34428 27344 34480 27353
rect 35072 27344 35124 27396
rect 36360 27412 36412 27464
rect 36636 27412 36688 27464
rect 37280 27412 37332 27464
rect 38200 27412 38252 27464
rect 32128 27276 32180 27328
rect 33232 27276 33284 27328
rect 33508 27276 33560 27328
rect 33692 27276 33744 27328
rect 33968 27276 34020 27328
rect 34704 27276 34756 27328
rect 34796 27319 34848 27328
rect 34796 27285 34805 27319
rect 34805 27285 34839 27319
rect 34839 27285 34848 27319
rect 34796 27276 34848 27285
rect 35532 27319 35584 27328
rect 35532 27285 35541 27319
rect 35541 27285 35575 27319
rect 35575 27285 35584 27319
rect 35532 27276 35584 27285
rect 38292 27387 38344 27396
rect 38292 27353 38301 27387
rect 38301 27353 38335 27387
rect 38335 27353 38344 27387
rect 38292 27344 38344 27353
rect 38476 27412 38528 27464
rect 38844 27412 38896 27464
rect 39856 27412 39908 27464
rect 41696 27412 41748 27464
rect 39396 27319 39448 27328
rect 39396 27285 39405 27319
rect 39405 27285 39439 27319
rect 39439 27285 39448 27319
rect 39396 27276 39448 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 5540 27072 5592 27124
rect 6000 27115 6052 27124
rect 6000 27081 6009 27115
rect 6009 27081 6043 27115
rect 6043 27081 6052 27115
rect 6000 27072 6052 27081
rect 7012 27072 7064 27124
rect 3056 27004 3108 27056
rect 3884 27004 3936 27056
rect 5908 27004 5960 27056
rect 6828 27004 6880 27056
rect 7748 27072 7800 27124
rect 7932 27072 7984 27124
rect 8300 27072 8352 27124
rect 8944 27072 8996 27124
rect 9128 27072 9180 27124
rect 9772 27072 9824 27124
rect 9864 27115 9916 27124
rect 9864 27081 9873 27115
rect 9873 27081 9907 27115
rect 9907 27081 9916 27115
rect 9864 27072 9916 27081
rect 10048 27072 10100 27124
rect 12348 27115 12400 27124
rect 12348 27081 12357 27115
rect 12357 27081 12391 27115
rect 12391 27081 12400 27115
rect 12348 27072 12400 27081
rect 12532 27072 12584 27124
rect 12808 27072 12860 27124
rect 12992 27072 13044 27124
rect 1400 26868 1452 26920
rect 1768 26911 1820 26920
rect 1768 26877 1777 26911
rect 1777 26877 1811 26911
rect 1811 26877 1820 26911
rect 1768 26868 1820 26877
rect 6092 26911 6144 26920
rect 6092 26877 6101 26911
rect 6101 26877 6135 26911
rect 6135 26877 6144 26911
rect 6092 26868 6144 26877
rect 7380 26868 7432 26920
rect 2872 26800 2924 26852
rect 7932 26979 7984 26988
rect 7932 26945 7941 26979
rect 7941 26945 7975 26979
rect 7975 26945 7984 26979
rect 7932 26936 7984 26945
rect 8116 26979 8168 26988
rect 8116 26945 8123 26979
rect 8123 26945 8168 26979
rect 8116 26936 8168 26945
rect 8300 26979 8352 26988
rect 8300 26945 8309 26979
rect 8309 26945 8343 26979
rect 8343 26945 8352 26979
rect 8300 26936 8352 26945
rect 8576 26936 8628 26988
rect 8852 26979 8904 26988
rect 8852 26945 8861 26979
rect 8861 26945 8895 26979
rect 8895 26945 8904 26979
rect 8852 26936 8904 26945
rect 9404 26979 9456 26988
rect 9404 26945 9411 26979
rect 9411 26945 9456 26979
rect 2412 26732 2464 26784
rect 3240 26775 3292 26784
rect 3240 26741 3249 26775
rect 3249 26741 3283 26775
rect 3283 26741 3292 26775
rect 3240 26732 3292 26741
rect 3516 26732 3568 26784
rect 4804 26732 4856 26784
rect 7840 26732 7892 26784
rect 8668 26732 8720 26784
rect 9036 26732 9088 26784
rect 9404 26936 9456 26945
rect 10692 27004 10744 27056
rect 11796 27004 11848 27056
rect 12072 27004 12124 27056
rect 9496 26800 9548 26852
rect 9680 26800 9732 26852
rect 9956 26979 10008 26988
rect 9956 26945 9965 26979
rect 9965 26945 9999 26979
rect 9999 26945 10008 26979
rect 9956 26936 10008 26945
rect 10048 26979 10100 26988
rect 10048 26945 10058 26979
rect 10058 26945 10092 26979
rect 10092 26945 10100 26979
rect 10048 26936 10100 26945
rect 10324 26979 10376 26988
rect 10324 26945 10333 26979
rect 10333 26945 10367 26979
rect 10367 26945 10376 26979
rect 10324 26936 10376 26945
rect 12532 26936 12584 26988
rect 14004 27072 14056 27124
rect 14556 27072 14608 27124
rect 14924 27115 14976 27124
rect 14924 27081 14933 27115
rect 14933 27081 14967 27115
rect 14967 27081 14976 27115
rect 14924 27072 14976 27081
rect 15752 27115 15804 27124
rect 15752 27081 15761 27115
rect 15761 27081 15795 27115
rect 15795 27081 15804 27115
rect 15752 27072 15804 27081
rect 15936 27072 15988 27124
rect 13728 27004 13780 27056
rect 11888 26911 11940 26920
rect 11888 26877 11897 26911
rect 11897 26877 11931 26911
rect 11931 26877 11940 26911
rect 11888 26868 11940 26877
rect 12440 26843 12492 26852
rect 12440 26809 12449 26843
rect 12449 26809 12483 26843
rect 12483 26809 12492 26843
rect 12440 26800 12492 26809
rect 13176 26979 13228 26988
rect 13176 26945 13185 26979
rect 13185 26945 13219 26979
rect 13219 26945 13228 26979
rect 13176 26936 13228 26945
rect 13176 26800 13228 26852
rect 13360 26800 13412 26852
rect 10784 26732 10836 26784
rect 13544 26936 13596 26988
rect 13820 26936 13872 26988
rect 14188 26979 14240 26988
rect 14188 26945 14197 26979
rect 14197 26945 14231 26979
rect 14231 26945 14240 26979
rect 14188 26936 14240 26945
rect 14372 26936 14424 26988
rect 14556 26936 14608 26988
rect 14096 26843 14148 26852
rect 14096 26809 14105 26843
rect 14105 26809 14139 26843
rect 14139 26809 14148 26843
rect 14096 26800 14148 26809
rect 15108 26979 15160 26988
rect 15108 26945 15117 26979
rect 15117 26945 15151 26979
rect 15151 26945 15160 26979
rect 15108 26936 15160 26945
rect 15292 26979 15344 26988
rect 15292 26945 15299 26979
rect 15299 26945 15344 26979
rect 15292 26936 15344 26945
rect 15384 26979 15436 26988
rect 15384 26945 15393 26979
rect 15393 26945 15427 26979
rect 15427 26945 15436 26979
rect 15384 26936 15436 26945
rect 15476 26979 15528 26988
rect 15476 26945 15485 26979
rect 15485 26945 15519 26979
rect 15519 26945 15528 26979
rect 15476 26936 15528 26945
rect 15568 26979 15620 26988
rect 16580 27072 16632 27124
rect 17960 27072 18012 27124
rect 15568 26945 15582 26979
rect 15582 26945 15616 26979
rect 15616 26945 15620 26979
rect 15568 26936 15620 26945
rect 13728 26775 13780 26784
rect 13728 26741 13737 26775
rect 13737 26741 13771 26775
rect 13771 26741 13780 26775
rect 13728 26732 13780 26741
rect 13912 26732 13964 26784
rect 15016 26800 15068 26852
rect 15384 26800 15436 26852
rect 16304 26843 16356 26852
rect 16304 26809 16313 26843
rect 16313 26809 16347 26843
rect 16347 26809 16356 26843
rect 16304 26800 16356 26809
rect 17592 26936 17644 26988
rect 19248 27072 19300 27124
rect 22100 27072 22152 27124
rect 22928 27072 22980 27124
rect 23388 27072 23440 27124
rect 23572 27072 23624 27124
rect 18696 26979 18748 26988
rect 18696 26945 18705 26979
rect 18705 26945 18739 26979
rect 18739 26945 18748 26979
rect 19984 27047 20036 27056
rect 19984 27013 19993 27047
rect 19993 27013 20027 27047
rect 20027 27013 20036 27047
rect 19984 27004 20036 27013
rect 20996 27004 21048 27056
rect 18696 26936 18748 26945
rect 19340 26979 19392 26988
rect 19340 26945 19349 26979
rect 19349 26945 19383 26979
rect 19383 26945 19392 26979
rect 19340 26936 19392 26945
rect 18328 26868 18380 26920
rect 22008 26979 22060 26988
rect 22008 26945 22017 26979
rect 22017 26945 22051 26979
rect 22051 26945 22060 26979
rect 22008 26936 22060 26945
rect 22836 26936 22888 26988
rect 28632 27072 28684 27124
rect 26608 27004 26660 27056
rect 29092 27004 29144 27056
rect 19616 26911 19668 26920
rect 19616 26877 19625 26911
rect 19625 26877 19659 26911
rect 19659 26877 19668 26911
rect 19616 26868 19668 26877
rect 21088 26868 21140 26920
rect 14464 26732 14516 26784
rect 16580 26732 16632 26784
rect 19248 26800 19300 26852
rect 25044 26936 25096 26988
rect 25136 26936 25188 26988
rect 26424 26936 26476 26988
rect 23572 26868 23624 26920
rect 24032 26868 24084 26920
rect 24768 26868 24820 26920
rect 28172 26936 28224 26988
rect 28540 26936 28592 26988
rect 30840 27072 30892 27124
rect 31116 27115 31168 27124
rect 31116 27081 31125 27115
rect 31125 27081 31159 27115
rect 31159 27081 31168 27115
rect 31116 27072 31168 27081
rect 31760 27072 31812 27124
rect 33416 27072 33468 27124
rect 33784 27072 33836 27124
rect 34888 27072 34940 27124
rect 31208 26936 31260 26988
rect 32036 26936 32088 26988
rect 32404 26936 32456 26988
rect 27160 26868 27212 26920
rect 28080 26868 28132 26920
rect 29828 26868 29880 26920
rect 30288 26868 30340 26920
rect 31668 26911 31720 26920
rect 31668 26877 31677 26911
rect 31677 26877 31711 26911
rect 31711 26877 31720 26911
rect 31668 26868 31720 26877
rect 32588 26868 32640 26920
rect 33324 26936 33376 26988
rect 33876 26979 33928 26988
rect 33876 26945 33885 26979
rect 33885 26945 33919 26979
rect 33919 26945 33928 26979
rect 33876 26936 33928 26945
rect 34244 26936 34296 26988
rect 34980 27004 35032 27056
rect 36084 27004 36136 27056
rect 36636 27004 36688 27056
rect 33692 26868 33744 26920
rect 35808 26936 35860 26988
rect 36452 26936 36504 26988
rect 37004 26936 37056 26988
rect 37372 26936 37424 26988
rect 37832 26936 37884 26988
rect 38292 27004 38344 27056
rect 39396 27072 39448 27124
rect 39488 27072 39540 27124
rect 40040 27004 40092 27056
rect 38108 26936 38160 26988
rect 27344 26843 27396 26852
rect 18880 26775 18932 26784
rect 18880 26741 18889 26775
rect 18889 26741 18923 26775
rect 18923 26741 18932 26775
rect 18880 26732 18932 26741
rect 20168 26732 20220 26784
rect 22100 26732 22152 26784
rect 22744 26732 22796 26784
rect 23204 26732 23256 26784
rect 24032 26775 24084 26784
rect 24032 26741 24041 26775
rect 24041 26741 24075 26775
rect 24075 26741 24084 26775
rect 24032 26732 24084 26741
rect 24216 26732 24268 26784
rect 24584 26732 24636 26784
rect 25136 26732 25188 26784
rect 27344 26809 27353 26843
rect 27353 26809 27387 26843
rect 27387 26809 27396 26843
rect 27344 26800 27396 26809
rect 26056 26732 26108 26784
rect 29276 26775 29328 26784
rect 29276 26741 29285 26775
rect 29285 26741 29319 26775
rect 29319 26741 29328 26775
rect 29276 26732 29328 26741
rect 29460 26732 29512 26784
rect 34428 26775 34480 26784
rect 34428 26741 34437 26775
rect 34437 26741 34471 26775
rect 34471 26741 34480 26775
rect 34428 26732 34480 26741
rect 34704 26800 34756 26852
rect 36544 26732 36596 26784
rect 37648 26732 37700 26784
rect 38844 26732 38896 26784
rect 39304 26732 39356 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 1768 26528 1820 26580
rect 5540 26571 5592 26580
rect 5540 26537 5549 26571
rect 5549 26537 5583 26571
rect 5583 26537 5592 26571
rect 5540 26528 5592 26537
rect 8852 26528 8904 26580
rect 6552 26460 6604 26512
rect 8300 26460 8352 26512
rect 8760 26460 8812 26512
rect 9680 26528 9732 26580
rect 3424 26435 3476 26444
rect 3424 26401 3433 26435
rect 3433 26401 3467 26435
rect 3467 26401 3476 26435
rect 3424 26392 3476 26401
rect 3240 26324 3292 26376
rect 4620 26392 4672 26444
rect 3792 26367 3844 26376
rect 3792 26333 3801 26367
rect 3801 26333 3835 26367
rect 3835 26333 3844 26367
rect 3792 26324 3844 26333
rect 3516 26256 3568 26308
rect 3976 26256 4028 26308
rect 3884 26188 3936 26240
rect 5816 26256 5868 26308
rect 8024 26367 8076 26376
rect 8024 26333 8031 26367
rect 8031 26333 8076 26367
rect 6368 26299 6420 26308
rect 6368 26265 6377 26299
rect 6377 26265 6411 26299
rect 6411 26265 6420 26299
rect 6368 26256 6420 26265
rect 6828 26256 6880 26308
rect 7012 26256 7064 26308
rect 8024 26324 8076 26333
rect 8576 26324 8628 26376
rect 7104 26188 7156 26240
rect 8944 26367 8996 26376
rect 8944 26333 8953 26367
rect 8953 26333 8987 26367
rect 8987 26333 8996 26367
rect 8944 26324 8996 26333
rect 9128 26367 9180 26376
rect 9128 26333 9135 26367
rect 9135 26333 9180 26367
rect 9128 26324 9180 26333
rect 10692 26528 10744 26580
rect 11336 26528 11388 26580
rect 9312 26299 9364 26308
rect 9312 26265 9321 26299
rect 9321 26265 9355 26299
rect 9355 26265 9364 26299
rect 9312 26256 9364 26265
rect 10968 26392 11020 26444
rect 10048 26256 10100 26308
rect 10416 26256 10468 26308
rect 9404 26188 9456 26240
rect 10692 26231 10744 26240
rect 10692 26197 10701 26231
rect 10701 26197 10735 26231
rect 10735 26197 10744 26231
rect 10692 26188 10744 26197
rect 11244 26367 11296 26376
rect 11244 26333 11253 26367
rect 11253 26333 11287 26367
rect 11287 26333 11296 26367
rect 11244 26324 11296 26333
rect 11428 26367 11480 26376
rect 11428 26333 11435 26367
rect 11435 26333 11480 26367
rect 11428 26324 11480 26333
rect 11520 26367 11572 26376
rect 11520 26333 11529 26367
rect 11529 26333 11563 26367
rect 11563 26333 11572 26367
rect 11520 26324 11572 26333
rect 11888 26571 11940 26580
rect 11888 26537 11897 26571
rect 11897 26537 11931 26571
rect 11931 26537 11940 26571
rect 11888 26528 11940 26537
rect 12440 26528 12492 26580
rect 13636 26528 13688 26580
rect 14464 26528 14516 26580
rect 16488 26528 16540 26580
rect 16672 26571 16724 26580
rect 16672 26537 16681 26571
rect 16681 26537 16715 26571
rect 16715 26537 16724 26571
rect 16672 26528 16724 26537
rect 16764 26528 16816 26580
rect 18880 26528 18932 26580
rect 19340 26571 19392 26580
rect 19340 26537 19349 26571
rect 19349 26537 19383 26571
rect 19383 26537 19392 26571
rect 19340 26528 19392 26537
rect 19432 26528 19484 26580
rect 11796 26324 11848 26376
rect 12532 26460 12584 26512
rect 14280 26392 14332 26444
rect 12624 26324 12676 26376
rect 12532 26256 12584 26308
rect 13268 26367 13320 26376
rect 13268 26333 13277 26367
rect 13277 26333 13311 26367
rect 13311 26333 13320 26367
rect 13268 26324 13320 26333
rect 13452 26324 13504 26376
rect 13544 26324 13596 26376
rect 16212 26324 16264 26376
rect 17040 26460 17092 26512
rect 19156 26460 19208 26512
rect 19616 26460 19668 26512
rect 20076 26528 20128 26580
rect 20352 26528 20404 26580
rect 20628 26528 20680 26580
rect 13912 26256 13964 26308
rect 14648 26256 14700 26308
rect 18144 26367 18196 26376
rect 18144 26333 18155 26367
rect 18155 26333 18189 26367
rect 18189 26333 18196 26367
rect 20444 26392 20496 26444
rect 20628 26392 20680 26444
rect 18144 26324 18196 26333
rect 18328 26367 18380 26376
rect 18328 26333 18337 26367
rect 18337 26333 18371 26367
rect 18371 26333 18380 26367
rect 18328 26324 18380 26333
rect 17592 26256 17644 26308
rect 12348 26188 12400 26240
rect 14924 26188 14976 26240
rect 15200 26188 15252 26240
rect 18236 26299 18288 26308
rect 18236 26265 18245 26299
rect 18245 26265 18279 26299
rect 18279 26265 18288 26299
rect 18236 26256 18288 26265
rect 18696 26324 18748 26376
rect 18880 26324 18932 26376
rect 19432 26324 19484 26376
rect 21548 26324 21600 26376
rect 21732 26367 21784 26376
rect 21732 26333 21741 26367
rect 21741 26333 21775 26367
rect 21775 26333 21784 26367
rect 21732 26324 21784 26333
rect 22744 26528 22796 26580
rect 22100 26460 22152 26512
rect 23664 26528 23716 26580
rect 23756 26528 23808 26580
rect 24032 26528 24084 26580
rect 24400 26528 24452 26580
rect 24584 26528 24636 26580
rect 25044 26528 25096 26580
rect 25320 26571 25372 26580
rect 25320 26537 25329 26571
rect 25329 26537 25363 26571
rect 25363 26537 25372 26571
rect 25320 26528 25372 26537
rect 26424 26528 26476 26580
rect 27804 26528 27856 26580
rect 28816 26528 28868 26580
rect 29368 26528 29420 26580
rect 30012 26571 30064 26580
rect 30012 26537 30021 26571
rect 30021 26537 30055 26571
rect 30055 26537 30064 26571
rect 30012 26528 30064 26537
rect 31668 26528 31720 26580
rect 22192 26367 22244 26376
rect 22192 26333 22201 26367
rect 22201 26333 22235 26367
rect 22235 26333 22244 26367
rect 22192 26324 22244 26333
rect 18880 26188 18932 26240
rect 19064 26188 19116 26240
rect 20904 26188 20956 26240
rect 21732 26188 21784 26240
rect 24216 26460 24268 26512
rect 23388 26392 23440 26444
rect 22744 26367 22796 26376
rect 22744 26333 22753 26367
rect 22753 26333 22787 26367
rect 22787 26333 22796 26367
rect 22744 26324 22796 26333
rect 23664 26324 23716 26376
rect 23756 26367 23808 26376
rect 23756 26333 23765 26367
rect 23765 26333 23799 26367
rect 23799 26333 23808 26367
rect 23756 26324 23808 26333
rect 24308 26324 24360 26376
rect 24768 26367 24820 26376
rect 24768 26333 24777 26367
rect 24777 26333 24811 26367
rect 24811 26333 24820 26367
rect 24768 26324 24820 26333
rect 24952 26324 25004 26376
rect 25136 26367 25188 26376
rect 25136 26333 25145 26367
rect 25145 26333 25179 26367
rect 25179 26333 25188 26367
rect 25136 26324 25188 26333
rect 25228 26367 25280 26376
rect 25228 26333 25237 26367
rect 25237 26333 25271 26367
rect 25271 26333 25280 26367
rect 25228 26324 25280 26333
rect 26148 26392 26200 26444
rect 26332 26367 26384 26376
rect 26332 26333 26341 26367
rect 26341 26333 26375 26367
rect 26375 26333 26384 26367
rect 26332 26324 26384 26333
rect 26700 26367 26752 26376
rect 26700 26333 26712 26367
rect 26712 26333 26746 26367
rect 26746 26333 26752 26367
rect 28908 26392 28960 26444
rect 26700 26324 26752 26333
rect 26976 26367 27028 26376
rect 26976 26333 26985 26367
rect 26985 26333 27019 26367
rect 27019 26333 27028 26367
rect 26976 26324 27028 26333
rect 27528 26367 27580 26376
rect 27528 26333 27537 26367
rect 27537 26333 27571 26367
rect 27571 26333 27580 26367
rect 27528 26324 27580 26333
rect 22100 26188 22152 26240
rect 22376 26188 22428 26240
rect 23940 26188 23992 26240
rect 24584 26188 24636 26240
rect 24768 26188 24820 26240
rect 25596 26256 25648 26308
rect 27804 26367 27856 26376
rect 27804 26333 27813 26367
rect 27813 26333 27847 26367
rect 27847 26333 27856 26367
rect 27804 26324 27856 26333
rect 30748 26460 30800 26512
rect 32036 26571 32088 26580
rect 32036 26537 32045 26571
rect 32045 26537 32079 26571
rect 32079 26537 32088 26571
rect 32036 26528 32088 26537
rect 33048 26528 33100 26580
rect 29276 26392 29328 26444
rect 29644 26435 29696 26444
rect 29644 26401 29653 26435
rect 29653 26401 29687 26435
rect 29687 26401 29696 26435
rect 29644 26392 29696 26401
rect 28632 26256 28684 26308
rect 29368 26299 29420 26308
rect 29368 26265 29377 26299
rect 29377 26265 29411 26299
rect 29411 26265 29420 26299
rect 29368 26256 29420 26265
rect 30472 26324 30524 26376
rect 32128 26392 32180 26444
rect 30840 26324 30892 26376
rect 31024 26324 31076 26376
rect 32036 26324 32088 26376
rect 32588 26324 32640 26376
rect 33508 26503 33560 26512
rect 33508 26469 33517 26503
rect 33517 26469 33551 26503
rect 33551 26469 33560 26503
rect 33508 26460 33560 26469
rect 32772 26324 32824 26376
rect 33232 26367 33284 26376
rect 33232 26333 33241 26367
rect 33241 26333 33275 26367
rect 33275 26333 33284 26367
rect 33232 26324 33284 26333
rect 33508 26324 33560 26376
rect 34060 26324 34112 26376
rect 37372 26528 37424 26580
rect 37556 26528 37608 26580
rect 38292 26528 38344 26580
rect 36544 26460 36596 26512
rect 34244 26392 34296 26444
rect 35992 26324 36044 26376
rect 36084 26367 36136 26376
rect 36084 26333 36093 26367
rect 36093 26333 36127 26367
rect 36127 26333 36136 26367
rect 36084 26324 36136 26333
rect 25964 26231 26016 26240
rect 25964 26197 25973 26231
rect 25973 26197 26007 26231
rect 26007 26197 26016 26231
rect 25964 26188 26016 26197
rect 27068 26188 27120 26240
rect 27344 26231 27396 26240
rect 27344 26197 27353 26231
rect 27353 26197 27387 26231
rect 27387 26197 27396 26231
rect 27344 26188 27396 26197
rect 27620 26188 27672 26240
rect 27896 26188 27948 26240
rect 27988 26188 28040 26240
rect 28448 26188 28500 26240
rect 29276 26188 29328 26240
rect 31760 26188 31812 26240
rect 32128 26188 32180 26240
rect 33692 26188 33744 26240
rect 37096 26256 37148 26308
rect 39212 26188 39264 26240
rect 39764 26256 39816 26308
rect 39948 26256 40000 26308
rect 40684 26299 40736 26308
rect 40684 26265 40693 26299
rect 40693 26265 40727 26299
rect 40727 26265 40736 26299
rect 40684 26256 40736 26265
rect 40500 26188 40552 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 5540 25984 5592 26036
rect 8944 25984 8996 26036
rect 11244 25984 11296 26036
rect 11520 25984 11572 26036
rect 12808 25984 12860 26036
rect 20444 25984 20496 26036
rect 2412 25916 2464 25968
rect 3792 25959 3844 25968
rect 3792 25925 3801 25959
rect 3801 25925 3835 25959
rect 3835 25925 3844 25959
rect 3792 25916 3844 25925
rect 2964 25891 3016 25900
rect 2964 25857 2973 25891
rect 2973 25857 3007 25891
rect 3007 25857 3016 25891
rect 2964 25848 3016 25857
rect 5448 25848 5500 25900
rect 9312 25916 9364 25968
rect 9588 25916 9640 25968
rect 13176 25916 13228 25968
rect 14096 25916 14148 25968
rect 18236 25916 18288 25968
rect 19156 25916 19208 25968
rect 20260 25916 20312 25968
rect 6920 25848 6972 25900
rect 3424 25712 3476 25764
rect 3884 25712 3936 25764
rect 6368 25780 6420 25832
rect 7104 25780 7156 25832
rect 7564 25780 7616 25832
rect 8116 25891 8168 25900
rect 8116 25857 8125 25891
rect 8125 25857 8159 25891
rect 8159 25857 8168 25891
rect 8116 25848 8168 25857
rect 9036 25848 9088 25900
rect 10416 25891 10468 25900
rect 10416 25857 10425 25891
rect 10425 25857 10459 25891
rect 10459 25857 10468 25891
rect 10416 25848 10468 25857
rect 8576 25780 8628 25832
rect 9588 25780 9640 25832
rect 10784 25891 10836 25900
rect 10784 25857 10793 25891
rect 10793 25857 10827 25891
rect 10827 25857 10836 25891
rect 10784 25848 10836 25857
rect 11612 25848 11664 25900
rect 13636 25848 13688 25900
rect 15200 25891 15252 25900
rect 15200 25857 15209 25891
rect 15209 25857 15243 25891
rect 15243 25857 15252 25891
rect 15200 25848 15252 25857
rect 16948 25891 17000 25900
rect 16948 25857 16957 25891
rect 16957 25857 16991 25891
rect 16991 25857 17000 25891
rect 16948 25848 17000 25857
rect 17592 25848 17644 25900
rect 19432 25891 19484 25900
rect 19432 25857 19441 25891
rect 19441 25857 19475 25891
rect 19475 25857 19484 25891
rect 19432 25848 19484 25857
rect 20076 25848 20128 25900
rect 19340 25780 19392 25832
rect 9220 25712 9272 25764
rect 20904 25848 20956 25900
rect 22008 25984 22060 26036
rect 22100 25984 22152 26036
rect 23572 25984 23624 26036
rect 23756 25984 23808 26036
rect 22284 25916 22336 25968
rect 22008 25780 22060 25832
rect 27436 25984 27488 26036
rect 28632 26027 28684 26036
rect 28632 25993 28641 26027
rect 28641 25993 28675 26027
rect 28675 25993 28684 26027
rect 28632 25984 28684 25993
rect 28724 25984 28776 26036
rect 26608 25916 26660 25968
rect 25412 25891 25464 25900
rect 25412 25857 25421 25891
rect 25421 25857 25455 25891
rect 25455 25857 25464 25891
rect 25412 25848 25464 25857
rect 25964 25848 26016 25900
rect 26056 25891 26108 25900
rect 26056 25857 26065 25891
rect 26065 25857 26099 25891
rect 26099 25857 26108 25891
rect 26056 25848 26108 25857
rect 26240 25891 26292 25900
rect 26240 25857 26249 25891
rect 26249 25857 26283 25891
rect 26283 25857 26292 25891
rect 26240 25848 26292 25857
rect 26884 25848 26936 25900
rect 27252 25916 27304 25968
rect 32036 25984 32088 26036
rect 34244 25984 34296 26036
rect 34336 25984 34388 26036
rect 27068 25848 27120 25900
rect 27344 25848 27396 25900
rect 35072 25916 35124 25968
rect 35532 25984 35584 26036
rect 37464 25984 37516 26036
rect 37740 25984 37792 26036
rect 39764 25984 39816 26036
rect 23020 25712 23072 25764
rect 24952 25712 25004 25764
rect 25872 25780 25924 25832
rect 4068 25644 4120 25696
rect 7196 25644 7248 25696
rect 9864 25644 9916 25696
rect 11796 25644 11848 25696
rect 15016 25687 15068 25696
rect 15016 25653 15025 25687
rect 15025 25653 15059 25687
rect 15059 25653 15068 25687
rect 15016 25644 15068 25653
rect 15752 25644 15804 25696
rect 18880 25644 18932 25696
rect 19340 25644 19392 25696
rect 20720 25644 20772 25696
rect 20996 25644 21048 25696
rect 21548 25644 21600 25696
rect 26056 25712 26108 25764
rect 27620 25780 27672 25832
rect 28448 25891 28500 25900
rect 28448 25857 28457 25891
rect 28457 25857 28491 25891
rect 28491 25857 28500 25891
rect 28448 25848 28500 25857
rect 29368 25891 29420 25900
rect 29368 25857 29377 25891
rect 29377 25857 29411 25891
rect 29411 25857 29420 25891
rect 29368 25848 29420 25857
rect 29920 25891 29972 25900
rect 29920 25857 29929 25891
rect 29929 25857 29963 25891
rect 29963 25857 29972 25891
rect 29920 25848 29972 25857
rect 30196 25891 30248 25900
rect 30196 25857 30205 25891
rect 30205 25857 30239 25891
rect 30239 25857 30248 25891
rect 30196 25848 30248 25857
rect 30564 25848 30616 25900
rect 31116 25848 31168 25900
rect 32036 25848 32088 25900
rect 33416 25848 33468 25900
rect 30380 25823 30432 25832
rect 30380 25789 30389 25823
rect 30389 25789 30423 25823
rect 30423 25789 30432 25823
rect 30380 25780 30432 25789
rect 33232 25780 33284 25832
rect 34796 25780 34848 25832
rect 35348 25780 35400 25832
rect 35808 25848 35860 25900
rect 37464 25848 37516 25900
rect 39212 25916 39264 25968
rect 40040 25916 40092 25968
rect 37832 25848 37884 25900
rect 38292 25848 38344 25900
rect 36084 25780 36136 25832
rect 39304 25823 39356 25832
rect 39304 25789 39313 25823
rect 39313 25789 39347 25823
rect 39347 25789 39356 25823
rect 39304 25780 39356 25789
rect 39580 25823 39632 25832
rect 39580 25789 39589 25823
rect 39589 25789 39623 25823
rect 39623 25789 39632 25823
rect 39580 25780 39632 25789
rect 35808 25712 35860 25764
rect 27436 25687 27488 25696
rect 27436 25653 27445 25687
rect 27445 25653 27479 25687
rect 27479 25653 27488 25687
rect 27436 25644 27488 25653
rect 27804 25687 27856 25696
rect 27804 25653 27813 25687
rect 27813 25653 27847 25687
rect 27847 25653 27856 25687
rect 27804 25644 27856 25653
rect 34796 25644 34848 25696
rect 36084 25644 36136 25696
rect 38292 25687 38344 25696
rect 38292 25653 38301 25687
rect 38301 25653 38335 25687
rect 38335 25653 38344 25687
rect 38292 25644 38344 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 3976 25440 4028 25492
rect 4068 25440 4120 25492
rect 5724 25440 5776 25492
rect 2412 25304 2464 25356
rect 3056 25236 3108 25288
rect 7380 25440 7432 25492
rect 7196 25347 7248 25356
rect 7196 25313 7205 25347
rect 7205 25313 7239 25347
rect 7239 25313 7248 25347
rect 7196 25304 7248 25313
rect 7564 25372 7616 25424
rect 9956 25440 10008 25492
rect 11888 25440 11940 25492
rect 13452 25440 13504 25492
rect 20260 25440 20312 25492
rect 20812 25440 20864 25492
rect 20904 25440 20956 25492
rect 11796 25415 11848 25424
rect 11796 25381 11805 25415
rect 11805 25381 11839 25415
rect 11839 25381 11848 25415
rect 11796 25372 11848 25381
rect 13912 25372 13964 25424
rect 14096 25372 14148 25424
rect 1676 25211 1728 25220
rect 1676 25177 1685 25211
rect 1685 25177 1719 25211
rect 1719 25177 1728 25211
rect 1676 25168 1728 25177
rect 7472 25236 7524 25288
rect 7288 25168 7340 25220
rect 3148 25143 3200 25152
rect 3148 25109 3157 25143
rect 3157 25109 3191 25143
rect 3191 25109 3200 25143
rect 3148 25100 3200 25109
rect 4068 25100 4120 25152
rect 6644 25143 6696 25152
rect 6644 25109 6653 25143
rect 6653 25109 6687 25143
rect 6687 25109 6696 25143
rect 6644 25100 6696 25109
rect 7472 25100 7524 25152
rect 9220 25279 9272 25288
rect 9220 25245 9229 25279
rect 9229 25245 9263 25279
rect 9263 25245 9272 25279
rect 9220 25236 9272 25245
rect 9404 25279 9456 25288
rect 9404 25245 9413 25279
rect 9413 25245 9447 25279
rect 9447 25245 9456 25279
rect 9404 25236 9456 25245
rect 9588 25279 9640 25288
rect 9588 25245 9597 25279
rect 9597 25245 9631 25279
rect 9631 25245 9640 25279
rect 9588 25236 9640 25245
rect 9772 25236 9824 25288
rect 10508 25279 10560 25288
rect 10508 25245 10517 25279
rect 10517 25245 10551 25279
rect 10551 25245 10560 25279
rect 10508 25236 10560 25245
rect 10784 25347 10836 25356
rect 10784 25313 10793 25347
rect 10793 25313 10827 25347
rect 10827 25313 10836 25347
rect 10784 25304 10836 25313
rect 11152 25304 11204 25356
rect 13544 25304 13596 25356
rect 14740 25347 14792 25356
rect 14740 25313 14749 25347
rect 14749 25313 14783 25347
rect 14783 25313 14792 25347
rect 14740 25304 14792 25313
rect 15016 25347 15068 25356
rect 15016 25313 15025 25347
rect 15025 25313 15059 25347
rect 15059 25313 15068 25347
rect 15016 25304 15068 25313
rect 9036 25168 9088 25220
rect 10232 25168 10284 25220
rect 11888 25236 11940 25288
rect 12072 25279 12124 25288
rect 12072 25245 12081 25279
rect 12081 25245 12115 25279
rect 12115 25245 12124 25279
rect 12072 25236 12124 25245
rect 12164 25279 12216 25288
rect 12164 25245 12173 25279
rect 12173 25245 12207 25279
rect 12207 25245 12216 25279
rect 12164 25236 12216 25245
rect 12348 25236 12400 25288
rect 12532 25236 12584 25288
rect 17132 25236 17184 25288
rect 19064 25304 19116 25356
rect 20444 25304 20496 25356
rect 20904 25304 20956 25356
rect 22560 25372 22612 25424
rect 25504 25440 25556 25492
rect 27804 25440 27856 25492
rect 29644 25440 29696 25492
rect 29920 25440 29972 25492
rect 31484 25483 31536 25492
rect 31484 25449 31493 25483
rect 31493 25449 31527 25483
rect 31527 25449 31536 25483
rect 31484 25440 31536 25449
rect 32128 25440 32180 25492
rect 32772 25483 32824 25492
rect 32772 25449 32781 25483
rect 32781 25449 32815 25483
rect 32815 25449 32824 25483
rect 32772 25440 32824 25449
rect 18052 25279 18104 25288
rect 18052 25245 18061 25279
rect 18061 25245 18095 25279
rect 18095 25245 18104 25279
rect 18052 25236 18104 25245
rect 19248 25236 19300 25288
rect 19984 25279 20036 25288
rect 19984 25245 19993 25279
rect 19993 25245 20027 25279
rect 20027 25245 20036 25279
rect 19984 25236 20036 25245
rect 11520 25100 11572 25152
rect 13544 25100 13596 25152
rect 16672 25211 16724 25220
rect 16672 25177 16681 25211
rect 16681 25177 16715 25211
rect 16715 25177 16724 25211
rect 16672 25168 16724 25177
rect 18512 25168 18564 25220
rect 20996 25236 21048 25288
rect 21824 25347 21876 25356
rect 21824 25313 21833 25347
rect 21833 25313 21867 25347
rect 21867 25313 21876 25347
rect 21824 25304 21876 25313
rect 15660 25100 15712 25152
rect 18144 25100 18196 25152
rect 20076 25100 20128 25152
rect 21548 25168 21600 25220
rect 22100 25236 22152 25288
rect 22744 25236 22796 25288
rect 25136 25279 25188 25288
rect 25136 25245 25145 25279
rect 25145 25245 25179 25279
rect 25179 25245 25188 25279
rect 25136 25236 25188 25245
rect 22008 25168 22060 25220
rect 23388 25168 23440 25220
rect 24492 25168 24544 25220
rect 22192 25100 22244 25152
rect 24952 25100 25004 25152
rect 25320 25236 25372 25288
rect 26976 25100 27028 25152
rect 27528 25304 27580 25356
rect 28724 25304 28776 25356
rect 27620 25279 27672 25288
rect 27620 25245 27629 25279
rect 27629 25245 27663 25279
rect 27663 25245 27672 25279
rect 27620 25236 27672 25245
rect 28908 25236 28960 25288
rect 29644 25236 29696 25288
rect 32496 25372 32548 25424
rect 34796 25440 34848 25492
rect 33968 25372 34020 25424
rect 27896 25168 27948 25220
rect 29920 25279 29972 25288
rect 29920 25245 29929 25279
rect 29929 25245 29963 25279
rect 29963 25245 29972 25279
rect 29920 25236 29972 25245
rect 30012 25279 30064 25288
rect 30012 25245 30021 25279
rect 30021 25245 30055 25279
rect 30055 25245 30064 25279
rect 30012 25236 30064 25245
rect 30380 25236 30432 25288
rect 30656 25279 30708 25288
rect 30656 25245 30665 25279
rect 30665 25245 30699 25279
rect 30699 25245 30708 25279
rect 30656 25236 30708 25245
rect 30840 25236 30892 25288
rect 33600 25304 33652 25356
rect 34244 25304 34296 25356
rect 30288 25168 30340 25220
rect 32036 25236 32088 25288
rect 32404 25236 32456 25288
rect 32680 25236 32732 25288
rect 32956 25279 33008 25288
rect 32956 25245 32965 25279
rect 32965 25245 32999 25279
rect 32999 25245 33008 25279
rect 32956 25236 33008 25245
rect 27804 25100 27856 25152
rect 31760 25168 31812 25220
rect 32496 25100 32548 25152
rect 32956 25100 33008 25152
rect 33324 25236 33376 25288
rect 34152 25279 34204 25288
rect 34152 25245 34161 25279
rect 34161 25245 34195 25279
rect 34195 25245 34204 25279
rect 36728 25440 36780 25492
rect 37556 25372 37608 25424
rect 37832 25483 37884 25492
rect 37832 25449 37841 25483
rect 37841 25449 37875 25483
rect 37875 25449 37884 25483
rect 37832 25440 37884 25449
rect 39580 25440 39632 25492
rect 40132 25440 40184 25492
rect 35808 25347 35860 25356
rect 35808 25313 35817 25347
rect 35817 25313 35851 25347
rect 35851 25313 35860 25347
rect 35808 25304 35860 25313
rect 34152 25236 34204 25245
rect 33600 25168 33652 25220
rect 36084 25279 36136 25288
rect 36084 25245 36087 25279
rect 36087 25245 36121 25279
rect 36121 25245 36136 25279
rect 36084 25236 36136 25245
rect 37004 25279 37056 25288
rect 37004 25245 37013 25279
rect 37013 25245 37047 25279
rect 37047 25245 37056 25279
rect 37004 25236 37056 25245
rect 37096 25236 37148 25288
rect 37372 25236 37424 25288
rect 38292 25304 38344 25356
rect 39764 25236 39816 25288
rect 40040 25279 40092 25288
rect 40040 25245 40049 25279
rect 40049 25245 40083 25279
rect 40083 25245 40092 25279
rect 40040 25236 40092 25245
rect 40500 25168 40552 25220
rect 36176 25100 36228 25152
rect 37096 25143 37148 25152
rect 37096 25109 37105 25143
rect 37105 25109 37139 25143
rect 37139 25109 37148 25143
rect 37096 25100 37148 25109
rect 37740 25100 37792 25152
rect 38108 25143 38160 25152
rect 38108 25109 38117 25143
rect 38117 25109 38151 25143
rect 38151 25109 38160 25143
rect 38108 25100 38160 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 1676 24896 1728 24948
rect 2872 24939 2924 24948
rect 2872 24905 2881 24939
rect 2881 24905 2915 24939
rect 2915 24905 2924 24939
rect 2872 24896 2924 24905
rect 3148 24896 3200 24948
rect 3976 24760 4028 24812
rect 5080 24896 5132 24948
rect 5632 24896 5684 24948
rect 5816 24939 5868 24948
rect 5816 24905 5825 24939
rect 5825 24905 5859 24939
rect 5859 24905 5868 24939
rect 5816 24896 5868 24905
rect 6644 24896 6696 24948
rect 7472 24896 7524 24948
rect 8116 24939 8168 24948
rect 8116 24905 8125 24939
rect 8125 24905 8159 24939
rect 8159 24905 8168 24939
rect 8116 24896 8168 24905
rect 3884 24692 3936 24744
rect 5080 24760 5132 24812
rect 5172 24760 5224 24812
rect 5540 24803 5592 24812
rect 5540 24769 5549 24803
rect 5549 24769 5583 24803
rect 5583 24769 5592 24803
rect 5540 24760 5592 24769
rect 5264 24735 5316 24744
rect 5264 24701 5273 24735
rect 5273 24701 5307 24735
rect 5307 24701 5316 24735
rect 5264 24692 5316 24701
rect 5632 24692 5684 24744
rect 7104 24828 7156 24880
rect 8024 24828 8076 24880
rect 9680 24896 9732 24948
rect 9772 24939 9824 24948
rect 9772 24905 9781 24939
rect 9781 24905 9815 24939
rect 9815 24905 9824 24939
rect 9772 24896 9824 24905
rect 12072 24896 12124 24948
rect 12256 24896 12308 24948
rect 13912 24896 13964 24948
rect 14832 24896 14884 24948
rect 15200 24896 15252 24948
rect 6368 24803 6420 24812
rect 6368 24769 6377 24803
rect 6377 24769 6411 24803
rect 6411 24769 6420 24803
rect 6368 24760 6420 24769
rect 8208 24803 8260 24812
rect 8208 24769 8217 24803
rect 8217 24769 8251 24803
rect 8251 24769 8260 24803
rect 8208 24760 8260 24769
rect 8300 24760 8352 24812
rect 8760 24760 8812 24812
rect 5908 24735 5960 24744
rect 5908 24701 5917 24735
rect 5917 24701 5951 24735
rect 5951 24701 5960 24735
rect 5908 24692 5960 24701
rect 4620 24624 4672 24676
rect 5172 24624 5224 24676
rect 12348 24828 12400 24880
rect 12808 24828 12860 24880
rect 10232 24760 10284 24812
rect 11152 24760 11204 24812
rect 9312 24735 9364 24744
rect 9312 24701 9321 24735
rect 9321 24701 9355 24735
rect 9355 24701 9364 24735
rect 9312 24692 9364 24701
rect 9220 24624 9272 24676
rect 8852 24599 8904 24608
rect 8852 24565 8861 24599
rect 8861 24565 8895 24599
rect 8895 24565 8904 24599
rect 8852 24556 8904 24565
rect 11980 24556 12032 24608
rect 12808 24556 12860 24608
rect 13268 24803 13320 24812
rect 13268 24769 13277 24803
rect 13277 24769 13311 24803
rect 13311 24769 13320 24803
rect 13268 24760 13320 24769
rect 13636 24828 13688 24880
rect 14280 24828 14332 24880
rect 14372 24828 14424 24880
rect 15660 24828 15712 24880
rect 13820 24803 13872 24812
rect 13820 24769 13829 24803
rect 13829 24769 13863 24803
rect 13863 24769 13872 24803
rect 13820 24760 13872 24769
rect 14464 24803 14516 24812
rect 14464 24769 14473 24803
rect 14473 24769 14507 24803
rect 14507 24769 14516 24803
rect 14464 24760 14516 24769
rect 14648 24803 14700 24812
rect 14648 24769 14657 24803
rect 14657 24769 14691 24803
rect 14691 24769 14700 24803
rect 14648 24760 14700 24769
rect 14740 24803 14792 24812
rect 14740 24769 14749 24803
rect 14749 24769 14783 24803
rect 14783 24769 14792 24803
rect 14740 24760 14792 24769
rect 13176 24624 13228 24676
rect 13268 24556 13320 24608
rect 13636 24624 13688 24676
rect 17040 24760 17092 24812
rect 19064 24896 19116 24948
rect 19248 24896 19300 24948
rect 22008 24939 22060 24948
rect 22008 24905 22017 24939
rect 22017 24905 22051 24939
rect 22051 24905 22060 24939
rect 22008 24896 22060 24905
rect 18052 24828 18104 24880
rect 15568 24692 15620 24744
rect 15752 24735 15804 24744
rect 15752 24701 15761 24735
rect 15761 24701 15795 24735
rect 15795 24701 15804 24735
rect 15752 24692 15804 24701
rect 15108 24556 15160 24608
rect 15476 24556 15528 24608
rect 17040 24556 17092 24608
rect 17316 24599 17368 24608
rect 17316 24565 17325 24599
rect 17325 24565 17359 24599
rect 17359 24565 17368 24599
rect 17316 24556 17368 24565
rect 17776 24624 17828 24676
rect 19248 24803 19300 24812
rect 19248 24769 19257 24803
rect 19257 24769 19291 24803
rect 19291 24769 19300 24803
rect 19248 24760 19300 24769
rect 19616 24828 19668 24880
rect 20260 24760 20312 24812
rect 20812 24760 20864 24812
rect 18512 24556 18564 24608
rect 18604 24599 18656 24608
rect 18604 24565 18613 24599
rect 18613 24565 18647 24599
rect 18647 24565 18656 24599
rect 18604 24556 18656 24565
rect 19800 24556 19852 24608
rect 21824 24871 21876 24880
rect 21824 24837 21833 24871
rect 21833 24837 21867 24871
rect 21867 24837 21876 24871
rect 21824 24828 21876 24837
rect 22100 24871 22152 24880
rect 22100 24837 22109 24871
rect 22109 24837 22143 24871
rect 22143 24837 22152 24871
rect 22100 24828 22152 24837
rect 22192 24871 22244 24880
rect 22192 24837 22201 24871
rect 22201 24837 22235 24871
rect 22235 24837 22244 24871
rect 22192 24828 22244 24837
rect 21548 24760 21600 24812
rect 23664 24896 23716 24948
rect 25504 24896 25556 24948
rect 26976 24939 27028 24948
rect 26976 24905 26985 24939
rect 26985 24905 27019 24939
rect 27019 24905 27028 24939
rect 26976 24896 27028 24905
rect 27620 24896 27672 24948
rect 22560 24803 22612 24812
rect 22560 24769 22569 24803
rect 22569 24769 22603 24803
rect 22603 24769 22612 24803
rect 22560 24760 22612 24769
rect 22468 24692 22520 24744
rect 27344 24828 27396 24880
rect 27436 24828 27488 24880
rect 22928 24803 22980 24812
rect 22928 24769 22937 24803
rect 22937 24769 22971 24803
rect 22971 24769 22980 24803
rect 22928 24760 22980 24769
rect 23020 24803 23072 24812
rect 23020 24769 23034 24803
rect 23034 24769 23068 24803
rect 23068 24769 23072 24803
rect 23020 24760 23072 24769
rect 26516 24760 26568 24812
rect 28080 24760 28132 24812
rect 24676 24692 24728 24744
rect 21272 24667 21324 24676
rect 21272 24633 21281 24667
rect 21281 24633 21315 24667
rect 21315 24633 21324 24667
rect 21272 24624 21324 24633
rect 28908 24896 28960 24948
rect 35348 24896 35400 24948
rect 29644 24828 29696 24880
rect 30012 24828 30064 24880
rect 28540 24803 28592 24812
rect 28540 24769 28549 24803
rect 28549 24769 28583 24803
rect 28583 24769 28592 24803
rect 28540 24760 28592 24769
rect 28632 24760 28684 24812
rect 28724 24760 28776 24812
rect 30932 24760 30984 24812
rect 32404 24828 32456 24880
rect 33968 24828 34020 24880
rect 34336 24828 34388 24880
rect 32864 24760 32916 24812
rect 33140 24760 33192 24812
rect 34060 24760 34112 24812
rect 35348 24803 35400 24812
rect 35348 24769 35381 24803
rect 35381 24769 35400 24803
rect 35348 24760 35400 24769
rect 40132 24828 40184 24880
rect 35624 24760 35676 24812
rect 30656 24692 30708 24744
rect 31208 24692 31260 24744
rect 32036 24692 32088 24744
rect 33416 24692 33468 24744
rect 34244 24692 34296 24744
rect 28448 24624 28500 24676
rect 36544 24760 36596 24812
rect 39028 24760 39080 24812
rect 36452 24692 36504 24744
rect 39304 24735 39356 24744
rect 39304 24701 39313 24735
rect 39313 24701 39347 24735
rect 39347 24701 39356 24735
rect 39304 24692 39356 24701
rect 39580 24735 39632 24744
rect 39580 24701 39589 24735
rect 39589 24701 39623 24735
rect 39623 24701 39632 24735
rect 39580 24692 39632 24701
rect 39948 24692 40000 24744
rect 21916 24556 21968 24608
rect 23020 24556 23072 24608
rect 23848 24556 23900 24608
rect 24492 24556 24544 24608
rect 25964 24556 26016 24608
rect 27252 24556 27304 24608
rect 28264 24556 28316 24608
rect 29644 24556 29696 24608
rect 30840 24556 30892 24608
rect 31300 24556 31352 24608
rect 32036 24556 32088 24608
rect 32128 24599 32180 24608
rect 32128 24565 32137 24599
rect 32137 24565 32171 24599
rect 32171 24565 32180 24599
rect 32128 24556 32180 24565
rect 32588 24599 32640 24608
rect 32588 24565 32597 24599
rect 32597 24565 32631 24599
rect 32631 24565 32640 24599
rect 32588 24556 32640 24565
rect 32864 24556 32916 24608
rect 33600 24556 33652 24608
rect 36176 24556 36228 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 4896 24395 4948 24404
rect 4896 24361 4905 24395
rect 4905 24361 4939 24395
rect 4939 24361 4948 24395
rect 4896 24352 4948 24361
rect 4988 24352 5040 24404
rect 5080 24352 5132 24404
rect 5632 24395 5684 24404
rect 5632 24361 5641 24395
rect 5641 24361 5675 24395
rect 5675 24361 5684 24395
rect 5632 24352 5684 24361
rect 6828 24352 6880 24404
rect 3884 24216 3936 24268
rect 4712 24148 4764 24200
rect 7748 24284 7800 24336
rect 9312 24352 9364 24404
rect 9496 24395 9548 24404
rect 9496 24361 9505 24395
rect 9505 24361 9539 24395
rect 9539 24361 9548 24395
rect 9496 24352 9548 24361
rect 5356 24148 5408 24200
rect 6460 24148 6512 24200
rect 7196 24216 7248 24268
rect 11152 24284 11204 24336
rect 12256 24352 12308 24404
rect 14004 24352 14056 24404
rect 14464 24352 14516 24404
rect 17316 24352 17368 24404
rect 17776 24352 17828 24404
rect 19340 24352 19392 24404
rect 19708 24352 19760 24404
rect 21272 24352 21324 24404
rect 21916 24352 21968 24404
rect 22560 24352 22612 24404
rect 23296 24352 23348 24404
rect 5264 24123 5316 24132
rect 5264 24089 5273 24123
rect 5273 24089 5307 24123
rect 5307 24089 5316 24123
rect 5264 24080 5316 24089
rect 5632 24123 5684 24132
rect 5632 24089 5641 24123
rect 5641 24089 5675 24123
rect 5675 24089 5684 24123
rect 5632 24080 5684 24089
rect 5724 24080 5776 24132
rect 6920 24080 6972 24132
rect 7196 24080 7248 24132
rect 7656 24123 7708 24132
rect 7656 24089 7665 24123
rect 7665 24089 7699 24123
rect 7699 24089 7708 24123
rect 7656 24080 7708 24089
rect 7840 24123 7892 24132
rect 7840 24089 7849 24123
rect 7849 24089 7883 24123
rect 7883 24089 7892 24123
rect 7840 24080 7892 24089
rect 2780 24055 2832 24064
rect 2780 24021 2789 24055
rect 2789 24021 2823 24055
rect 2823 24021 2832 24055
rect 2780 24012 2832 24021
rect 4252 24055 4304 24064
rect 4252 24021 4261 24055
rect 4261 24021 4295 24055
rect 4295 24021 4304 24055
rect 4252 24012 4304 24021
rect 5816 24055 5868 24064
rect 5816 24021 5825 24055
rect 5825 24021 5859 24055
rect 5859 24021 5868 24055
rect 8116 24148 8168 24200
rect 8300 24123 8352 24132
rect 8300 24089 8309 24123
rect 8309 24089 8343 24123
rect 8343 24089 8352 24123
rect 8300 24080 8352 24089
rect 8668 24148 8720 24200
rect 9036 24148 9088 24200
rect 9956 24216 10008 24268
rect 11796 24216 11848 24268
rect 12532 24284 12584 24336
rect 12900 24327 12952 24336
rect 12900 24293 12909 24327
rect 12909 24293 12943 24327
rect 12943 24293 12952 24327
rect 12900 24284 12952 24293
rect 13176 24284 13228 24336
rect 12808 24259 12860 24268
rect 12808 24225 12817 24259
rect 12817 24225 12851 24259
rect 12851 24225 12860 24259
rect 12808 24216 12860 24225
rect 9588 24148 9640 24200
rect 10232 24148 10284 24200
rect 11980 24191 12032 24200
rect 11980 24157 11989 24191
rect 11989 24157 12023 24191
rect 12023 24157 12032 24191
rect 11980 24148 12032 24157
rect 12348 24191 12400 24200
rect 12348 24157 12357 24191
rect 12357 24157 12391 24191
rect 12391 24157 12400 24191
rect 12348 24148 12400 24157
rect 13636 24284 13688 24336
rect 15200 24284 15252 24336
rect 13360 24148 13412 24200
rect 8760 24080 8812 24132
rect 14372 24148 14424 24200
rect 20904 24284 20956 24336
rect 21364 24284 21416 24336
rect 16212 24148 16264 24200
rect 16488 24148 16540 24200
rect 20628 24216 20680 24268
rect 21732 24216 21784 24268
rect 18144 24148 18196 24200
rect 18328 24191 18380 24200
rect 18328 24157 18337 24191
rect 18337 24157 18371 24191
rect 18371 24157 18380 24191
rect 18328 24148 18380 24157
rect 14004 24080 14056 24132
rect 14648 24080 14700 24132
rect 5816 24012 5868 24021
rect 12992 24012 13044 24064
rect 15384 24012 15436 24064
rect 15844 24055 15896 24064
rect 15844 24021 15853 24055
rect 15853 24021 15887 24055
rect 15887 24021 15896 24055
rect 15844 24012 15896 24021
rect 18052 24080 18104 24132
rect 19984 24148 20036 24200
rect 22468 24148 22520 24200
rect 19800 24080 19852 24132
rect 22744 24148 22796 24200
rect 23296 24259 23348 24268
rect 23296 24225 23305 24259
rect 23305 24225 23339 24259
rect 23339 24225 23348 24259
rect 23296 24216 23348 24225
rect 23020 24148 23072 24200
rect 24400 24395 24452 24404
rect 24400 24361 24409 24395
rect 24409 24361 24443 24395
rect 24443 24361 24452 24395
rect 24400 24352 24452 24361
rect 24952 24395 25004 24404
rect 24952 24361 24961 24395
rect 24961 24361 24995 24395
rect 24995 24361 25004 24395
rect 24952 24352 25004 24361
rect 25136 24352 25188 24404
rect 25412 24352 25464 24404
rect 27436 24352 27488 24404
rect 28540 24352 28592 24404
rect 28816 24352 28868 24404
rect 29644 24352 29696 24404
rect 30012 24352 30064 24404
rect 31484 24395 31536 24404
rect 31484 24361 31493 24395
rect 31493 24361 31527 24395
rect 31527 24361 31536 24395
rect 31484 24352 31536 24361
rect 31852 24352 31904 24404
rect 32496 24352 32548 24404
rect 33600 24352 33652 24404
rect 35348 24352 35400 24404
rect 35532 24352 35584 24404
rect 38292 24352 38344 24404
rect 39580 24352 39632 24404
rect 27620 24284 27672 24336
rect 28264 24284 28316 24336
rect 30840 24284 30892 24336
rect 32220 24284 32272 24336
rect 33508 24327 33560 24336
rect 33508 24293 33517 24327
rect 33517 24293 33551 24327
rect 33551 24293 33560 24327
rect 33508 24284 33560 24293
rect 33876 24284 33928 24336
rect 34152 24284 34204 24336
rect 24584 24259 24636 24268
rect 24584 24225 24593 24259
rect 24593 24225 24627 24259
rect 24627 24225 24636 24259
rect 24584 24216 24636 24225
rect 25964 24216 26016 24268
rect 28724 24216 28776 24268
rect 17500 24012 17552 24064
rect 17684 24012 17736 24064
rect 20260 24055 20312 24064
rect 20260 24021 20269 24055
rect 20269 24021 20303 24055
rect 20303 24021 20312 24055
rect 20260 24012 20312 24021
rect 23296 24080 23348 24132
rect 23664 24123 23716 24132
rect 23664 24089 23673 24123
rect 23673 24089 23707 24123
rect 23707 24089 23716 24123
rect 23664 24080 23716 24089
rect 23848 24055 23900 24064
rect 23848 24021 23873 24055
rect 23873 24021 23900 24055
rect 24400 24123 24452 24132
rect 24400 24089 24409 24123
rect 24409 24089 24443 24123
rect 24443 24089 24452 24123
rect 24400 24080 24452 24089
rect 24676 24191 24728 24200
rect 24676 24157 24685 24191
rect 24685 24157 24719 24191
rect 24719 24157 24728 24191
rect 24676 24148 24728 24157
rect 24952 24148 25004 24200
rect 25228 24080 25280 24132
rect 25320 24080 25372 24132
rect 25504 24123 25556 24132
rect 25504 24089 25513 24123
rect 25513 24089 25547 24123
rect 25547 24089 25556 24123
rect 25504 24080 25556 24089
rect 25688 24123 25740 24132
rect 25688 24089 25713 24123
rect 25713 24089 25740 24123
rect 25688 24080 25740 24089
rect 26056 24080 26108 24132
rect 26976 24148 27028 24200
rect 27528 24148 27580 24200
rect 27620 24191 27672 24200
rect 27620 24157 27629 24191
rect 27629 24157 27663 24191
rect 27663 24157 27672 24191
rect 27620 24148 27672 24157
rect 27896 24148 27948 24200
rect 28172 24148 28224 24200
rect 28264 24191 28316 24200
rect 28264 24157 28273 24191
rect 28273 24157 28307 24191
rect 28307 24157 28316 24191
rect 28264 24148 28316 24157
rect 28448 24148 28500 24200
rect 29460 24148 29512 24200
rect 29736 24148 29788 24200
rect 29092 24080 29144 24132
rect 30104 24191 30156 24200
rect 30104 24157 30113 24191
rect 30113 24157 30147 24191
rect 30147 24157 30156 24191
rect 30104 24148 30156 24157
rect 30288 24148 30340 24200
rect 30380 24148 30432 24200
rect 30840 24148 30892 24200
rect 23848 24012 23900 24021
rect 26148 24012 26200 24064
rect 26700 24012 26752 24064
rect 27252 24012 27304 24064
rect 27344 24012 27396 24064
rect 28356 24012 28408 24064
rect 31300 24123 31352 24132
rect 31300 24089 31309 24123
rect 31309 24089 31343 24123
rect 31343 24089 31352 24123
rect 31300 24080 31352 24089
rect 31484 24191 31536 24200
rect 31484 24157 31493 24191
rect 31493 24157 31527 24191
rect 31527 24157 31536 24191
rect 31484 24148 31536 24157
rect 33324 24259 33376 24268
rect 33324 24225 33333 24259
rect 33333 24225 33367 24259
rect 33367 24225 33376 24259
rect 33324 24216 33376 24225
rect 32864 24148 32916 24200
rect 29920 24012 29972 24064
rect 30104 24012 30156 24064
rect 30380 24012 30432 24064
rect 32496 24012 32548 24064
rect 33232 24012 33284 24064
rect 33968 24191 34020 24200
rect 33968 24157 33977 24191
rect 33977 24157 34011 24191
rect 34011 24157 34020 24191
rect 37556 24259 37608 24268
rect 37556 24225 37565 24259
rect 37565 24225 37599 24259
rect 37599 24225 37608 24259
rect 37556 24216 37608 24225
rect 33968 24148 34020 24157
rect 34428 24080 34480 24132
rect 37280 24148 37332 24200
rect 37740 24148 37792 24200
rect 37832 24148 37884 24200
rect 38384 24148 38436 24200
rect 40316 24191 40368 24200
rect 40316 24157 40325 24191
rect 40325 24157 40359 24191
rect 40359 24157 40368 24191
rect 40316 24148 40368 24157
rect 35164 24080 35216 24132
rect 36728 24080 36780 24132
rect 38660 24080 38712 24132
rect 35992 24012 36044 24064
rect 37372 24055 37424 24064
rect 37372 24021 37381 24055
rect 37381 24021 37415 24055
rect 37415 24021 37424 24055
rect 37372 24012 37424 24021
rect 38476 24012 38528 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 2780 23808 2832 23860
rect 3056 23808 3108 23860
rect 4068 23808 4120 23860
rect 5816 23808 5868 23860
rect 7196 23851 7248 23860
rect 7196 23817 7205 23851
rect 7205 23817 7239 23851
rect 7239 23817 7248 23851
rect 7196 23808 7248 23817
rect 4252 23740 4304 23792
rect 5264 23740 5316 23792
rect 5540 23740 5592 23792
rect 2412 23647 2464 23656
rect 2412 23613 2421 23647
rect 2421 23613 2455 23647
rect 2455 23613 2464 23647
rect 2412 23604 2464 23613
rect 7380 23715 7432 23724
rect 7380 23681 7389 23715
rect 7389 23681 7423 23715
rect 7423 23681 7432 23715
rect 7380 23672 7432 23681
rect 8852 23808 8904 23860
rect 9496 23808 9548 23860
rect 9956 23808 10008 23860
rect 11060 23808 11112 23860
rect 13084 23808 13136 23860
rect 13636 23808 13688 23860
rect 8484 23672 8536 23724
rect 9036 23715 9088 23724
rect 9036 23681 9045 23715
rect 9045 23681 9079 23715
rect 9079 23681 9088 23715
rect 9036 23672 9088 23681
rect 9404 23715 9456 23724
rect 9404 23681 9413 23715
rect 9413 23681 9447 23715
rect 9447 23681 9456 23715
rect 9404 23672 9456 23681
rect 9588 23672 9640 23724
rect 9680 23672 9732 23724
rect 10508 23672 10560 23724
rect 14556 23783 14608 23792
rect 14556 23749 14565 23783
rect 14565 23749 14599 23783
rect 14599 23749 14608 23783
rect 14556 23740 14608 23749
rect 7472 23579 7524 23588
rect 7472 23545 7481 23579
rect 7481 23545 7515 23579
rect 7515 23545 7524 23579
rect 7472 23536 7524 23545
rect 9496 23536 9548 23588
rect 7104 23468 7156 23520
rect 12992 23715 13044 23724
rect 12992 23681 13001 23715
rect 13001 23681 13035 23715
rect 13035 23681 13044 23715
rect 12992 23672 13044 23681
rect 13084 23715 13136 23724
rect 13084 23681 13105 23715
rect 13105 23681 13136 23715
rect 13084 23672 13136 23681
rect 14372 23672 14424 23724
rect 14464 23715 14516 23724
rect 14464 23681 14473 23715
rect 14473 23681 14507 23715
rect 14507 23681 14516 23715
rect 14464 23672 14516 23681
rect 15016 23808 15068 23860
rect 11244 23604 11296 23656
rect 12164 23536 12216 23588
rect 13820 23536 13872 23588
rect 15384 23740 15436 23792
rect 15660 23740 15712 23792
rect 15108 23715 15160 23724
rect 15108 23681 15117 23715
rect 15117 23681 15151 23715
rect 15151 23681 15160 23715
rect 15108 23672 15160 23681
rect 15476 23715 15528 23724
rect 15476 23681 15485 23715
rect 15485 23681 15519 23715
rect 15519 23681 15528 23715
rect 15476 23672 15528 23681
rect 15844 23715 15896 23724
rect 15844 23681 15853 23715
rect 15853 23681 15887 23715
rect 15887 23681 15896 23715
rect 15844 23672 15896 23681
rect 16580 23672 16632 23724
rect 17316 23808 17368 23860
rect 18328 23851 18380 23860
rect 17684 23672 17736 23724
rect 18328 23817 18337 23851
rect 18337 23817 18371 23851
rect 18371 23817 18380 23851
rect 18328 23808 18380 23817
rect 18604 23808 18656 23860
rect 20168 23808 20220 23860
rect 20444 23808 20496 23860
rect 20720 23851 20772 23860
rect 20720 23817 20729 23851
rect 20729 23817 20763 23851
rect 20763 23817 20772 23851
rect 20720 23808 20772 23817
rect 21272 23808 21324 23860
rect 21456 23808 21508 23860
rect 21732 23808 21784 23860
rect 22928 23808 22980 23860
rect 21824 23740 21876 23792
rect 12716 23468 12768 23520
rect 17500 23536 17552 23588
rect 17776 23579 17828 23588
rect 17776 23545 17785 23579
rect 17785 23545 17819 23579
rect 17819 23545 17828 23579
rect 17776 23536 17828 23545
rect 17960 23579 18012 23588
rect 17960 23545 17969 23579
rect 17969 23545 18003 23579
rect 18003 23545 18012 23579
rect 17960 23536 18012 23545
rect 20168 23536 20220 23588
rect 21180 23715 21232 23724
rect 21180 23681 21189 23715
rect 21189 23681 21223 23715
rect 21223 23681 21232 23715
rect 21180 23672 21232 23681
rect 21364 23715 21416 23724
rect 21364 23681 21373 23715
rect 21373 23681 21407 23715
rect 21407 23681 21416 23715
rect 21364 23672 21416 23681
rect 23480 23740 23532 23792
rect 25228 23808 25280 23860
rect 26608 23808 26660 23860
rect 20720 23604 20772 23656
rect 22468 23647 22520 23656
rect 22468 23613 22477 23647
rect 22477 23613 22511 23647
rect 22511 23613 22520 23647
rect 22468 23604 22520 23613
rect 23848 23672 23900 23724
rect 24492 23672 24544 23724
rect 24584 23715 24636 23724
rect 24584 23681 24593 23715
rect 24593 23681 24627 23715
rect 24627 23681 24636 23715
rect 24584 23672 24636 23681
rect 24860 23715 24912 23724
rect 24860 23681 24869 23715
rect 24869 23681 24903 23715
rect 24903 23681 24912 23715
rect 24860 23672 24912 23681
rect 26240 23783 26292 23792
rect 26240 23749 26249 23783
rect 26249 23749 26283 23783
rect 26283 23749 26292 23783
rect 26240 23740 26292 23749
rect 25044 23715 25096 23724
rect 25044 23681 25058 23715
rect 25058 23681 25092 23715
rect 25092 23681 25096 23715
rect 25044 23672 25096 23681
rect 25412 23672 25464 23724
rect 26700 23740 26752 23792
rect 25320 23604 25372 23656
rect 25964 23604 26016 23656
rect 26608 23715 26660 23724
rect 26608 23681 26617 23715
rect 26617 23681 26651 23715
rect 26651 23681 26660 23715
rect 26608 23672 26660 23681
rect 17224 23511 17276 23520
rect 17224 23477 17233 23511
rect 17233 23477 17267 23511
rect 17267 23477 17276 23511
rect 17224 23468 17276 23477
rect 18144 23468 18196 23520
rect 20260 23511 20312 23520
rect 20260 23477 20269 23511
rect 20269 23477 20303 23511
rect 20303 23477 20312 23511
rect 20260 23468 20312 23477
rect 20996 23536 21048 23588
rect 21548 23468 21600 23520
rect 22376 23511 22428 23520
rect 22376 23477 22385 23511
rect 22385 23477 22419 23511
rect 22419 23477 22428 23511
rect 22376 23468 22428 23477
rect 23480 23536 23532 23588
rect 23756 23468 23808 23520
rect 25780 23468 25832 23520
rect 26332 23536 26384 23588
rect 26884 23468 26936 23520
rect 28172 23808 28224 23860
rect 28264 23808 28316 23860
rect 31300 23808 31352 23860
rect 31668 23808 31720 23860
rect 32588 23808 32640 23860
rect 32680 23808 32732 23860
rect 34060 23808 34112 23860
rect 28080 23740 28132 23792
rect 28448 23740 28500 23792
rect 28816 23740 28868 23792
rect 27712 23672 27764 23724
rect 28172 23672 28224 23724
rect 28908 23672 28960 23724
rect 29000 23715 29052 23724
rect 29000 23681 29009 23715
rect 29009 23681 29043 23715
rect 29043 23681 29052 23715
rect 29000 23672 29052 23681
rect 29368 23672 29420 23724
rect 29460 23672 29512 23724
rect 29644 23672 29696 23724
rect 30104 23672 30156 23724
rect 30196 23672 30248 23724
rect 28264 23604 28316 23656
rect 27712 23536 27764 23588
rect 31208 23715 31260 23724
rect 31208 23681 31217 23715
rect 31217 23681 31251 23715
rect 31251 23681 31260 23715
rect 31208 23672 31260 23681
rect 31300 23715 31352 23724
rect 31300 23681 31309 23715
rect 31309 23681 31343 23715
rect 31343 23681 31352 23715
rect 31300 23672 31352 23681
rect 27436 23468 27488 23520
rect 27988 23468 28040 23520
rect 28356 23468 28408 23520
rect 32404 23604 32456 23656
rect 29736 23511 29788 23520
rect 29736 23477 29745 23511
rect 29745 23477 29779 23511
rect 29779 23477 29788 23511
rect 29736 23468 29788 23477
rect 31208 23536 31260 23588
rect 32588 23672 32640 23724
rect 32956 23715 33008 23724
rect 32956 23681 32965 23715
rect 32965 23681 32999 23715
rect 32999 23681 33008 23715
rect 32956 23672 33008 23681
rect 33692 23672 33744 23724
rect 33876 23672 33928 23724
rect 34520 23740 34572 23792
rect 32588 23536 32640 23588
rect 32680 23536 32732 23588
rect 35164 23715 35216 23724
rect 35164 23681 35173 23715
rect 35173 23681 35207 23715
rect 35207 23681 35216 23715
rect 35164 23672 35216 23681
rect 37832 23808 37884 23860
rect 38016 23808 38068 23860
rect 35532 23604 35584 23656
rect 36452 23647 36504 23656
rect 36452 23613 36461 23647
rect 36461 23613 36495 23647
rect 36495 23613 36504 23647
rect 36452 23604 36504 23613
rect 37464 23672 37516 23724
rect 34060 23468 34112 23520
rect 34428 23468 34480 23520
rect 37556 23579 37608 23588
rect 37556 23545 37565 23579
rect 37565 23545 37599 23579
rect 37599 23545 37608 23579
rect 37556 23536 37608 23545
rect 38292 23672 38344 23724
rect 38384 23672 38436 23724
rect 38752 23783 38804 23792
rect 38752 23749 38761 23783
rect 38761 23749 38795 23783
rect 38795 23749 38804 23783
rect 38752 23740 38804 23749
rect 39120 23808 39172 23860
rect 38476 23604 38528 23656
rect 38936 23715 38988 23724
rect 38936 23681 38945 23715
rect 38945 23681 38979 23715
rect 38979 23681 38988 23715
rect 38936 23672 38988 23681
rect 36544 23468 36596 23520
rect 37004 23468 37056 23520
rect 39120 23579 39172 23588
rect 39120 23545 39129 23579
rect 39129 23545 39163 23579
rect 39163 23545 39172 23579
rect 39120 23536 39172 23545
rect 37740 23511 37792 23520
rect 37740 23477 37749 23511
rect 37749 23477 37783 23511
rect 37783 23477 37792 23511
rect 37740 23468 37792 23477
rect 38752 23468 38804 23520
rect 39580 23715 39632 23724
rect 39580 23681 39589 23715
rect 39589 23681 39623 23715
rect 39623 23681 39632 23715
rect 39580 23672 39632 23681
rect 39764 23511 39816 23520
rect 39764 23477 39773 23511
rect 39773 23477 39807 23511
rect 39807 23477 39816 23511
rect 39764 23468 39816 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 5080 23264 5132 23316
rect 7104 23264 7156 23316
rect 7472 23264 7524 23316
rect 8116 23264 8168 23316
rect 3148 23239 3200 23248
rect 3148 23205 3157 23239
rect 3157 23205 3191 23239
rect 3191 23205 3200 23239
rect 3148 23196 3200 23205
rect 2412 23128 2464 23180
rect 3056 23060 3108 23112
rect 5080 23103 5132 23112
rect 5080 23069 5089 23103
rect 5089 23069 5123 23103
rect 5123 23069 5132 23103
rect 5080 23060 5132 23069
rect 1676 23035 1728 23044
rect 1676 23001 1685 23035
rect 1685 23001 1719 23035
rect 1719 23001 1728 23035
rect 1676 22992 1728 23001
rect 9404 23196 9456 23248
rect 5264 23103 5316 23112
rect 5264 23069 5273 23103
rect 5273 23069 5307 23103
rect 5307 23069 5316 23103
rect 5264 23060 5316 23069
rect 6000 23060 6052 23112
rect 7104 23060 7156 23112
rect 7472 23103 7524 23112
rect 7472 23069 7481 23103
rect 7481 23069 7515 23103
rect 7515 23069 7524 23103
rect 7472 23060 7524 23069
rect 7932 23060 7984 23112
rect 8576 23060 8628 23112
rect 8852 23060 8904 23112
rect 10600 23128 10652 23180
rect 8116 22992 8168 23044
rect 10508 23060 10560 23112
rect 4804 22924 4856 22976
rect 9496 22924 9548 22976
rect 9588 22924 9640 22976
rect 11980 23307 12032 23316
rect 11980 23273 11989 23307
rect 11989 23273 12023 23307
rect 12023 23273 12032 23307
rect 11980 23264 12032 23273
rect 14464 23264 14516 23316
rect 15844 23264 15896 23316
rect 17684 23264 17736 23316
rect 22192 23264 22244 23316
rect 22744 23264 22796 23316
rect 23940 23264 23992 23316
rect 26424 23264 26476 23316
rect 26884 23264 26936 23316
rect 27344 23264 27396 23316
rect 27620 23264 27672 23316
rect 30012 23264 30064 23316
rect 39856 23264 39908 23316
rect 40224 23264 40276 23316
rect 40316 23307 40368 23316
rect 40316 23273 40325 23307
rect 40325 23273 40359 23307
rect 40359 23273 40368 23307
rect 40316 23264 40368 23273
rect 14004 23128 14056 23180
rect 17500 23196 17552 23248
rect 11612 22992 11664 23044
rect 11152 22924 11204 22976
rect 11244 22924 11296 22976
rect 11980 23060 12032 23112
rect 12348 22992 12400 23044
rect 13360 22924 13412 22976
rect 14648 23103 14700 23112
rect 14648 23069 14657 23103
rect 14657 23069 14691 23103
rect 14691 23069 14700 23103
rect 16120 23128 16172 23180
rect 16304 23128 16356 23180
rect 19340 23128 19392 23180
rect 14648 23060 14700 23069
rect 14832 22992 14884 23044
rect 15200 22992 15252 23044
rect 15752 23103 15804 23112
rect 15752 23069 15761 23103
rect 15761 23069 15795 23103
rect 15795 23069 15804 23103
rect 15752 23060 15804 23069
rect 15936 23103 15988 23112
rect 15936 23069 15945 23103
rect 15945 23069 15979 23103
rect 15979 23069 15988 23103
rect 15936 23060 15988 23069
rect 17316 23060 17368 23112
rect 17408 23103 17460 23112
rect 17408 23069 17417 23103
rect 17417 23069 17451 23103
rect 17451 23069 17460 23103
rect 17408 23060 17460 23069
rect 18052 23060 18104 23112
rect 18328 23060 18380 23112
rect 20536 23060 20588 23112
rect 16488 22992 16540 23044
rect 16672 22992 16724 23044
rect 17224 22992 17276 23044
rect 18696 22992 18748 23044
rect 21180 23171 21232 23180
rect 21180 23137 21189 23171
rect 21189 23137 21223 23171
rect 21223 23137 21232 23171
rect 21180 23128 21232 23137
rect 24676 23196 24728 23248
rect 22928 23128 22980 23180
rect 29460 23196 29512 23248
rect 29828 23196 29880 23248
rect 30196 23196 30248 23248
rect 32680 23196 32732 23248
rect 25044 23128 25096 23180
rect 14556 22924 14608 22976
rect 16212 22924 16264 22976
rect 17408 22924 17460 22976
rect 18052 22967 18104 22976
rect 18052 22933 18061 22967
rect 18061 22933 18095 22967
rect 18095 22933 18104 22967
rect 18052 22924 18104 22933
rect 20720 22967 20772 22976
rect 20720 22933 20729 22967
rect 20729 22933 20763 22967
rect 20763 22933 20772 22967
rect 20720 22924 20772 22933
rect 21456 23060 21508 23112
rect 21548 23060 21600 23112
rect 21272 23035 21324 23044
rect 21272 23001 21281 23035
rect 21281 23001 21315 23035
rect 21315 23001 21324 23035
rect 21272 22992 21324 23001
rect 23388 23103 23440 23112
rect 23388 23069 23397 23103
rect 23397 23069 23431 23103
rect 23431 23069 23440 23103
rect 23388 23060 23440 23069
rect 26516 23128 26568 23180
rect 26056 23103 26108 23112
rect 26056 23069 26065 23103
rect 26065 23069 26099 23103
rect 26099 23069 26108 23103
rect 26056 23060 26108 23069
rect 26884 23103 26936 23112
rect 26884 23069 26893 23103
rect 26893 23069 26927 23103
rect 26927 23069 26936 23103
rect 26884 23060 26936 23069
rect 27252 23103 27304 23112
rect 27252 23069 27261 23103
rect 27261 23069 27295 23103
rect 27295 23069 27304 23103
rect 27252 23060 27304 23069
rect 27620 23060 27672 23112
rect 27896 23103 27948 23112
rect 27896 23069 27905 23103
rect 27905 23069 27939 23103
rect 27939 23069 27948 23103
rect 27896 23060 27948 23069
rect 28356 23060 28408 23112
rect 25504 22992 25556 23044
rect 28540 23060 28592 23112
rect 30380 23060 30432 23112
rect 31668 23103 31720 23112
rect 31668 23069 31677 23103
rect 31677 23069 31711 23103
rect 31711 23069 31720 23103
rect 31668 23060 31720 23069
rect 31760 23103 31812 23112
rect 31760 23069 31769 23103
rect 31769 23069 31803 23103
rect 31803 23069 31812 23103
rect 31760 23060 31812 23069
rect 32588 23128 32640 23180
rect 32864 23128 32916 23180
rect 36176 23171 36228 23180
rect 36176 23137 36185 23171
rect 36185 23137 36219 23171
rect 36219 23137 36228 23171
rect 36176 23128 36228 23137
rect 32036 23060 32088 23112
rect 22836 22924 22888 22976
rect 23572 22924 23624 22976
rect 24860 22924 24912 22976
rect 26884 22924 26936 22976
rect 28080 22967 28132 22976
rect 28080 22933 28089 22967
rect 28089 22933 28123 22967
rect 28123 22933 28132 22967
rect 28080 22924 28132 22933
rect 30564 22924 30616 22976
rect 31852 22967 31904 22976
rect 31852 22933 31861 22967
rect 31861 22933 31895 22967
rect 31895 22933 31904 22967
rect 31852 22924 31904 22933
rect 32220 22992 32272 23044
rect 33232 23060 33284 23112
rect 32956 22992 33008 23044
rect 32680 22924 32732 22976
rect 34428 23103 34480 23112
rect 34428 23069 34437 23103
rect 34437 23069 34471 23103
rect 34471 23069 34480 23103
rect 34428 23060 34480 23069
rect 36268 23103 36320 23112
rect 36268 23069 36277 23103
rect 36277 23069 36311 23103
rect 36311 23069 36320 23103
rect 36268 23060 36320 23069
rect 37188 23060 37240 23112
rect 38568 23060 38620 23112
rect 39028 23196 39080 23248
rect 34520 22992 34572 23044
rect 35808 22992 35860 23044
rect 36636 23035 36688 23044
rect 36636 23001 36645 23035
rect 36645 23001 36679 23035
rect 36679 23001 36688 23035
rect 36636 22992 36688 23001
rect 38752 22992 38804 23044
rect 33508 22924 33560 22976
rect 37280 22924 37332 22976
rect 37464 22924 37516 22976
rect 39580 23060 39632 23112
rect 39948 23035 40000 23044
rect 39948 23001 39957 23035
rect 39957 23001 39991 23035
rect 39991 23001 40000 23035
rect 39948 22992 40000 23001
rect 40592 22992 40644 23044
rect 39212 22967 39264 22976
rect 39212 22933 39221 22967
rect 39221 22933 39255 22967
rect 39255 22933 39264 22967
rect 39212 22924 39264 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 1676 22720 1728 22772
rect 2872 22763 2924 22772
rect 2872 22729 2881 22763
rect 2881 22729 2915 22763
rect 2915 22729 2924 22763
rect 2872 22720 2924 22729
rect 3148 22720 3200 22772
rect 5908 22763 5960 22772
rect 5908 22729 5917 22763
rect 5917 22729 5951 22763
rect 5951 22729 5960 22763
rect 5908 22720 5960 22729
rect 7472 22720 7524 22772
rect 11888 22720 11940 22772
rect 5816 22652 5868 22704
rect 7288 22652 7340 22704
rect 9128 22652 9180 22704
rect 6368 22584 6420 22636
rect 8208 22584 8260 22636
rect 4160 22559 4212 22568
rect 4160 22525 4169 22559
rect 4169 22525 4203 22559
rect 4203 22525 4212 22559
rect 4160 22516 4212 22525
rect 4528 22516 4580 22568
rect 7196 22516 7248 22568
rect 9404 22516 9456 22568
rect 9496 22516 9548 22568
rect 9772 22584 9824 22636
rect 10048 22584 10100 22636
rect 12072 22584 12124 22636
rect 12164 22627 12216 22636
rect 12164 22593 12173 22627
rect 12173 22593 12207 22627
rect 12207 22593 12216 22627
rect 12164 22584 12216 22593
rect 12532 22627 12584 22636
rect 12532 22593 12541 22627
rect 12541 22593 12575 22627
rect 12575 22593 12584 22627
rect 12532 22584 12584 22593
rect 12716 22627 12768 22636
rect 12716 22593 12725 22627
rect 12725 22593 12759 22627
rect 12759 22593 12768 22627
rect 12716 22584 12768 22593
rect 9588 22448 9640 22500
rect 12440 22516 12492 22568
rect 13728 22627 13780 22636
rect 13728 22593 13737 22627
rect 13737 22593 13771 22627
rect 13771 22593 13780 22627
rect 13728 22584 13780 22593
rect 14096 22584 14148 22636
rect 14740 22627 14792 22636
rect 14740 22593 14749 22627
rect 14749 22593 14783 22627
rect 14783 22593 14792 22627
rect 14740 22584 14792 22593
rect 15016 22584 15068 22636
rect 15476 22652 15528 22704
rect 16028 22652 16080 22704
rect 16488 22763 16540 22772
rect 16488 22729 16497 22763
rect 16497 22729 16531 22763
rect 16531 22729 16540 22763
rect 16488 22720 16540 22729
rect 15660 22627 15712 22636
rect 15660 22593 15669 22627
rect 15669 22593 15703 22627
rect 15703 22593 15712 22627
rect 15660 22584 15712 22593
rect 15844 22584 15896 22636
rect 15936 22627 15988 22636
rect 15936 22593 15945 22627
rect 15945 22593 15979 22627
rect 15979 22593 15988 22627
rect 15936 22584 15988 22593
rect 11704 22448 11756 22500
rect 3148 22380 3200 22432
rect 8392 22423 8444 22432
rect 8392 22389 8401 22423
rect 8401 22389 8435 22423
rect 8435 22389 8444 22423
rect 8392 22380 8444 22389
rect 10784 22380 10836 22432
rect 13912 22448 13964 22500
rect 14188 22380 14240 22432
rect 14924 22448 14976 22500
rect 15752 22448 15804 22500
rect 16764 22652 16816 22704
rect 16672 22584 16724 22636
rect 17040 22720 17092 22772
rect 17316 22720 17368 22772
rect 20168 22720 20220 22772
rect 21456 22720 21508 22772
rect 18052 22652 18104 22704
rect 18144 22652 18196 22704
rect 19892 22652 19944 22704
rect 21548 22652 21600 22704
rect 22100 22652 22152 22704
rect 22928 22720 22980 22772
rect 23664 22720 23716 22772
rect 16304 22516 16356 22568
rect 16488 22516 16540 22568
rect 17224 22627 17276 22636
rect 17224 22593 17233 22627
rect 17233 22593 17267 22627
rect 17267 22593 17276 22627
rect 17224 22584 17276 22593
rect 17408 22584 17460 22636
rect 18880 22584 18932 22636
rect 21272 22584 21324 22636
rect 23020 22652 23072 22704
rect 18420 22559 18472 22568
rect 18420 22525 18429 22559
rect 18429 22525 18463 22559
rect 18463 22525 18472 22559
rect 18420 22516 18472 22525
rect 18696 22516 18748 22568
rect 20720 22516 20772 22568
rect 21364 22516 21416 22568
rect 22836 22584 22888 22636
rect 24216 22652 24268 22704
rect 24676 22720 24728 22772
rect 27528 22720 27580 22772
rect 24492 22652 24544 22704
rect 25044 22652 25096 22704
rect 24032 22627 24084 22636
rect 24032 22593 24041 22627
rect 24041 22593 24075 22627
rect 24075 22593 24084 22627
rect 24032 22584 24084 22593
rect 30840 22720 30892 22772
rect 31760 22720 31812 22772
rect 32496 22720 32548 22772
rect 34888 22720 34940 22772
rect 28448 22695 28500 22704
rect 28448 22661 28457 22695
rect 28457 22661 28491 22695
rect 28491 22661 28500 22695
rect 28448 22652 28500 22661
rect 28264 22627 28316 22636
rect 28264 22593 28273 22627
rect 28273 22593 28307 22627
rect 28307 22593 28316 22627
rect 28264 22584 28316 22593
rect 28632 22584 28684 22636
rect 24492 22516 24544 22568
rect 25596 22516 25648 22568
rect 26240 22516 26292 22568
rect 16212 22423 16264 22432
rect 16212 22389 16221 22423
rect 16221 22389 16255 22423
rect 16255 22389 16264 22423
rect 16212 22380 16264 22389
rect 16764 22380 16816 22432
rect 17224 22380 17276 22432
rect 17408 22380 17460 22432
rect 23020 22448 23072 22500
rect 23848 22448 23900 22500
rect 23940 22448 23992 22500
rect 28724 22516 28776 22568
rect 20812 22380 20864 22432
rect 21272 22380 21324 22432
rect 22100 22423 22152 22432
rect 22100 22389 22109 22423
rect 22109 22389 22143 22423
rect 22143 22389 22152 22423
rect 22100 22380 22152 22389
rect 22192 22380 22244 22432
rect 22744 22380 22796 22432
rect 24216 22423 24268 22432
rect 24216 22389 24225 22423
rect 24225 22389 24259 22423
rect 24259 22389 24268 22423
rect 24216 22380 24268 22389
rect 29184 22584 29236 22636
rect 29644 22627 29696 22636
rect 29644 22593 29653 22627
rect 29653 22593 29687 22627
rect 29687 22593 29696 22627
rect 29644 22584 29696 22593
rect 29460 22559 29512 22568
rect 29460 22525 29469 22559
rect 29469 22525 29503 22559
rect 29503 22525 29512 22559
rect 29460 22516 29512 22525
rect 31208 22652 31260 22704
rect 31668 22652 31720 22704
rect 32220 22652 32272 22704
rect 34060 22652 34112 22704
rect 37464 22720 37516 22772
rect 39948 22720 40000 22772
rect 36636 22652 36688 22704
rect 38660 22652 38712 22704
rect 38844 22695 38896 22704
rect 38844 22661 38853 22695
rect 38853 22661 38887 22695
rect 38887 22661 38896 22695
rect 38844 22652 38896 22661
rect 30196 22584 30248 22636
rect 30012 22448 30064 22500
rect 30380 22584 30432 22636
rect 30656 22584 30708 22636
rect 30748 22584 30800 22636
rect 30932 22584 30984 22636
rect 31392 22584 31444 22636
rect 30472 22491 30524 22500
rect 30472 22457 30481 22491
rect 30481 22457 30515 22491
rect 30515 22457 30524 22491
rect 30472 22448 30524 22457
rect 30196 22380 30248 22432
rect 30656 22380 30708 22432
rect 31024 22516 31076 22568
rect 31576 22627 31628 22636
rect 31576 22593 31585 22627
rect 31585 22593 31619 22627
rect 31619 22593 31628 22627
rect 31576 22584 31628 22593
rect 31852 22584 31904 22636
rect 32128 22584 32180 22636
rect 32680 22627 32732 22636
rect 32680 22593 32689 22627
rect 32689 22593 32723 22627
rect 32723 22593 32732 22627
rect 32680 22584 32732 22593
rect 33232 22584 33284 22636
rect 34520 22584 34572 22636
rect 35348 22584 35400 22636
rect 33876 22516 33928 22568
rect 35808 22584 35860 22636
rect 35532 22516 35584 22568
rect 31024 22380 31076 22432
rect 32496 22423 32548 22432
rect 32496 22389 32505 22423
rect 32505 22389 32539 22423
rect 32539 22389 32548 22423
rect 32496 22380 32548 22389
rect 33232 22448 33284 22500
rect 33784 22448 33836 22500
rect 34428 22448 34480 22500
rect 36360 22627 36412 22636
rect 36360 22593 36369 22627
rect 36369 22593 36403 22627
rect 36403 22593 36412 22627
rect 36360 22584 36412 22593
rect 38568 22627 38620 22636
rect 38568 22593 38578 22627
rect 38578 22593 38612 22627
rect 38612 22593 38620 22627
rect 38568 22584 38620 22593
rect 39028 22584 39080 22636
rect 39120 22516 39172 22568
rect 39396 22627 39448 22636
rect 39396 22593 39405 22627
rect 39405 22593 39439 22627
rect 39439 22593 39448 22627
rect 39396 22584 39448 22593
rect 39488 22559 39540 22568
rect 39488 22525 39497 22559
rect 39497 22525 39531 22559
rect 39531 22525 39540 22559
rect 39488 22516 39540 22525
rect 38844 22448 38896 22500
rect 40684 22516 40736 22568
rect 35348 22380 35400 22432
rect 37832 22380 37884 22432
rect 39120 22423 39172 22432
rect 39120 22389 39129 22423
rect 39129 22389 39163 22423
rect 39163 22389 39172 22423
rect 39120 22380 39172 22389
rect 39212 22380 39264 22432
rect 39856 22380 39908 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 4620 22176 4672 22228
rect 5816 22219 5868 22228
rect 5816 22185 5825 22219
rect 5825 22185 5859 22219
rect 5859 22185 5868 22219
rect 5816 22176 5868 22185
rect 6092 22176 6144 22228
rect 7196 22219 7248 22228
rect 7196 22185 7205 22219
rect 7205 22185 7239 22219
rect 7239 22185 7248 22219
rect 7196 22176 7248 22185
rect 9220 22176 9272 22228
rect 11428 22176 11480 22228
rect 12164 22176 12216 22228
rect 12716 22176 12768 22228
rect 13820 22176 13872 22228
rect 14740 22219 14792 22228
rect 14740 22185 14749 22219
rect 14749 22185 14783 22219
rect 14783 22185 14792 22219
rect 14740 22176 14792 22185
rect 3148 22108 3200 22160
rect 5448 22083 5500 22092
rect 5448 22049 5457 22083
rect 5457 22049 5491 22083
rect 5491 22049 5500 22083
rect 5448 22040 5500 22049
rect 5908 22040 5960 22092
rect 7104 22040 7156 22092
rect 7472 22040 7524 22092
rect 4620 21904 4672 21956
rect 2504 21879 2556 21888
rect 2504 21845 2513 21879
rect 2513 21845 2547 21879
rect 2547 21845 2556 21879
rect 2504 21836 2556 21845
rect 2872 21879 2924 21888
rect 2872 21845 2881 21879
rect 2881 21845 2915 21879
rect 2915 21845 2924 21879
rect 2872 21836 2924 21845
rect 3148 21836 3200 21888
rect 8392 21972 8444 22024
rect 8852 21972 8904 22024
rect 9772 22108 9824 22160
rect 10140 22040 10192 22092
rect 10692 22040 10744 22092
rect 9312 22015 9364 22024
rect 9312 21981 9321 22015
rect 9321 21981 9355 22015
rect 9355 21981 9364 22015
rect 9312 21972 9364 21981
rect 9588 21972 9640 22024
rect 9772 22015 9824 22024
rect 9772 21981 9781 22015
rect 9781 21981 9815 22015
rect 9815 21981 9824 22015
rect 9772 21972 9824 21981
rect 10048 22015 10100 22024
rect 10048 21981 10057 22015
rect 10057 21981 10091 22015
rect 10091 21981 10100 22015
rect 10048 21972 10100 21981
rect 4988 21836 5040 21888
rect 5356 21904 5408 21956
rect 5632 21836 5684 21888
rect 5816 21904 5868 21956
rect 7288 21836 7340 21888
rect 9680 21879 9732 21888
rect 9680 21845 9689 21879
rect 9689 21845 9723 21879
rect 9723 21845 9732 21879
rect 9680 21836 9732 21845
rect 10600 22015 10652 22024
rect 10600 21981 10609 22015
rect 10609 21981 10643 22015
rect 10643 21981 10652 22015
rect 10600 21972 10652 21981
rect 10692 21904 10744 21956
rect 10876 22015 10928 22024
rect 10876 21981 10885 22015
rect 10885 21981 10919 22015
rect 10919 21981 10928 22015
rect 10876 21972 10928 21981
rect 11244 22040 11296 22092
rect 11980 22015 12032 22024
rect 11980 21981 11989 22015
rect 11989 21981 12023 22015
rect 12023 21981 12032 22015
rect 11980 21972 12032 21981
rect 12164 22015 12216 22024
rect 12164 21981 12171 22015
rect 12171 21981 12216 22015
rect 12164 21972 12216 21981
rect 12808 22108 12860 22160
rect 13084 22108 13136 22160
rect 12440 22015 12492 22024
rect 12440 21981 12454 22015
rect 12454 21981 12488 22015
rect 12488 21981 12492 22015
rect 12440 21972 12492 21981
rect 11152 21947 11204 21956
rect 11152 21913 11161 21947
rect 11161 21913 11195 21947
rect 11195 21913 11204 21947
rect 11152 21904 11204 21913
rect 11244 21947 11296 21956
rect 11244 21913 11253 21947
rect 11253 21913 11287 21947
rect 11287 21913 11296 21947
rect 11244 21904 11296 21913
rect 10416 21836 10468 21888
rect 11520 21879 11572 21888
rect 11520 21845 11529 21879
rect 11529 21845 11563 21879
rect 11563 21845 11572 21879
rect 11520 21836 11572 21845
rect 11888 21904 11940 21956
rect 13728 22108 13780 22160
rect 21640 22176 21692 22228
rect 22008 22176 22060 22228
rect 22284 22176 22336 22228
rect 29092 22176 29144 22228
rect 29276 22176 29328 22228
rect 29460 22176 29512 22228
rect 30472 22176 30524 22228
rect 30656 22176 30708 22228
rect 30840 22176 30892 22228
rect 31208 22176 31260 22228
rect 31576 22176 31628 22228
rect 35532 22176 35584 22228
rect 35808 22176 35860 22228
rect 39396 22176 39448 22228
rect 19340 22108 19392 22160
rect 12900 21836 12952 21888
rect 13084 21947 13136 21956
rect 13084 21913 13093 21947
rect 13093 21913 13127 21947
rect 13127 21913 13136 21947
rect 13084 21904 13136 21913
rect 13360 21904 13412 21956
rect 14096 22015 14148 22024
rect 14096 21981 14105 22015
rect 14105 21981 14139 22015
rect 14139 21981 14148 22015
rect 14096 21972 14148 21981
rect 17408 22083 17460 22092
rect 17408 22049 17417 22083
rect 17417 22049 17451 22083
rect 17451 22049 17460 22083
rect 17408 22040 17460 22049
rect 17316 21972 17368 22024
rect 17776 22015 17828 22024
rect 17776 21981 17785 22015
rect 17785 21981 17819 22015
rect 17819 21981 17828 22015
rect 17776 21972 17828 21981
rect 17960 22015 18012 22024
rect 17960 21981 17969 22015
rect 17969 21981 18003 22015
rect 18003 21981 18012 22015
rect 17960 21972 18012 21981
rect 18052 22015 18104 22024
rect 18052 21981 18061 22015
rect 18061 21981 18095 22015
rect 18095 21981 18104 22015
rect 18052 21972 18104 21981
rect 18420 21972 18472 22024
rect 18512 22015 18564 22024
rect 18512 21981 18521 22015
rect 18521 21981 18555 22015
rect 18555 21981 18564 22015
rect 18512 21972 18564 21981
rect 18696 21972 18748 22024
rect 18880 22015 18932 22024
rect 18880 21981 18889 22015
rect 18889 21981 18923 22015
rect 18923 21981 18932 22015
rect 18880 21972 18932 21981
rect 19892 22040 19944 22092
rect 13912 21879 13964 21888
rect 13912 21845 13921 21879
rect 13921 21845 13955 21879
rect 13955 21845 13964 21879
rect 13912 21836 13964 21845
rect 14280 21904 14332 21956
rect 14464 21947 14516 21956
rect 14464 21913 14473 21947
rect 14473 21913 14507 21947
rect 14507 21913 14516 21947
rect 14464 21904 14516 21913
rect 16488 21904 16540 21956
rect 17408 21904 17460 21956
rect 19156 21904 19208 21956
rect 20628 21972 20680 22024
rect 20168 21947 20220 21956
rect 20168 21913 20177 21947
rect 20177 21913 20211 21947
rect 20211 21913 20220 21947
rect 20168 21904 20220 21913
rect 19984 21836 20036 21888
rect 20444 21836 20496 21888
rect 20996 21972 21048 22024
rect 22100 22108 22152 22160
rect 23020 22108 23072 22160
rect 23204 22108 23256 22160
rect 24124 22108 24176 22160
rect 24860 22108 24912 22160
rect 25320 22151 25372 22160
rect 25320 22117 25329 22151
rect 25329 22117 25363 22151
rect 25363 22117 25372 22151
rect 25320 22108 25372 22117
rect 21824 21972 21876 22024
rect 22468 21972 22520 22024
rect 22836 21972 22888 22024
rect 23296 21972 23348 22024
rect 23940 22015 23992 22024
rect 23940 21981 23949 22015
rect 23949 21981 23983 22015
rect 23983 21981 23992 22015
rect 23940 21972 23992 21981
rect 24400 21972 24452 22024
rect 25504 22108 25556 22160
rect 26056 22108 26108 22160
rect 27068 22108 27120 22160
rect 20996 21836 21048 21888
rect 23572 21904 23624 21956
rect 23848 21904 23900 21956
rect 25228 21904 25280 21956
rect 21548 21836 21600 21888
rect 21640 21879 21692 21888
rect 21640 21845 21649 21879
rect 21649 21845 21683 21879
rect 21683 21845 21692 21879
rect 21640 21836 21692 21845
rect 21732 21836 21784 21888
rect 22008 21836 22060 21888
rect 22468 21879 22520 21888
rect 22468 21845 22477 21879
rect 22477 21845 22511 21879
rect 22511 21845 22520 21879
rect 22468 21836 22520 21845
rect 23020 21836 23072 21888
rect 24400 21879 24452 21888
rect 24400 21845 24409 21879
rect 24409 21845 24443 21879
rect 24443 21845 24452 21879
rect 24400 21836 24452 21845
rect 25596 21836 25648 21888
rect 25780 22015 25832 22024
rect 25780 21981 25789 22015
rect 25789 21981 25823 22015
rect 25823 21981 25832 22015
rect 25780 21972 25832 21981
rect 25964 22015 26016 22024
rect 25964 21981 25973 22015
rect 25973 21981 26007 22015
rect 26007 21981 26016 22015
rect 25964 21972 26016 21981
rect 26332 21972 26384 22024
rect 26424 21972 26476 22024
rect 29552 22108 29604 22160
rect 29276 22040 29328 22092
rect 27068 22015 27120 22024
rect 27068 21981 27077 22015
rect 27077 21981 27111 22015
rect 27111 21981 27120 22015
rect 27068 21972 27120 21981
rect 26056 21904 26108 21956
rect 27344 21972 27396 22024
rect 27436 21904 27488 21956
rect 27620 21947 27672 21956
rect 27620 21913 27629 21947
rect 27629 21913 27663 21947
rect 27663 21913 27672 21947
rect 27620 21904 27672 21913
rect 27988 22015 28040 22024
rect 27988 21981 27997 22015
rect 27997 21981 28031 22015
rect 28031 21981 28040 22015
rect 27988 21972 28040 21981
rect 28264 22015 28316 22024
rect 28264 21981 28273 22015
rect 28273 21981 28307 22015
rect 28307 21981 28316 22015
rect 28264 21972 28316 21981
rect 28540 22015 28592 22024
rect 28540 21981 28549 22015
rect 28549 21981 28583 22015
rect 28583 21981 28592 22015
rect 28540 21972 28592 21981
rect 28632 22015 28684 22024
rect 28632 21981 28641 22015
rect 28641 21981 28675 22015
rect 28675 21981 28684 22015
rect 28632 21972 28684 21981
rect 30932 22040 30984 22092
rect 32036 22108 32088 22160
rect 33324 22108 33376 22160
rect 28724 21904 28776 21956
rect 29092 21904 29144 21956
rect 30104 21972 30156 22024
rect 30380 21972 30432 22024
rect 31576 22015 31628 22024
rect 31576 21981 31585 22015
rect 31585 21981 31619 22015
rect 31619 21981 31628 22015
rect 31576 21972 31628 21981
rect 32680 21972 32732 22024
rect 33876 22015 33928 22024
rect 33876 21981 33885 22015
rect 33885 21981 33919 22015
rect 33919 21981 33928 22015
rect 33876 21972 33928 21981
rect 34336 22015 34388 22024
rect 34336 21981 34345 22015
rect 34345 21981 34379 22015
rect 34379 21981 34388 22015
rect 34336 21972 34388 21981
rect 28080 21879 28132 21888
rect 28080 21845 28089 21879
rect 28089 21845 28123 21879
rect 28123 21845 28132 21879
rect 28080 21836 28132 21845
rect 29552 21836 29604 21888
rect 30656 21904 30708 21956
rect 33324 21904 33376 21956
rect 33968 21947 34020 21956
rect 33968 21913 33977 21947
rect 33977 21913 34011 21947
rect 34011 21913 34020 21947
rect 33968 21904 34020 21913
rect 31300 21836 31352 21888
rect 31944 21836 31996 21888
rect 34520 21836 34572 21888
rect 36360 21836 36412 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 2504 21632 2556 21684
rect 3240 21564 3292 21616
rect 5632 21632 5684 21684
rect 7656 21632 7708 21684
rect 8208 21632 8260 21684
rect 5172 21564 5224 21616
rect 5448 21564 5500 21616
rect 2688 21471 2740 21480
rect 2688 21437 2697 21471
rect 2697 21437 2731 21471
rect 2731 21437 2740 21471
rect 2688 21428 2740 21437
rect 4068 21360 4120 21412
rect 7564 21496 7616 21548
rect 9220 21632 9272 21684
rect 9312 21632 9364 21684
rect 9772 21632 9824 21684
rect 11428 21632 11480 21684
rect 11520 21632 11572 21684
rect 8484 21564 8536 21616
rect 8852 21539 8904 21548
rect 8852 21505 8861 21539
rect 8861 21505 8895 21539
rect 8895 21505 8904 21539
rect 8852 21496 8904 21505
rect 1860 21335 1912 21344
rect 1860 21301 1869 21335
rect 1869 21301 1903 21335
rect 1903 21301 1912 21335
rect 1860 21292 1912 21301
rect 2688 21292 2740 21344
rect 4160 21292 4212 21344
rect 5908 21292 5960 21344
rect 6276 21292 6328 21344
rect 6920 21360 6972 21412
rect 9588 21496 9640 21548
rect 9680 21496 9732 21548
rect 10876 21564 10928 21616
rect 10416 21539 10468 21548
rect 10416 21505 10425 21539
rect 10425 21505 10459 21539
rect 10459 21505 10468 21539
rect 10416 21496 10468 21505
rect 10508 21539 10560 21548
rect 10508 21505 10517 21539
rect 10517 21505 10551 21539
rect 10551 21505 10560 21539
rect 10508 21496 10560 21505
rect 10692 21496 10744 21548
rect 13912 21564 13964 21616
rect 14004 21496 14056 21548
rect 14280 21496 14332 21548
rect 11612 21428 11664 21480
rect 12072 21428 12124 21480
rect 15752 21632 15804 21684
rect 16396 21632 16448 21684
rect 17776 21632 17828 21684
rect 19064 21632 19116 21684
rect 19524 21632 19576 21684
rect 20996 21632 21048 21684
rect 15660 21564 15712 21616
rect 17960 21496 18012 21548
rect 15384 21428 15436 21480
rect 15476 21471 15528 21480
rect 15476 21437 15485 21471
rect 15485 21437 15519 21471
rect 15519 21437 15528 21471
rect 15476 21428 15528 21437
rect 15752 21471 15804 21480
rect 15752 21437 15761 21471
rect 15761 21437 15795 21471
rect 15795 21437 15804 21471
rect 15752 21428 15804 21437
rect 19340 21564 19392 21616
rect 20168 21564 20220 21616
rect 18972 21539 19024 21548
rect 18972 21505 18981 21539
rect 18981 21505 19015 21539
rect 19015 21505 19024 21539
rect 18972 21496 19024 21505
rect 19432 21496 19484 21548
rect 20720 21564 20772 21616
rect 21180 21632 21232 21684
rect 22928 21632 22980 21684
rect 23848 21632 23900 21684
rect 24400 21632 24452 21684
rect 27160 21632 27212 21684
rect 27436 21632 27488 21684
rect 28632 21632 28684 21684
rect 29184 21632 29236 21684
rect 29736 21632 29788 21684
rect 30840 21632 30892 21684
rect 34060 21632 34112 21684
rect 8852 21292 8904 21344
rect 11980 21360 12032 21412
rect 12992 21360 13044 21412
rect 13636 21403 13688 21412
rect 13636 21369 13645 21403
rect 13645 21369 13679 21403
rect 13679 21369 13688 21403
rect 13636 21360 13688 21369
rect 18512 21428 18564 21480
rect 19064 21360 19116 21412
rect 13820 21292 13872 21344
rect 14464 21292 14516 21344
rect 15752 21292 15804 21344
rect 16120 21335 16172 21344
rect 16120 21301 16129 21335
rect 16129 21301 16163 21335
rect 16163 21301 16172 21335
rect 16120 21292 16172 21301
rect 19248 21292 19300 21344
rect 20076 21292 20128 21344
rect 20720 21428 20772 21480
rect 21272 21539 21324 21548
rect 21272 21505 21281 21539
rect 21281 21505 21315 21539
rect 21315 21505 21324 21539
rect 21272 21496 21324 21505
rect 21824 21539 21876 21548
rect 21824 21505 21833 21539
rect 21833 21505 21867 21539
rect 21867 21505 21876 21539
rect 21824 21496 21876 21505
rect 20444 21360 20496 21412
rect 23572 21564 23624 21616
rect 22192 21539 22244 21548
rect 22192 21505 22201 21539
rect 22201 21505 22235 21539
rect 22235 21505 22244 21539
rect 22192 21496 22244 21505
rect 22744 21496 22796 21548
rect 23848 21496 23900 21548
rect 25964 21564 26016 21616
rect 25412 21496 25464 21548
rect 21640 21292 21692 21344
rect 22744 21360 22796 21412
rect 23020 21360 23072 21412
rect 24400 21428 24452 21480
rect 25504 21428 25556 21480
rect 24860 21360 24912 21412
rect 27068 21564 27120 21616
rect 26332 21428 26384 21480
rect 26700 21428 26752 21480
rect 23940 21292 23992 21344
rect 24216 21335 24268 21344
rect 24216 21301 24225 21335
rect 24225 21301 24259 21335
rect 24259 21301 24268 21335
rect 24216 21292 24268 21301
rect 24400 21335 24452 21344
rect 24400 21301 24409 21335
rect 24409 21301 24443 21335
rect 24443 21301 24452 21335
rect 24400 21292 24452 21301
rect 25044 21292 25096 21344
rect 25780 21292 25832 21344
rect 27068 21292 27120 21344
rect 27804 21564 27856 21616
rect 27988 21564 28040 21616
rect 27712 21496 27764 21548
rect 28080 21539 28132 21548
rect 28080 21505 28089 21539
rect 28089 21505 28123 21539
rect 28123 21505 28132 21539
rect 28080 21496 28132 21505
rect 28540 21496 28592 21548
rect 34336 21564 34388 21616
rect 34704 21564 34756 21616
rect 35348 21607 35400 21616
rect 35348 21573 35357 21607
rect 35357 21573 35391 21607
rect 35391 21573 35400 21607
rect 35348 21564 35400 21573
rect 36360 21632 36412 21684
rect 38016 21632 38068 21684
rect 39028 21632 39080 21684
rect 39948 21632 40000 21684
rect 40868 21675 40920 21684
rect 40868 21641 40877 21675
rect 40877 21641 40911 21675
rect 40911 21641 40920 21675
rect 40868 21632 40920 21641
rect 30104 21496 30156 21548
rect 31392 21496 31444 21548
rect 33140 21496 33192 21548
rect 36636 21564 36688 21616
rect 37280 21607 37332 21616
rect 37280 21573 37289 21607
rect 37289 21573 37323 21607
rect 37323 21573 37332 21607
rect 37280 21564 37332 21573
rect 28264 21428 28316 21480
rect 31760 21428 31812 21480
rect 28448 21360 28500 21412
rect 29460 21360 29512 21412
rect 31116 21360 31168 21412
rect 31300 21360 31352 21412
rect 31392 21360 31444 21412
rect 27804 21292 27856 21344
rect 28908 21335 28960 21344
rect 28908 21301 28917 21335
rect 28917 21301 28951 21335
rect 28951 21301 28960 21335
rect 28908 21292 28960 21301
rect 35348 21428 35400 21480
rect 35624 21428 35676 21480
rect 37464 21496 37516 21548
rect 38844 21496 38896 21548
rect 41420 21496 41472 21548
rect 37372 21471 37424 21480
rect 37372 21437 37381 21471
rect 37381 21437 37415 21471
rect 37415 21437 37424 21471
rect 37372 21428 37424 21437
rect 38660 21428 38712 21480
rect 38476 21360 38528 21412
rect 35440 21292 35492 21344
rect 35532 21292 35584 21344
rect 37648 21292 37700 21344
rect 37832 21292 37884 21344
rect 38568 21292 38620 21344
rect 39212 21292 39264 21344
rect 39304 21335 39356 21344
rect 39304 21301 39313 21335
rect 39313 21301 39347 21335
rect 39347 21301 39356 21335
rect 39304 21292 39356 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1860 21088 1912 21140
rect 3240 21088 3292 21140
rect 1400 20995 1452 21004
rect 1400 20961 1409 20995
rect 1409 20961 1443 20995
rect 1443 20961 1452 20995
rect 1400 20952 1452 20961
rect 2688 20952 2740 21004
rect 3148 20995 3200 21004
rect 3148 20961 3157 20995
rect 3157 20961 3191 20995
rect 3191 20961 3200 20995
rect 3148 20952 3200 20961
rect 3056 20816 3108 20868
rect 4068 20952 4120 21004
rect 7656 21131 7708 21140
rect 7656 21097 7665 21131
rect 7665 21097 7699 21131
rect 7699 21097 7708 21131
rect 7656 21088 7708 21097
rect 10508 21088 10560 21140
rect 11520 21088 11572 21140
rect 14556 21131 14608 21140
rect 14556 21097 14565 21131
rect 14565 21097 14599 21131
rect 14599 21097 14608 21131
rect 14556 21088 14608 21097
rect 7932 21020 7984 21072
rect 5172 20884 5224 20936
rect 5356 20884 5408 20936
rect 5908 20995 5960 21004
rect 5908 20961 5917 20995
rect 5917 20961 5951 20995
rect 5951 20961 5960 20995
rect 5908 20952 5960 20961
rect 6276 20952 6328 21004
rect 9404 20952 9456 21004
rect 15568 21088 15620 21140
rect 15476 21020 15528 21072
rect 16856 21088 16908 21140
rect 17684 21088 17736 21140
rect 18972 21088 19024 21140
rect 20076 21088 20128 21140
rect 21732 21088 21784 21140
rect 21916 21088 21968 21140
rect 15752 21020 15804 21072
rect 16028 21020 16080 21072
rect 16212 21020 16264 21072
rect 23204 21020 23256 21072
rect 24216 21088 24268 21140
rect 24400 21088 24452 21140
rect 27344 21088 27396 21140
rect 27528 21088 27580 21140
rect 28172 21088 28224 21140
rect 30932 21131 30984 21140
rect 30932 21097 30941 21131
rect 30941 21097 30975 21131
rect 30975 21097 30984 21131
rect 30932 21088 30984 21097
rect 31760 21088 31812 21140
rect 32496 21088 32548 21140
rect 32864 21088 32916 21140
rect 36084 21088 36136 21140
rect 36268 21088 36320 21140
rect 36728 21088 36780 21140
rect 36912 21088 36964 21140
rect 15384 20952 15436 21004
rect 5816 20884 5868 20936
rect 7288 20884 7340 20936
rect 10876 20884 10928 20936
rect 11336 20884 11388 20936
rect 12440 20884 12492 20936
rect 16856 20884 16908 20936
rect 19156 20952 19208 21004
rect 19432 20952 19484 21004
rect 20260 20952 20312 21004
rect 21824 20952 21876 21004
rect 22100 20952 22152 21004
rect 22284 20952 22336 21004
rect 4712 20748 4764 20800
rect 5080 20748 5132 20800
rect 5632 20748 5684 20800
rect 6000 20748 6052 20800
rect 7748 20748 7800 20800
rect 8392 20748 8444 20800
rect 10968 20748 11020 20800
rect 11888 20748 11940 20800
rect 12164 20748 12216 20800
rect 15660 20816 15712 20868
rect 16212 20816 16264 20868
rect 16672 20859 16724 20868
rect 16672 20825 16681 20859
rect 16681 20825 16715 20859
rect 16715 20825 16724 20859
rect 16672 20816 16724 20825
rect 15752 20748 15804 20800
rect 19248 20927 19300 20936
rect 19248 20893 19257 20927
rect 19257 20893 19291 20927
rect 19291 20893 19300 20927
rect 19248 20884 19300 20893
rect 20628 20884 20680 20936
rect 22008 20884 22060 20936
rect 22376 20816 22428 20868
rect 22928 20927 22980 20936
rect 22928 20893 22937 20927
rect 22937 20893 22971 20927
rect 22971 20893 22980 20927
rect 22928 20884 22980 20893
rect 23112 20884 23164 20936
rect 23664 20952 23716 21004
rect 24860 20952 24912 21004
rect 25780 20952 25832 21004
rect 23940 20884 23992 20936
rect 26516 20884 26568 20936
rect 27988 20952 28040 21004
rect 30196 20952 30248 21004
rect 27068 20884 27120 20936
rect 29828 20927 29880 20936
rect 29828 20893 29837 20927
rect 29837 20893 29871 20927
rect 29871 20893 29880 20927
rect 29828 20884 29880 20893
rect 30288 20884 30340 20936
rect 30380 20884 30432 20936
rect 30656 20884 30708 20936
rect 17132 20748 17184 20800
rect 21640 20791 21692 20800
rect 21640 20757 21649 20791
rect 21649 20757 21683 20791
rect 21683 20757 21692 20791
rect 21640 20748 21692 20757
rect 22468 20748 22520 20800
rect 24952 20748 25004 20800
rect 29644 20791 29696 20800
rect 29644 20757 29653 20791
rect 29653 20757 29687 20791
rect 29687 20757 29696 20791
rect 29644 20748 29696 20757
rect 30932 20884 30984 20936
rect 31208 20884 31260 20936
rect 31116 20748 31168 20800
rect 31576 20859 31628 20868
rect 31576 20825 31585 20859
rect 31585 20825 31619 20859
rect 31619 20825 31628 20859
rect 31576 20816 31628 20825
rect 31944 20816 31996 20868
rect 31392 20748 31444 20800
rect 32496 20927 32548 20936
rect 32496 20893 32505 20927
rect 32505 20893 32539 20927
rect 32539 20893 32548 20927
rect 32496 20884 32548 20893
rect 32220 20816 32272 20868
rect 32588 20748 32640 20800
rect 33140 20884 33192 20936
rect 37280 21020 37332 21072
rect 37464 21020 37516 21072
rect 38568 21088 38620 21140
rect 39212 21088 39264 21140
rect 38292 21020 38344 21072
rect 35440 20884 35492 20936
rect 35532 20927 35584 20936
rect 35532 20893 35541 20927
rect 35541 20893 35575 20927
rect 35575 20893 35584 20927
rect 35532 20884 35584 20893
rect 34704 20816 34756 20868
rect 32864 20748 32916 20800
rect 33416 20748 33468 20800
rect 33876 20748 33928 20800
rect 34520 20748 34572 20800
rect 35900 20927 35952 20936
rect 35900 20893 35909 20927
rect 35909 20893 35943 20927
rect 35943 20893 35952 20927
rect 35900 20884 35952 20893
rect 36360 20884 36412 20936
rect 36728 20884 36780 20936
rect 35716 20816 35768 20868
rect 37188 20816 37240 20868
rect 37464 20927 37516 20936
rect 37464 20893 37474 20927
rect 37474 20893 37508 20927
rect 37508 20893 37516 20927
rect 37464 20884 37516 20893
rect 37740 20927 37792 20936
rect 37740 20893 37749 20927
rect 37749 20893 37783 20927
rect 37783 20893 37792 20927
rect 37740 20884 37792 20893
rect 38016 20884 38068 20936
rect 36636 20748 36688 20800
rect 38936 20995 38988 21004
rect 38936 20961 38945 20995
rect 38945 20961 38979 20995
rect 38979 20961 38988 20995
rect 38936 20952 38988 20961
rect 39488 20952 39540 21004
rect 39764 20952 39816 21004
rect 39672 20884 39724 20936
rect 39856 20927 39908 20936
rect 39856 20893 39865 20927
rect 39865 20893 39899 20927
rect 39899 20893 39908 20927
rect 39856 20884 39908 20893
rect 38016 20791 38068 20800
rect 38016 20757 38025 20791
rect 38025 20757 38059 20791
rect 38059 20757 38068 20791
rect 38016 20748 38068 20757
rect 39212 20791 39264 20800
rect 39212 20757 39221 20791
rect 39221 20757 39255 20791
rect 39255 20757 39264 20791
rect 39212 20748 39264 20757
rect 40776 20791 40828 20800
rect 40776 20757 40785 20791
rect 40785 20757 40819 20791
rect 40819 20757 40828 20791
rect 40776 20748 40828 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 5816 20587 5868 20596
rect 5816 20553 5825 20587
rect 5825 20553 5859 20587
rect 5859 20553 5868 20587
rect 5816 20544 5868 20553
rect 7656 20544 7708 20596
rect 2964 20476 3016 20528
rect 5908 20476 5960 20528
rect 6828 20476 6880 20528
rect 2596 20408 2648 20460
rect 4988 20408 5040 20460
rect 2688 20340 2740 20392
rect 3424 20204 3476 20256
rect 3608 20204 3660 20256
rect 5356 20408 5408 20460
rect 6000 20408 6052 20460
rect 6920 20340 6972 20392
rect 7656 20451 7708 20460
rect 7656 20417 7665 20451
rect 7665 20417 7699 20451
rect 7699 20417 7708 20451
rect 7656 20408 7708 20417
rect 7748 20408 7800 20460
rect 8024 20451 8076 20460
rect 8024 20417 8033 20451
rect 8033 20417 8067 20451
rect 8067 20417 8076 20451
rect 8024 20408 8076 20417
rect 9864 20587 9916 20596
rect 9864 20553 9873 20587
rect 9873 20553 9907 20587
rect 9907 20553 9916 20587
rect 9864 20544 9916 20553
rect 10324 20544 10376 20596
rect 10968 20544 11020 20596
rect 9956 20476 10008 20528
rect 9220 20451 9272 20460
rect 9220 20417 9229 20451
rect 9229 20417 9263 20451
rect 9263 20417 9272 20451
rect 9220 20408 9272 20417
rect 10508 20408 10560 20460
rect 12348 20544 12400 20596
rect 7748 20272 7800 20324
rect 8024 20272 8076 20324
rect 9864 20340 9916 20392
rect 11796 20408 11848 20460
rect 13084 20476 13136 20528
rect 13912 20476 13964 20528
rect 14832 20587 14884 20596
rect 14832 20553 14841 20587
rect 14841 20553 14875 20587
rect 14875 20553 14884 20587
rect 14832 20544 14884 20553
rect 15936 20544 15988 20596
rect 19984 20544 20036 20596
rect 22928 20544 22980 20596
rect 25228 20544 25280 20596
rect 25964 20544 26016 20596
rect 26608 20544 26660 20596
rect 15660 20519 15712 20528
rect 11704 20340 11756 20392
rect 12164 20451 12216 20460
rect 12164 20417 12173 20451
rect 12173 20417 12207 20451
rect 12207 20417 12216 20451
rect 12164 20408 12216 20417
rect 12348 20408 12400 20460
rect 12716 20451 12768 20460
rect 12716 20417 12725 20451
rect 12725 20417 12759 20451
rect 12759 20417 12768 20451
rect 12716 20408 12768 20417
rect 15660 20485 15669 20519
rect 15669 20485 15703 20519
rect 15703 20485 15712 20519
rect 15660 20476 15712 20485
rect 15752 20476 15804 20528
rect 16672 20476 16724 20528
rect 19432 20476 19484 20528
rect 20076 20476 20128 20528
rect 15384 20408 15436 20460
rect 15476 20451 15528 20460
rect 15476 20417 15485 20451
rect 15485 20417 15519 20451
rect 15519 20417 15528 20451
rect 15476 20408 15528 20417
rect 21456 20476 21508 20528
rect 26148 20476 26200 20528
rect 26240 20476 26292 20528
rect 16120 20451 16172 20460
rect 16120 20417 16129 20451
rect 16129 20417 16163 20451
rect 16163 20417 16172 20451
rect 16120 20408 16172 20417
rect 17408 20451 17460 20460
rect 17408 20417 17417 20451
rect 17417 20417 17451 20451
rect 17451 20417 17460 20451
rect 17408 20408 17460 20417
rect 20444 20408 20496 20460
rect 8208 20247 8260 20256
rect 8208 20213 8217 20247
rect 8217 20213 8251 20247
rect 8251 20213 8260 20247
rect 8208 20204 8260 20213
rect 8576 20247 8628 20256
rect 8576 20213 8585 20247
rect 8585 20213 8619 20247
rect 8619 20213 8628 20247
rect 8576 20204 8628 20213
rect 10416 20204 10468 20256
rect 10600 20247 10652 20256
rect 10600 20213 10609 20247
rect 10609 20213 10643 20247
rect 10643 20213 10652 20247
rect 10600 20204 10652 20213
rect 11612 20204 11664 20256
rect 11796 20204 11848 20256
rect 12624 20272 12676 20324
rect 12532 20247 12584 20256
rect 12532 20213 12541 20247
rect 12541 20213 12575 20247
rect 12575 20213 12584 20247
rect 12532 20204 12584 20213
rect 13084 20383 13136 20392
rect 13084 20349 13093 20383
rect 13093 20349 13127 20383
rect 13127 20349 13136 20383
rect 13084 20340 13136 20349
rect 13360 20383 13412 20392
rect 13360 20349 13369 20383
rect 13369 20349 13403 20383
rect 13403 20349 13412 20383
rect 13360 20340 13412 20349
rect 15844 20340 15896 20392
rect 19064 20340 19116 20392
rect 20168 20340 20220 20392
rect 20996 20340 21048 20392
rect 21088 20340 21140 20392
rect 23296 20408 23348 20460
rect 23572 20408 23624 20460
rect 24400 20408 24452 20460
rect 27436 20451 27488 20460
rect 27436 20417 27445 20451
rect 27445 20417 27479 20451
rect 27479 20417 27488 20451
rect 27436 20408 27488 20417
rect 28172 20519 28224 20528
rect 28172 20485 28181 20519
rect 28181 20485 28215 20519
rect 28215 20485 28224 20519
rect 28172 20476 28224 20485
rect 28356 20519 28408 20528
rect 28356 20485 28381 20519
rect 28381 20485 28408 20519
rect 35624 20544 35676 20596
rect 37464 20544 37516 20596
rect 38936 20544 38988 20596
rect 39212 20544 39264 20596
rect 40040 20544 40092 20596
rect 28356 20476 28408 20485
rect 30012 20476 30064 20528
rect 15016 20272 15068 20324
rect 16396 20272 16448 20324
rect 19340 20272 19392 20324
rect 19984 20315 20036 20324
rect 19984 20281 19993 20315
rect 19993 20281 20027 20315
rect 20027 20281 20036 20315
rect 19984 20272 20036 20281
rect 26884 20340 26936 20392
rect 23480 20272 23532 20324
rect 26240 20272 26292 20324
rect 15200 20204 15252 20256
rect 16304 20204 16356 20256
rect 16856 20247 16908 20256
rect 16856 20213 16865 20247
rect 16865 20213 16899 20247
rect 16899 20213 16908 20247
rect 16856 20204 16908 20213
rect 17224 20247 17276 20256
rect 17224 20213 17233 20247
rect 17233 20213 17267 20247
rect 17267 20213 17276 20247
rect 17224 20204 17276 20213
rect 20260 20204 20312 20256
rect 20904 20204 20956 20256
rect 22376 20204 22428 20256
rect 23020 20204 23072 20256
rect 26056 20204 26108 20256
rect 31576 20451 31628 20460
rect 31576 20417 31585 20451
rect 31585 20417 31619 20451
rect 31619 20417 31628 20451
rect 31576 20408 31628 20417
rect 27620 20272 27672 20324
rect 31300 20340 31352 20392
rect 31392 20383 31444 20392
rect 31392 20349 31401 20383
rect 31401 20349 31435 20383
rect 31435 20349 31444 20383
rect 32036 20476 32088 20528
rect 33416 20476 33468 20528
rect 31392 20340 31444 20349
rect 34060 20340 34112 20392
rect 37372 20408 37424 20460
rect 27896 20272 27948 20324
rect 28448 20272 28500 20324
rect 34152 20272 34204 20324
rect 27804 20247 27856 20256
rect 27804 20213 27813 20247
rect 27813 20213 27847 20247
rect 27847 20213 27856 20247
rect 27804 20204 27856 20213
rect 29000 20204 29052 20256
rect 29276 20204 29328 20256
rect 29552 20204 29604 20256
rect 29828 20204 29880 20256
rect 30656 20204 30708 20256
rect 31484 20204 31536 20256
rect 31576 20204 31628 20256
rect 33416 20204 33468 20256
rect 33784 20204 33836 20256
rect 36084 20204 36136 20256
rect 36544 20204 36596 20256
rect 37372 20204 37424 20256
rect 37556 20451 37608 20460
rect 37556 20417 37565 20451
rect 37565 20417 37599 20451
rect 37599 20417 37608 20451
rect 37556 20408 37608 20417
rect 39764 20408 39816 20460
rect 41236 20408 41288 20460
rect 38844 20340 38896 20392
rect 39580 20204 39632 20256
rect 40776 20204 40828 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 3608 20000 3660 20052
rect 3976 20000 4028 20052
rect 1400 19907 1452 19916
rect 1400 19873 1409 19907
rect 1409 19873 1443 19907
rect 1443 19873 1452 19907
rect 1400 19864 1452 19873
rect 3792 19932 3844 19984
rect 5724 20000 5776 20052
rect 5816 20000 5868 20052
rect 3976 19839 4028 19848
rect 3976 19805 3985 19839
rect 3985 19805 4019 19839
rect 4019 19805 4028 19839
rect 3976 19796 4028 19805
rect 4252 19839 4304 19848
rect 4252 19805 4261 19839
rect 4261 19805 4295 19839
rect 4295 19805 4304 19839
rect 4252 19796 4304 19805
rect 8208 20000 8260 20052
rect 8300 20000 8352 20052
rect 8484 20000 8536 20052
rect 8024 19932 8076 19984
rect 10232 19932 10284 19984
rect 1676 19771 1728 19780
rect 1676 19737 1685 19771
rect 1685 19737 1719 19771
rect 1719 19737 1728 19771
rect 1676 19728 1728 19737
rect 3056 19728 3108 19780
rect 4436 19728 4488 19780
rect 5080 19839 5132 19848
rect 5080 19805 5090 19839
rect 5090 19805 5124 19839
rect 5124 19805 5132 19839
rect 5080 19796 5132 19805
rect 5724 19796 5776 19848
rect 7840 19839 7892 19848
rect 7840 19805 7850 19839
rect 7850 19805 7884 19839
rect 7884 19805 7892 19839
rect 7840 19796 7892 19805
rect 3608 19660 3660 19712
rect 5172 19660 5224 19712
rect 5356 19771 5408 19780
rect 5356 19737 5365 19771
rect 5365 19737 5399 19771
rect 5399 19737 5408 19771
rect 5356 19728 5408 19737
rect 5816 19728 5868 19780
rect 7012 19728 7064 19780
rect 8484 19796 8536 19848
rect 8760 19796 8812 19848
rect 9036 19839 9088 19848
rect 9036 19805 9045 19839
rect 9045 19805 9079 19839
rect 9079 19805 9088 19839
rect 9036 19796 9088 19805
rect 9404 19839 9456 19848
rect 9404 19805 9413 19839
rect 9413 19805 9447 19839
rect 9447 19805 9456 19839
rect 9404 19796 9456 19805
rect 9588 19796 9640 19848
rect 6828 19660 6880 19712
rect 8116 19771 8168 19780
rect 8116 19737 8125 19771
rect 8125 19737 8159 19771
rect 8159 19737 8168 19771
rect 8116 19728 8168 19737
rect 8944 19728 8996 19780
rect 9496 19660 9548 19712
rect 10416 19907 10468 19916
rect 10416 19873 10425 19907
rect 10425 19873 10459 19907
rect 10459 19873 10468 19907
rect 10416 19864 10468 19873
rect 9956 19796 10008 19848
rect 11060 19932 11112 19984
rect 13084 20000 13136 20052
rect 13360 20000 13412 20052
rect 17224 20043 17276 20052
rect 17224 20009 17254 20043
rect 17254 20009 17276 20043
rect 17224 20000 17276 20009
rect 17316 20000 17368 20052
rect 12532 19864 12584 19916
rect 10784 19796 10836 19848
rect 11520 19839 11572 19848
rect 11520 19805 11529 19839
rect 11529 19805 11563 19839
rect 11563 19805 11572 19839
rect 11520 19796 11572 19805
rect 14740 19907 14792 19916
rect 14740 19873 14749 19907
rect 14749 19873 14783 19907
rect 14783 19873 14792 19907
rect 14740 19864 14792 19873
rect 14832 19864 14884 19916
rect 17868 19864 17920 19916
rect 19064 19932 19116 19984
rect 19708 19975 19760 19984
rect 19708 19941 19717 19975
rect 19717 19941 19751 19975
rect 19751 19941 19760 19975
rect 19708 19932 19760 19941
rect 21456 20000 21508 20052
rect 22192 20000 22244 20052
rect 24676 20000 24728 20052
rect 19340 19864 19392 19916
rect 20168 19864 20220 19916
rect 20628 19864 20680 19916
rect 27620 19932 27672 19984
rect 28172 20043 28224 20052
rect 28172 20009 28181 20043
rect 28181 20009 28215 20043
rect 28215 20009 28224 20043
rect 28172 20000 28224 20009
rect 28908 20000 28960 20052
rect 30656 20000 30708 20052
rect 31024 20000 31076 20052
rect 34060 20000 34112 20052
rect 34336 20000 34388 20052
rect 34612 20000 34664 20052
rect 20812 19864 20864 19916
rect 24768 19864 24820 19916
rect 15200 19839 15252 19848
rect 15200 19805 15209 19839
rect 15209 19805 15243 19839
rect 15243 19805 15252 19839
rect 15200 19796 15252 19805
rect 16028 19796 16080 19848
rect 19616 19839 19668 19848
rect 19616 19805 19625 19839
rect 19625 19805 19659 19839
rect 19659 19805 19668 19839
rect 19616 19796 19668 19805
rect 13912 19728 13964 19780
rect 16948 19728 17000 19780
rect 20996 19796 21048 19848
rect 22284 19796 22336 19848
rect 23848 19839 23900 19848
rect 23848 19805 23857 19839
rect 23857 19805 23891 19839
rect 23891 19805 23900 19839
rect 23848 19796 23900 19805
rect 24032 19796 24084 19848
rect 25780 19864 25832 19916
rect 25136 19839 25188 19848
rect 25136 19805 25143 19839
rect 25143 19805 25188 19839
rect 25136 19796 25188 19805
rect 25596 19796 25648 19848
rect 25872 19796 25924 19848
rect 11796 19660 11848 19712
rect 13360 19703 13412 19712
rect 13360 19669 13369 19703
rect 13369 19669 13403 19703
rect 13403 19669 13412 19703
rect 13360 19660 13412 19669
rect 14372 19660 14424 19712
rect 14556 19660 14608 19712
rect 15752 19660 15804 19712
rect 17960 19660 18012 19712
rect 18144 19660 18196 19712
rect 23940 19728 23992 19780
rect 19432 19703 19484 19712
rect 19432 19669 19441 19703
rect 19441 19669 19475 19703
rect 19475 19669 19484 19703
rect 19432 19660 19484 19669
rect 20444 19703 20496 19712
rect 20444 19669 20453 19703
rect 20453 19669 20487 19703
rect 20487 19669 20496 19703
rect 20444 19660 20496 19669
rect 20536 19660 20588 19712
rect 20720 19660 20772 19712
rect 23020 19660 23072 19712
rect 23388 19703 23440 19712
rect 23388 19669 23397 19703
rect 23397 19669 23431 19703
rect 23431 19669 23440 19703
rect 23388 19660 23440 19669
rect 27528 19728 27580 19780
rect 28448 19796 28500 19848
rect 28816 19796 28868 19848
rect 29000 19932 29052 19984
rect 29368 19839 29420 19848
rect 29368 19805 29389 19839
rect 29389 19805 29420 19839
rect 29368 19796 29420 19805
rect 25412 19660 25464 19712
rect 27436 19660 27488 19712
rect 27712 19660 27764 19712
rect 28356 19660 28408 19712
rect 29276 19728 29328 19780
rect 29552 19975 29604 19984
rect 29552 19941 29561 19975
rect 29561 19941 29595 19975
rect 29595 19941 29604 19975
rect 29552 19932 29604 19941
rect 30012 19932 30064 19984
rect 33784 19932 33836 19984
rect 29828 19839 29880 19848
rect 29828 19805 29837 19839
rect 29837 19805 29871 19839
rect 29871 19805 29880 19839
rect 29828 19796 29880 19805
rect 29920 19839 29972 19848
rect 29920 19805 29929 19839
rect 29929 19805 29963 19839
rect 29963 19805 29972 19839
rect 29920 19796 29972 19805
rect 30380 19864 30432 19916
rect 31300 19864 31352 19916
rect 31392 19864 31444 19916
rect 30840 19796 30892 19848
rect 31484 19839 31536 19848
rect 31484 19805 31493 19839
rect 31493 19805 31527 19839
rect 31527 19805 31536 19839
rect 31484 19796 31536 19805
rect 31576 19771 31628 19780
rect 31576 19737 31585 19771
rect 31585 19737 31619 19771
rect 31619 19737 31628 19771
rect 31576 19728 31628 19737
rect 33416 19864 33468 19916
rect 34060 19907 34112 19916
rect 34060 19873 34069 19907
rect 34069 19873 34103 19907
rect 34103 19873 34112 19907
rect 34060 19864 34112 19873
rect 34152 19907 34204 19916
rect 34152 19873 34161 19907
rect 34161 19873 34195 19907
rect 34195 19873 34204 19907
rect 34152 19864 34204 19873
rect 32036 19796 32088 19848
rect 32220 19796 32272 19848
rect 32772 19796 32824 19848
rect 33784 19839 33836 19848
rect 33784 19805 33793 19839
rect 33793 19805 33827 19839
rect 33827 19805 33836 19839
rect 33784 19796 33836 19805
rect 33876 19796 33928 19848
rect 34336 19839 34388 19848
rect 34336 19805 34345 19839
rect 34345 19805 34379 19839
rect 34379 19805 34388 19839
rect 34336 19796 34388 19805
rect 34520 19796 34572 19848
rect 35440 19796 35492 19848
rect 35900 19796 35952 19848
rect 40500 19796 40552 19848
rect 33416 19771 33468 19780
rect 33416 19737 33425 19771
rect 33425 19737 33459 19771
rect 33459 19737 33468 19771
rect 33416 19728 33468 19737
rect 29828 19660 29880 19712
rect 30012 19660 30064 19712
rect 30656 19660 30708 19712
rect 32220 19660 32272 19712
rect 33140 19703 33192 19712
rect 33140 19669 33149 19703
rect 33149 19669 33183 19703
rect 33183 19669 33192 19703
rect 33140 19660 33192 19669
rect 33324 19660 33376 19712
rect 34060 19728 34112 19780
rect 34152 19728 34204 19780
rect 38844 19728 38896 19780
rect 39488 19728 39540 19780
rect 37924 19660 37976 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 1676 19456 1728 19508
rect 2596 19499 2648 19508
rect 2596 19465 2605 19499
rect 2605 19465 2639 19499
rect 2639 19465 2648 19499
rect 2596 19456 2648 19465
rect 2780 19320 2832 19372
rect 3424 19456 3476 19508
rect 4620 19456 4672 19508
rect 5080 19456 5132 19508
rect 5540 19499 5592 19508
rect 5540 19465 5549 19499
rect 5549 19465 5583 19499
rect 5583 19465 5592 19499
rect 5540 19456 5592 19465
rect 7012 19456 7064 19508
rect 8576 19456 8628 19508
rect 8760 19456 8812 19508
rect 9404 19456 9456 19508
rect 3608 19388 3660 19440
rect 4436 19320 4488 19372
rect 4712 19320 4764 19372
rect 8300 19388 8352 19440
rect 4068 19252 4120 19304
rect 5172 19363 5224 19372
rect 5172 19329 5181 19363
rect 5181 19329 5215 19363
rect 5215 19329 5224 19363
rect 5172 19320 5224 19329
rect 2872 19116 2924 19168
rect 3884 19116 3936 19168
rect 5632 19320 5684 19372
rect 5724 19320 5776 19372
rect 7564 19320 7616 19372
rect 5632 19184 5684 19236
rect 5816 19184 5868 19236
rect 6828 19184 6880 19236
rect 6920 19159 6972 19168
rect 6920 19125 6929 19159
rect 6929 19125 6963 19159
rect 6963 19125 6972 19159
rect 6920 19116 6972 19125
rect 8024 19184 8076 19236
rect 9496 19320 9548 19372
rect 9956 19456 10008 19508
rect 12716 19456 12768 19508
rect 13728 19456 13780 19508
rect 10140 19388 10192 19440
rect 11060 19388 11112 19440
rect 12348 19388 12400 19440
rect 14556 19388 14608 19440
rect 8944 19252 8996 19304
rect 9864 19252 9916 19304
rect 9956 19252 10008 19304
rect 10784 19295 10836 19304
rect 10784 19261 10793 19295
rect 10793 19261 10827 19295
rect 10827 19261 10836 19295
rect 10784 19252 10836 19261
rect 12532 19363 12584 19372
rect 12532 19329 12541 19363
rect 12541 19329 12575 19363
rect 12575 19329 12584 19363
rect 12532 19320 12584 19329
rect 13360 19320 13412 19372
rect 12716 19252 12768 19304
rect 14740 19320 14792 19372
rect 16856 19456 16908 19508
rect 17408 19456 17460 19508
rect 17868 19456 17920 19508
rect 24584 19456 24636 19508
rect 25136 19456 25188 19508
rect 25596 19456 25648 19508
rect 16028 19388 16080 19440
rect 16396 19388 16448 19440
rect 14464 19252 14516 19304
rect 15752 19363 15804 19372
rect 15752 19329 15761 19363
rect 15761 19329 15795 19363
rect 15795 19329 15804 19363
rect 15752 19320 15804 19329
rect 17316 19363 17368 19372
rect 17316 19329 17325 19363
rect 17325 19329 17359 19363
rect 17359 19329 17368 19363
rect 17316 19320 17368 19329
rect 17592 19388 17644 19440
rect 18144 19388 18196 19440
rect 18236 19431 18288 19440
rect 18236 19397 18245 19431
rect 18245 19397 18279 19431
rect 18279 19397 18288 19431
rect 18236 19388 18288 19397
rect 20168 19388 20220 19440
rect 20536 19388 20588 19440
rect 21732 19388 21784 19440
rect 20720 19320 20772 19372
rect 22192 19320 22244 19372
rect 22376 19388 22428 19440
rect 12900 19184 12952 19236
rect 13728 19184 13780 19236
rect 14648 19184 14700 19236
rect 15108 19184 15160 19236
rect 19064 19252 19116 19304
rect 19156 19295 19208 19304
rect 19156 19261 19165 19295
rect 19165 19261 19199 19295
rect 19199 19261 19208 19295
rect 19156 19252 19208 19261
rect 19432 19252 19484 19304
rect 21548 19252 21600 19304
rect 22376 19295 22428 19304
rect 22376 19261 22385 19295
rect 22385 19261 22419 19295
rect 22419 19261 22428 19295
rect 22376 19252 22428 19261
rect 23204 19320 23256 19372
rect 24032 19388 24084 19440
rect 24308 19388 24360 19440
rect 24676 19431 24728 19440
rect 24676 19397 24685 19431
rect 24685 19397 24719 19431
rect 24719 19397 24728 19431
rect 24676 19388 24728 19397
rect 25228 19431 25280 19440
rect 25228 19397 25237 19431
rect 25237 19397 25271 19431
rect 25271 19397 25280 19431
rect 25228 19388 25280 19397
rect 25688 19388 25740 19440
rect 25964 19388 26016 19440
rect 27712 19456 27764 19508
rect 27896 19456 27948 19508
rect 29552 19456 29604 19508
rect 23572 19320 23624 19372
rect 23664 19363 23716 19372
rect 23664 19329 23673 19363
rect 23673 19329 23707 19363
rect 23707 19329 23716 19363
rect 23664 19320 23716 19329
rect 23848 19320 23900 19372
rect 24400 19363 24452 19372
rect 24400 19329 24409 19363
rect 24409 19329 24443 19363
rect 24443 19329 24452 19363
rect 24400 19320 24452 19329
rect 20628 19184 20680 19236
rect 9404 19116 9456 19168
rect 12072 19116 12124 19168
rect 15568 19116 15620 19168
rect 16580 19116 16632 19168
rect 17224 19116 17276 19168
rect 18144 19116 18196 19168
rect 19064 19159 19116 19168
rect 19064 19125 19073 19159
rect 19073 19125 19107 19159
rect 19107 19125 19116 19159
rect 19064 19116 19116 19125
rect 21180 19116 21232 19168
rect 22560 19116 22612 19168
rect 23204 19159 23256 19168
rect 23204 19125 23213 19159
rect 23213 19125 23247 19159
rect 23247 19125 23256 19159
rect 23204 19116 23256 19125
rect 24584 19184 24636 19236
rect 24860 19295 24912 19304
rect 24860 19261 24869 19295
rect 24869 19261 24903 19295
rect 24903 19261 24912 19295
rect 24860 19252 24912 19261
rect 25136 19320 25188 19372
rect 25596 19363 25648 19372
rect 25596 19329 25605 19363
rect 25605 19329 25639 19363
rect 25639 19329 25648 19363
rect 25596 19320 25648 19329
rect 25412 19252 25464 19304
rect 26056 19320 26108 19372
rect 26148 19252 26200 19304
rect 26516 19363 26568 19372
rect 26516 19329 26525 19363
rect 26525 19329 26559 19363
rect 26559 19329 26568 19363
rect 26516 19320 26568 19329
rect 26608 19320 26660 19372
rect 24952 19116 25004 19168
rect 25136 19116 25188 19168
rect 25780 19116 25832 19168
rect 26884 19252 26936 19304
rect 28172 19431 28224 19440
rect 28172 19397 28181 19431
rect 28181 19397 28215 19431
rect 28215 19397 28224 19431
rect 28172 19388 28224 19397
rect 29920 19456 29972 19508
rect 30380 19456 30432 19508
rect 27712 19320 27764 19372
rect 27896 19320 27948 19372
rect 27344 19252 27396 19304
rect 28080 19252 28132 19304
rect 29092 19320 29144 19372
rect 30472 19388 30524 19440
rect 33140 19456 33192 19508
rect 39672 19456 39724 19508
rect 40132 19456 40184 19508
rect 30932 19320 30984 19372
rect 33600 19388 33652 19440
rect 33416 19320 33468 19372
rect 34152 19388 34204 19440
rect 34612 19388 34664 19440
rect 35624 19388 35676 19440
rect 39120 19388 39172 19440
rect 33784 19320 33836 19372
rect 35716 19320 35768 19372
rect 39580 19363 39632 19372
rect 39580 19329 39589 19363
rect 39589 19329 39623 19363
rect 39623 19329 39632 19363
rect 39580 19320 39632 19329
rect 39672 19363 39724 19372
rect 39672 19329 39681 19363
rect 39681 19329 39715 19363
rect 39715 19329 39724 19363
rect 39672 19320 39724 19329
rect 26608 19184 26660 19236
rect 31116 19295 31168 19304
rect 31116 19261 31125 19295
rect 31125 19261 31159 19295
rect 31159 19261 31168 19295
rect 31116 19252 31168 19261
rect 32956 19252 33008 19304
rect 33508 19252 33560 19304
rect 38752 19252 38804 19304
rect 39120 19252 39172 19304
rect 30748 19184 30800 19236
rect 27712 19159 27764 19168
rect 27712 19125 27721 19159
rect 27721 19125 27755 19159
rect 27755 19125 27764 19159
rect 27712 19116 27764 19125
rect 30932 19159 30984 19168
rect 30932 19125 30941 19159
rect 30941 19125 30975 19159
rect 30975 19125 30984 19159
rect 30932 19116 30984 19125
rect 31576 19184 31628 19236
rect 37372 19184 37424 19236
rect 32956 19116 33008 19168
rect 33140 19116 33192 19168
rect 37740 19116 37792 19168
rect 39304 19116 39356 19168
rect 39856 19159 39908 19168
rect 39856 19125 39865 19159
rect 39865 19125 39899 19159
rect 39899 19125 39908 19159
rect 39856 19116 39908 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 3976 18912 4028 18964
rect 5724 18912 5776 18964
rect 7380 18912 7432 18964
rect 7840 18955 7892 18964
rect 7840 18921 7849 18955
rect 7849 18921 7883 18955
rect 7883 18921 7892 18955
rect 7840 18912 7892 18921
rect 8300 18912 8352 18964
rect 8760 18912 8812 18964
rect 2872 18776 2924 18828
rect 5080 18776 5132 18828
rect 4436 18708 4488 18760
rect 5540 18708 5592 18760
rect 5632 18751 5684 18760
rect 5632 18717 5641 18751
rect 5641 18717 5675 18751
rect 5675 18717 5684 18751
rect 5632 18708 5684 18717
rect 12164 18912 12216 18964
rect 12808 18912 12860 18964
rect 15936 18912 15988 18964
rect 17960 18912 18012 18964
rect 18788 18912 18840 18964
rect 14832 18844 14884 18896
rect 10600 18776 10652 18828
rect 6000 18708 6052 18760
rect 9956 18708 10008 18760
rect 11612 18708 11664 18760
rect 12716 18776 12768 18828
rect 16856 18776 16908 18828
rect 19156 18844 19208 18896
rect 12164 18751 12216 18760
rect 12164 18717 12174 18751
rect 12174 18717 12208 18751
rect 12208 18717 12216 18751
rect 12164 18708 12216 18717
rect 12348 18751 12400 18760
rect 12348 18717 12357 18751
rect 12357 18717 12391 18751
rect 12391 18717 12400 18751
rect 12348 18708 12400 18717
rect 12900 18708 12952 18760
rect 20628 18776 20680 18828
rect 20904 18776 20956 18828
rect 20996 18776 21048 18828
rect 21180 18819 21232 18828
rect 21180 18785 21189 18819
rect 21189 18785 21223 18819
rect 21223 18785 21232 18819
rect 21180 18776 21232 18785
rect 17960 18708 18012 18760
rect 18328 18708 18380 18760
rect 21088 18708 21140 18760
rect 21456 18955 21508 18964
rect 21456 18921 21465 18955
rect 21465 18921 21499 18955
rect 21499 18921 21508 18955
rect 21456 18912 21508 18921
rect 23204 18912 23256 18964
rect 23756 18912 23808 18964
rect 24584 18912 24636 18964
rect 25596 18912 25648 18964
rect 25688 18912 25740 18964
rect 26608 18912 26660 18964
rect 30932 18912 30984 18964
rect 31576 18912 31628 18964
rect 31668 18912 31720 18964
rect 32496 18912 32548 18964
rect 22008 18819 22060 18828
rect 22008 18785 22017 18819
rect 22017 18785 22051 18819
rect 22051 18785 22060 18819
rect 22008 18776 22060 18785
rect 22836 18819 22888 18828
rect 22836 18785 22845 18819
rect 22845 18785 22879 18819
rect 22879 18785 22888 18819
rect 22836 18776 22888 18785
rect 4804 18572 4856 18624
rect 6184 18572 6236 18624
rect 7104 18572 7156 18624
rect 7288 18572 7340 18624
rect 9312 18572 9364 18624
rect 12256 18572 12308 18624
rect 18604 18683 18656 18692
rect 18604 18649 18613 18683
rect 18613 18649 18647 18683
rect 18647 18649 18656 18683
rect 18604 18640 18656 18649
rect 14740 18572 14792 18624
rect 18696 18615 18748 18624
rect 18696 18581 18705 18615
rect 18705 18581 18739 18615
rect 18739 18581 18748 18615
rect 18696 18572 18748 18581
rect 20536 18615 20588 18624
rect 20536 18581 20551 18615
rect 20551 18581 20585 18615
rect 20585 18581 20588 18615
rect 20536 18572 20588 18581
rect 21548 18615 21600 18624
rect 21548 18581 21557 18615
rect 21557 18581 21591 18615
rect 21591 18581 21600 18615
rect 21548 18572 21600 18581
rect 21732 18572 21784 18624
rect 23388 18708 23440 18760
rect 23480 18708 23532 18760
rect 22192 18640 22244 18692
rect 23756 18640 23808 18692
rect 23296 18572 23348 18624
rect 23388 18615 23440 18624
rect 23388 18581 23397 18615
rect 23397 18581 23431 18615
rect 23431 18581 23440 18615
rect 23388 18572 23440 18581
rect 24768 18708 24820 18760
rect 25136 18751 25188 18760
rect 25136 18717 25145 18751
rect 25145 18717 25179 18751
rect 25179 18717 25188 18751
rect 25136 18708 25188 18717
rect 25320 18683 25372 18692
rect 25320 18649 25329 18683
rect 25329 18649 25363 18683
rect 25363 18649 25372 18683
rect 25320 18640 25372 18649
rect 25504 18640 25556 18692
rect 26056 18751 26108 18760
rect 32680 18844 32732 18896
rect 34060 18912 34112 18964
rect 35440 18912 35492 18964
rect 32588 18776 32640 18828
rect 26056 18717 26070 18751
rect 26070 18717 26104 18751
rect 26104 18717 26108 18751
rect 26056 18708 26108 18717
rect 25872 18683 25924 18692
rect 25872 18649 25881 18683
rect 25881 18649 25915 18683
rect 25915 18649 25924 18683
rect 25872 18640 25924 18649
rect 26148 18640 26200 18692
rect 26332 18683 26384 18692
rect 26332 18649 26341 18683
rect 26341 18649 26375 18683
rect 26375 18649 26384 18683
rect 26332 18640 26384 18649
rect 26516 18615 26568 18624
rect 26516 18581 26541 18615
rect 26541 18581 26568 18615
rect 26516 18572 26568 18581
rect 27344 18572 27396 18624
rect 31392 18572 31444 18624
rect 31760 18751 31812 18760
rect 31760 18717 31795 18751
rect 31795 18717 31812 18751
rect 31760 18708 31812 18717
rect 32772 18708 32824 18760
rect 33140 18751 33192 18760
rect 33140 18717 33149 18751
rect 33149 18717 33183 18751
rect 33183 18717 33192 18751
rect 33140 18708 33192 18717
rect 34428 18776 34480 18828
rect 34888 18776 34940 18828
rect 31668 18572 31720 18624
rect 33416 18640 33468 18692
rect 34060 18708 34112 18760
rect 34704 18708 34756 18760
rect 35716 18751 35768 18760
rect 35716 18717 35725 18751
rect 35725 18717 35759 18751
rect 35759 18717 35768 18751
rect 35716 18708 35768 18717
rect 35808 18751 35860 18760
rect 35808 18717 35817 18751
rect 35817 18717 35851 18751
rect 35851 18717 35860 18751
rect 35808 18708 35860 18717
rect 36636 18887 36688 18896
rect 36636 18853 36645 18887
rect 36645 18853 36679 18887
rect 36679 18853 36688 18887
rect 36636 18844 36688 18853
rect 37280 18912 37332 18964
rect 37832 18955 37884 18964
rect 37832 18921 37841 18955
rect 37841 18921 37875 18955
rect 37875 18921 37884 18955
rect 37832 18912 37884 18921
rect 38016 18912 38068 18964
rect 39856 18912 39908 18964
rect 38292 18844 38344 18896
rect 37556 18776 37608 18828
rect 33692 18683 33744 18692
rect 33692 18649 33701 18683
rect 33701 18649 33735 18683
rect 33735 18649 33744 18683
rect 33692 18640 33744 18649
rect 32496 18572 32548 18624
rect 33140 18572 33192 18624
rect 33508 18572 33560 18624
rect 35164 18640 35216 18692
rect 36360 18640 36412 18692
rect 37372 18708 37424 18760
rect 37924 18708 37976 18760
rect 37280 18640 37332 18692
rect 38108 18640 38160 18692
rect 38752 18751 38804 18760
rect 38752 18717 38761 18751
rect 38761 18717 38795 18751
rect 38795 18717 38804 18751
rect 38752 18708 38804 18717
rect 39028 18640 39080 18692
rect 40224 18955 40276 18964
rect 40224 18921 40233 18955
rect 40233 18921 40267 18955
rect 40267 18921 40276 18955
rect 40224 18912 40276 18921
rect 36452 18572 36504 18624
rect 38200 18615 38252 18624
rect 38200 18581 38209 18615
rect 38209 18581 38243 18615
rect 38243 18581 38252 18615
rect 38200 18572 38252 18581
rect 40040 18572 40092 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 4068 18232 4120 18284
rect 6920 18368 6972 18420
rect 7104 18411 7156 18420
rect 7104 18377 7113 18411
rect 7113 18377 7147 18411
rect 7147 18377 7156 18411
rect 7104 18368 7156 18377
rect 9772 18368 9824 18420
rect 10416 18368 10468 18420
rect 14464 18411 14516 18420
rect 14464 18377 14473 18411
rect 14473 18377 14507 18411
rect 14507 18377 14516 18411
rect 14464 18368 14516 18377
rect 2964 18207 3016 18216
rect 2964 18173 2973 18207
rect 2973 18173 3007 18207
rect 3007 18173 3016 18207
rect 2964 18164 3016 18173
rect 3424 18207 3476 18216
rect 3424 18173 3433 18207
rect 3433 18173 3467 18207
rect 3467 18173 3476 18207
rect 3424 18164 3476 18173
rect 5264 18164 5316 18216
rect 4436 18096 4488 18148
rect 5632 18164 5684 18216
rect 8392 18232 8444 18284
rect 9220 18207 9272 18216
rect 9220 18173 9229 18207
rect 9229 18173 9263 18207
rect 9263 18173 9272 18207
rect 9220 18164 9272 18173
rect 9404 18207 9456 18216
rect 9404 18173 9413 18207
rect 9413 18173 9447 18207
rect 9447 18173 9456 18207
rect 14372 18232 14424 18284
rect 16028 18368 16080 18420
rect 16948 18368 17000 18420
rect 18512 18368 18564 18420
rect 18604 18368 18656 18420
rect 20628 18368 20680 18420
rect 21548 18368 21600 18420
rect 24124 18368 24176 18420
rect 26516 18368 26568 18420
rect 27344 18368 27396 18420
rect 15476 18232 15528 18284
rect 15936 18232 15988 18284
rect 16028 18275 16080 18284
rect 16028 18241 16037 18275
rect 16037 18241 16071 18275
rect 16071 18241 16080 18275
rect 16028 18232 16080 18241
rect 16304 18275 16356 18284
rect 16304 18241 16313 18275
rect 16313 18241 16347 18275
rect 16347 18241 16356 18275
rect 16304 18232 16356 18241
rect 9404 18164 9456 18173
rect 14740 18207 14792 18216
rect 14740 18173 14749 18207
rect 14749 18173 14783 18207
rect 14783 18173 14792 18207
rect 14740 18164 14792 18173
rect 15568 18164 15620 18216
rect 17224 18232 17276 18284
rect 17776 18232 17828 18284
rect 18236 18275 18288 18284
rect 18236 18241 18245 18275
rect 18245 18241 18279 18275
rect 18279 18241 18288 18275
rect 18236 18232 18288 18241
rect 19064 18232 19116 18284
rect 19340 18275 19392 18284
rect 19340 18241 19349 18275
rect 19349 18241 19383 18275
rect 19383 18241 19392 18275
rect 19340 18232 19392 18241
rect 12440 18096 12492 18148
rect 16488 18096 16540 18148
rect 17132 18207 17184 18216
rect 17132 18173 17141 18207
rect 17141 18173 17175 18207
rect 17175 18173 17184 18207
rect 17132 18164 17184 18173
rect 18972 18164 19024 18216
rect 19432 18207 19484 18216
rect 19432 18173 19441 18207
rect 19441 18173 19475 18207
rect 19475 18173 19484 18207
rect 19432 18164 19484 18173
rect 23296 18300 23348 18352
rect 23756 18232 23808 18284
rect 24400 18232 24452 18284
rect 27896 18232 27948 18284
rect 30472 18368 30524 18420
rect 20904 18096 20956 18148
rect 21548 18096 21600 18148
rect 2504 18071 2556 18080
rect 2504 18037 2513 18071
rect 2513 18037 2547 18071
rect 2547 18037 2556 18071
rect 2504 18028 2556 18037
rect 4712 18071 4764 18080
rect 4712 18037 4721 18071
rect 4721 18037 4755 18071
rect 4755 18037 4764 18071
rect 4712 18028 4764 18037
rect 8760 18071 8812 18080
rect 8760 18037 8769 18071
rect 8769 18037 8803 18071
rect 8803 18037 8812 18071
rect 8760 18028 8812 18037
rect 14096 18071 14148 18080
rect 14096 18037 14105 18071
rect 14105 18037 14139 18071
rect 14139 18037 14148 18071
rect 14096 18028 14148 18037
rect 15752 18071 15804 18080
rect 15752 18037 15761 18071
rect 15761 18037 15795 18071
rect 15795 18037 15804 18071
rect 15752 18028 15804 18037
rect 16580 18028 16632 18080
rect 16672 18071 16724 18080
rect 16672 18037 16681 18071
rect 16681 18037 16715 18071
rect 16715 18037 16724 18071
rect 16672 18028 16724 18037
rect 17776 18028 17828 18080
rect 18604 18028 18656 18080
rect 18972 18071 19024 18080
rect 18972 18037 18981 18071
rect 18981 18037 19015 18071
rect 19015 18037 19024 18071
rect 18972 18028 19024 18037
rect 19616 18028 19668 18080
rect 30012 18207 30064 18216
rect 30012 18173 30021 18207
rect 30021 18173 30055 18207
rect 30055 18173 30064 18207
rect 30012 18164 30064 18173
rect 30104 18207 30156 18216
rect 30104 18173 30113 18207
rect 30113 18173 30147 18207
rect 30147 18173 30156 18207
rect 30104 18164 30156 18173
rect 30656 18275 30708 18284
rect 30656 18241 30665 18275
rect 30665 18241 30699 18275
rect 30699 18241 30708 18275
rect 30656 18232 30708 18241
rect 30748 18232 30800 18284
rect 31852 18368 31904 18420
rect 32680 18368 32732 18420
rect 35164 18368 35216 18420
rect 33048 18300 33100 18352
rect 31392 18275 31444 18284
rect 31392 18241 31401 18275
rect 31401 18241 31435 18275
rect 31435 18241 31444 18275
rect 31392 18232 31444 18241
rect 32772 18232 32824 18284
rect 33508 18300 33560 18352
rect 33968 18300 34020 18352
rect 33416 18232 33468 18284
rect 34520 18232 34572 18284
rect 34888 18275 34940 18284
rect 34888 18241 34897 18275
rect 34897 18241 34931 18275
rect 34931 18241 34940 18275
rect 34888 18232 34940 18241
rect 36176 18300 36228 18352
rect 34060 18164 34112 18216
rect 35256 18275 35308 18284
rect 35256 18241 35265 18275
rect 35265 18241 35299 18275
rect 35299 18241 35308 18275
rect 35256 18232 35308 18241
rect 23940 18096 23992 18148
rect 24860 18096 24912 18148
rect 26148 18096 26200 18148
rect 30380 18096 30432 18148
rect 30564 18139 30616 18148
rect 30564 18105 30573 18139
rect 30573 18105 30607 18139
rect 30607 18105 30616 18139
rect 35900 18232 35952 18284
rect 36544 18232 36596 18284
rect 37648 18343 37700 18352
rect 37648 18309 37657 18343
rect 37657 18309 37691 18343
rect 37691 18309 37700 18343
rect 37648 18300 37700 18309
rect 30564 18096 30616 18105
rect 29736 18028 29788 18080
rect 30012 18028 30064 18080
rect 30472 18028 30524 18080
rect 30656 18028 30708 18080
rect 31116 18028 31168 18080
rect 33048 18028 33100 18080
rect 33876 18028 33928 18080
rect 36452 18096 36504 18148
rect 37648 18164 37700 18216
rect 38200 18368 38252 18420
rect 41328 18368 41380 18420
rect 41512 18368 41564 18420
rect 37924 18275 37976 18284
rect 37924 18241 37933 18275
rect 37933 18241 37967 18275
rect 37967 18241 37976 18275
rect 37924 18232 37976 18241
rect 38108 18232 38160 18284
rect 39580 18232 39632 18284
rect 40316 18232 40368 18284
rect 40500 18275 40552 18284
rect 40500 18241 40509 18275
rect 40509 18241 40543 18275
rect 40543 18241 40552 18275
rect 40500 18232 40552 18241
rect 40132 18207 40184 18216
rect 40132 18173 40141 18207
rect 40141 18173 40175 18207
rect 40175 18173 40184 18207
rect 40132 18164 40184 18173
rect 41696 18164 41748 18216
rect 39028 18096 39080 18148
rect 39580 18096 39632 18148
rect 36636 18028 36688 18080
rect 37096 18028 37148 18080
rect 38108 18071 38160 18080
rect 38108 18037 38117 18071
rect 38117 18037 38151 18071
rect 38151 18037 38160 18071
rect 38108 18028 38160 18037
rect 39764 18071 39816 18080
rect 39764 18037 39773 18071
rect 39773 18037 39807 18071
rect 39807 18037 39816 18071
rect 39764 18028 39816 18037
rect 40040 18071 40092 18080
rect 40040 18037 40049 18071
rect 40049 18037 40083 18071
rect 40083 18037 40092 18071
rect 40040 18028 40092 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 6000 17824 6052 17876
rect 6368 17824 6420 17876
rect 3424 17756 3476 17808
rect 5632 17756 5684 17808
rect 4620 17688 4672 17740
rect 6552 17756 6604 17808
rect 9680 17756 9732 17808
rect 8024 17688 8076 17740
rect 9956 17731 10008 17740
rect 9956 17697 9965 17731
rect 9965 17697 9999 17731
rect 9999 17697 10008 17731
rect 9956 17688 10008 17697
rect 5632 17620 5684 17672
rect 6092 17620 6144 17672
rect 8116 17620 8168 17672
rect 8760 17663 8812 17672
rect 8760 17629 8769 17663
rect 8769 17629 8803 17663
rect 8803 17629 8812 17663
rect 8760 17620 8812 17629
rect 9128 17620 9180 17672
rect 9588 17620 9640 17672
rect 13176 17824 13228 17876
rect 13912 17824 13964 17876
rect 15292 17824 15344 17876
rect 15476 17824 15528 17876
rect 16672 17824 16724 17876
rect 18328 17824 18380 17876
rect 18880 17824 18932 17876
rect 19340 17824 19392 17876
rect 21456 17824 21508 17876
rect 24492 17824 24544 17876
rect 24584 17824 24636 17876
rect 24768 17824 24820 17876
rect 29644 17824 29696 17876
rect 36636 17824 36688 17876
rect 37924 17867 37976 17876
rect 37924 17833 37933 17867
rect 37933 17833 37967 17867
rect 37967 17833 37976 17867
rect 37924 17824 37976 17833
rect 38844 17867 38896 17876
rect 38844 17833 38853 17867
rect 38853 17833 38887 17867
rect 38887 17833 38896 17867
rect 38844 17824 38896 17833
rect 12164 17756 12216 17808
rect 12440 17731 12492 17740
rect 12440 17697 12449 17731
rect 12449 17697 12483 17731
rect 12483 17697 12492 17731
rect 12440 17688 12492 17697
rect 18052 17756 18104 17808
rect 18696 17756 18748 17808
rect 20628 17756 20680 17808
rect 12532 17620 12584 17672
rect 14188 17688 14240 17740
rect 17868 17688 17920 17740
rect 18328 17731 18380 17740
rect 18328 17697 18337 17731
rect 18337 17697 18371 17731
rect 18371 17697 18380 17731
rect 18328 17688 18380 17697
rect 19248 17688 19300 17740
rect 1676 17595 1728 17604
rect 1676 17561 1685 17595
rect 1685 17561 1719 17595
rect 1719 17561 1728 17595
rect 1676 17552 1728 17561
rect 3424 17552 3476 17604
rect 10232 17595 10284 17604
rect 10232 17561 10241 17595
rect 10241 17561 10275 17595
rect 10275 17561 10284 17595
rect 10232 17552 10284 17561
rect 11244 17552 11296 17604
rect 11612 17552 11664 17604
rect 4712 17484 4764 17536
rect 8484 17527 8536 17536
rect 8484 17493 8493 17527
rect 8493 17493 8527 17527
rect 8527 17493 8536 17527
rect 8484 17484 8536 17493
rect 8576 17527 8628 17536
rect 8576 17493 8585 17527
rect 8585 17493 8619 17527
rect 8619 17493 8628 17527
rect 8576 17484 8628 17493
rect 11796 17527 11848 17536
rect 11796 17493 11805 17527
rect 11805 17493 11839 17527
rect 11839 17493 11848 17527
rect 11796 17484 11848 17493
rect 13544 17663 13596 17672
rect 13544 17629 13553 17663
rect 13553 17629 13587 17663
rect 13587 17629 13596 17663
rect 13544 17620 13596 17629
rect 14096 17620 14148 17672
rect 15292 17620 15344 17672
rect 17224 17620 17276 17672
rect 17776 17663 17828 17672
rect 17776 17629 17785 17663
rect 17785 17629 17819 17663
rect 17819 17629 17828 17663
rect 17776 17620 17828 17629
rect 18052 17663 18104 17672
rect 18052 17629 18061 17663
rect 18061 17629 18095 17663
rect 18095 17629 18104 17663
rect 18052 17620 18104 17629
rect 14096 17527 14148 17536
rect 14096 17493 14105 17527
rect 14105 17493 14139 17527
rect 14139 17493 14148 17527
rect 14096 17484 14148 17493
rect 15292 17484 15344 17536
rect 17592 17595 17644 17604
rect 17592 17561 17601 17595
rect 17601 17561 17635 17595
rect 17635 17561 17644 17595
rect 17592 17552 17644 17561
rect 16672 17484 16724 17536
rect 17960 17527 18012 17536
rect 17960 17493 17969 17527
rect 17969 17493 18003 17527
rect 18003 17493 18012 17527
rect 17960 17484 18012 17493
rect 18236 17484 18288 17536
rect 18512 17663 18564 17672
rect 18512 17629 18521 17663
rect 18521 17629 18555 17663
rect 18555 17629 18564 17663
rect 18512 17620 18564 17629
rect 18880 17620 18932 17672
rect 19156 17620 19208 17672
rect 19616 17731 19668 17740
rect 19616 17697 19625 17731
rect 19625 17697 19659 17731
rect 19659 17697 19668 17731
rect 19616 17688 19668 17697
rect 23572 17688 23624 17740
rect 24124 17688 24176 17740
rect 18696 17484 18748 17536
rect 21456 17620 21508 17672
rect 22008 17620 22060 17672
rect 23756 17620 23808 17672
rect 25228 17688 25280 17740
rect 26056 17756 26108 17808
rect 24952 17620 25004 17672
rect 25504 17620 25556 17672
rect 21180 17552 21232 17604
rect 22836 17552 22888 17604
rect 26332 17688 26384 17740
rect 27712 17731 27764 17740
rect 27712 17697 27721 17731
rect 27721 17697 27755 17731
rect 27755 17697 27764 17731
rect 27712 17688 27764 17697
rect 29000 17688 29052 17740
rect 29276 17688 29328 17740
rect 31576 17799 31628 17808
rect 31576 17765 31585 17799
rect 31585 17765 31619 17799
rect 31619 17765 31628 17799
rect 31576 17756 31628 17765
rect 32588 17756 32640 17808
rect 33784 17756 33836 17808
rect 27804 17663 27856 17672
rect 27804 17629 27813 17663
rect 27813 17629 27847 17663
rect 27847 17629 27856 17663
rect 27804 17620 27856 17629
rect 28264 17663 28316 17672
rect 28264 17629 28273 17663
rect 28273 17629 28307 17663
rect 28307 17629 28316 17663
rect 28264 17620 28316 17629
rect 28540 17663 28592 17672
rect 28540 17629 28549 17663
rect 28549 17629 28583 17663
rect 28583 17629 28592 17663
rect 28540 17620 28592 17629
rect 27528 17595 27580 17604
rect 27528 17561 27537 17595
rect 27537 17561 27571 17595
rect 27571 17561 27580 17595
rect 27528 17552 27580 17561
rect 21272 17484 21324 17536
rect 23480 17484 23532 17536
rect 24124 17484 24176 17536
rect 26148 17484 26200 17536
rect 29552 17552 29604 17604
rect 29644 17552 29696 17604
rect 30380 17663 30432 17672
rect 30380 17629 30389 17663
rect 30389 17629 30423 17663
rect 30423 17629 30432 17663
rect 30380 17620 30432 17629
rect 30472 17620 30524 17672
rect 31024 17620 31076 17672
rect 31760 17620 31812 17672
rect 33692 17663 33744 17672
rect 33692 17629 33701 17663
rect 33701 17629 33735 17663
rect 33735 17629 33744 17663
rect 33692 17620 33744 17629
rect 33784 17663 33836 17672
rect 33784 17629 33794 17663
rect 33794 17629 33828 17663
rect 33828 17629 33836 17663
rect 34244 17756 34296 17808
rect 36360 17756 36412 17808
rect 39672 17867 39724 17876
rect 39672 17833 39681 17867
rect 39681 17833 39715 17867
rect 39715 17833 39724 17867
rect 39672 17824 39724 17833
rect 40132 17756 40184 17808
rect 33784 17620 33836 17629
rect 33600 17552 33652 17604
rect 33508 17484 33560 17536
rect 33876 17484 33928 17536
rect 34336 17620 34388 17672
rect 35440 17663 35492 17672
rect 35440 17629 35449 17663
rect 35449 17629 35483 17663
rect 35483 17629 35492 17663
rect 35440 17620 35492 17629
rect 37556 17731 37608 17740
rect 37556 17697 37565 17731
rect 37565 17697 37599 17731
rect 37599 17697 37608 17731
rect 37556 17688 37608 17697
rect 38016 17688 38068 17740
rect 35348 17552 35400 17604
rect 35716 17484 35768 17536
rect 35808 17484 35860 17536
rect 36912 17620 36964 17672
rect 37740 17663 37792 17672
rect 37740 17629 37749 17663
rect 37749 17629 37783 17663
rect 37783 17629 37792 17663
rect 37740 17620 37792 17629
rect 39028 17620 39080 17672
rect 38200 17552 38252 17604
rect 36544 17484 36596 17536
rect 40408 17688 40460 17740
rect 39580 17620 39632 17672
rect 39396 17484 39448 17536
rect 40040 17484 40092 17536
rect 41604 17484 41656 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 1676 17280 1728 17332
rect 2504 17280 2556 17332
rect 8484 17280 8536 17332
rect 8576 17280 8628 17332
rect 9772 17323 9824 17332
rect 9772 17289 9781 17323
rect 9781 17289 9815 17323
rect 9815 17289 9824 17323
rect 9772 17280 9824 17289
rect 10232 17280 10284 17332
rect 2964 17212 3016 17264
rect 3976 17212 4028 17264
rect 6000 17144 6052 17196
rect 9312 17212 9364 17264
rect 8024 17187 8076 17196
rect 3884 17076 3936 17128
rect 8024 17153 8033 17187
rect 8033 17153 8067 17187
rect 8067 17153 8076 17187
rect 8024 17144 8076 17153
rect 9680 17144 9732 17196
rect 7564 17119 7616 17128
rect 7564 17085 7573 17119
rect 7573 17085 7607 17119
rect 7607 17085 7616 17119
rect 7564 17076 7616 17085
rect 2136 16940 2188 16992
rect 3332 16940 3384 16992
rect 4068 16940 4120 16992
rect 6644 16940 6696 16992
rect 6828 16940 6880 16992
rect 11796 17280 11848 17332
rect 12532 17280 12584 17332
rect 14096 17280 14148 17332
rect 14464 17280 14516 17332
rect 16304 17323 16356 17332
rect 16304 17289 16313 17323
rect 16313 17289 16347 17323
rect 16347 17289 16356 17323
rect 16304 17280 16356 17289
rect 16580 17280 16632 17332
rect 13728 17212 13780 17264
rect 13912 17212 13964 17264
rect 16488 17212 16540 17264
rect 16672 17212 16724 17264
rect 15292 17144 15344 17196
rect 16396 17144 16448 17196
rect 17868 17212 17920 17264
rect 18696 17280 18748 17332
rect 19340 17212 19392 17264
rect 12072 17119 12124 17128
rect 12072 17085 12081 17119
rect 12081 17085 12115 17119
rect 12115 17085 12124 17119
rect 12072 17076 12124 17085
rect 12256 17076 12308 17128
rect 13176 17119 13228 17128
rect 13176 17085 13185 17119
rect 13185 17085 13219 17119
rect 13219 17085 13228 17119
rect 13176 17076 13228 17085
rect 10692 17008 10744 17060
rect 17224 17119 17276 17128
rect 17224 17085 17233 17119
rect 17233 17085 17267 17119
rect 17267 17085 17276 17119
rect 17224 17076 17276 17085
rect 18236 17076 18288 17128
rect 18512 17076 18564 17128
rect 20628 17255 20680 17264
rect 20628 17221 20637 17255
rect 20637 17221 20671 17255
rect 20671 17221 20680 17255
rect 20628 17212 20680 17221
rect 23756 17280 23808 17332
rect 24584 17280 24636 17332
rect 26148 17280 26200 17332
rect 26700 17323 26752 17332
rect 26700 17289 26709 17323
rect 26709 17289 26743 17323
rect 26743 17289 26752 17323
rect 26700 17280 26752 17289
rect 23204 17212 23256 17264
rect 23572 17212 23624 17264
rect 20812 17144 20864 17196
rect 21272 17187 21324 17196
rect 21272 17153 21281 17187
rect 21281 17153 21315 17187
rect 21315 17153 21324 17187
rect 21272 17144 21324 17153
rect 21640 17144 21692 17196
rect 21364 17119 21416 17128
rect 21364 17085 21373 17119
rect 21373 17085 21407 17119
rect 21407 17085 21416 17119
rect 21364 17076 21416 17085
rect 21456 17076 21508 17128
rect 22652 17144 22704 17196
rect 22744 17187 22796 17196
rect 22744 17153 22753 17187
rect 22753 17153 22787 17187
rect 22787 17153 22796 17187
rect 22744 17144 22796 17153
rect 23020 17187 23072 17196
rect 23020 17153 23029 17187
rect 23029 17153 23063 17187
rect 23063 17153 23072 17187
rect 23020 17144 23072 17153
rect 23388 17144 23440 17196
rect 9680 16940 9732 16992
rect 10784 16940 10836 16992
rect 11152 16940 11204 16992
rect 15844 16983 15896 16992
rect 15844 16949 15853 16983
rect 15853 16949 15887 16983
rect 15887 16949 15896 16983
rect 15844 16940 15896 16949
rect 17132 16940 17184 16992
rect 17868 16940 17920 16992
rect 19340 16940 19392 16992
rect 20168 16940 20220 16992
rect 20628 16940 20680 16992
rect 22192 16940 22244 16992
rect 22560 16983 22612 16992
rect 22560 16949 22569 16983
rect 22569 16949 22603 16983
rect 22603 16949 22612 16983
rect 22560 16940 22612 16949
rect 24124 17144 24176 17196
rect 24492 17187 24544 17196
rect 24492 17153 24501 17187
rect 24501 17153 24535 17187
rect 24535 17153 24544 17187
rect 24492 17144 24544 17153
rect 24584 17144 24636 17196
rect 25780 17076 25832 17128
rect 26332 17076 26384 17128
rect 26516 17187 26568 17196
rect 26516 17153 26525 17187
rect 26525 17153 26559 17187
rect 26559 17153 26568 17187
rect 26516 17144 26568 17153
rect 27160 17144 27212 17196
rect 27528 17280 27580 17332
rect 27344 17187 27396 17196
rect 27344 17153 27353 17187
rect 27353 17153 27387 17187
rect 27387 17153 27396 17187
rect 27344 17144 27396 17153
rect 27896 17212 27948 17264
rect 28080 17144 28132 17196
rect 28816 17280 28868 17332
rect 29644 17280 29696 17332
rect 30012 17323 30064 17332
rect 30012 17289 30021 17323
rect 30021 17289 30055 17323
rect 30055 17289 30064 17323
rect 30012 17280 30064 17289
rect 32956 17280 33008 17332
rect 36084 17280 36136 17332
rect 39948 17280 40000 17332
rect 40500 17280 40552 17332
rect 29184 17212 29236 17264
rect 35900 17212 35952 17264
rect 39764 17212 39816 17264
rect 28632 17187 28684 17196
rect 28632 17153 28641 17187
rect 28641 17153 28675 17187
rect 28675 17153 28684 17187
rect 28632 17144 28684 17153
rect 27252 17076 27304 17128
rect 28172 17076 28224 17128
rect 23664 17008 23716 17060
rect 23756 17008 23808 17060
rect 23940 16983 23992 16992
rect 23940 16949 23949 16983
rect 23949 16949 23983 16983
rect 23983 16949 23992 16983
rect 23940 16940 23992 16949
rect 26240 16940 26292 16992
rect 26516 16940 26568 16992
rect 27528 16983 27580 16992
rect 27528 16949 27537 16983
rect 27537 16949 27571 16983
rect 27571 16949 27580 16983
rect 27528 16940 27580 16949
rect 27620 16983 27672 16992
rect 27620 16949 27629 16983
rect 27629 16949 27663 16983
rect 27663 16949 27672 16983
rect 27620 16940 27672 16949
rect 29000 17144 29052 17196
rect 29828 17076 29880 17128
rect 28632 16940 28684 16992
rect 28908 17051 28960 17060
rect 28908 17017 28917 17051
rect 28917 17017 28951 17051
rect 28951 17017 28960 17051
rect 28908 17008 28960 17017
rect 29276 17008 29328 17060
rect 29092 16940 29144 16992
rect 29460 16983 29512 16992
rect 29460 16949 29469 16983
rect 29469 16949 29503 16983
rect 29503 16949 29512 16983
rect 30196 17144 30248 17196
rect 33416 17119 33468 17128
rect 33416 17085 33425 17119
rect 33425 17085 33459 17119
rect 33459 17085 33468 17119
rect 33416 17076 33468 17085
rect 32588 17008 32640 17060
rect 34060 17144 34112 17196
rect 35624 17144 35676 17196
rect 33784 17119 33836 17128
rect 33784 17085 33793 17119
rect 33793 17085 33827 17119
rect 33827 17085 33836 17119
rect 33784 17076 33836 17085
rect 40040 17144 40092 17196
rect 39948 17076 40000 17128
rect 35900 17008 35952 17060
rect 40224 17144 40276 17196
rect 29460 16940 29512 16949
rect 31760 16940 31812 16992
rect 32220 16940 32272 16992
rect 33508 16940 33560 16992
rect 33968 16940 34020 16992
rect 37372 16940 37424 16992
rect 39580 16940 39632 16992
rect 39672 16983 39724 16992
rect 39672 16949 39681 16983
rect 39681 16949 39715 16983
rect 39715 16949 39724 16983
rect 39672 16940 39724 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 3516 16736 3568 16788
rect 3884 16736 3936 16788
rect 4068 16736 4120 16788
rect 2136 16600 2188 16652
rect 4804 16643 4856 16652
rect 4804 16609 4813 16643
rect 4813 16609 4847 16643
rect 4847 16609 4856 16643
rect 4804 16600 4856 16609
rect 6736 16736 6788 16788
rect 8116 16736 8168 16788
rect 9680 16736 9732 16788
rect 5356 16600 5408 16652
rect 6276 16643 6328 16652
rect 6276 16609 6285 16643
rect 6285 16609 6319 16643
rect 6319 16609 6328 16643
rect 6276 16600 6328 16609
rect 6644 16600 6696 16652
rect 12256 16736 12308 16788
rect 12072 16668 12124 16720
rect 14740 16736 14792 16788
rect 20720 16736 20772 16788
rect 21824 16736 21876 16788
rect 22652 16736 22704 16788
rect 23664 16779 23716 16788
rect 23664 16745 23673 16779
rect 23673 16745 23707 16779
rect 23707 16745 23716 16779
rect 23664 16736 23716 16745
rect 24492 16736 24544 16788
rect 25780 16736 25832 16788
rect 28724 16779 28776 16788
rect 28724 16745 28733 16779
rect 28733 16745 28767 16779
rect 28767 16745 28776 16779
rect 28724 16736 28776 16745
rect 32220 16736 32272 16788
rect 13176 16668 13228 16720
rect 9956 16600 10008 16652
rect 10784 16600 10836 16652
rect 19892 16668 19944 16720
rect 20812 16668 20864 16720
rect 22284 16668 22336 16720
rect 16580 16600 16632 16652
rect 3424 16464 3476 16516
rect 4068 16396 4120 16448
rect 5080 16396 5132 16448
rect 5448 16396 5500 16448
rect 6092 16575 6144 16584
rect 6092 16541 6101 16575
rect 6101 16541 6135 16575
rect 6135 16541 6144 16575
rect 6092 16532 6144 16541
rect 9036 16532 9088 16584
rect 9496 16532 9548 16584
rect 13912 16575 13964 16584
rect 13912 16541 13921 16575
rect 13921 16541 13955 16575
rect 13955 16541 13964 16575
rect 13912 16532 13964 16541
rect 18144 16532 18196 16584
rect 19248 16532 19300 16584
rect 20076 16600 20128 16652
rect 21640 16643 21692 16652
rect 21640 16609 21649 16643
rect 21649 16609 21683 16643
rect 21683 16609 21692 16643
rect 21640 16600 21692 16609
rect 21916 16643 21968 16652
rect 21916 16609 21925 16643
rect 21925 16609 21959 16643
rect 21959 16609 21968 16643
rect 27620 16668 27672 16720
rect 34336 16779 34388 16788
rect 34336 16745 34345 16779
rect 34345 16745 34379 16779
rect 34379 16745 34388 16779
rect 34336 16736 34388 16745
rect 34520 16779 34572 16788
rect 34520 16745 34529 16779
rect 34529 16745 34563 16779
rect 34563 16745 34572 16779
rect 34520 16736 34572 16745
rect 34796 16736 34848 16788
rect 35440 16736 35492 16788
rect 35624 16736 35676 16788
rect 37372 16736 37424 16788
rect 37740 16736 37792 16788
rect 38660 16736 38712 16788
rect 39948 16736 40000 16788
rect 21916 16600 21968 16609
rect 20628 16532 20680 16584
rect 11244 16464 11296 16516
rect 8116 16396 8168 16448
rect 8944 16439 8996 16448
rect 8944 16405 8953 16439
rect 8953 16405 8987 16439
rect 8987 16405 8996 16439
rect 8944 16396 8996 16405
rect 9220 16396 9272 16448
rect 9312 16439 9364 16448
rect 9312 16405 9321 16439
rect 9321 16405 9355 16439
rect 9355 16405 9364 16439
rect 9312 16396 9364 16405
rect 14648 16464 14700 16516
rect 18420 16464 18472 16516
rect 18972 16464 19024 16516
rect 17684 16396 17736 16448
rect 20720 16396 20772 16448
rect 21548 16575 21600 16584
rect 21548 16541 21557 16575
rect 21557 16541 21591 16575
rect 21591 16541 21600 16575
rect 21548 16532 21600 16541
rect 21456 16464 21508 16516
rect 22928 16532 22980 16584
rect 23480 16575 23532 16584
rect 23480 16541 23489 16575
rect 23489 16541 23523 16575
rect 23523 16541 23532 16575
rect 23480 16532 23532 16541
rect 25044 16575 25096 16584
rect 25044 16541 25053 16575
rect 25053 16541 25087 16575
rect 25087 16541 25096 16575
rect 25044 16532 25096 16541
rect 25228 16575 25280 16584
rect 25228 16541 25235 16575
rect 25235 16541 25280 16575
rect 25228 16532 25280 16541
rect 25504 16575 25556 16584
rect 25504 16541 25518 16575
rect 25518 16541 25552 16575
rect 25552 16541 25556 16575
rect 25504 16532 25556 16541
rect 25688 16532 25740 16584
rect 25872 16575 25924 16584
rect 25872 16541 25882 16575
rect 25882 16541 25916 16575
rect 25916 16541 25924 16575
rect 28632 16600 28684 16652
rect 25872 16532 25924 16541
rect 23572 16464 23624 16516
rect 23756 16464 23808 16516
rect 22008 16396 22060 16448
rect 22100 16396 22152 16448
rect 24860 16396 24912 16448
rect 26056 16507 26108 16516
rect 26056 16473 26065 16507
rect 26065 16473 26099 16507
rect 26099 16473 26108 16507
rect 26056 16464 26108 16473
rect 25780 16396 25832 16448
rect 25872 16396 25924 16448
rect 26332 16464 26384 16516
rect 31576 16575 31628 16584
rect 31576 16541 31611 16575
rect 31611 16541 31628 16575
rect 31576 16532 31628 16541
rect 31852 16532 31904 16584
rect 33048 16600 33100 16652
rect 33416 16643 33468 16652
rect 33416 16609 33425 16643
rect 33425 16609 33459 16643
rect 33459 16609 33468 16643
rect 33416 16600 33468 16609
rect 33508 16600 33560 16652
rect 33784 16600 33836 16652
rect 34152 16600 34204 16652
rect 29460 16464 29512 16516
rect 31208 16464 31260 16516
rect 27344 16396 27396 16448
rect 27804 16396 27856 16448
rect 30380 16396 30432 16448
rect 31116 16439 31168 16448
rect 31116 16405 31125 16439
rect 31125 16405 31159 16439
rect 31159 16405 31168 16439
rect 31116 16396 31168 16405
rect 31944 16464 31996 16516
rect 32220 16396 32272 16448
rect 32680 16464 32732 16516
rect 33416 16464 33468 16516
rect 34060 16396 34112 16448
rect 34428 16464 34480 16516
rect 34520 16464 34572 16516
rect 35164 16507 35216 16516
rect 35164 16473 35173 16507
rect 35173 16473 35207 16507
rect 35207 16473 35216 16507
rect 35164 16464 35216 16473
rect 35256 16507 35308 16516
rect 35256 16473 35265 16507
rect 35265 16473 35299 16507
rect 35299 16473 35308 16507
rect 35256 16464 35308 16473
rect 35348 16507 35400 16516
rect 35348 16473 35383 16507
rect 35383 16473 35400 16507
rect 35348 16464 35400 16473
rect 36084 16600 36136 16652
rect 40132 16668 40184 16720
rect 37372 16532 37424 16584
rect 37464 16575 37516 16584
rect 37464 16541 37473 16575
rect 37473 16541 37507 16575
rect 37507 16541 37516 16575
rect 37464 16532 37516 16541
rect 39212 16532 39264 16584
rect 40684 16532 40736 16584
rect 39304 16464 39356 16516
rect 36360 16396 36412 16448
rect 38384 16396 38436 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 5356 16192 5408 16244
rect 6092 16192 6144 16244
rect 9588 16192 9640 16244
rect 9680 16192 9732 16244
rect 5080 16124 5132 16176
rect 5632 16124 5684 16176
rect 9036 16124 9088 16176
rect 11244 16124 11296 16176
rect 3516 16099 3568 16108
rect 3516 16065 3525 16099
rect 3525 16065 3559 16099
rect 3559 16065 3568 16099
rect 3516 16056 3568 16065
rect 8024 16099 8076 16108
rect 8024 16065 8033 16099
rect 8033 16065 8067 16099
rect 8067 16065 8076 16099
rect 8024 16056 8076 16065
rect 3792 16031 3844 16040
rect 3792 15997 3801 16031
rect 3801 15997 3835 16031
rect 3835 15997 3844 16031
rect 3792 15988 3844 15997
rect 5264 15988 5316 16040
rect 6184 15988 6236 16040
rect 6828 15988 6880 16040
rect 8300 16031 8352 16040
rect 8300 15997 8309 16031
rect 8309 15997 8343 16031
rect 8343 15997 8352 16031
rect 8300 15988 8352 15997
rect 9036 15988 9088 16040
rect 10048 16056 10100 16108
rect 13084 16124 13136 16176
rect 13912 16192 13964 16244
rect 14648 16192 14700 16244
rect 17960 16192 18012 16244
rect 18788 16192 18840 16244
rect 13360 16099 13412 16108
rect 13360 16065 13369 16099
rect 13369 16065 13403 16099
rect 13403 16065 13412 16099
rect 13360 16056 13412 16065
rect 13544 16099 13596 16108
rect 13544 16065 13553 16099
rect 13553 16065 13587 16099
rect 13587 16065 13596 16099
rect 13544 16056 13596 16065
rect 14188 16056 14240 16108
rect 14556 16031 14608 16040
rect 14556 15997 14565 16031
rect 14565 15997 14599 16031
rect 14599 15997 14608 16031
rect 14556 15988 14608 15997
rect 14740 16031 14792 16040
rect 14740 15997 14749 16031
rect 14749 15997 14783 16031
rect 14783 15997 14792 16031
rect 14740 15988 14792 15997
rect 16948 16056 17000 16108
rect 17868 16056 17920 16108
rect 18052 16056 18104 16108
rect 16120 15988 16172 16040
rect 18420 16124 18472 16176
rect 21916 16192 21968 16244
rect 18236 16099 18288 16108
rect 18236 16065 18245 16099
rect 18245 16065 18279 16099
rect 18279 16065 18288 16099
rect 21456 16124 21508 16176
rect 23756 16192 23808 16244
rect 25228 16192 25280 16244
rect 24676 16124 24728 16176
rect 28540 16192 28592 16244
rect 33416 16192 33468 16244
rect 34612 16192 34664 16244
rect 34980 16192 35032 16244
rect 35440 16192 35492 16244
rect 37280 16192 37332 16244
rect 37556 16192 37608 16244
rect 18236 16056 18288 16065
rect 18512 16031 18564 16040
rect 18512 15997 18521 16031
rect 18521 15997 18555 16031
rect 18555 15997 18564 16031
rect 18512 15988 18564 15997
rect 18972 16056 19024 16108
rect 19248 16056 19300 16108
rect 20628 16056 20680 16108
rect 25044 16056 25096 16108
rect 25504 16056 25556 16108
rect 26700 16124 26752 16176
rect 28356 16124 28408 16176
rect 31116 16124 31168 16176
rect 31484 16124 31536 16176
rect 32864 16124 32916 16176
rect 34520 16124 34572 16176
rect 7840 15852 7892 15904
rect 12716 15895 12768 15904
rect 12716 15861 12725 15895
rect 12725 15861 12759 15895
rect 12759 15861 12768 15895
rect 12716 15852 12768 15861
rect 12900 15895 12952 15904
rect 12900 15861 12909 15895
rect 12909 15861 12943 15895
rect 12943 15861 12952 15895
rect 12900 15852 12952 15861
rect 16212 15895 16264 15904
rect 16212 15861 16221 15895
rect 16221 15861 16255 15895
rect 16255 15861 16264 15895
rect 16212 15852 16264 15861
rect 17408 15852 17460 15904
rect 17500 15852 17552 15904
rect 18512 15852 18564 15904
rect 19156 15963 19208 15972
rect 19156 15929 19165 15963
rect 19165 15929 19199 15963
rect 19199 15929 19208 15963
rect 19156 15920 19208 15929
rect 22008 15920 22060 15972
rect 22560 15920 22612 15972
rect 25320 15988 25372 16040
rect 25412 15988 25464 16040
rect 25688 16031 25740 16040
rect 25688 15997 25697 16031
rect 25697 15997 25731 16031
rect 25731 15997 25740 16031
rect 25688 15988 25740 15997
rect 25044 15920 25096 15972
rect 25872 15920 25924 15972
rect 26608 16056 26660 16108
rect 28632 16056 28684 16108
rect 30380 16056 30432 16108
rect 30932 16056 30984 16108
rect 31392 16099 31444 16108
rect 31392 16065 31401 16099
rect 31401 16065 31435 16099
rect 31435 16065 31444 16099
rect 31392 16056 31444 16065
rect 34428 16056 34480 16108
rect 35256 16124 35308 16176
rect 35624 16167 35676 16176
rect 39488 16192 39540 16244
rect 35624 16133 35659 16167
rect 35659 16133 35676 16167
rect 35624 16124 35676 16133
rect 35164 16056 35216 16108
rect 26332 15988 26384 16040
rect 28724 15988 28776 16040
rect 35440 16099 35492 16108
rect 35440 16065 35449 16099
rect 35449 16065 35483 16099
rect 35483 16065 35492 16099
rect 35440 16056 35492 16065
rect 26240 15920 26292 15972
rect 26792 15920 26844 15972
rect 35624 15988 35676 16040
rect 36084 16056 36136 16108
rect 36268 16056 36320 16108
rect 36544 16056 36596 16108
rect 37464 16056 37516 16108
rect 39028 16056 39080 16108
rect 39396 16056 39448 16108
rect 39580 15988 39632 16040
rect 39856 15920 39908 15972
rect 23940 15852 23992 15904
rect 24216 15895 24268 15904
rect 24216 15861 24225 15895
rect 24225 15861 24259 15895
rect 24259 15861 24268 15895
rect 24216 15852 24268 15861
rect 24308 15852 24360 15904
rect 30288 15852 30340 15904
rect 37372 15852 37424 15904
rect 37556 15895 37608 15904
rect 37556 15861 37565 15895
rect 37565 15861 37599 15895
rect 37599 15861 37608 15895
rect 37556 15852 37608 15861
rect 38660 15852 38712 15904
rect 39212 15895 39264 15904
rect 39212 15861 39221 15895
rect 39221 15861 39255 15895
rect 39255 15861 39264 15895
rect 39212 15852 39264 15861
rect 39672 15895 39724 15904
rect 39672 15861 39681 15895
rect 39681 15861 39715 15895
rect 39715 15861 39724 15895
rect 39672 15852 39724 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 3792 15648 3844 15700
rect 5448 15648 5500 15700
rect 6184 15648 6236 15700
rect 8300 15648 8352 15700
rect 8944 15648 8996 15700
rect 12716 15648 12768 15700
rect 12900 15648 12952 15700
rect 3332 15555 3384 15564
rect 3332 15521 3341 15555
rect 3341 15521 3375 15555
rect 3375 15521 3384 15555
rect 3332 15512 3384 15521
rect 3516 15512 3568 15564
rect 3700 15444 3752 15496
rect 4160 15487 4212 15496
rect 4160 15453 4169 15487
rect 4169 15453 4203 15487
rect 4203 15453 4212 15487
rect 4160 15444 4212 15453
rect 6276 15444 6328 15496
rect 7840 15487 7892 15496
rect 7840 15453 7849 15487
rect 7849 15453 7883 15487
rect 7883 15453 7892 15487
rect 7840 15444 7892 15453
rect 8116 15487 8168 15496
rect 8116 15453 8125 15487
rect 8125 15453 8159 15487
rect 8159 15453 8168 15487
rect 8116 15444 8168 15453
rect 8392 15444 8444 15496
rect 11612 15512 11664 15564
rect 17224 15648 17276 15700
rect 17960 15648 18012 15700
rect 18052 15648 18104 15700
rect 13268 15580 13320 15632
rect 13728 15580 13780 15632
rect 15200 15580 15252 15632
rect 3240 15376 3292 15428
rect 5632 15376 5684 15428
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 2044 15351 2096 15360
rect 2044 15317 2053 15351
rect 2053 15317 2087 15351
rect 2087 15317 2096 15351
rect 2044 15308 2096 15317
rect 2780 15308 2832 15360
rect 4068 15308 4120 15360
rect 8760 15376 8812 15428
rect 10968 15376 11020 15428
rect 11520 15376 11572 15428
rect 12900 15376 12952 15428
rect 18788 15580 18840 15632
rect 20720 15648 20772 15700
rect 22100 15648 22152 15700
rect 22744 15648 22796 15700
rect 23848 15648 23900 15700
rect 21456 15580 21508 15632
rect 15292 15444 15344 15496
rect 9956 15308 10008 15360
rect 10784 15351 10836 15360
rect 10784 15317 10793 15351
rect 10793 15317 10827 15351
rect 10827 15317 10836 15351
rect 10784 15308 10836 15317
rect 11060 15308 11112 15360
rect 14280 15308 14332 15360
rect 14464 15308 14516 15360
rect 15752 15376 15804 15428
rect 18144 15487 18196 15496
rect 18144 15453 18153 15487
rect 18153 15453 18187 15487
rect 18187 15453 18196 15487
rect 18144 15444 18196 15453
rect 18696 15444 18748 15496
rect 16856 15351 16908 15360
rect 16856 15317 16865 15351
rect 16865 15317 16899 15351
rect 16899 15317 16908 15351
rect 16856 15308 16908 15317
rect 17408 15376 17460 15428
rect 17868 15376 17920 15428
rect 21180 15444 21232 15496
rect 20720 15376 20772 15428
rect 21640 15444 21692 15496
rect 24216 15580 24268 15632
rect 25688 15648 25740 15700
rect 26884 15691 26936 15700
rect 26884 15657 26893 15691
rect 26893 15657 26927 15691
rect 26927 15657 26936 15691
rect 26884 15648 26936 15657
rect 30104 15648 30156 15700
rect 30288 15691 30340 15700
rect 30288 15657 30297 15691
rect 30297 15657 30331 15691
rect 30331 15657 30340 15691
rect 30288 15648 30340 15657
rect 32220 15648 32272 15700
rect 37464 15648 37516 15700
rect 39028 15648 39080 15700
rect 39672 15648 39724 15700
rect 39856 15691 39908 15700
rect 39856 15657 39865 15691
rect 39865 15657 39899 15691
rect 39899 15657 39908 15691
rect 39856 15648 39908 15657
rect 40592 15648 40644 15700
rect 22192 15487 22244 15496
rect 22192 15453 22201 15487
rect 22201 15453 22235 15487
rect 22235 15453 22244 15487
rect 22192 15444 22244 15453
rect 22652 15444 22704 15496
rect 24032 15444 24084 15496
rect 24400 15444 24452 15496
rect 25780 15444 25832 15496
rect 25964 15444 26016 15496
rect 26148 15555 26200 15564
rect 26148 15521 26157 15555
rect 26157 15521 26191 15555
rect 26191 15521 26200 15555
rect 26148 15512 26200 15521
rect 26240 15512 26292 15564
rect 26608 15444 26660 15496
rect 19156 15308 19208 15360
rect 19432 15308 19484 15360
rect 21180 15308 21232 15360
rect 21548 15351 21600 15360
rect 21548 15317 21557 15351
rect 21557 15317 21591 15351
rect 21591 15317 21600 15351
rect 21548 15308 21600 15317
rect 21732 15308 21784 15360
rect 23664 15351 23716 15360
rect 23664 15317 23673 15351
rect 23673 15317 23707 15351
rect 23707 15317 23716 15351
rect 23664 15308 23716 15317
rect 26148 15376 26200 15428
rect 26792 15487 26844 15496
rect 26792 15453 26801 15487
rect 26801 15453 26835 15487
rect 26835 15453 26844 15487
rect 26792 15444 26844 15453
rect 26976 15555 27028 15564
rect 26976 15521 26985 15555
rect 26985 15521 27019 15555
rect 27019 15521 27028 15555
rect 26976 15512 27028 15521
rect 30196 15623 30248 15632
rect 30196 15589 30205 15623
rect 30205 15589 30239 15623
rect 30239 15589 30248 15623
rect 30196 15580 30248 15589
rect 34520 15580 34572 15632
rect 27252 15444 27304 15496
rect 30104 15487 30156 15496
rect 30104 15453 30113 15487
rect 30113 15453 30147 15487
rect 30147 15453 30156 15487
rect 30104 15444 30156 15453
rect 30380 15444 30432 15496
rect 37188 15512 37240 15564
rect 30840 15444 30892 15496
rect 31760 15444 31812 15496
rect 32588 15487 32640 15496
rect 32588 15453 32597 15487
rect 32597 15453 32631 15487
rect 32631 15453 32640 15487
rect 32588 15444 32640 15453
rect 33600 15444 33652 15496
rect 35624 15487 35676 15496
rect 35624 15453 35633 15487
rect 35633 15453 35667 15487
rect 35667 15453 35676 15487
rect 35624 15444 35676 15453
rect 31208 15376 31260 15428
rect 34060 15376 34112 15428
rect 35348 15376 35400 15428
rect 26332 15308 26384 15360
rect 26884 15308 26936 15360
rect 29736 15308 29788 15360
rect 30196 15308 30248 15360
rect 31668 15308 31720 15360
rect 32312 15308 32364 15360
rect 34244 15308 34296 15360
rect 34612 15308 34664 15360
rect 35624 15308 35676 15360
rect 35900 15376 35952 15428
rect 36084 15376 36136 15428
rect 37004 15444 37056 15496
rect 37464 15487 37516 15496
rect 37464 15453 37471 15487
rect 37471 15453 37516 15487
rect 37464 15444 37516 15453
rect 38936 15444 38988 15496
rect 39764 15512 39816 15564
rect 38384 15376 38436 15428
rect 37188 15308 37240 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 2044 15104 2096 15156
rect 3700 15104 3752 15156
rect 3976 15104 4028 15156
rect 3148 15036 3200 15088
rect 5632 15036 5684 15088
rect 8024 15104 8076 15156
rect 10784 15104 10836 15156
rect 10968 15147 11020 15156
rect 10968 15113 10977 15147
rect 10977 15113 11011 15147
rect 11011 15113 11020 15147
rect 10968 15104 11020 15113
rect 11428 15104 11480 15156
rect 12900 15147 12952 15156
rect 12900 15113 12909 15147
rect 12909 15113 12943 15147
rect 12943 15113 12952 15147
rect 12900 15104 12952 15113
rect 15292 15147 15344 15156
rect 15292 15113 15301 15147
rect 15301 15113 15335 15147
rect 15335 15113 15344 15147
rect 15292 15104 15344 15113
rect 15844 15104 15896 15156
rect 19616 15104 19668 15156
rect 13636 15036 13688 15088
rect 8392 15011 8444 15020
rect 8392 14977 8401 15011
rect 8401 14977 8435 15011
rect 8435 14977 8444 15011
rect 8392 14968 8444 14977
rect 8484 15011 8536 15020
rect 8484 14977 8493 15011
rect 8493 14977 8527 15011
rect 8527 14977 8536 15011
rect 8484 14968 8536 14977
rect 6276 14900 6328 14952
rect 1584 14764 1636 14816
rect 6736 14900 6788 14952
rect 9128 14832 9180 14884
rect 11060 15011 11112 15020
rect 11060 14977 11069 15011
rect 11069 14977 11103 15011
rect 11103 14977 11112 15011
rect 11060 14968 11112 14977
rect 10784 14900 10836 14952
rect 11152 14943 11204 14952
rect 11152 14909 11161 14943
rect 11161 14909 11195 14943
rect 11195 14909 11204 14943
rect 11152 14900 11204 14909
rect 12440 14900 12492 14952
rect 6644 14764 6696 14816
rect 8576 14807 8628 14816
rect 8576 14773 8585 14807
rect 8585 14773 8619 14807
rect 8619 14773 8628 14807
rect 8576 14764 8628 14773
rect 9404 14764 9456 14816
rect 10600 14807 10652 14816
rect 10600 14773 10609 14807
rect 10609 14773 10643 14807
rect 10643 14773 10652 14807
rect 10600 14764 10652 14773
rect 11060 14764 11112 14816
rect 11428 14764 11480 14816
rect 12900 14764 12952 14816
rect 14464 14968 14516 15020
rect 15108 15036 15160 15088
rect 16120 15079 16172 15088
rect 16120 15045 16129 15079
rect 16129 15045 16163 15079
rect 16163 15045 16172 15079
rect 16120 15036 16172 15045
rect 16856 15036 16908 15088
rect 17224 15036 17276 15088
rect 18328 15036 18380 15088
rect 18788 15036 18840 15088
rect 15016 14968 15068 15020
rect 16580 14968 16632 15020
rect 14004 14900 14056 14952
rect 15568 14943 15620 14952
rect 15568 14909 15577 14943
rect 15577 14909 15611 14943
rect 15611 14909 15620 14943
rect 15568 14900 15620 14909
rect 16304 14900 16356 14952
rect 16948 14900 17000 14952
rect 17316 14900 17368 14952
rect 19432 15036 19484 15088
rect 20168 15104 20220 15156
rect 21272 15104 21324 15156
rect 20352 15036 20404 15088
rect 19524 15011 19576 15020
rect 19524 14977 19533 15011
rect 19533 14977 19567 15011
rect 19567 14977 19576 15011
rect 19524 14968 19576 14977
rect 20904 15036 20956 15088
rect 20812 14968 20864 15020
rect 22008 15104 22060 15156
rect 22192 15104 22244 15156
rect 23664 15104 23716 15156
rect 26240 15104 26292 15156
rect 26792 15104 26844 15156
rect 27068 15104 27120 15156
rect 28448 15147 28500 15156
rect 28448 15113 28457 15147
rect 28457 15113 28491 15147
rect 28491 15113 28500 15147
rect 28448 15104 28500 15113
rect 29276 15104 29328 15156
rect 32220 15104 32272 15156
rect 32404 15104 32456 15156
rect 21824 15036 21876 15088
rect 13360 14764 13412 14816
rect 16488 14764 16540 14816
rect 17316 14764 17368 14816
rect 17592 14764 17644 14816
rect 18696 14832 18748 14884
rect 18328 14764 18380 14816
rect 19248 14832 19300 14884
rect 22008 15011 22060 15020
rect 22008 14977 22017 15011
rect 22017 14977 22051 15011
rect 22051 14977 22060 15011
rect 22008 14968 22060 14977
rect 22744 14968 22796 15020
rect 23664 14968 23716 15020
rect 23940 14968 23992 15020
rect 25964 15036 26016 15088
rect 24308 14968 24360 15020
rect 24400 14968 24452 15020
rect 26240 14968 26292 15020
rect 19340 14807 19392 14816
rect 19340 14773 19349 14807
rect 19349 14773 19383 14807
rect 19383 14773 19392 14807
rect 19340 14764 19392 14773
rect 19432 14764 19484 14816
rect 20536 14764 20588 14816
rect 21640 14832 21692 14884
rect 25136 14900 25188 14952
rect 25964 14900 26016 14952
rect 24676 14832 24728 14884
rect 26516 14900 26568 14952
rect 27896 15011 27948 15020
rect 27896 14977 27905 15011
rect 27905 14977 27939 15011
rect 27939 14977 27948 15011
rect 27896 14968 27948 14977
rect 28264 15079 28316 15088
rect 28264 15045 28273 15079
rect 28273 15045 28307 15079
rect 28307 15045 28316 15079
rect 28264 15036 28316 15045
rect 28908 14968 28960 15020
rect 29644 14968 29696 15020
rect 29828 15036 29880 15088
rect 31576 14968 31628 15020
rect 31852 14968 31904 15020
rect 33232 15036 33284 15088
rect 38660 15104 38712 15156
rect 38752 15104 38804 15156
rect 26148 14832 26200 14884
rect 27160 14832 27212 14884
rect 27344 14875 27396 14884
rect 27344 14841 27353 14875
rect 27353 14841 27387 14875
rect 27387 14841 27396 14875
rect 27344 14832 27396 14841
rect 27620 14832 27672 14884
rect 22008 14764 22060 14816
rect 22284 14807 22336 14816
rect 22284 14773 22293 14807
rect 22293 14773 22327 14807
rect 22327 14773 22336 14807
rect 22284 14764 22336 14773
rect 22560 14807 22612 14816
rect 22560 14773 22569 14807
rect 22569 14773 22603 14807
rect 22603 14773 22612 14807
rect 22560 14764 22612 14773
rect 23296 14807 23348 14816
rect 23296 14773 23305 14807
rect 23305 14773 23339 14807
rect 23339 14773 23348 14807
rect 23296 14764 23348 14773
rect 23572 14807 23624 14816
rect 23572 14773 23581 14807
rect 23581 14773 23615 14807
rect 23615 14773 23624 14807
rect 23572 14764 23624 14773
rect 23664 14807 23716 14816
rect 23664 14773 23673 14807
rect 23673 14773 23707 14807
rect 23707 14773 23716 14807
rect 23664 14764 23716 14773
rect 23756 14764 23808 14816
rect 24124 14807 24176 14816
rect 24124 14773 24133 14807
rect 24133 14773 24167 14807
rect 24167 14773 24176 14807
rect 24124 14764 24176 14773
rect 24308 14764 24360 14816
rect 29460 14900 29512 14952
rect 29920 14900 29972 14952
rect 30932 14900 30984 14952
rect 29092 14832 29144 14884
rect 29184 14875 29236 14884
rect 29184 14841 29193 14875
rect 29193 14841 29227 14875
rect 29227 14841 29236 14875
rect 29184 14832 29236 14841
rect 31668 14832 31720 14884
rect 31760 14832 31812 14884
rect 32220 14832 32272 14884
rect 32864 14968 32916 15020
rect 32772 14943 32824 14952
rect 32772 14909 32781 14943
rect 32781 14909 32815 14943
rect 32815 14909 32824 14943
rect 32772 14900 32824 14909
rect 32680 14832 32732 14884
rect 33600 14968 33652 15020
rect 33876 15011 33928 15020
rect 33876 14977 33890 15011
rect 33890 14977 33924 15011
rect 33924 14977 33928 15011
rect 33876 14968 33928 14977
rect 34244 14968 34296 15020
rect 35256 14968 35308 15020
rect 37648 14968 37700 15020
rect 38108 14968 38160 15020
rect 38384 15036 38436 15088
rect 38568 15079 38620 15088
rect 38568 15045 38577 15079
rect 38577 15045 38611 15079
rect 38611 15045 38620 15079
rect 38568 15036 38620 15045
rect 34428 14900 34480 14952
rect 35716 14900 35768 14952
rect 38936 14968 38988 15020
rect 39396 14968 39448 15020
rect 38476 14900 38528 14952
rect 28356 14764 28408 14816
rect 29920 14764 29972 14816
rect 32036 14764 32088 14816
rect 33140 14764 33192 14816
rect 34428 14764 34480 14816
rect 37004 14764 37056 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 4068 14560 4120 14612
rect 8484 14560 8536 14612
rect 3240 14424 3292 14476
rect 14648 14492 14700 14544
rect 14924 14560 14976 14612
rect 16028 14560 16080 14612
rect 16488 14560 16540 14612
rect 16948 14560 17000 14612
rect 17684 14560 17736 14612
rect 17960 14560 18012 14612
rect 18144 14560 18196 14612
rect 15568 14492 15620 14544
rect 17500 14492 17552 14544
rect 19432 14492 19484 14544
rect 19616 14603 19668 14612
rect 19616 14569 19625 14603
rect 19625 14569 19659 14603
rect 19659 14569 19668 14603
rect 19616 14560 19668 14569
rect 20628 14560 20680 14612
rect 23664 14560 23716 14612
rect 25780 14603 25832 14612
rect 25780 14569 25789 14603
rect 25789 14569 25823 14603
rect 25823 14569 25832 14603
rect 25780 14560 25832 14569
rect 26884 14560 26936 14612
rect 19800 14492 19852 14544
rect 19984 14492 20036 14544
rect 21272 14492 21324 14544
rect 6276 14424 6328 14476
rect 7932 14424 7984 14476
rect 9220 14424 9272 14476
rect 10600 14356 10652 14408
rect 10968 14467 11020 14476
rect 10968 14433 10977 14467
rect 10977 14433 11011 14467
rect 11011 14433 11020 14467
rect 10968 14424 11020 14433
rect 12440 14424 12492 14476
rect 7840 14288 7892 14340
rect 9864 14288 9916 14340
rect 10876 14288 10928 14340
rect 11060 14288 11112 14340
rect 12256 14288 12308 14340
rect 14280 14356 14332 14408
rect 2780 14220 2832 14272
rect 7656 14263 7708 14272
rect 7656 14229 7665 14263
rect 7665 14229 7699 14263
rect 7699 14229 7708 14263
rect 7656 14220 7708 14229
rect 9036 14220 9088 14272
rect 11980 14263 12032 14272
rect 11980 14229 11989 14263
rect 11989 14229 12023 14263
rect 12023 14229 12032 14263
rect 14924 14356 14976 14408
rect 11980 14220 12032 14229
rect 17408 14356 17460 14408
rect 17592 14331 17644 14340
rect 17592 14297 17601 14331
rect 17601 14297 17635 14331
rect 17635 14297 17644 14331
rect 17592 14288 17644 14297
rect 17960 14356 18012 14408
rect 22560 14492 22612 14544
rect 23572 14492 23624 14544
rect 24308 14492 24360 14544
rect 24400 14535 24452 14544
rect 24400 14501 24409 14535
rect 24409 14501 24443 14535
rect 24443 14501 24452 14535
rect 24400 14492 24452 14501
rect 18420 14356 18472 14408
rect 18880 14356 18932 14408
rect 19248 14356 19300 14408
rect 19432 14288 19484 14340
rect 20352 14356 20404 14408
rect 20536 14399 20588 14408
rect 20536 14365 20545 14399
rect 20545 14365 20579 14399
rect 20579 14365 20588 14399
rect 20536 14356 20588 14365
rect 15292 14263 15344 14272
rect 15292 14229 15301 14263
rect 15301 14229 15335 14263
rect 15335 14229 15344 14263
rect 15292 14220 15344 14229
rect 17408 14263 17460 14272
rect 17408 14229 17417 14263
rect 17417 14229 17451 14263
rect 17451 14229 17460 14263
rect 17408 14220 17460 14229
rect 17960 14263 18012 14272
rect 17960 14229 17969 14263
rect 17969 14229 18003 14263
rect 18003 14229 18012 14263
rect 17960 14220 18012 14229
rect 18420 14220 18472 14272
rect 18696 14220 18748 14272
rect 19064 14220 19116 14272
rect 20720 14288 20772 14340
rect 23756 14424 23808 14476
rect 24124 14424 24176 14476
rect 23296 14356 23348 14408
rect 27068 14560 27120 14612
rect 27436 14603 27488 14612
rect 27436 14569 27445 14603
rect 27445 14569 27479 14603
rect 27479 14569 27488 14603
rect 27436 14560 27488 14569
rect 27896 14560 27948 14612
rect 29184 14560 29236 14612
rect 30656 14560 30708 14612
rect 22744 14288 22796 14340
rect 24676 14399 24728 14408
rect 24676 14365 24685 14399
rect 24685 14365 24719 14399
rect 24719 14365 24728 14399
rect 24676 14356 24728 14365
rect 24952 14356 25004 14408
rect 24492 14288 24544 14340
rect 24768 14288 24820 14340
rect 25228 14288 25280 14340
rect 25504 14399 25556 14408
rect 25504 14365 25513 14399
rect 25513 14365 25547 14399
rect 25547 14365 25556 14399
rect 25504 14356 25556 14365
rect 25780 14356 25832 14408
rect 25964 14399 26016 14408
rect 25964 14365 25973 14399
rect 25973 14365 26007 14399
rect 26007 14365 26016 14399
rect 25964 14356 26016 14365
rect 28264 14492 28316 14544
rect 27896 14424 27948 14476
rect 27712 14356 27764 14408
rect 31484 14492 31536 14544
rect 33692 14560 33744 14612
rect 35992 14560 36044 14612
rect 36268 14560 36320 14612
rect 37096 14560 37148 14612
rect 38200 14560 38252 14612
rect 38660 14603 38712 14612
rect 38660 14569 38669 14603
rect 38669 14569 38703 14603
rect 38703 14569 38712 14603
rect 38660 14560 38712 14569
rect 39764 14560 39816 14612
rect 31944 14535 31996 14544
rect 31944 14501 31953 14535
rect 31953 14501 31987 14535
rect 31987 14501 31996 14535
rect 31944 14492 31996 14501
rect 40316 14603 40368 14612
rect 40316 14569 40325 14603
rect 40325 14569 40359 14603
rect 40359 14569 40368 14603
rect 40316 14560 40368 14569
rect 30380 14356 30432 14408
rect 30840 14399 30892 14408
rect 30840 14365 30849 14399
rect 30849 14365 30883 14399
rect 30883 14365 30892 14399
rect 30840 14356 30892 14365
rect 30932 14399 30984 14408
rect 30932 14365 30941 14399
rect 30941 14365 30975 14399
rect 30975 14365 30984 14399
rect 30932 14356 30984 14365
rect 31024 14399 31076 14408
rect 31024 14365 31033 14399
rect 31033 14365 31067 14399
rect 31067 14365 31076 14399
rect 31024 14356 31076 14365
rect 31300 14399 31352 14408
rect 31300 14365 31309 14399
rect 31309 14365 31343 14399
rect 31343 14365 31352 14399
rect 31300 14356 31352 14365
rect 31484 14399 31536 14408
rect 31484 14365 31491 14399
rect 31491 14365 31536 14399
rect 31484 14356 31536 14365
rect 31576 14399 31628 14408
rect 31576 14365 31585 14399
rect 31585 14365 31619 14399
rect 31619 14365 31628 14399
rect 31576 14356 31628 14365
rect 31668 14399 31720 14408
rect 31668 14365 31677 14399
rect 31677 14365 31711 14399
rect 31711 14365 31720 14399
rect 31668 14356 31720 14365
rect 32404 14356 32456 14408
rect 32496 14356 32548 14408
rect 33416 14356 33468 14408
rect 34336 14424 34388 14476
rect 34612 14424 34664 14476
rect 34244 14356 34296 14408
rect 26700 14288 26752 14340
rect 23020 14263 23072 14272
rect 23020 14229 23029 14263
rect 23029 14229 23063 14263
rect 23063 14229 23072 14263
rect 23020 14220 23072 14229
rect 25412 14220 25464 14272
rect 25872 14220 25924 14272
rect 27436 14263 27488 14272
rect 27436 14229 27445 14263
rect 27445 14229 27479 14263
rect 27479 14229 27488 14263
rect 27436 14220 27488 14229
rect 27804 14288 27856 14340
rect 30564 14288 30616 14340
rect 33692 14331 33744 14340
rect 33692 14297 33701 14331
rect 33701 14297 33735 14331
rect 33735 14297 33744 14331
rect 33692 14288 33744 14297
rect 34428 14288 34480 14340
rect 35440 14356 35492 14408
rect 38752 14467 38804 14476
rect 38752 14433 38761 14467
rect 38761 14433 38795 14467
rect 38795 14433 38804 14467
rect 38752 14424 38804 14433
rect 39948 14467 40000 14476
rect 39948 14433 39957 14467
rect 39957 14433 39991 14467
rect 39991 14433 40000 14467
rect 39948 14424 40000 14433
rect 36912 14399 36964 14408
rect 36912 14365 36921 14399
rect 36921 14365 36955 14399
rect 36955 14365 36964 14399
rect 36912 14356 36964 14365
rect 37004 14356 37056 14408
rect 37832 14356 37884 14408
rect 38844 14399 38896 14408
rect 38844 14365 38853 14399
rect 38853 14365 38887 14399
rect 38887 14365 38896 14399
rect 38844 14356 38896 14365
rect 39212 14356 39264 14408
rect 40040 14356 40092 14408
rect 35072 14331 35124 14340
rect 35072 14297 35081 14331
rect 35081 14297 35115 14331
rect 35115 14297 35124 14331
rect 35072 14288 35124 14297
rect 35164 14331 35216 14340
rect 35164 14297 35199 14331
rect 35199 14297 35216 14331
rect 35164 14288 35216 14297
rect 35532 14288 35584 14340
rect 35624 14288 35676 14340
rect 35992 14288 36044 14340
rect 28172 14220 28224 14272
rect 28540 14220 28592 14272
rect 28908 14220 28960 14272
rect 30196 14220 30248 14272
rect 31300 14220 31352 14272
rect 32128 14220 32180 14272
rect 32772 14220 32824 14272
rect 33600 14220 33652 14272
rect 33968 14220 34020 14272
rect 34704 14263 34756 14272
rect 34704 14229 34713 14263
rect 34713 14229 34747 14263
rect 34747 14229 34756 14263
rect 34704 14220 34756 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 1584 14016 1636 14068
rect 3516 14016 3568 14068
rect 6736 14016 6788 14068
rect 7656 14016 7708 14068
rect 3148 13948 3200 14000
rect 3240 13948 3292 14000
rect 1768 13855 1820 13864
rect 1768 13821 1777 13855
rect 1777 13821 1811 13855
rect 1811 13821 1820 13855
rect 1768 13812 1820 13821
rect 5632 13948 5684 14000
rect 5356 13923 5408 13932
rect 5356 13889 5365 13923
rect 5365 13889 5399 13923
rect 5399 13889 5408 13923
rect 5356 13880 5408 13889
rect 3700 13855 3752 13864
rect 3700 13821 3709 13855
rect 3709 13821 3743 13855
rect 3743 13821 3752 13855
rect 3700 13812 3752 13821
rect 6552 13923 6604 13932
rect 6552 13889 6561 13923
rect 6561 13889 6595 13923
rect 6595 13889 6604 13923
rect 6552 13880 6604 13889
rect 6736 13923 6788 13932
rect 6736 13889 6745 13923
rect 6745 13889 6779 13923
rect 6779 13889 6788 13923
rect 6736 13880 6788 13889
rect 7840 13880 7892 13932
rect 7932 13923 7984 13932
rect 7932 13889 7941 13923
rect 7941 13889 7975 13923
rect 7975 13889 7984 13923
rect 7932 13880 7984 13889
rect 8852 13991 8904 14000
rect 8852 13957 8861 13991
rect 8861 13957 8895 13991
rect 8895 13957 8904 13991
rect 8852 13948 8904 13957
rect 9036 13948 9088 14000
rect 9864 14016 9916 14068
rect 12348 13948 12400 14000
rect 13176 13948 13228 14000
rect 16580 13948 16632 14000
rect 7104 13812 7156 13864
rect 9128 13880 9180 13932
rect 8576 13812 8628 13864
rect 9220 13812 9272 13864
rect 9404 13923 9456 13932
rect 9404 13889 9413 13923
rect 9413 13889 9447 13923
rect 9447 13889 9456 13923
rect 9404 13880 9456 13889
rect 12164 13880 12216 13932
rect 9496 13812 9548 13864
rect 12808 13923 12860 13932
rect 12808 13889 12817 13923
rect 12817 13889 12851 13923
rect 12851 13889 12860 13923
rect 12808 13880 12860 13889
rect 12992 13923 13044 13932
rect 12992 13889 13001 13923
rect 13001 13889 13035 13923
rect 13035 13889 13044 13923
rect 12992 13880 13044 13889
rect 16764 13880 16816 13932
rect 17684 13923 17736 13932
rect 17684 13889 17693 13923
rect 17693 13889 17727 13923
rect 17727 13889 17736 13923
rect 17684 13880 17736 13889
rect 13084 13812 13136 13864
rect 5540 13744 5592 13796
rect 7288 13744 7340 13796
rect 6000 13719 6052 13728
rect 6000 13685 6009 13719
rect 6009 13685 6043 13719
rect 6043 13685 6052 13719
rect 6000 13676 6052 13685
rect 6828 13676 6880 13728
rect 7012 13676 7064 13728
rect 8484 13676 8536 13728
rect 8668 13744 8720 13796
rect 12072 13744 12124 13796
rect 18144 13880 18196 13932
rect 19340 14016 19392 14068
rect 20720 14016 20772 14068
rect 22008 14016 22060 14068
rect 24952 14016 25004 14068
rect 25780 14059 25832 14068
rect 25780 14025 25789 14059
rect 25789 14025 25823 14059
rect 25823 14025 25832 14059
rect 25780 14016 25832 14025
rect 19800 13923 19852 13932
rect 19800 13889 19809 13923
rect 19809 13889 19843 13923
rect 19843 13889 19852 13923
rect 19800 13880 19852 13889
rect 19984 13880 20036 13932
rect 22836 13948 22888 14000
rect 25044 13948 25096 14000
rect 18328 13855 18380 13864
rect 17316 13744 17368 13796
rect 18328 13821 18337 13855
rect 18337 13821 18371 13855
rect 18371 13821 18380 13855
rect 18328 13812 18380 13821
rect 19708 13812 19760 13864
rect 25596 13880 25648 13932
rect 25780 13880 25832 13932
rect 27344 14016 27396 14068
rect 27712 14059 27764 14068
rect 27712 14025 27721 14059
rect 27721 14025 27755 14059
rect 27755 14025 27764 14059
rect 27712 14016 27764 14025
rect 27804 14016 27856 14068
rect 28080 14016 28132 14068
rect 28448 14016 28500 14068
rect 29368 14016 29420 14068
rect 29920 14059 29972 14068
rect 29920 14025 29929 14059
rect 29929 14025 29963 14059
rect 29963 14025 29972 14059
rect 29920 14016 29972 14025
rect 30472 14016 30524 14068
rect 31392 14016 31444 14068
rect 26516 13880 26568 13932
rect 26976 13923 27028 13932
rect 26976 13889 26985 13923
rect 26985 13889 27019 13923
rect 27019 13889 27028 13923
rect 26976 13880 27028 13889
rect 27068 13880 27120 13932
rect 18696 13744 18748 13796
rect 10232 13676 10284 13728
rect 13544 13676 13596 13728
rect 14832 13676 14884 13728
rect 18052 13676 18104 13728
rect 20812 13744 20864 13796
rect 25228 13744 25280 13796
rect 19064 13719 19116 13728
rect 19064 13685 19073 13719
rect 19073 13685 19107 13719
rect 19107 13685 19116 13719
rect 19064 13676 19116 13685
rect 19432 13676 19484 13728
rect 26424 13787 26476 13796
rect 26424 13753 26433 13787
rect 26433 13753 26467 13787
rect 26467 13753 26476 13787
rect 26424 13744 26476 13753
rect 26608 13744 26660 13796
rect 26792 13744 26844 13796
rect 27620 13812 27672 13864
rect 27712 13812 27764 13864
rect 28172 13923 28224 13932
rect 28172 13889 28181 13923
rect 28181 13889 28215 13923
rect 28215 13889 28224 13923
rect 28172 13880 28224 13889
rect 28908 13880 28960 13932
rect 29736 13880 29788 13932
rect 29920 13880 29972 13932
rect 31024 13923 31076 13932
rect 31024 13889 31033 13923
rect 31033 13889 31067 13923
rect 31067 13889 31076 13923
rect 31024 13880 31076 13889
rect 30012 13855 30064 13864
rect 30012 13821 30021 13855
rect 30021 13821 30055 13855
rect 30055 13821 30064 13855
rect 30012 13812 30064 13821
rect 32036 13948 32088 14000
rect 32588 14059 32640 14068
rect 32588 14025 32597 14059
rect 32597 14025 32631 14059
rect 32631 14025 32640 14059
rect 32588 14016 32640 14025
rect 33784 13948 33836 14000
rect 34704 14016 34756 14068
rect 31760 13880 31812 13932
rect 32680 13880 32732 13932
rect 33140 13880 33192 13932
rect 30104 13744 30156 13796
rect 32864 13812 32916 13864
rect 37188 14016 37240 14068
rect 37556 13991 37608 14000
rect 37556 13957 37565 13991
rect 37565 13957 37599 13991
rect 37599 13957 37608 13991
rect 37556 13948 37608 13957
rect 35164 13880 35216 13932
rect 32496 13744 32548 13796
rect 33232 13744 33284 13796
rect 34152 13744 34204 13796
rect 34428 13744 34480 13796
rect 35716 13812 35768 13864
rect 35992 13923 36044 13932
rect 35992 13889 36001 13923
rect 36001 13889 36035 13923
rect 36035 13889 36044 13923
rect 35992 13880 36044 13889
rect 36084 13923 36136 13932
rect 36084 13889 36119 13923
rect 36119 13889 36136 13923
rect 36084 13880 36136 13889
rect 36268 13923 36320 13932
rect 36268 13889 36277 13923
rect 36277 13889 36311 13923
rect 36311 13889 36320 13923
rect 36268 13880 36320 13889
rect 36912 13880 36964 13932
rect 37280 13923 37332 13932
rect 37280 13889 37289 13923
rect 37289 13889 37323 13923
rect 37323 13889 37332 13923
rect 37280 13880 37332 13889
rect 37832 14059 37884 14068
rect 37832 14025 37841 14059
rect 37841 14025 37875 14059
rect 37875 14025 37884 14059
rect 37832 14016 37884 14025
rect 39488 13880 39540 13932
rect 38936 13812 38988 13864
rect 39120 13812 39172 13864
rect 28172 13676 28224 13728
rect 32128 13719 32180 13728
rect 32128 13685 32137 13719
rect 32137 13685 32171 13719
rect 32171 13685 32180 13719
rect 32128 13676 32180 13685
rect 34520 13719 34572 13728
rect 34520 13685 34529 13719
rect 34529 13685 34563 13719
rect 34563 13685 34572 13719
rect 34520 13676 34572 13685
rect 36452 13744 36504 13796
rect 36728 13744 36780 13796
rect 37004 13744 37056 13796
rect 35624 13719 35676 13728
rect 35624 13685 35633 13719
rect 35633 13685 35667 13719
rect 35667 13685 35676 13719
rect 35624 13676 35676 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 1768 13472 1820 13524
rect 3700 13472 3752 13524
rect 6552 13472 6604 13524
rect 6828 13472 6880 13524
rect 8300 13472 8352 13524
rect 10784 13472 10836 13524
rect 14648 13472 14700 13524
rect 2780 13268 2832 13320
rect 6092 13404 6144 13456
rect 6736 13404 6788 13456
rect 5264 13311 5316 13320
rect 5264 13277 5273 13311
rect 5273 13277 5307 13311
rect 5307 13277 5316 13311
rect 5264 13268 5316 13277
rect 5448 13311 5500 13320
rect 5448 13277 5457 13311
rect 5457 13277 5491 13311
rect 5491 13277 5500 13311
rect 5448 13268 5500 13277
rect 5540 13268 5592 13320
rect 6000 13268 6052 13320
rect 6460 13268 6512 13320
rect 7012 13268 7064 13320
rect 7932 13404 7984 13456
rect 8116 13404 8168 13456
rect 10416 13404 10468 13456
rect 7656 13311 7708 13320
rect 7656 13277 7665 13311
rect 7665 13277 7699 13311
rect 7699 13277 7708 13311
rect 7656 13268 7708 13277
rect 8852 13336 8904 13388
rect 8116 13268 8168 13320
rect 8668 13268 8720 13320
rect 8944 13311 8996 13320
rect 8944 13277 8953 13311
rect 8953 13277 8987 13311
rect 8987 13277 8996 13311
rect 8944 13268 8996 13277
rect 9404 13336 9456 13388
rect 10600 13379 10652 13388
rect 10600 13345 10609 13379
rect 10609 13345 10643 13379
rect 10643 13345 10652 13379
rect 10600 13336 10652 13345
rect 7380 13243 7432 13252
rect 7380 13209 7389 13243
rect 7389 13209 7423 13243
rect 7423 13209 7432 13243
rect 7380 13200 7432 13209
rect 6736 13175 6788 13184
rect 6736 13141 6745 13175
rect 6745 13141 6779 13175
rect 6779 13141 6788 13175
rect 6736 13132 6788 13141
rect 7196 13175 7248 13184
rect 7196 13141 7205 13175
rect 7205 13141 7239 13175
rect 7239 13141 7248 13175
rect 7196 13132 7248 13141
rect 8024 13175 8076 13184
rect 8024 13141 8033 13175
rect 8033 13141 8067 13175
rect 8067 13141 8076 13175
rect 8024 13132 8076 13141
rect 8392 13243 8444 13252
rect 8392 13209 8401 13243
rect 8401 13209 8435 13243
rect 8435 13209 8444 13243
rect 8392 13200 8444 13209
rect 8484 13243 8536 13252
rect 8484 13209 8493 13243
rect 8493 13209 8527 13243
rect 8527 13209 8536 13243
rect 8484 13200 8536 13209
rect 9404 13200 9456 13252
rect 9864 13268 9916 13320
rect 11060 13311 11112 13320
rect 11060 13277 11069 13311
rect 11069 13277 11103 13311
rect 11103 13277 11112 13311
rect 11060 13268 11112 13277
rect 11152 13268 11204 13320
rect 11888 13268 11940 13320
rect 11980 13311 12032 13320
rect 11980 13277 11989 13311
rect 11989 13277 12023 13311
rect 12023 13277 12032 13311
rect 11980 13268 12032 13277
rect 12164 13268 12216 13320
rect 9036 13132 9088 13184
rect 9496 13132 9548 13184
rect 9680 13132 9732 13184
rect 10508 13175 10560 13184
rect 10508 13141 10517 13175
rect 10517 13141 10551 13175
rect 10551 13141 10560 13175
rect 10508 13132 10560 13141
rect 10600 13132 10652 13184
rect 11980 13132 12032 13184
rect 12164 13132 12216 13184
rect 12532 13311 12584 13320
rect 12532 13277 12541 13311
rect 12541 13277 12575 13311
rect 12575 13277 12584 13311
rect 12532 13268 12584 13277
rect 12992 13404 13044 13456
rect 16028 13472 16080 13524
rect 16396 13515 16448 13524
rect 16396 13481 16405 13515
rect 16405 13481 16439 13515
rect 16439 13481 16448 13515
rect 16396 13472 16448 13481
rect 13084 13379 13136 13388
rect 13084 13345 13093 13379
rect 13093 13345 13127 13379
rect 13127 13345 13136 13379
rect 13084 13336 13136 13345
rect 12808 13200 12860 13252
rect 13176 13311 13228 13320
rect 13176 13277 13185 13311
rect 13185 13277 13219 13311
rect 13219 13277 13228 13311
rect 13176 13268 13228 13277
rect 15292 13404 15344 13456
rect 17224 13472 17276 13524
rect 13636 13200 13688 13252
rect 14004 13200 14056 13252
rect 14096 13200 14148 13252
rect 14188 13200 14240 13252
rect 16672 13336 16724 13388
rect 15660 13311 15712 13320
rect 15660 13277 15669 13311
rect 15669 13277 15703 13311
rect 15703 13277 15712 13311
rect 15660 13268 15712 13277
rect 20812 13404 20864 13456
rect 17408 13336 17460 13388
rect 19984 13336 20036 13388
rect 12624 13132 12676 13184
rect 14280 13132 14332 13184
rect 15384 13175 15436 13184
rect 15384 13141 15393 13175
rect 15393 13141 15427 13175
rect 15427 13141 15436 13175
rect 15384 13132 15436 13141
rect 17592 13268 17644 13320
rect 17684 13268 17736 13320
rect 18144 13268 18196 13320
rect 19708 13268 19760 13320
rect 20812 13243 20864 13252
rect 20812 13209 20821 13243
rect 20821 13209 20855 13243
rect 20855 13209 20864 13243
rect 20812 13200 20864 13209
rect 15844 13132 15896 13184
rect 17684 13175 17736 13184
rect 17684 13141 17693 13175
rect 17693 13141 17727 13175
rect 17727 13141 17736 13175
rect 17684 13132 17736 13141
rect 22192 13404 22244 13456
rect 23020 13472 23072 13524
rect 26976 13472 27028 13524
rect 27712 13472 27764 13524
rect 28172 13472 28224 13524
rect 29368 13472 29420 13524
rect 32864 13472 32916 13524
rect 34612 13472 34664 13524
rect 35808 13515 35860 13524
rect 35808 13481 35817 13515
rect 35817 13481 35851 13515
rect 35851 13481 35860 13515
rect 35808 13472 35860 13481
rect 37924 13472 37976 13524
rect 39856 13515 39908 13524
rect 39856 13481 39865 13515
rect 39865 13481 39899 13515
rect 39899 13481 39908 13515
rect 39856 13472 39908 13481
rect 40040 13472 40092 13524
rect 26792 13404 26844 13456
rect 31484 13404 31536 13456
rect 33232 13404 33284 13456
rect 21272 13268 21324 13320
rect 32680 13336 32732 13388
rect 33876 13336 33928 13388
rect 22192 13243 22244 13252
rect 22192 13209 22201 13243
rect 22201 13209 22235 13243
rect 22235 13209 22244 13243
rect 22192 13200 22244 13209
rect 21180 13175 21232 13184
rect 21180 13141 21189 13175
rect 21189 13141 21223 13175
rect 21223 13141 21232 13175
rect 21180 13132 21232 13141
rect 22744 13268 22796 13320
rect 22376 13200 22428 13252
rect 26240 13268 26292 13320
rect 27436 13268 27488 13320
rect 27896 13268 27948 13320
rect 29736 13268 29788 13320
rect 33968 13311 34020 13320
rect 33968 13277 33977 13311
rect 33977 13277 34011 13311
rect 34011 13277 34020 13311
rect 33968 13268 34020 13277
rect 34060 13268 34112 13320
rect 35256 13336 35308 13388
rect 36360 13404 36412 13456
rect 35440 13268 35492 13320
rect 27068 13243 27120 13252
rect 27068 13209 27077 13243
rect 27077 13209 27111 13243
rect 27111 13209 27120 13243
rect 27068 13200 27120 13209
rect 27252 13200 27304 13252
rect 27528 13200 27580 13252
rect 32312 13243 32364 13252
rect 32312 13209 32321 13243
rect 32321 13209 32355 13243
rect 32355 13209 32364 13243
rect 32312 13200 32364 13209
rect 33324 13200 33376 13252
rect 34888 13200 34940 13252
rect 35808 13268 35860 13320
rect 36452 13268 36504 13320
rect 22836 13132 22888 13184
rect 28080 13132 28132 13184
rect 31852 13132 31904 13184
rect 32220 13132 32272 13184
rect 33784 13132 33836 13184
rect 34520 13175 34572 13184
rect 34520 13141 34529 13175
rect 34529 13141 34563 13175
rect 34563 13141 34572 13175
rect 34520 13132 34572 13141
rect 35992 13132 36044 13184
rect 36636 13175 36688 13184
rect 36636 13141 36645 13175
rect 36645 13141 36679 13175
rect 36679 13141 36688 13175
rect 36636 13132 36688 13141
rect 38844 13336 38896 13388
rect 37280 13311 37332 13320
rect 37280 13277 37289 13311
rect 37289 13277 37323 13311
rect 37323 13277 37332 13311
rect 37280 13268 37332 13277
rect 37188 13200 37240 13252
rect 37648 13311 37700 13320
rect 37648 13277 37657 13311
rect 37657 13277 37691 13311
rect 37691 13277 37700 13311
rect 37648 13268 37700 13277
rect 37832 13268 37884 13320
rect 38108 13268 38160 13320
rect 39028 13311 39080 13320
rect 39028 13277 39037 13311
rect 39037 13277 39071 13311
rect 39071 13277 39080 13311
rect 39028 13268 39080 13277
rect 39488 13336 39540 13388
rect 38660 13200 38712 13252
rect 38844 13200 38896 13252
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 7012 12928 7064 12980
rect 7196 12928 7248 12980
rect 8392 12928 8444 12980
rect 6460 12860 6512 12912
rect 9128 12928 9180 12980
rect 9864 12928 9916 12980
rect 10416 12971 10468 12980
rect 10416 12937 10425 12971
rect 10425 12937 10459 12971
rect 10459 12937 10468 12971
rect 10416 12928 10468 12937
rect 10508 12928 10560 12980
rect 12624 12928 12676 12980
rect 14004 12928 14056 12980
rect 17500 12928 17552 12980
rect 22284 12971 22336 12980
rect 22284 12937 22293 12971
rect 22293 12937 22327 12971
rect 22327 12937 22336 12971
rect 22284 12928 22336 12937
rect 24308 12971 24360 12980
rect 24308 12937 24317 12971
rect 24317 12937 24351 12971
rect 24351 12937 24360 12971
rect 24308 12928 24360 12937
rect 6368 12835 6420 12844
rect 6368 12801 6377 12835
rect 6377 12801 6411 12835
rect 6411 12801 6420 12835
rect 6368 12792 6420 12801
rect 6736 12835 6788 12844
rect 6736 12801 6745 12835
rect 6745 12801 6779 12835
rect 6779 12801 6788 12835
rect 6736 12792 6788 12801
rect 7196 12792 7248 12844
rect 7748 12792 7800 12844
rect 8300 12792 8352 12844
rect 8576 12835 8628 12844
rect 8576 12801 8593 12835
rect 8593 12801 8627 12835
rect 8627 12801 8628 12835
rect 8576 12792 8628 12801
rect 7104 12724 7156 12776
rect 9220 12860 9272 12912
rect 10784 12860 10836 12912
rect 9036 12835 9088 12844
rect 9036 12801 9045 12835
rect 9045 12801 9079 12835
rect 9079 12801 9088 12835
rect 9036 12792 9088 12801
rect 9680 12792 9732 12844
rect 10048 12835 10100 12844
rect 10048 12801 10057 12835
rect 10057 12801 10091 12835
rect 10091 12801 10100 12835
rect 10048 12792 10100 12801
rect 10232 12792 10284 12844
rect 4620 12656 4672 12708
rect 6736 12588 6788 12640
rect 7380 12699 7432 12708
rect 7380 12665 7389 12699
rect 7389 12665 7423 12699
rect 7423 12665 7432 12699
rect 7380 12656 7432 12665
rect 9864 12588 9916 12640
rect 10232 12588 10284 12640
rect 10508 12724 10560 12776
rect 10784 12724 10836 12776
rect 11796 12835 11848 12844
rect 11796 12801 11805 12835
rect 11805 12801 11839 12835
rect 11839 12801 11848 12835
rect 11796 12792 11848 12801
rect 12164 12792 12216 12844
rect 12348 12792 12400 12844
rect 14096 12792 14148 12844
rect 14188 12792 14240 12844
rect 14280 12835 14332 12844
rect 14280 12801 14289 12835
rect 14289 12801 14323 12835
rect 14323 12801 14332 12835
rect 14280 12792 14332 12801
rect 11336 12724 11388 12776
rect 11612 12699 11664 12708
rect 11612 12665 11621 12699
rect 11621 12665 11655 12699
rect 11655 12665 11664 12699
rect 11612 12656 11664 12665
rect 12072 12767 12124 12776
rect 12072 12733 12081 12767
rect 12081 12733 12115 12767
rect 12115 12733 12124 12767
rect 12072 12724 12124 12733
rect 14648 12792 14700 12844
rect 15016 12792 15068 12844
rect 15292 12903 15344 12912
rect 15292 12869 15301 12903
rect 15301 12869 15335 12903
rect 15335 12869 15344 12903
rect 15292 12860 15344 12869
rect 15568 12792 15620 12844
rect 15936 12835 15988 12844
rect 15936 12801 15971 12835
rect 15971 12801 15988 12835
rect 15936 12792 15988 12801
rect 16120 12835 16172 12844
rect 16120 12801 16129 12835
rect 16129 12801 16163 12835
rect 16163 12801 16172 12835
rect 16120 12792 16172 12801
rect 15108 12656 15160 12708
rect 15844 12724 15896 12776
rect 18788 12860 18840 12912
rect 17500 12792 17552 12844
rect 17316 12724 17368 12776
rect 17868 12835 17920 12844
rect 17868 12801 17877 12835
rect 17877 12801 17911 12835
rect 17911 12801 17920 12835
rect 17868 12792 17920 12801
rect 17960 12792 18012 12844
rect 18052 12792 18104 12844
rect 18604 12835 18656 12844
rect 18604 12801 18613 12835
rect 18613 12801 18647 12835
rect 18647 12801 18656 12835
rect 18604 12792 18656 12801
rect 18696 12835 18748 12844
rect 18696 12801 18705 12835
rect 18705 12801 18739 12835
rect 18739 12801 18748 12835
rect 18696 12792 18748 12801
rect 22468 12860 22520 12912
rect 23940 12903 23992 12912
rect 23940 12869 23949 12903
rect 23949 12869 23983 12903
rect 23983 12869 23992 12903
rect 23940 12860 23992 12869
rect 24032 12860 24084 12912
rect 24584 12903 24636 12912
rect 21364 12792 21416 12844
rect 22192 12792 22244 12844
rect 12992 12588 13044 12640
rect 14372 12588 14424 12640
rect 15292 12588 15344 12640
rect 19616 12724 19668 12776
rect 23480 12724 23532 12776
rect 18972 12656 19024 12708
rect 24584 12869 24593 12903
rect 24593 12869 24627 12903
rect 24627 12869 24636 12903
rect 24584 12860 24636 12869
rect 26608 12928 26660 12980
rect 27896 12860 27948 12912
rect 29736 12928 29788 12980
rect 30288 12928 30340 12980
rect 31760 12928 31812 12980
rect 32128 12928 32180 12980
rect 32588 12928 32640 12980
rect 32956 12928 33008 12980
rect 33048 12928 33100 12980
rect 30104 12860 30156 12912
rect 31668 12860 31720 12912
rect 32496 12860 32548 12912
rect 32680 12860 32732 12912
rect 24860 12792 24912 12844
rect 25136 12792 25188 12844
rect 25872 12724 25924 12776
rect 26240 12792 26292 12844
rect 27712 12792 27764 12844
rect 29092 12792 29144 12844
rect 29828 12835 29880 12844
rect 29828 12801 29834 12835
rect 29834 12801 29868 12835
rect 29868 12801 29880 12835
rect 29828 12792 29880 12801
rect 26700 12724 26752 12776
rect 27620 12724 27672 12776
rect 30104 12724 30156 12776
rect 31300 12724 31352 12776
rect 32864 12792 32916 12844
rect 32680 12724 32732 12776
rect 33140 12792 33192 12844
rect 19064 12588 19116 12640
rect 21916 12631 21968 12640
rect 21916 12597 21925 12631
rect 21925 12597 21959 12631
rect 21959 12597 21968 12631
rect 21916 12588 21968 12597
rect 23296 12588 23348 12640
rect 32956 12656 33008 12708
rect 33784 12835 33836 12844
rect 33784 12801 33793 12835
rect 33793 12801 33827 12835
rect 33827 12801 33836 12835
rect 33784 12792 33836 12801
rect 34060 12835 34112 12844
rect 34060 12801 34069 12835
rect 34069 12801 34103 12835
rect 34103 12801 34112 12835
rect 34060 12792 34112 12801
rect 34152 12835 34204 12844
rect 34152 12801 34161 12835
rect 34161 12801 34195 12835
rect 34195 12801 34204 12835
rect 34152 12792 34204 12801
rect 34152 12656 34204 12708
rect 23848 12588 23900 12640
rect 24124 12631 24176 12640
rect 24124 12597 24133 12631
rect 24133 12597 24167 12631
rect 24167 12597 24176 12631
rect 24124 12588 24176 12597
rect 24952 12631 25004 12640
rect 24952 12597 24961 12631
rect 24961 12597 24995 12631
rect 24995 12597 25004 12631
rect 24952 12588 25004 12597
rect 25412 12588 25464 12640
rect 32312 12588 32364 12640
rect 33876 12588 33928 12640
rect 34888 12971 34940 12980
rect 34888 12937 34897 12971
rect 34897 12937 34931 12971
rect 34931 12937 34940 12971
rect 34888 12928 34940 12937
rect 35624 12928 35676 12980
rect 35900 12928 35952 12980
rect 36176 12928 36228 12980
rect 38200 12928 38252 12980
rect 39856 12928 39908 12980
rect 38936 12860 38988 12912
rect 39120 12903 39172 12912
rect 39120 12869 39129 12903
rect 39129 12869 39163 12903
rect 39163 12869 39172 12903
rect 39120 12860 39172 12869
rect 36544 12835 36596 12844
rect 36544 12801 36553 12835
rect 36553 12801 36587 12835
rect 36587 12801 36596 12835
rect 36544 12792 36596 12801
rect 38844 12835 38896 12844
rect 38844 12801 38853 12835
rect 38853 12801 38887 12835
rect 38887 12801 38896 12835
rect 38844 12792 38896 12801
rect 34520 12767 34572 12776
rect 34520 12733 34529 12767
rect 34529 12733 34563 12767
rect 34563 12733 34572 12767
rect 34520 12724 34572 12733
rect 38660 12724 38712 12776
rect 39396 12792 39448 12844
rect 35256 12656 35308 12708
rect 38936 12656 38988 12708
rect 39488 12656 39540 12708
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 6460 12384 6512 12436
rect 8208 12384 8260 12436
rect 11060 12384 11112 12436
rect 4344 12180 4396 12232
rect 4896 12316 4948 12368
rect 7380 12316 7432 12368
rect 15108 12384 15160 12436
rect 15384 12384 15436 12436
rect 17224 12384 17276 12436
rect 18144 12384 18196 12436
rect 18972 12427 19024 12436
rect 18972 12393 18981 12427
rect 18981 12393 19015 12427
rect 19015 12393 19024 12427
rect 18972 12384 19024 12393
rect 19340 12384 19392 12436
rect 14740 12316 14792 12368
rect 14832 12316 14884 12368
rect 5264 12248 5316 12300
rect 6368 12248 6420 12300
rect 7288 12248 7340 12300
rect 4804 12223 4856 12232
rect 4804 12189 4813 12223
rect 4813 12189 4847 12223
rect 4847 12189 4856 12223
rect 4804 12180 4856 12189
rect 4896 12223 4948 12232
rect 4896 12189 4905 12223
rect 4905 12189 4939 12223
rect 4939 12189 4948 12223
rect 4896 12180 4948 12189
rect 4988 12223 5040 12232
rect 4988 12189 4997 12223
rect 4997 12189 5031 12223
rect 5031 12189 5040 12223
rect 4988 12180 5040 12189
rect 5356 12180 5408 12232
rect 3976 12044 4028 12096
rect 4344 12044 4396 12096
rect 5448 12044 5500 12096
rect 5632 12112 5684 12164
rect 5908 12223 5960 12232
rect 5908 12189 5917 12223
rect 5917 12189 5951 12223
rect 5951 12189 5960 12223
rect 5908 12180 5960 12189
rect 6644 12155 6696 12164
rect 6644 12121 6653 12155
rect 6653 12121 6687 12155
rect 6687 12121 6696 12155
rect 6644 12112 6696 12121
rect 7012 12112 7064 12164
rect 9036 12223 9088 12232
rect 9036 12189 9045 12223
rect 9045 12189 9079 12223
rect 9079 12189 9088 12223
rect 9036 12180 9088 12189
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 11152 12248 11204 12300
rect 16580 12248 16632 12300
rect 19616 12427 19668 12436
rect 19616 12393 19625 12427
rect 19625 12393 19659 12427
rect 19659 12393 19668 12427
rect 19616 12384 19668 12393
rect 20076 12384 20128 12436
rect 23480 12427 23532 12436
rect 23480 12393 23489 12427
rect 23489 12393 23523 12427
rect 23523 12393 23532 12427
rect 23480 12384 23532 12393
rect 10692 12223 10744 12232
rect 10692 12189 10701 12223
rect 10701 12189 10735 12223
rect 10735 12189 10744 12223
rect 10692 12180 10744 12189
rect 14280 12223 14332 12232
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 14464 12223 14516 12232
rect 14464 12189 14473 12223
rect 14473 12189 14507 12223
rect 14507 12189 14516 12223
rect 14464 12180 14516 12189
rect 15108 12223 15160 12232
rect 15108 12189 15117 12223
rect 15117 12189 15151 12223
rect 15151 12189 15160 12223
rect 15108 12180 15160 12189
rect 15752 12180 15804 12232
rect 17132 12180 17184 12232
rect 17316 12223 17368 12232
rect 17316 12189 17325 12223
rect 17325 12189 17359 12223
rect 17359 12189 17368 12223
rect 17316 12180 17368 12189
rect 17500 12223 17552 12232
rect 17500 12189 17509 12223
rect 17509 12189 17543 12223
rect 17543 12189 17552 12223
rect 17500 12180 17552 12189
rect 18788 12223 18840 12232
rect 18788 12189 18797 12223
rect 18797 12189 18831 12223
rect 18831 12189 18840 12223
rect 18788 12180 18840 12189
rect 11152 12112 11204 12164
rect 12716 12112 12768 12164
rect 13084 12112 13136 12164
rect 13728 12112 13780 12164
rect 5816 12044 5868 12096
rect 6368 12044 6420 12096
rect 7288 12087 7340 12096
rect 7288 12053 7297 12087
rect 7297 12053 7331 12087
rect 7331 12053 7340 12087
rect 7288 12044 7340 12053
rect 13820 12044 13872 12096
rect 14096 12112 14148 12164
rect 18604 12087 18656 12096
rect 18604 12053 18613 12087
rect 18613 12053 18647 12087
rect 18647 12053 18656 12087
rect 18604 12044 18656 12053
rect 19064 12223 19116 12232
rect 19064 12189 19073 12223
rect 19073 12189 19107 12223
rect 19107 12189 19116 12223
rect 19064 12180 19116 12189
rect 23940 12384 23992 12436
rect 24860 12384 24912 12436
rect 25596 12384 25648 12436
rect 25872 12427 25924 12436
rect 25872 12393 25881 12427
rect 25881 12393 25915 12427
rect 25915 12393 25924 12427
rect 25872 12384 25924 12393
rect 26056 12427 26108 12436
rect 26056 12393 26065 12427
rect 26065 12393 26099 12427
rect 26099 12393 26108 12427
rect 26056 12384 26108 12393
rect 26608 12427 26660 12436
rect 26608 12393 26617 12427
rect 26617 12393 26651 12427
rect 26651 12393 26660 12427
rect 26608 12384 26660 12393
rect 26884 12384 26936 12436
rect 21088 12248 21140 12300
rect 21364 12291 21416 12300
rect 21364 12257 21373 12291
rect 21373 12257 21407 12291
rect 21407 12257 21416 12291
rect 21364 12248 21416 12257
rect 21548 12291 21600 12300
rect 21548 12257 21557 12291
rect 21557 12257 21591 12291
rect 21591 12257 21600 12291
rect 21548 12248 21600 12257
rect 21916 12291 21968 12300
rect 21916 12257 21925 12291
rect 21925 12257 21959 12291
rect 21959 12257 21968 12291
rect 21916 12248 21968 12257
rect 23480 12248 23532 12300
rect 23848 12291 23900 12300
rect 23848 12257 23857 12291
rect 23857 12257 23891 12291
rect 23891 12257 23900 12291
rect 23848 12248 23900 12257
rect 24032 12248 24084 12300
rect 20260 12180 20312 12232
rect 23296 12180 23348 12232
rect 23664 12223 23716 12232
rect 23664 12189 23673 12223
rect 23673 12189 23707 12223
rect 23707 12189 23716 12223
rect 23664 12180 23716 12189
rect 24400 12180 24452 12232
rect 25596 12223 25648 12232
rect 25596 12189 25605 12223
rect 25605 12189 25639 12223
rect 25639 12189 25648 12223
rect 25596 12180 25648 12189
rect 26056 12248 26108 12300
rect 25872 12223 25924 12232
rect 25872 12189 25881 12223
rect 25881 12189 25915 12223
rect 25915 12189 25924 12223
rect 25872 12180 25924 12189
rect 19984 12044 20036 12096
rect 20904 12087 20956 12096
rect 20904 12053 20913 12087
rect 20913 12053 20947 12087
rect 20947 12053 20956 12087
rect 20904 12044 20956 12053
rect 21364 12044 21416 12096
rect 23112 12044 23164 12096
rect 25688 12112 25740 12164
rect 26056 12112 26108 12164
rect 26332 12223 26384 12232
rect 26332 12189 26341 12223
rect 26341 12189 26375 12223
rect 26375 12189 26384 12223
rect 26332 12180 26384 12189
rect 26608 12180 26660 12232
rect 26976 12223 27028 12232
rect 26976 12189 26985 12223
rect 26985 12189 27019 12223
rect 27019 12189 27028 12223
rect 26976 12180 27028 12189
rect 27068 12180 27120 12232
rect 28632 12248 28684 12300
rect 27528 12223 27580 12232
rect 27528 12189 27537 12223
rect 27537 12189 27571 12223
rect 27571 12189 27580 12223
rect 27528 12180 27580 12189
rect 27620 12223 27672 12232
rect 27620 12189 27629 12223
rect 27629 12189 27663 12223
rect 27663 12189 27672 12223
rect 27620 12180 27672 12189
rect 27712 12180 27764 12232
rect 28080 12180 28132 12232
rect 29368 12180 29420 12232
rect 29920 12180 29972 12232
rect 31576 12384 31628 12436
rect 31024 12359 31076 12368
rect 31024 12325 31033 12359
rect 31033 12325 31067 12359
rect 31067 12325 31076 12359
rect 31024 12316 31076 12325
rect 32312 12384 32364 12436
rect 33048 12384 33100 12436
rect 33508 12384 33560 12436
rect 37188 12384 37240 12436
rect 38108 12384 38160 12436
rect 30380 12291 30432 12300
rect 30380 12257 30389 12291
rect 30389 12257 30423 12291
rect 30423 12257 30432 12291
rect 30380 12248 30432 12257
rect 30472 12223 30524 12232
rect 24676 12044 24728 12096
rect 29736 12112 29788 12164
rect 26516 12044 26568 12096
rect 27068 12044 27120 12096
rect 27896 12044 27948 12096
rect 30472 12189 30481 12223
rect 30481 12189 30515 12223
rect 30515 12189 30524 12223
rect 30472 12180 30524 12189
rect 31576 12223 31628 12232
rect 31576 12189 31585 12223
rect 31585 12189 31619 12223
rect 31619 12189 31628 12223
rect 31576 12180 31628 12189
rect 32312 12291 32364 12300
rect 32312 12257 32321 12291
rect 32321 12257 32355 12291
rect 32355 12257 32364 12291
rect 32312 12248 32364 12257
rect 30288 12112 30340 12164
rect 31208 12112 31260 12164
rect 31392 12112 31444 12164
rect 32588 12180 32640 12232
rect 33140 12316 33192 12368
rect 39028 12316 39080 12368
rect 33692 12248 33744 12300
rect 35256 12248 35308 12300
rect 36452 12248 36504 12300
rect 37004 12248 37056 12300
rect 30380 12044 30432 12096
rect 30656 12087 30708 12096
rect 30656 12053 30665 12087
rect 30665 12053 30699 12087
rect 30699 12053 30708 12087
rect 30656 12044 30708 12053
rect 30932 12044 30984 12096
rect 32496 12112 32548 12164
rect 32772 12155 32824 12164
rect 32772 12121 32781 12155
rect 32781 12121 32815 12155
rect 32815 12121 32824 12155
rect 32772 12112 32824 12121
rect 33140 12155 33192 12164
rect 33140 12121 33149 12155
rect 33149 12121 33183 12155
rect 33183 12121 33192 12155
rect 33140 12112 33192 12121
rect 34060 12223 34112 12232
rect 34060 12189 34069 12223
rect 34069 12189 34103 12223
rect 34103 12189 34112 12223
rect 34060 12180 34112 12189
rect 34336 12180 34388 12232
rect 35808 12180 35860 12232
rect 36268 12180 36320 12232
rect 33600 12112 33652 12164
rect 37188 12112 37240 12164
rect 34520 12044 34572 12096
rect 36268 12044 36320 12096
rect 36820 12044 36872 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 3976 11840 4028 11892
rect 4804 11840 4856 11892
rect 5816 11883 5868 11892
rect 5816 11849 5825 11883
rect 5825 11849 5859 11883
rect 5859 11849 5868 11883
rect 5816 11840 5868 11849
rect 6736 11840 6788 11892
rect 7288 11840 7340 11892
rect 8116 11883 8168 11892
rect 8116 11849 8125 11883
rect 8125 11849 8159 11883
rect 8159 11849 8168 11883
rect 8116 11840 8168 11849
rect 9128 11840 9180 11892
rect 10232 11840 10284 11892
rect 11336 11840 11388 11892
rect 12716 11840 12768 11892
rect 18604 11840 18656 11892
rect 940 11704 992 11756
rect 1676 11679 1728 11688
rect 1676 11645 1685 11679
rect 1685 11645 1719 11679
rect 1719 11645 1728 11679
rect 1676 11636 1728 11645
rect 5632 11704 5684 11756
rect 4436 11636 4488 11688
rect 4804 11636 4856 11688
rect 6184 11704 6236 11756
rect 8300 11772 8352 11824
rect 8208 11747 8260 11756
rect 8208 11713 8217 11747
rect 8217 11713 8251 11747
rect 8251 11713 8260 11747
rect 8208 11704 8260 11713
rect 5356 11568 5408 11620
rect 5264 11500 5316 11552
rect 6828 11679 6880 11688
rect 6828 11645 6837 11679
rect 6837 11645 6871 11679
rect 6871 11645 6880 11679
rect 6828 11636 6880 11645
rect 7564 11636 7616 11688
rect 12532 11772 12584 11824
rect 14096 11772 14148 11824
rect 14740 11772 14792 11824
rect 20904 11840 20956 11892
rect 23664 11840 23716 11892
rect 19340 11772 19392 11824
rect 20168 11772 20220 11824
rect 10876 11747 10928 11756
rect 10876 11713 10885 11747
rect 10885 11713 10919 11747
rect 10919 11713 10928 11747
rect 10876 11704 10928 11713
rect 11060 11747 11112 11756
rect 11060 11713 11069 11747
rect 11069 11713 11103 11747
rect 11103 11713 11112 11747
rect 11060 11704 11112 11713
rect 13820 11704 13872 11756
rect 15108 11704 15160 11756
rect 16580 11704 16632 11756
rect 17408 11704 17460 11756
rect 25780 11840 25832 11892
rect 23756 11704 23808 11756
rect 25596 11772 25648 11824
rect 14832 11636 14884 11688
rect 5540 11568 5592 11620
rect 13728 11568 13780 11620
rect 15568 11568 15620 11620
rect 16304 11568 16356 11620
rect 16856 11568 16908 11620
rect 18328 11568 18380 11620
rect 10232 11500 10284 11552
rect 10324 11500 10376 11552
rect 16396 11500 16448 11552
rect 17500 11500 17552 11552
rect 21824 11568 21876 11620
rect 20260 11500 20312 11552
rect 23480 11636 23532 11688
rect 24952 11704 25004 11756
rect 24032 11568 24084 11620
rect 25964 11636 26016 11688
rect 26792 11840 26844 11892
rect 26884 11840 26936 11892
rect 30564 11840 30616 11892
rect 30656 11840 30708 11892
rect 31208 11840 31260 11892
rect 31300 11883 31352 11892
rect 31300 11849 31309 11883
rect 31309 11849 31343 11883
rect 31343 11849 31352 11883
rect 31300 11840 31352 11849
rect 31392 11840 31444 11892
rect 32312 11840 32364 11892
rect 26608 11772 26660 11824
rect 26424 11704 26476 11756
rect 26516 11636 26568 11688
rect 25872 11500 25924 11552
rect 29736 11772 29788 11824
rect 26700 11747 26752 11756
rect 26700 11713 26709 11747
rect 26709 11713 26743 11747
rect 26743 11713 26752 11747
rect 26700 11704 26752 11713
rect 27252 11747 27304 11756
rect 27252 11713 27261 11747
rect 27261 11713 27295 11747
rect 27295 11713 27304 11747
rect 27252 11704 27304 11713
rect 27344 11704 27396 11756
rect 29000 11747 29052 11756
rect 29000 11713 29009 11747
rect 29009 11713 29043 11747
rect 29043 11713 29052 11747
rect 29368 11747 29420 11756
rect 29000 11704 29052 11713
rect 29368 11713 29377 11747
rect 29377 11713 29411 11747
rect 29411 11713 29420 11747
rect 29368 11704 29420 11713
rect 26792 11636 26844 11688
rect 29276 11679 29328 11688
rect 29276 11645 29285 11679
rect 29285 11645 29319 11679
rect 29319 11645 29328 11679
rect 29276 11636 29328 11645
rect 30104 11704 30156 11756
rect 30288 11772 30340 11824
rect 30564 11704 30616 11756
rect 29920 11636 29972 11688
rect 30748 11704 30800 11756
rect 32036 11772 32088 11824
rect 34888 11772 34940 11824
rect 35072 11815 35124 11824
rect 35072 11781 35081 11815
rect 35081 11781 35115 11815
rect 35115 11781 35124 11815
rect 35072 11772 35124 11781
rect 35256 11772 35308 11824
rect 35992 11815 36044 11824
rect 35992 11781 36001 11815
rect 36001 11781 36035 11815
rect 36035 11781 36044 11815
rect 35992 11772 36044 11781
rect 33876 11704 33928 11756
rect 29736 11568 29788 11620
rect 31576 11636 31628 11688
rect 33784 11636 33836 11688
rect 34152 11636 34204 11688
rect 34428 11636 34480 11688
rect 35716 11747 35768 11756
rect 35716 11713 35726 11747
rect 35726 11713 35760 11747
rect 35760 11713 35768 11747
rect 35716 11704 35768 11713
rect 36084 11747 36136 11756
rect 36084 11713 36098 11747
rect 36098 11713 36132 11747
rect 36132 11713 36136 11747
rect 36084 11704 36136 11713
rect 36636 11840 36688 11892
rect 36820 11840 36872 11892
rect 37464 11840 37516 11892
rect 36636 11704 36688 11756
rect 39396 11772 39448 11824
rect 32404 11568 32456 11620
rect 33140 11568 33192 11620
rect 27160 11543 27212 11552
rect 27160 11509 27169 11543
rect 27169 11509 27203 11543
rect 27203 11509 27212 11543
rect 27160 11500 27212 11509
rect 27620 11500 27672 11552
rect 29368 11500 29420 11552
rect 30380 11500 30432 11552
rect 30656 11500 30708 11552
rect 34060 11500 34112 11552
rect 34520 11500 34572 11552
rect 37740 11636 37792 11688
rect 38844 11568 38896 11620
rect 39120 11636 39172 11688
rect 39672 11747 39724 11756
rect 39672 11713 39681 11747
rect 39681 11713 39715 11747
rect 39715 11713 39724 11747
rect 39672 11704 39724 11713
rect 41236 11840 41288 11892
rect 39856 11747 39908 11756
rect 39856 11713 39865 11747
rect 39865 11713 39899 11747
rect 39899 11713 39908 11747
rect 39856 11704 39908 11713
rect 40132 11747 40184 11756
rect 40132 11713 40141 11747
rect 40141 11713 40175 11747
rect 40175 11713 40184 11747
rect 40132 11704 40184 11713
rect 40040 11679 40092 11688
rect 40040 11645 40049 11679
rect 40049 11645 40083 11679
rect 40083 11645 40092 11679
rect 40040 11636 40092 11645
rect 36360 11500 36412 11552
rect 39212 11500 39264 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1676 11296 1728 11348
rect 4988 11296 5040 11348
rect 6184 11339 6236 11348
rect 6184 11305 6193 11339
rect 6193 11305 6227 11339
rect 6227 11305 6236 11339
rect 6184 11296 6236 11305
rect 6368 11339 6420 11348
rect 6368 11305 6377 11339
rect 6377 11305 6411 11339
rect 6411 11305 6420 11339
rect 6368 11296 6420 11305
rect 7656 11296 7708 11348
rect 8116 11296 8168 11348
rect 8300 11296 8352 11348
rect 12256 11296 12308 11348
rect 7932 11228 7984 11280
rect 6460 11135 6512 11144
rect 6460 11101 6469 11135
rect 6469 11101 6503 11135
rect 6503 11101 6512 11135
rect 6460 11092 6512 11101
rect 5264 10956 5316 11008
rect 7104 10956 7156 11008
rect 7196 10956 7248 11008
rect 10140 11160 10192 11212
rect 10692 11160 10744 11212
rect 10968 11203 11020 11212
rect 10968 11169 10977 11203
rect 10977 11169 11011 11203
rect 11011 11169 11020 11203
rect 10968 11160 11020 11169
rect 12900 11228 12952 11280
rect 7656 11024 7708 11076
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 8576 11092 8628 11144
rect 9956 11092 10008 11144
rect 10324 11092 10376 11144
rect 12164 11160 12216 11212
rect 12256 11203 12308 11212
rect 12256 11169 12265 11203
rect 12265 11169 12299 11203
rect 12299 11169 12308 11203
rect 12256 11160 12308 11169
rect 14556 11296 14608 11348
rect 12440 11135 12492 11144
rect 12440 11101 12449 11135
rect 12449 11101 12483 11135
rect 12483 11101 12492 11135
rect 12440 11092 12492 11101
rect 12532 11092 12584 11144
rect 15568 11160 15620 11212
rect 15936 11296 15988 11348
rect 16120 11296 16172 11348
rect 21364 11339 21416 11348
rect 21364 11305 21373 11339
rect 21373 11305 21407 11339
rect 21407 11305 21416 11339
rect 21364 11296 21416 11305
rect 26056 11296 26108 11348
rect 26792 11296 26844 11348
rect 27528 11296 27580 11348
rect 22100 11228 22152 11280
rect 8116 10956 8168 11008
rect 11612 11067 11664 11076
rect 11612 11033 11621 11067
rect 11621 11033 11655 11067
rect 11655 11033 11664 11067
rect 11612 11024 11664 11033
rect 11888 11024 11940 11076
rect 16304 11092 16356 11144
rect 17408 11160 17460 11212
rect 17500 11203 17552 11212
rect 17500 11169 17509 11203
rect 17509 11169 17543 11203
rect 17543 11169 17552 11203
rect 17500 11160 17552 11169
rect 17776 11160 17828 11212
rect 18604 11160 18656 11212
rect 20260 11160 20312 11212
rect 29000 11228 29052 11280
rect 30840 11271 30892 11280
rect 30840 11237 30849 11271
rect 30849 11237 30883 11271
rect 30883 11237 30892 11271
rect 30840 11228 30892 11237
rect 31024 11339 31076 11348
rect 31024 11305 31033 11339
rect 31033 11305 31067 11339
rect 31067 11305 31076 11339
rect 31024 11296 31076 11305
rect 36084 11296 36136 11348
rect 36176 11296 36228 11348
rect 38660 11296 38712 11348
rect 39120 11296 39172 11348
rect 39304 11339 39356 11348
rect 39304 11305 39313 11339
rect 39313 11305 39347 11339
rect 39347 11305 39356 11339
rect 39304 11296 39356 11305
rect 33508 11228 33560 11280
rect 25872 11160 25924 11212
rect 22376 11092 22428 11144
rect 22652 11135 22704 11144
rect 22652 11101 22661 11135
rect 22661 11101 22695 11135
rect 22695 11101 22704 11135
rect 22652 11092 22704 11101
rect 23112 11135 23164 11144
rect 23112 11101 23121 11135
rect 23121 11101 23155 11135
rect 23155 11101 23164 11135
rect 23112 11092 23164 11101
rect 9864 10956 9916 11008
rect 10416 10999 10468 11008
rect 10416 10965 10425 10999
rect 10425 10965 10459 10999
rect 10459 10965 10468 10999
rect 10416 10956 10468 10965
rect 11244 10999 11296 11008
rect 11244 10965 11253 10999
rect 11253 10965 11287 10999
rect 11287 10965 11296 10999
rect 11244 10956 11296 10965
rect 12624 10999 12676 11008
rect 12624 10965 12633 10999
rect 12633 10965 12667 10999
rect 12667 10965 12676 10999
rect 12624 10956 12676 10965
rect 17132 11024 17184 11076
rect 22468 11024 22520 11076
rect 13820 10956 13872 11008
rect 16304 10999 16356 11008
rect 16304 10965 16313 10999
rect 16313 10965 16347 10999
rect 16347 10965 16356 10999
rect 16304 10956 16356 10965
rect 17040 10999 17092 11008
rect 17040 10965 17049 10999
rect 17049 10965 17083 10999
rect 17083 10965 17092 10999
rect 17040 10956 17092 10965
rect 17316 10956 17368 11008
rect 21456 10956 21508 11008
rect 25964 11024 26016 11076
rect 26700 11024 26752 11076
rect 27160 11024 27212 11076
rect 31484 11092 31536 11144
rect 32956 11203 33008 11212
rect 32956 11169 32965 11203
rect 32965 11169 32999 11203
rect 32999 11169 33008 11203
rect 32956 11160 33008 11169
rect 36360 11271 36412 11280
rect 36360 11237 36369 11271
rect 36369 11237 36403 11271
rect 36403 11237 36412 11271
rect 36360 11228 36412 11237
rect 36636 11228 36688 11280
rect 37648 11228 37700 11280
rect 30196 11024 30248 11076
rect 30564 11067 30616 11076
rect 30564 11033 30573 11067
rect 30573 11033 30607 11067
rect 30607 11033 30616 11067
rect 30564 11024 30616 11033
rect 31668 11024 31720 11076
rect 32036 11092 32088 11144
rect 33600 11135 33652 11144
rect 33600 11101 33609 11135
rect 33609 11101 33643 11135
rect 33643 11101 33652 11135
rect 33600 11092 33652 11101
rect 33876 11160 33928 11212
rect 35440 11160 35492 11212
rect 25136 10956 25188 11008
rect 29184 10956 29236 11008
rect 29552 10956 29604 11008
rect 31208 10956 31260 11008
rect 32956 10956 33008 11008
rect 33140 10956 33192 11008
rect 33324 11067 33376 11076
rect 33324 11033 33333 11067
rect 33333 11033 33367 11067
rect 33367 11033 33376 11067
rect 33324 11024 33376 11033
rect 34060 11092 34112 11144
rect 35164 11092 35216 11144
rect 36084 11135 36136 11144
rect 36084 11101 36093 11135
rect 36093 11101 36127 11135
rect 36127 11101 36136 11135
rect 36084 11092 36136 11101
rect 36176 11135 36228 11144
rect 36176 11101 36185 11135
rect 36185 11101 36219 11135
rect 36219 11101 36228 11135
rect 36176 11092 36228 11101
rect 36360 11092 36412 11144
rect 36820 11092 36872 11144
rect 35992 11067 36044 11076
rect 35992 11033 36001 11067
rect 36001 11033 36035 11067
rect 36035 11033 36044 11067
rect 35992 11024 36044 11033
rect 37188 11024 37240 11076
rect 37556 11092 37608 11144
rect 38384 11092 38436 11144
rect 38752 11135 38804 11144
rect 38752 11101 38762 11135
rect 38762 11101 38796 11135
rect 38796 11101 38804 11135
rect 38752 11092 38804 11101
rect 39948 11228 40000 11280
rect 39120 11135 39172 11144
rect 39120 11101 39134 11135
rect 39134 11101 39168 11135
rect 39168 11101 39172 11135
rect 39120 11092 39172 11101
rect 36636 10956 36688 11008
rect 36820 10999 36872 11008
rect 36820 10965 36829 10999
rect 36829 10965 36863 10999
rect 36863 10965 36872 10999
rect 36820 10956 36872 10965
rect 37096 10956 37148 11008
rect 39028 10956 39080 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 6460 10795 6512 10804
rect 6460 10761 6469 10795
rect 6469 10761 6503 10795
rect 6503 10761 6512 10795
rect 6460 10752 6512 10761
rect 7104 10795 7156 10804
rect 7104 10761 7113 10795
rect 7113 10761 7147 10795
rect 7147 10761 7156 10795
rect 7104 10752 7156 10761
rect 7932 10752 7984 10804
rect 11244 10752 11296 10804
rect 11980 10795 12032 10804
rect 11980 10761 11989 10795
rect 11989 10761 12023 10795
rect 12023 10761 12032 10795
rect 11980 10752 12032 10761
rect 12164 10752 12216 10804
rect 16488 10752 16540 10804
rect 17960 10752 18012 10804
rect 19340 10752 19392 10804
rect 20904 10752 20956 10804
rect 6920 10659 6972 10668
rect 6920 10625 6929 10659
rect 6929 10625 6963 10659
rect 6963 10625 6972 10659
rect 6920 10616 6972 10625
rect 7196 10659 7248 10668
rect 7196 10625 7205 10659
rect 7205 10625 7239 10659
rect 7239 10625 7248 10659
rect 7196 10616 7248 10625
rect 8484 10616 8536 10668
rect 10876 10684 10928 10736
rect 8668 10616 8720 10668
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 8208 10548 8260 10600
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 9404 10616 9456 10668
rect 9496 10659 9548 10668
rect 9496 10625 9505 10659
rect 9505 10625 9539 10659
rect 9539 10625 9548 10659
rect 9496 10616 9548 10625
rect 9956 10659 10008 10668
rect 9956 10625 9965 10659
rect 9965 10625 9999 10659
rect 9999 10625 10008 10659
rect 9956 10616 10008 10625
rect 10140 10616 10192 10668
rect 10324 10548 10376 10600
rect 16856 10684 16908 10736
rect 17040 10684 17092 10736
rect 17684 10727 17736 10736
rect 17684 10693 17693 10727
rect 17693 10693 17727 10727
rect 17727 10693 17736 10727
rect 17684 10684 17736 10693
rect 18972 10684 19024 10736
rect 19064 10684 19116 10736
rect 20720 10684 20772 10736
rect 10416 10480 10468 10532
rect 12624 10548 12676 10600
rect 12992 10659 13044 10668
rect 12992 10625 13001 10659
rect 13001 10625 13035 10659
rect 13035 10625 13044 10659
rect 12992 10616 13044 10625
rect 17408 10659 17460 10668
rect 17408 10625 17417 10659
rect 17417 10625 17451 10659
rect 17451 10625 17460 10659
rect 17408 10616 17460 10625
rect 18696 10616 18748 10668
rect 19984 10616 20036 10668
rect 26240 10616 26292 10668
rect 26700 10616 26752 10668
rect 19156 10591 19208 10600
rect 15660 10480 15712 10532
rect 19156 10557 19165 10591
rect 19165 10557 19199 10591
rect 19199 10557 19208 10591
rect 19156 10548 19208 10557
rect 19340 10591 19392 10600
rect 19340 10557 19349 10591
rect 19349 10557 19383 10591
rect 19383 10557 19392 10591
rect 19340 10548 19392 10557
rect 20260 10548 20312 10600
rect 23572 10548 23624 10600
rect 21456 10480 21508 10532
rect 4804 10412 4856 10464
rect 5356 10412 5408 10464
rect 8392 10455 8444 10464
rect 8392 10421 8401 10455
rect 8401 10421 8435 10455
rect 8435 10421 8444 10455
rect 8392 10412 8444 10421
rect 10232 10412 10284 10464
rect 12900 10455 12952 10464
rect 12900 10421 12909 10455
rect 12909 10421 12943 10455
rect 12943 10421 12952 10455
rect 12900 10412 12952 10421
rect 16120 10412 16172 10464
rect 19984 10455 20036 10464
rect 19984 10421 19993 10455
rect 19993 10421 20027 10455
rect 20027 10421 20036 10455
rect 19984 10412 20036 10421
rect 21640 10412 21692 10464
rect 23756 10412 23808 10464
rect 23848 10455 23900 10464
rect 23848 10421 23857 10455
rect 23857 10421 23891 10455
rect 23891 10421 23900 10455
rect 23848 10412 23900 10421
rect 25136 10412 25188 10464
rect 26424 10412 26476 10464
rect 30472 10752 30524 10804
rect 31760 10795 31812 10804
rect 31760 10761 31769 10795
rect 31769 10761 31803 10795
rect 31803 10761 31812 10795
rect 31760 10752 31812 10761
rect 27436 10659 27488 10668
rect 27436 10625 27445 10659
rect 27445 10625 27479 10659
rect 27479 10625 27488 10659
rect 27436 10616 27488 10625
rect 28724 10616 28776 10668
rect 32404 10684 32456 10736
rect 32772 10727 32824 10736
rect 32772 10693 32797 10727
rect 32797 10693 32824 10727
rect 33048 10752 33100 10804
rect 34428 10752 34480 10804
rect 40960 10752 41012 10804
rect 32772 10684 32824 10693
rect 35900 10684 35952 10736
rect 29184 10616 29236 10668
rect 29552 10659 29604 10668
rect 29552 10625 29561 10659
rect 29561 10625 29595 10659
rect 29595 10625 29604 10659
rect 29552 10616 29604 10625
rect 29644 10616 29696 10668
rect 30104 10616 30156 10668
rect 30196 10659 30248 10668
rect 30196 10625 30205 10659
rect 30205 10625 30239 10659
rect 30239 10625 30248 10659
rect 30196 10616 30248 10625
rect 30840 10616 30892 10668
rect 31484 10616 31536 10668
rect 31208 10548 31260 10600
rect 32036 10616 32088 10668
rect 32956 10616 33008 10668
rect 33508 10616 33560 10668
rect 33784 10659 33836 10668
rect 33784 10625 33793 10659
rect 33793 10625 33827 10659
rect 33827 10625 33836 10659
rect 33784 10616 33836 10625
rect 36084 10616 36136 10668
rect 37648 10659 37700 10668
rect 37648 10625 37657 10659
rect 37657 10625 37691 10659
rect 37691 10625 37700 10659
rect 37648 10616 37700 10625
rect 31024 10480 31076 10532
rect 34060 10548 34112 10600
rect 35440 10548 35492 10600
rect 36360 10548 36412 10600
rect 37556 10548 37608 10600
rect 32128 10480 32180 10532
rect 28448 10412 28500 10464
rect 29552 10412 29604 10464
rect 29920 10412 29972 10464
rect 30564 10412 30616 10464
rect 32680 10412 32732 10464
rect 37832 10455 37884 10464
rect 37832 10421 37841 10455
rect 37841 10421 37875 10455
rect 37875 10421 37884 10455
rect 37832 10412 37884 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 4804 10208 4856 10260
rect 8392 10208 8444 10260
rect 8484 10208 8536 10260
rect 11428 10208 11480 10260
rect 17500 10208 17552 10260
rect 19340 10208 19392 10260
rect 20444 10251 20496 10260
rect 20444 10217 20453 10251
rect 20453 10217 20487 10251
rect 20487 10217 20496 10251
rect 20444 10208 20496 10217
rect 20812 10208 20864 10260
rect 21456 10251 21508 10260
rect 21456 10217 21465 10251
rect 21465 10217 21499 10251
rect 21499 10217 21508 10251
rect 21456 10208 21508 10217
rect 22192 10208 22244 10260
rect 22376 10251 22428 10260
rect 22376 10217 22385 10251
rect 22385 10217 22419 10251
rect 22419 10217 22428 10251
rect 22376 10208 22428 10217
rect 22560 10208 22612 10260
rect 23848 10208 23900 10260
rect 24492 10208 24544 10260
rect 26240 10208 26292 10260
rect 26516 10208 26568 10260
rect 26976 10208 27028 10260
rect 27436 10208 27488 10260
rect 28724 10208 28776 10260
rect 30196 10208 30248 10260
rect 31484 10208 31536 10260
rect 32680 10208 32732 10260
rect 37832 10208 37884 10260
rect 39856 10208 39908 10260
rect 7748 10140 7800 10192
rect 6000 10072 6052 10124
rect 8760 10140 8812 10192
rect 13636 10140 13688 10192
rect 16028 10183 16080 10192
rect 16028 10149 16037 10183
rect 16037 10149 16071 10183
rect 16071 10149 16080 10183
rect 16028 10140 16080 10149
rect 22100 10183 22152 10192
rect 22100 10149 22109 10183
rect 22109 10149 22143 10183
rect 22143 10149 22152 10183
rect 22100 10140 22152 10149
rect 4896 9979 4948 9988
rect 4896 9945 4926 9979
rect 4926 9945 4948 9979
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 9312 10072 9364 10124
rect 8852 10004 8904 10056
rect 9772 10072 9824 10124
rect 10232 10072 10284 10124
rect 4896 9936 4948 9945
rect 5264 9936 5316 9988
rect 5356 9979 5408 9988
rect 5356 9945 5365 9979
rect 5365 9945 5399 9979
rect 5399 9945 5408 9979
rect 5356 9936 5408 9945
rect 9864 10004 9916 10056
rect 12624 10004 12676 10056
rect 14188 10004 14240 10056
rect 13820 9936 13872 9988
rect 15936 9936 15988 9988
rect 5724 9868 5776 9920
rect 9588 9911 9640 9920
rect 9588 9877 9597 9911
rect 9597 9877 9631 9911
rect 9631 9877 9640 9911
rect 9588 9868 9640 9877
rect 9864 9868 9916 9920
rect 12164 9911 12216 9920
rect 12164 9877 12173 9911
rect 12173 9877 12207 9911
rect 12207 9877 12216 9911
rect 12164 9868 12216 9877
rect 13912 9911 13964 9920
rect 13912 9877 13921 9911
rect 13921 9877 13955 9911
rect 13955 9877 13964 9911
rect 13912 9868 13964 9877
rect 14004 9868 14056 9920
rect 15844 9868 15896 9920
rect 16304 10072 16356 10124
rect 16120 10047 16172 10056
rect 16120 10013 16129 10047
rect 16129 10013 16163 10047
rect 16163 10013 16172 10047
rect 16120 10004 16172 10013
rect 16856 10072 16908 10124
rect 20168 10072 20220 10124
rect 19156 10004 19208 10056
rect 20996 10072 21048 10124
rect 21180 10004 21232 10056
rect 21640 10004 21692 10056
rect 22008 10004 22060 10056
rect 23388 10183 23440 10192
rect 23388 10149 23397 10183
rect 23397 10149 23431 10183
rect 23431 10149 23440 10183
rect 23388 10140 23440 10149
rect 25228 10072 25280 10124
rect 27068 10115 27120 10124
rect 27068 10081 27077 10115
rect 27077 10081 27111 10115
rect 27111 10081 27120 10115
rect 27068 10072 27120 10081
rect 28540 10072 28592 10124
rect 29276 10072 29328 10124
rect 31852 10140 31904 10192
rect 32496 10140 32548 10192
rect 22560 10047 22612 10056
rect 22560 10013 22569 10047
rect 22569 10013 22603 10047
rect 22603 10013 22612 10047
rect 22560 10004 22612 10013
rect 23112 10004 23164 10056
rect 23572 10047 23624 10056
rect 23572 10013 23581 10047
rect 23581 10013 23615 10047
rect 23615 10013 23624 10047
rect 23572 10004 23624 10013
rect 20904 9936 20956 9988
rect 21272 9936 21324 9988
rect 26792 10047 26844 10056
rect 26792 10013 26801 10047
rect 26801 10013 26835 10047
rect 26835 10013 26844 10047
rect 26792 10004 26844 10013
rect 27620 10004 27672 10056
rect 24952 9936 25004 9988
rect 25136 9936 25188 9988
rect 29736 10004 29788 10056
rect 30472 10072 30524 10124
rect 31024 10072 31076 10124
rect 32404 10072 32456 10124
rect 31300 10004 31352 10056
rect 31576 10047 31628 10056
rect 31576 10013 31585 10047
rect 31585 10013 31619 10047
rect 31619 10013 31628 10047
rect 31576 10004 31628 10013
rect 16948 9868 17000 9920
rect 24124 9868 24176 9920
rect 26424 9911 26476 9920
rect 26424 9877 26433 9911
rect 26433 9877 26467 9911
rect 26467 9877 26476 9911
rect 26424 9868 26476 9877
rect 27068 9868 27120 9920
rect 27988 9868 28040 9920
rect 28080 9868 28132 9920
rect 32128 10004 32180 10056
rect 38200 10115 38252 10124
rect 38200 10081 38209 10115
rect 38209 10081 38243 10115
rect 38243 10081 38252 10115
rect 38200 10072 38252 10081
rect 33508 10047 33560 10056
rect 33508 10013 33517 10047
rect 33517 10013 33551 10047
rect 33551 10013 33560 10047
rect 33508 10004 33560 10013
rect 38108 10047 38160 10056
rect 38108 10013 38117 10047
rect 38117 10013 38151 10047
rect 38151 10013 38160 10047
rect 38108 10004 38160 10013
rect 38384 10047 38436 10056
rect 38384 10013 38393 10047
rect 38393 10013 38427 10047
rect 38427 10013 38436 10047
rect 38384 10004 38436 10013
rect 28448 9868 28500 9920
rect 29000 9868 29052 9920
rect 30288 9868 30340 9920
rect 31852 9868 31904 9920
rect 32036 9868 32088 9920
rect 32312 9868 32364 9920
rect 33140 9868 33192 9920
rect 33692 9911 33744 9920
rect 33692 9877 33701 9911
rect 33701 9877 33735 9911
rect 33735 9877 33744 9911
rect 33692 9868 33744 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 8668 9664 8720 9716
rect 9404 9664 9456 9716
rect 5080 9528 5132 9580
rect 5448 9528 5500 9580
rect 5724 9528 5776 9580
rect 6000 9571 6052 9580
rect 6000 9537 6009 9571
rect 6009 9537 6043 9571
rect 6043 9537 6052 9571
rect 6000 9528 6052 9537
rect 7656 9596 7708 9648
rect 7840 9596 7892 9648
rect 8944 9596 8996 9648
rect 6552 9571 6604 9580
rect 6552 9537 6561 9571
rect 6561 9537 6595 9571
rect 6595 9537 6604 9571
rect 6552 9528 6604 9537
rect 6920 9528 6972 9580
rect 7564 9571 7616 9580
rect 7564 9537 7573 9571
rect 7573 9537 7607 9571
rect 7607 9537 7616 9571
rect 7564 9528 7616 9537
rect 7748 9571 7800 9580
rect 7748 9537 7757 9571
rect 7757 9537 7791 9571
rect 7791 9537 7800 9571
rect 7748 9528 7800 9537
rect 9128 9596 9180 9648
rect 9588 9596 9640 9648
rect 9772 9596 9824 9648
rect 9864 9639 9916 9648
rect 9864 9605 9873 9639
rect 9873 9605 9907 9639
rect 9907 9605 9916 9639
rect 9864 9596 9916 9605
rect 9496 9528 9548 9580
rect 9956 9528 10008 9580
rect 5264 9392 5316 9444
rect 7564 9392 7616 9444
rect 7932 9392 7984 9444
rect 12900 9664 12952 9716
rect 11888 9596 11940 9648
rect 11060 9460 11112 9512
rect 11244 9460 11296 9512
rect 11336 9460 11388 9512
rect 12532 9528 12584 9580
rect 12716 9571 12768 9580
rect 12716 9537 12725 9571
rect 12725 9537 12759 9571
rect 12759 9537 12768 9571
rect 12716 9528 12768 9537
rect 13820 9571 13872 9580
rect 13820 9537 13829 9571
rect 13829 9537 13863 9571
rect 13863 9537 13872 9571
rect 13820 9528 13872 9537
rect 13912 9528 13964 9580
rect 14188 9528 14240 9580
rect 16120 9664 16172 9716
rect 20720 9664 20772 9716
rect 15844 9528 15896 9580
rect 19432 9596 19484 9648
rect 19800 9596 19852 9648
rect 19984 9596 20036 9648
rect 16120 9571 16172 9580
rect 16120 9537 16129 9571
rect 16129 9537 16163 9571
rect 16163 9537 16172 9571
rect 16120 9528 16172 9537
rect 9588 9435 9640 9444
rect 9588 9401 9597 9435
rect 9597 9401 9631 9435
rect 9631 9401 9640 9435
rect 9588 9392 9640 9401
rect 9864 9392 9916 9444
rect 6184 9367 6236 9376
rect 6184 9333 6193 9367
rect 6193 9333 6227 9367
rect 6227 9333 6236 9367
rect 6184 9324 6236 9333
rect 8024 9324 8076 9376
rect 9220 9324 9272 9376
rect 11428 9324 11480 9376
rect 12164 9324 12216 9376
rect 12256 9367 12308 9376
rect 12256 9333 12265 9367
rect 12265 9333 12299 9367
rect 12299 9333 12308 9367
rect 12256 9324 12308 9333
rect 13176 9367 13228 9376
rect 13176 9333 13185 9367
rect 13185 9333 13219 9367
rect 13219 9333 13228 9367
rect 13176 9324 13228 9333
rect 16580 9460 16632 9512
rect 16856 9571 16908 9580
rect 16856 9537 16865 9571
rect 16865 9537 16899 9571
rect 16899 9537 16908 9571
rect 16856 9528 16908 9537
rect 16948 9571 17000 9580
rect 16948 9537 16957 9571
rect 16957 9537 16991 9571
rect 16991 9537 17000 9571
rect 16948 9528 17000 9537
rect 17132 9571 17184 9580
rect 17132 9537 17141 9571
rect 17141 9537 17175 9571
rect 17175 9537 17184 9571
rect 17132 9528 17184 9537
rect 13728 9392 13780 9444
rect 16948 9392 17000 9444
rect 15200 9324 15252 9376
rect 16396 9324 16448 9376
rect 16488 9324 16540 9376
rect 19156 9571 19208 9580
rect 19156 9537 19165 9571
rect 19165 9537 19199 9571
rect 19199 9537 19208 9571
rect 19156 9528 19208 9537
rect 21180 9596 21232 9648
rect 23112 9664 23164 9716
rect 24860 9664 24912 9716
rect 25136 9664 25188 9716
rect 25964 9707 26016 9716
rect 25964 9673 25973 9707
rect 25973 9673 26007 9707
rect 26007 9673 26016 9707
rect 25964 9664 26016 9673
rect 22008 9571 22060 9580
rect 22008 9537 22017 9571
rect 22017 9537 22051 9571
rect 22051 9537 22060 9571
rect 22008 9528 22060 9537
rect 22192 9571 22244 9580
rect 22192 9537 22201 9571
rect 22201 9537 22235 9571
rect 22235 9537 22244 9571
rect 22192 9528 22244 9537
rect 21824 9460 21876 9512
rect 19432 9324 19484 9376
rect 19708 9324 19760 9376
rect 22560 9460 22612 9512
rect 24124 9460 24176 9512
rect 24216 9503 24268 9512
rect 24216 9469 24225 9503
rect 24225 9469 24259 9503
rect 24259 9469 24268 9503
rect 24216 9460 24268 9469
rect 24492 9503 24544 9512
rect 24492 9469 24501 9503
rect 24501 9469 24535 9503
rect 24535 9469 24544 9503
rect 24492 9460 24544 9469
rect 24952 9460 25004 9512
rect 26056 9571 26108 9580
rect 26056 9537 26065 9571
rect 26065 9537 26099 9571
rect 26099 9537 26108 9571
rect 26056 9528 26108 9537
rect 26332 9639 26384 9648
rect 26332 9605 26341 9639
rect 26341 9605 26375 9639
rect 26375 9605 26384 9639
rect 26332 9596 26384 9605
rect 31484 9664 31536 9716
rect 33140 9664 33192 9716
rect 33600 9664 33652 9716
rect 30380 9596 30432 9648
rect 31576 9596 31628 9648
rect 27160 9528 27212 9580
rect 27252 9571 27304 9580
rect 27252 9537 27261 9571
rect 27261 9537 27295 9571
rect 27295 9537 27304 9571
rect 27252 9528 27304 9537
rect 30104 9528 30156 9580
rect 27528 9460 27580 9512
rect 27344 9392 27396 9444
rect 28356 9460 28408 9512
rect 29644 9460 29696 9512
rect 31852 9528 31904 9580
rect 33508 9596 33560 9648
rect 33968 9639 34020 9648
rect 33968 9605 33977 9639
rect 33977 9605 34011 9639
rect 34011 9605 34020 9639
rect 33968 9596 34020 9605
rect 31392 9460 31444 9512
rect 27620 9367 27672 9376
rect 27620 9333 27629 9367
rect 27629 9333 27663 9367
rect 27663 9333 27672 9367
rect 27620 9324 27672 9333
rect 27896 9324 27948 9376
rect 32036 9324 32088 9376
rect 33416 9528 33468 9580
rect 32772 9460 32824 9512
rect 33876 9571 33928 9580
rect 33876 9537 33885 9571
rect 33885 9537 33919 9571
rect 33919 9537 33928 9571
rect 33876 9528 33928 9537
rect 34244 9596 34296 9648
rect 34520 9596 34572 9648
rect 34428 9571 34480 9580
rect 34428 9537 34437 9571
rect 34437 9537 34471 9571
rect 34471 9537 34480 9571
rect 34428 9528 34480 9537
rect 35716 9596 35768 9648
rect 38936 9596 38988 9648
rect 39580 9596 39632 9648
rect 32312 9392 32364 9444
rect 33508 9392 33560 9444
rect 33968 9392 34020 9444
rect 34244 9435 34296 9444
rect 34244 9401 34253 9435
rect 34253 9401 34287 9435
rect 34287 9401 34296 9435
rect 34244 9392 34296 9401
rect 35256 9503 35308 9512
rect 35256 9469 35265 9503
rect 35265 9469 35299 9503
rect 35299 9469 35308 9503
rect 35256 9460 35308 9469
rect 35348 9460 35400 9512
rect 34612 9392 34664 9444
rect 34796 9324 34848 9376
rect 35992 9324 36044 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 6184 9120 6236 9172
rect 6552 9163 6604 9172
rect 6552 9129 6561 9163
rect 6561 9129 6595 9163
rect 6595 9129 6604 9163
rect 6552 9120 6604 9129
rect 6920 9120 6972 9172
rect 7656 9120 7708 9172
rect 8024 9163 8076 9172
rect 8024 9129 8033 9163
rect 8033 9129 8067 9163
rect 8067 9129 8076 9163
rect 8024 9120 8076 9129
rect 5448 9052 5500 9104
rect 7196 9052 7248 9104
rect 9588 9120 9640 9172
rect 11612 9120 11664 9172
rect 12256 9120 12308 9172
rect 13176 9120 13228 9172
rect 13820 9120 13872 9172
rect 16488 9120 16540 9172
rect 16580 9120 16632 9172
rect 16856 9120 16908 9172
rect 19156 9120 19208 9172
rect 20812 9163 20864 9172
rect 20812 9129 20821 9163
rect 20821 9129 20855 9163
rect 20855 9129 20864 9163
rect 20812 9120 20864 9129
rect 21824 9120 21876 9172
rect 24492 9120 24544 9172
rect 4068 8916 4120 8968
rect 6644 8984 6696 9036
rect 7104 8916 7156 8968
rect 6552 8848 6604 8900
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 11520 9095 11572 9104
rect 11520 9061 11529 9095
rect 11529 9061 11563 9095
rect 11563 9061 11572 9095
rect 11520 9052 11572 9061
rect 11244 9027 11296 9036
rect 11244 8993 11253 9027
rect 11253 8993 11287 9027
rect 11287 8993 11296 9027
rect 11244 8984 11296 8993
rect 13544 9052 13596 9104
rect 15200 9052 15252 9104
rect 16120 9052 16172 9104
rect 7104 8780 7156 8832
rect 7656 8780 7708 8832
rect 8024 8848 8076 8900
rect 9312 8959 9364 8968
rect 9312 8925 9321 8959
rect 9321 8925 9355 8959
rect 9355 8925 9364 8959
rect 9312 8916 9364 8925
rect 9772 8959 9824 8968
rect 9772 8925 9781 8959
rect 9781 8925 9815 8959
rect 9815 8925 9824 8959
rect 9772 8916 9824 8925
rect 9864 8916 9916 8968
rect 11060 8916 11112 8968
rect 11428 8916 11480 8968
rect 11520 8916 11572 8968
rect 11796 8916 11848 8968
rect 8944 8780 8996 8832
rect 9496 8848 9548 8900
rect 11336 8848 11388 8900
rect 11980 8959 12032 8968
rect 11980 8925 11989 8959
rect 11989 8925 12023 8959
rect 12023 8925 12032 8959
rect 11980 8916 12032 8925
rect 12072 8959 12124 8968
rect 12072 8925 12081 8959
rect 12081 8925 12115 8959
rect 12115 8925 12124 8959
rect 12072 8916 12124 8925
rect 12164 8959 12216 8968
rect 12164 8925 12173 8959
rect 12173 8925 12207 8959
rect 12207 8925 12216 8959
rect 12164 8916 12216 8925
rect 14004 8916 14056 8968
rect 14096 8823 14148 8832
rect 14096 8789 14105 8823
rect 14105 8789 14139 8823
rect 14139 8789 14148 8823
rect 14096 8780 14148 8789
rect 15292 8916 15344 8968
rect 16028 8984 16080 9036
rect 16212 8959 16264 8968
rect 16212 8925 16221 8959
rect 16221 8925 16255 8959
rect 16255 8925 16264 8959
rect 16212 8916 16264 8925
rect 21272 9052 21324 9104
rect 19340 8984 19392 9036
rect 19708 8984 19760 9036
rect 20996 8984 21048 9036
rect 22100 8984 22152 9036
rect 23756 9027 23808 9036
rect 23756 8993 23765 9027
rect 23765 8993 23799 9027
rect 23799 8993 23808 9027
rect 23756 8984 23808 8993
rect 18972 8916 19024 8968
rect 19064 8916 19116 8968
rect 26424 9120 26476 9172
rect 27620 9120 27672 9172
rect 27896 9120 27948 9172
rect 30288 9120 30340 9172
rect 30564 9163 30616 9172
rect 30564 9129 30573 9163
rect 30573 9129 30607 9163
rect 30607 9129 30616 9163
rect 30564 9120 30616 9129
rect 32680 9120 32732 9172
rect 33416 9120 33468 9172
rect 33508 9163 33560 9172
rect 33508 9129 33517 9163
rect 33517 9129 33551 9163
rect 33551 9129 33560 9163
rect 33508 9120 33560 9129
rect 34428 9120 34480 9172
rect 35992 9163 36044 9172
rect 35992 9129 36001 9163
rect 36001 9129 36035 9163
rect 36035 9129 36044 9163
rect 35992 9120 36044 9129
rect 37464 9163 37516 9172
rect 37464 9129 37473 9163
rect 37473 9129 37507 9163
rect 37507 9129 37516 9163
rect 37464 9120 37516 9129
rect 25228 8984 25280 9036
rect 28080 9095 28132 9104
rect 28080 9061 28089 9095
rect 28089 9061 28123 9095
rect 28123 9061 28132 9095
rect 28080 9052 28132 9061
rect 17592 8891 17644 8900
rect 17592 8857 17601 8891
rect 17601 8857 17635 8891
rect 17635 8857 17644 8891
rect 17592 8848 17644 8857
rect 14832 8780 14884 8832
rect 18972 8780 19024 8832
rect 19248 8780 19300 8832
rect 21916 8848 21968 8900
rect 22100 8848 22152 8900
rect 22560 8848 22612 8900
rect 27344 8848 27396 8900
rect 28264 8984 28316 9036
rect 29552 9052 29604 9104
rect 21088 8780 21140 8832
rect 27252 8780 27304 8832
rect 28540 8891 28592 8900
rect 28540 8857 28549 8891
rect 28549 8857 28583 8891
rect 28583 8857 28592 8891
rect 28540 8848 28592 8857
rect 29736 8916 29788 8968
rect 29920 8959 29972 8968
rect 29920 8925 29929 8959
rect 29929 8925 29963 8959
rect 29963 8925 29972 8959
rect 29920 8916 29972 8925
rect 30104 9027 30156 9036
rect 30104 8993 30113 9027
rect 30113 8993 30147 9027
rect 30147 8993 30156 9027
rect 30104 8984 30156 8993
rect 30196 8984 30248 9036
rect 30472 8984 30524 9036
rect 31668 9052 31720 9104
rect 31852 8916 31904 8968
rect 32036 8916 32088 8968
rect 28632 8780 28684 8832
rect 30196 8891 30248 8900
rect 30196 8857 30205 8891
rect 30205 8857 30239 8891
rect 30239 8857 30248 8891
rect 30196 8848 30248 8857
rect 30288 8848 30340 8900
rect 30472 8848 30524 8900
rect 34060 9052 34112 9104
rect 34336 9052 34388 9104
rect 32312 8959 32364 8968
rect 32312 8925 32321 8959
rect 32321 8925 32355 8959
rect 32355 8925 32364 8959
rect 32312 8916 32364 8925
rect 33048 8916 33100 8968
rect 34244 8984 34296 9036
rect 33692 8916 33744 8968
rect 33784 8848 33836 8900
rect 37372 8984 37424 9036
rect 34612 8916 34664 8968
rect 35808 8959 35860 8968
rect 35808 8925 35817 8959
rect 35817 8925 35851 8959
rect 35851 8925 35860 8959
rect 35808 8916 35860 8925
rect 32220 8823 32272 8832
rect 32220 8789 32229 8823
rect 32229 8789 32263 8823
rect 32263 8789 32272 8823
rect 32220 8780 32272 8789
rect 33692 8780 33744 8832
rect 35992 8848 36044 8900
rect 37832 8916 37884 8968
rect 37924 8959 37976 8968
rect 37924 8925 37933 8959
rect 37933 8925 37967 8959
rect 37967 8925 37976 8959
rect 37924 8916 37976 8925
rect 38936 8916 38988 8968
rect 34336 8823 34388 8832
rect 34336 8789 34345 8823
rect 34345 8789 34379 8823
rect 34379 8789 34388 8823
rect 34336 8780 34388 8789
rect 34428 8780 34480 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 8944 8576 8996 8628
rect 9036 8576 9088 8628
rect 11336 8576 11388 8628
rect 11980 8576 12032 8628
rect 12716 8576 12768 8628
rect 13728 8576 13780 8628
rect 17592 8576 17644 8628
rect 19248 8576 19300 8628
rect 19432 8576 19484 8628
rect 27160 8576 27212 8628
rect 28632 8576 28684 8628
rect 28724 8576 28776 8628
rect 30472 8576 30524 8628
rect 9128 8483 9180 8492
rect 9128 8449 9137 8483
rect 9137 8449 9171 8483
rect 9171 8449 9180 8483
rect 9128 8440 9180 8449
rect 11520 8440 11572 8492
rect 11612 8440 11664 8492
rect 11980 8483 12032 8492
rect 11980 8449 11989 8483
rect 11989 8449 12023 8483
rect 12023 8449 12032 8483
rect 11980 8440 12032 8449
rect 12164 8483 12216 8492
rect 12164 8449 12173 8483
rect 12173 8449 12207 8483
rect 12207 8449 12216 8483
rect 12164 8440 12216 8449
rect 14372 8508 14424 8560
rect 16764 8508 16816 8560
rect 17316 8551 17368 8560
rect 17316 8517 17325 8551
rect 17325 8517 17359 8551
rect 17359 8517 17368 8551
rect 17316 8508 17368 8517
rect 13544 8483 13596 8492
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 13728 8440 13780 8492
rect 15108 8440 15160 8492
rect 15292 8440 15344 8492
rect 16028 8483 16080 8492
rect 16028 8449 16037 8483
rect 16037 8449 16071 8483
rect 16071 8449 16080 8483
rect 16028 8440 16080 8449
rect 16212 8440 16264 8492
rect 7564 8304 7616 8356
rect 6092 8236 6144 8288
rect 8300 8236 8352 8288
rect 9128 8236 9180 8288
rect 9772 8304 9824 8356
rect 11336 8304 11388 8356
rect 11152 8236 11204 8288
rect 12164 8304 12216 8356
rect 16304 8415 16356 8424
rect 16304 8381 16313 8415
rect 16313 8381 16347 8415
rect 16347 8381 16356 8415
rect 16304 8372 16356 8381
rect 16396 8372 16448 8424
rect 19984 8508 20036 8560
rect 27252 8508 27304 8560
rect 28356 8508 28408 8560
rect 19524 8483 19576 8492
rect 19524 8449 19533 8483
rect 19533 8449 19567 8483
rect 19567 8449 19576 8483
rect 19524 8440 19576 8449
rect 20076 8440 20128 8492
rect 18328 8372 18380 8424
rect 26976 8415 27028 8424
rect 26976 8381 26985 8415
rect 26985 8381 27019 8415
rect 27019 8381 27028 8415
rect 26976 8372 27028 8381
rect 28080 8483 28132 8492
rect 28080 8449 28089 8483
rect 28089 8449 28123 8483
rect 28123 8449 28132 8483
rect 28080 8440 28132 8449
rect 28356 8415 28408 8424
rect 28356 8381 28365 8415
rect 28365 8381 28399 8415
rect 28399 8381 28408 8415
rect 28356 8372 28408 8381
rect 28632 8483 28684 8492
rect 28632 8449 28641 8483
rect 28641 8449 28675 8483
rect 28675 8449 28684 8483
rect 28632 8440 28684 8449
rect 29460 8440 29512 8492
rect 29644 8440 29696 8492
rect 31392 8483 31444 8492
rect 31392 8449 31401 8483
rect 31401 8449 31435 8483
rect 31435 8449 31444 8483
rect 31392 8440 31444 8449
rect 31668 8483 31720 8492
rect 31668 8449 31677 8483
rect 31677 8449 31711 8483
rect 31711 8449 31720 8483
rect 31668 8440 31720 8449
rect 32036 8508 32088 8560
rect 31208 8372 31260 8424
rect 32220 8440 32272 8492
rect 33508 8576 33560 8628
rect 33692 8619 33744 8628
rect 33692 8585 33701 8619
rect 33701 8585 33735 8619
rect 33735 8585 33744 8619
rect 33692 8576 33744 8585
rect 35808 8576 35860 8628
rect 37924 8576 37976 8628
rect 34428 8508 34480 8560
rect 34520 8508 34572 8560
rect 35900 8508 35952 8560
rect 32036 8372 32088 8424
rect 33048 8415 33100 8424
rect 33048 8381 33057 8415
rect 33057 8381 33091 8415
rect 33091 8381 33100 8415
rect 33048 8372 33100 8381
rect 11796 8236 11848 8288
rect 16672 8279 16724 8288
rect 16672 8245 16681 8279
rect 16681 8245 16715 8279
rect 16715 8245 16724 8279
rect 16672 8236 16724 8245
rect 18604 8236 18656 8288
rect 20628 8236 20680 8288
rect 27436 8236 27488 8288
rect 27712 8279 27764 8288
rect 27712 8245 27721 8279
rect 27721 8245 27755 8279
rect 27755 8245 27764 8279
rect 27712 8236 27764 8245
rect 28080 8236 28132 8288
rect 28632 8236 28684 8288
rect 30012 8304 30064 8356
rect 30288 8236 30340 8288
rect 31668 8304 31720 8356
rect 33232 8304 33284 8356
rect 34244 8483 34296 8492
rect 34244 8449 34253 8483
rect 34253 8449 34287 8483
rect 34287 8449 34296 8483
rect 34244 8440 34296 8449
rect 35348 8440 35400 8492
rect 37464 8483 37516 8492
rect 37464 8449 37473 8483
rect 37473 8449 37507 8483
rect 37507 8449 37516 8483
rect 37464 8440 37516 8449
rect 37556 8483 37608 8492
rect 37556 8449 37565 8483
rect 37565 8449 37599 8483
rect 37599 8449 37608 8483
rect 37556 8440 37608 8449
rect 38108 8483 38160 8492
rect 38108 8449 38117 8483
rect 38117 8449 38151 8483
rect 38151 8449 38160 8483
rect 38108 8440 38160 8449
rect 38384 8483 38436 8492
rect 38384 8449 38393 8483
rect 38393 8449 38427 8483
rect 38427 8449 38436 8483
rect 38384 8440 38436 8449
rect 33968 8372 34020 8424
rect 34796 8372 34848 8424
rect 38200 8372 38252 8424
rect 41144 8304 41196 8356
rect 32772 8236 32824 8288
rect 33876 8236 33928 8288
rect 34336 8279 34388 8288
rect 34336 8245 34345 8279
rect 34345 8245 34379 8279
rect 34379 8245 34388 8279
rect 34336 8236 34388 8245
rect 35716 8236 35768 8288
rect 41052 8236 41104 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 7564 8032 7616 8084
rect 7748 8032 7800 8084
rect 8116 8032 8168 8084
rect 7472 7964 7524 8016
rect 8208 7964 8260 8016
rect 11060 8007 11112 8016
rect 11060 7973 11069 8007
rect 11069 7973 11103 8007
rect 11103 7973 11112 8007
rect 11060 7964 11112 7973
rect 8024 7896 8076 7948
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 11152 7828 11204 7880
rect 940 7760 992 7812
rect 8392 7803 8444 7812
rect 8392 7769 8401 7803
rect 8401 7769 8435 7803
rect 8435 7769 8444 7803
rect 8392 7760 8444 7769
rect 8668 7760 8720 7812
rect 11796 7828 11848 7880
rect 11888 7871 11940 7880
rect 11888 7837 11897 7871
rect 11897 7837 11931 7871
rect 11931 7837 11940 7871
rect 11888 7828 11940 7837
rect 12072 7828 12124 7880
rect 18972 8032 19024 8084
rect 12716 7964 12768 8016
rect 12716 7828 12768 7880
rect 13544 7964 13596 8016
rect 12256 7760 12308 7812
rect 19432 7896 19484 7948
rect 20260 8032 20312 8084
rect 20812 8032 20864 8084
rect 23572 7964 23624 8016
rect 26976 8032 27028 8084
rect 29552 8032 29604 8084
rect 29828 8032 29880 8084
rect 30932 8032 30984 8084
rect 27712 7964 27764 8016
rect 32404 8032 32456 8084
rect 34060 8032 34112 8084
rect 38384 8032 38436 8084
rect 21824 7896 21876 7948
rect 24216 7896 24268 7948
rect 14004 7828 14056 7880
rect 17776 7828 17828 7880
rect 18880 7828 18932 7880
rect 18696 7760 18748 7812
rect 8116 7735 8168 7744
rect 8116 7701 8125 7735
rect 8125 7701 8159 7735
rect 8159 7701 8168 7735
rect 8116 7692 8168 7701
rect 11428 7735 11480 7744
rect 11428 7701 11437 7735
rect 11437 7701 11471 7735
rect 11471 7701 11480 7735
rect 11428 7692 11480 7701
rect 11520 7692 11572 7744
rect 11704 7692 11756 7744
rect 15476 7692 15528 7744
rect 16212 7692 16264 7744
rect 23388 7828 23440 7880
rect 32036 7964 32088 8016
rect 29736 7896 29788 7948
rect 20260 7803 20312 7812
rect 20260 7769 20269 7803
rect 20269 7769 20303 7803
rect 20303 7769 20312 7803
rect 20260 7760 20312 7769
rect 20720 7760 20772 7812
rect 21916 7803 21968 7812
rect 20904 7692 20956 7744
rect 21916 7769 21925 7803
rect 21925 7769 21959 7803
rect 21959 7769 21968 7803
rect 21916 7760 21968 7769
rect 29276 7828 29328 7880
rect 30104 7828 30156 7880
rect 31576 7828 31628 7880
rect 34888 7828 34940 7880
rect 34980 7828 35032 7880
rect 23572 7735 23624 7744
rect 23572 7701 23581 7735
rect 23581 7701 23615 7735
rect 23615 7701 23624 7735
rect 23572 7692 23624 7701
rect 24952 7760 25004 7812
rect 26056 7760 26108 7812
rect 27160 7760 27212 7812
rect 29460 7760 29512 7812
rect 29552 7803 29604 7812
rect 29552 7769 29561 7803
rect 29561 7769 29595 7803
rect 29595 7769 29604 7803
rect 29552 7760 29604 7769
rect 29736 7803 29788 7812
rect 29736 7769 29745 7803
rect 29745 7769 29779 7803
rect 29779 7769 29788 7803
rect 29736 7760 29788 7769
rect 30472 7760 30524 7812
rect 33784 7760 33836 7812
rect 35072 7803 35124 7812
rect 35072 7769 35081 7803
rect 35081 7769 35115 7803
rect 35115 7769 35124 7803
rect 35072 7760 35124 7769
rect 28356 7692 28408 7744
rect 29092 7692 29144 7744
rect 30196 7692 30248 7744
rect 30656 7692 30708 7744
rect 32128 7692 32180 7744
rect 34704 7692 34756 7744
rect 34980 7735 35032 7744
rect 34980 7701 34995 7735
rect 34995 7701 35029 7735
rect 35029 7701 35032 7735
rect 34980 7692 35032 7701
rect 35348 7692 35400 7744
rect 35992 7828 36044 7880
rect 37464 7896 37516 7948
rect 37556 7896 37608 7948
rect 35716 7803 35768 7812
rect 35716 7769 35725 7803
rect 35725 7769 35759 7803
rect 35759 7769 35768 7803
rect 35716 7760 35768 7769
rect 35808 7760 35860 7812
rect 36084 7692 36136 7744
rect 40776 7692 40828 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 7840 7488 7892 7540
rect 8116 7488 8168 7540
rect 8668 7488 8720 7540
rect 7196 7420 7248 7472
rect 7748 7395 7800 7404
rect 7748 7361 7757 7395
rect 7757 7361 7791 7395
rect 7791 7361 7800 7395
rect 7748 7352 7800 7361
rect 7840 7395 7892 7404
rect 7840 7361 7849 7395
rect 7849 7361 7883 7395
rect 7883 7361 7892 7395
rect 7840 7352 7892 7361
rect 8300 7352 8352 7404
rect 8392 7395 8444 7404
rect 8392 7361 8401 7395
rect 8401 7361 8435 7395
rect 8435 7361 8444 7395
rect 8392 7352 8444 7361
rect 8484 7352 8536 7404
rect 9128 7463 9180 7472
rect 9128 7429 9137 7463
rect 9137 7429 9171 7463
rect 9171 7429 9180 7463
rect 9128 7420 9180 7429
rect 7564 7284 7616 7336
rect 8208 7284 8260 7336
rect 8852 7284 8904 7336
rect 11796 7488 11848 7540
rect 11520 7420 11572 7472
rect 11704 7352 11756 7404
rect 11612 7216 11664 7268
rect 11888 7284 11940 7336
rect 12256 7395 12308 7404
rect 12256 7361 12265 7395
rect 12265 7361 12299 7395
rect 12299 7361 12308 7395
rect 12256 7352 12308 7361
rect 14096 7488 14148 7540
rect 12716 7463 12768 7472
rect 12716 7429 12725 7463
rect 12725 7429 12759 7463
rect 12759 7429 12768 7463
rect 12716 7420 12768 7429
rect 14004 7463 14056 7472
rect 14004 7429 14013 7463
rect 14013 7429 14047 7463
rect 14047 7429 14056 7463
rect 14004 7420 14056 7429
rect 12532 7352 12584 7404
rect 7380 7148 7432 7200
rect 7472 7191 7524 7200
rect 7472 7157 7481 7191
rect 7481 7157 7515 7191
rect 7515 7157 7524 7191
rect 7472 7148 7524 7157
rect 7748 7148 7800 7200
rect 8484 7148 8536 7200
rect 12808 7284 12860 7336
rect 14372 7352 14424 7404
rect 14832 7352 14884 7404
rect 16028 7488 16080 7540
rect 15016 7284 15068 7336
rect 13820 7216 13872 7268
rect 15476 7352 15528 7404
rect 15384 7327 15436 7336
rect 15384 7293 15393 7327
rect 15393 7293 15427 7327
rect 15427 7293 15436 7327
rect 15384 7284 15436 7293
rect 15844 7327 15896 7336
rect 15844 7293 15854 7327
rect 15854 7293 15888 7327
rect 15888 7293 15896 7327
rect 15844 7284 15896 7293
rect 16028 7352 16080 7404
rect 16212 7395 16264 7404
rect 16212 7361 16221 7395
rect 16221 7361 16255 7395
rect 16255 7361 16264 7395
rect 16212 7352 16264 7361
rect 16672 7352 16724 7404
rect 19340 7488 19392 7540
rect 20260 7488 20312 7540
rect 18696 7420 18748 7472
rect 18880 7420 18932 7472
rect 20352 7420 20404 7472
rect 20812 7352 20864 7404
rect 23572 7488 23624 7540
rect 24124 7488 24176 7540
rect 25780 7488 25832 7540
rect 22100 7395 22152 7404
rect 22100 7361 22109 7395
rect 22109 7361 22143 7395
rect 22143 7361 22152 7395
rect 22100 7352 22152 7361
rect 26148 7420 26200 7472
rect 24860 7352 24912 7404
rect 25228 7352 25280 7404
rect 27160 7463 27212 7472
rect 27160 7429 27169 7463
rect 27169 7429 27203 7463
rect 27203 7429 27212 7463
rect 27160 7420 27212 7429
rect 28356 7420 28408 7472
rect 19432 7284 19484 7336
rect 15476 7191 15528 7200
rect 15476 7157 15485 7191
rect 15485 7157 15519 7191
rect 15519 7157 15528 7191
rect 15476 7148 15528 7157
rect 15568 7148 15620 7200
rect 16304 7191 16356 7200
rect 16304 7157 16313 7191
rect 16313 7157 16347 7191
rect 16347 7157 16356 7191
rect 16304 7148 16356 7157
rect 26792 7284 26844 7336
rect 27436 7352 27488 7404
rect 27620 7395 27672 7404
rect 27620 7361 27629 7395
rect 27629 7361 27663 7395
rect 27663 7361 27672 7395
rect 27620 7352 27672 7361
rect 29552 7420 29604 7472
rect 28632 7284 28684 7336
rect 29184 7395 29236 7404
rect 29184 7361 29193 7395
rect 29193 7361 29227 7395
rect 29227 7361 29236 7395
rect 29184 7352 29236 7361
rect 29276 7352 29328 7404
rect 29460 7352 29512 7404
rect 29828 7352 29880 7404
rect 29920 7395 29972 7404
rect 29920 7361 29929 7395
rect 29929 7361 29963 7395
rect 29963 7361 29972 7395
rect 29920 7352 29972 7361
rect 30288 7352 30340 7404
rect 29092 7327 29144 7336
rect 29092 7293 29101 7327
rect 29101 7293 29135 7327
rect 29135 7293 29144 7327
rect 29092 7284 29144 7293
rect 27252 7148 27304 7200
rect 27528 7191 27580 7200
rect 27528 7157 27537 7191
rect 27537 7157 27571 7191
rect 27571 7157 27580 7191
rect 27528 7148 27580 7157
rect 28632 7191 28684 7200
rect 28632 7157 28641 7191
rect 28641 7157 28675 7191
rect 28675 7157 28684 7191
rect 28632 7148 28684 7157
rect 28908 7148 28960 7200
rect 30472 7352 30524 7404
rect 30656 7352 30708 7404
rect 30932 7352 30984 7404
rect 31208 7352 31260 7404
rect 31576 7463 31628 7472
rect 31576 7429 31585 7463
rect 31585 7429 31619 7463
rect 31619 7429 31628 7463
rect 31576 7420 31628 7429
rect 31668 7352 31720 7404
rect 32036 7420 32088 7472
rect 32128 7420 32180 7472
rect 32496 7463 32548 7472
rect 32496 7429 32505 7463
rect 32505 7429 32539 7463
rect 32539 7429 32548 7463
rect 32496 7420 32548 7429
rect 34336 7488 34388 7540
rect 35072 7488 35124 7540
rect 32036 7284 32088 7336
rect 32772 7395 32824 7404
rect 32772 7361 32781 7395
rect 32781 7361 32815 7395
rect 32815 7361 32824 7395
rect 32772 7352 32824 7361
rect 33692 7420 33744 7472
rect 33140 7352 33192 7404
rect 33232 7352 33284 7404
rect 33416 7395 33468 7404
rect 33416 7361 33425 7395
rect 33425 7361 33459 7395
rect 33459 7361 33468 7395
rect 33416 7352 33468 7361
rect 33876 7352 33928 7404
rect 34980 7420 35032 7472
rect 35348 7463 35400 7472
rect 35348 7429 35357 7463
rect 35357 7429 35391 7463
rect 35391 7429 35400 7463
rect 35348 7420 35400 7429
rect 29644 7216 29696 7268
rect 30380 7259 30432 7268
rect 30380 7225 30389 7259
rect 30389 7225 30423 7259
rect 30423 7225 30432 7259
rect 30380 7216 30432 7225
rect 30748 7148 30800 7200
rect 31208 7148 31260 7200
rect 31300 7191 31352 7200
rect 31300 7157 31309 7191
rect 31309 7157 31343 7191
rect 31343 7157 31352 7191
rect 31300 7148 31352 7157
rect 34888 7352 34940 7404
rect 35164 7352 35216 7404
rect 35256 7352 35308 7404
rect 34888 7216 34940 7268
rect 34980 7216 35032 7268
rect 35716 7488 35768 7540
rect 36176 7531 36228 7540
rect 36176 7497 36185 7531
rect 36185 7497 36219 7531
rect 36219 7497 36228 7531
rect 36176 7488 36228 7497
rect 36452 7488 36504 7540
rect 36912 7488 36964 7540
rect 35992 7463 36044 7472
rect 35992 7429 36001 7463
rect 36001 7429 36035 7463
rect 36035 7429 36044 7463
rect 35992 7420 36044 7429
rect 35716 7352 35768 7404
rect 36452 7395 36504 7404
rect 36452 7361 36461 7395
rect 36461 7361 36495 7395
rect 36495 7361 36504 7395
rect 36452 7352 36504 7361
rect 32128 7191 32180 7200
rect 32128 7157 32137 7191
rect 32137 7157 32171 7191
rect 32171 7157 32180 7191
rect 32128 7148 32180 7157
rect 32312 7148 32364 7200
rect 32404 7148 32456 7200
rect 33784 7148 33836 7200
rect 34796 7148 34848 7200
rect 35716 7259 35768 7268
rect 35716 7225 35725 7259
rect 35725 7225 35759 7259
rect 35759 7225 35768 7259
rect 35716 7216 35768 7225
rect 35624 7148 35676 7200
rect 35900 7148 35952 7200
rect 36544 7191 36596 7200
rect 36544 7157 36553 7191
rect 36553 7157 36587 7191
rect 36587 7157 36596 7191
rect 36544 7148 36596 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 7564 6944 7616 6996
rect 11428 6944 11480 6996
rect 12624 6944 12676 6996
rect 12808 6944 12860 6996
rect 1860 6740 1912 6792
rect 4068 6740 4120 6792
rect 5172 6783 5224 6792
rect 5172 6749 5181 6783
rect 5181 6749 5215 6783
rect 5215 6749 5224 6783
rect 5172 6740 5224 6749
rect 6552 6740 6604 6792
rect 8208 6876 8260 6928
rect 10324 6876 10376 6928
rect 7288 6740 7340 6792
rect 7472 6740 7524 6792
rect 8484 6783 8536 6792
rect 8484 6749 8493 6783
rect 8493 6749 8527 6783
rect 8527 6749 8536 6783
rect 8484 6740 8536 6749
rect 8668 6783 8720 6792
rect 8668 6749 8677 6783
rect 8677 6749 8711 6783
rect 8711 6749 8720 6783
rect 8668 6740 8720 6749
rect 8852 6740 8904 6792
rect 9680 6740 9732 6792
rect 11244 6740 11296 6792
rect 11336 6783 11388 6792
rect 11336 6749 11345 6783
rect 11345 6749 11379 6783
rect 11379 6749 11388 6783
rect 11336 6740 11388 6749
rect 11520 6783 11572 6792
rect 11520 6749 11527 6783
rect 11527 6749 11572 6783
rect 11520 6740 11572 6749
rect 15476 6944 15528 6996
rect 27528 6944 27580 6996
rect 27620 6944 27672 6996
rect 28172 6944 28224 6996
rect 27712 6876 27764 6928
rect 28632 6876 28684 6928
rect 29184 6944 29236 6996
rect 29644 6876 29696 6928
rect 32036 6944 32088 6996
rect 32220 6987 32272 6996
rect 32220 6953 32229 6987
rect 32229 6953 32263 6987
rect 32263 6953 32272 6987
rect 32220 6944 32272 6953
rect 32312 6944 32364 6996
rect 31668 6876 31720 6928
rect 14280 6808 14332 6860
rect 15016 6851 15068 6860
rect 15016 6817 15025 6851
rect 15025 6817 15059 6851
rect 15059 6817 15068 6851
rect 15016 6808 15068 6817
rect 16304 6808 16356 6860
rect 17316 6808 17368 6860
rect 18420 6851 18472 6860
rect 18420 6817 18429 6851
rect 18429 6817 18463 6851
rect 18463 6817 18472 6851
rect 18420 6808 18472 6817
rect 19064 6808 19116 6860
rect 20904 6808 20956 6860
rect 5540 6672 5592 6724
rect 7380 6672 7432 6724
rect 7656 6647 7708 6656
rect 7656 6613 7665 6647
rect 7665 6613 7699 6647
rect 7699 6613 7708 6647
rect 7656 6604 7708 6613
rect 7932 6604 7984 6656
rect 10968 6672 11020 6724
rect 11704 6715 11756 6724
rect 11704 6681 11713 6715
rect 11713 6681 11747 6715
rect 11747 6681 11756 6715
rect 11704 6672 11756 6681
rect 8392 6647 8444 6656
rect 8392 6613 8401 6647
rect 8401 6613 8435 6647
rect 8435 6613 8444 6647
rect 8392 6604 8444 6613
rect 11152 6604 11204 6656
rect 12072 6715 12124 6724
rect 12072 6681 12081 6715
rect 12081 6681 12115 6715
rect 12115 6681 12124 6715
rect 12072 6672 12124 6681
rect 12256 6672 12308 6724
rect 11980 6647 12032 6656
rect 11980 6613 11989 6647
rect 11989 6613 12023 6647
rect 12023 6613 12032 6647
rect 11980 6604 12032 6613
rect 13636 6783 13688 6792
rect 12992 6715 13044 6724
rect 12992 6681 13022 6715
rect 13022 6681 13044 6715
rect 13636 6749 13645 6783
rect 13645 6749 13679 6783
rect 13679 6749 13688 6783
rect 13636 6740 13688 6749
rect 13728 6783 13780 6792
rect 13728 6749 13737 6783
rect 13737 6749 13771 6783
rect 13771 6749 13780 6783
rect 13728 6740 13780 6749
rect 14004 6740 14056 6792
rect 12992 6672 13044 6681
rect 13544 6672 13596 6724
rect 17500 6740 17552 6792
rect 17868 6672 17920 6724
rect 18052 6740 18104 6792
rect 19432 6783 19484 6792
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 21088 6740 21140 6792
rect 21824 6851 21876 6860
rect 21824 6817 21833 6851
rect 21833 6817 21867 6851
rect 21867 6817 21876 6851
rect 21824 6808 21876 6817
rect 26056 6851 26108 6860
rect 26056 6817 26065 6851
rect 26065 6817 26099 6851
rect 26099 6817 26108 6851
rect 26056 6808 26108 6817
rect 26792 6808 26844 6860
rect 30380 6851 30432 6860
rect 30380 6817 30389 6851
rect 30389 6817 30423 6851
rect 30423 6817 30432 6851
rect 30380 6808 30432 6817
rect 31484 6808 31536 6860
rect 32128 6808 32180 6860
rect 32496 6876 32548 6928
rect 33508 6876 33560 6928
rect 24492 6740 24544 6792
rect 13820 6604 13872 6656
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 14556 6647 14608 6656
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14556 6604 14608 6613
rect 15292 6647 15344 6656
rect 15292 6613 15301 6647
rect 15301 6613 15335 6647
rect 15335 6613 15344 6647
rect 15292 6604 15344 6613
rect 18696 6604 18748 6656
rect 20444 6604 20496 6656
rect 22560 6672 22612 6724
rect 23848 6715 23900 6724
rect 23848 6681 23857 6715
rect 23857 6681 23891 6715
rect 23891 6681 23900 6715
rect 23848 6672 23900 6681
rect 25780 6672 25832 6724
rect 27436 6740 27488 6792
rect 28724 6740 28776 6792
rect 28908 6740 28960 6792
rect 26240 6672 26292 6724
rect 22376 6604 22428 6656
rect 26700 6604 26752 6656
rect 29276 6740 29328 6792
rect 29460 6740 29512 6792
rect 29644 6672 29696 6724
rect 30288 6740 30340 6792
rect 30656 6740 30708 6792
rect 31300 6740 31352 6792
rect 29000 6647 29052 6656
rect 29000 6613 29009 6647
rect 29009 6613 29043 6647
rect 29043 6613 29052 6647
rect 29000 6604 29052 6613
rect 32404 6740 32456 6792
rect 32496 6783 32548 6792
rect 32496 6749 32505 6783
rect 32505 6749 32539 6783
rect 32539 6749 32548 6783
rect 32496 6740 32548 6749
rect 31576 6647 31628 6656
rect 31576 6613 31585 6647
rect 31585 6613 31619 6647
rect 31619 6613 31628 6647
rect 31576 6604 31628 6613
rect 33048 6672 33100 6724
rect 32496 6604 32548 6656
rect 32680 6647 32732 6656
rect 32680 6613 32689 6647
rect 32689 6613 32723 6647
rect 32723 6613 32732 6647
rect 32680 6604 32732 6613
rect 33324 6783 33376 6792
rect 33324 6749 33333 6783
rect 33333 6749 33367 6783
rect 33367 6749 33376 6783
rect 33324 6740 33376 6749
rect 34152 6944 34204 6996
rect 34336 6944 34388 6996
rect 34704 6944 34756 6996
rect 36452 6944 36504 6996
rect 36544 6876 36596 6928
rect 34612 6808 34664 6860
rect 33968 6783 34020 6792
rect 33968 6749 33977 6783
rect 33977 6749 34011 6783
rect 34011 6749 34020 6783
rect 33968 6740 34020 6749
rect 34152 6783 34204 6792
rect 34152 6749 34161 6783
rect 34161 6749 34195 6783
rect 34195 6749 34204 6783
rect 34152 6740 34204 6749
rect 34428 6783 34480 6792
rect 34428 6749 34437 6783
rect 34437 6749 34471 6783
rect 34471 6749 34480 6783
rect 34428 6740 34480 6749
rect 33232 6672 33284 6724
rect 33876 6672 33928 6724
rect 34336 6672 34388 6724
rect 34980 6740 35032 6792
rect 35624 6808 35676 6860
rect 35348 6740 35400 6792
rect 35808 6740 35860 6792
rect 35532 6647 35584 6656
rect 35532 6613 35541 6647
rect 35541 6613 35575 6647
rect 35575 6613 35584 6647
rect 35532 6604 35584 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 5540 6443 5592 6452
rect 5540 6409 5549 6443
rect 5549 6409 5583 6443
rect 5583 6409 5592 6443
rect 5540 6400 5592 6409
rect 5172 6264 5224 6316
rect 7656 6400 7708 6452
rect 8392 6400 8444 6452
rect 10048 6400 10100 6452
rect 10876 6443 10928 6452
rect 10876 6409 10885 6443
rect 10885 6409 10919 6443
rect 10919 6409 10928 6443
rect 10876 6400 10928 6409
rect 11520 6443 11572 6452
rect 11520 6409 11529 6443
rect 11529 6409 11563 6443
rect 11563 6409 11572 6443
rect 11520 6400 11572 6409
rect 11704 6400 11756 6452
rect 12072 6400 12124 6452
rect 12808 6400 12860 6452
rect 13636 6400 13688 6452
rect 14556 6400 14608 6452
rect 15292 6400 15344 6452
rect 19432 6400 19484 6452
rect 20444 6400 20496 6452
rect 20628 6443 20680 6452
rect 20628 6409 20637 6443
rect 20637 6409 20671 6443
rect 20671 6409 20680 6443
rect 20628 6400 20680 6409
rect 7932 6332 7984 6384
rect 10324 6375 10376 6384
rect 10324 6341 10333 6375
rect 10333 6341 10367 6375
rect 10367 6341 10376 6375
rect 10324 6332 10376 6341
rect 9680 6264 9732 6316
rect 6276 6196 6328 6248
rect 6828 6196 6880 6248
rect 8116 6196 8168 6248
rect 8668 6196 8720 6248
rect 11152 6332 11204 6384
rect 12348 6332 12400 6384
rect 11060 6264 11112 6316
rect 11796 6264 11848 6316
rect 12992 6264 13044 6316
rect 11612 6196 11664 6248
rect 12256 6196 12308 6248
rect 14372 6264 14424 6316
rect 17960 6332 18012 6384
rect 19064 6332 19116 6384
rect 19340 6332 19392 6384
rect 20076 6264 20128 6316
rect 18972 6239 19024 6248
rect 18972 6205 18981 6239
rect 18981 6205 19015 6239
rect 19015 6205 19024 6239
rect 18972 6196 19024 6205
rect 22376 6375 22428 6384
rect 22376 6341 22385 6375
rect 22385 6341 22419 6375
rect 22419 6341 22428 6375
rect 22376 6332 22428 6341
rect 10416 6103 10468 6112
rect 10416 6069 10425 6103
rect 10425 6069 10459 6103
rect 10459 6069 10468 6103
rect 10416 6060 10468 6069
rect 12164 6060 12216 6112
rect 12808 6060 12860 6112
rect 13452 6128 13504 6180
rect 18052 6128 18104 6180
rect 20812 6239 20864 6248
rect 20812 6205 20821 6239
rect 20821 6205 20855 6239
rect 20855 6205 20864 6239
rect 20812 6196 20864 6205
rect 14096 6060 14148 6112
rect 18972 6060 19024 6112
rect 20260 6060 20312 6112
rect 22284 6307 22336 6316
rect 22284 6273 22293 6307
rect 22293 6273 22327 6307
rect 22327 6273 22336 6307
rect 22284 6264 22336 6273
rect 23848 6332 23900 6384
rect 25228 6332 25280 6384
rect 26240 6443 26292 6452
rect 26240 6409 26249 6443
rect 26249 6409 26283 6443
rect 26283 6409 26292 6443
rect 26240 6400 26292 6409
rect 26700 6443 26752 6452
rect 26700 6409 26709 6443
rect 26709 6409 26743 6443
rect 26743 6409 26752 6443
rect 26700 6400 26752 6409
rect 29000 6332 29052 6384
rect 29552 6375 29604 6384
rect 29552 6341 29561 6375
rect 29561 6341 29595 6375
rect 29595 6341 29604 6375
rect 29552 6332 29604 6341
rect 33692 6375 33744 6384
rect 33692 6341 33701 6375
rect 33701 6341 33735 6375
rect 33735 6341 33744 6375
rect 33692 6332 33744 6341
rect 34428 6400 34480 6452
rect 40960 6332 41012 6384
rect 24492 6307 24544 6316
rect 24492 6273 24501 6307
rect 24501 6273 24535 6307
rect 24535 6273 24544 6307
rect 24492 6264 24544 6273
rect 27528 6264 27580 6316
rect 29184 6264 29236 6316
rect 29644 6305 29696 6316
rect 29644 6271 29653 6305
rect 29653 6271 29687 6305
rect 29687 6271 29696 6305
rect 29644 6264 29696 6271
rect 31300 6264 31352 6316
rect 32220 6264 32272 6316
rect 20996 6103 21048 6112
rect 20996 6069 21005 6103
rect 21005 6069 21039 6103
rect 21039 6069 21048 6103
rect 20996 6060 21048 6069
rect 21088 6060 21140 6112
rect 22008 6060 22060 6112
rect 28724 6060 28776 6112
rect 30840 6060 30892 6112
rect 33600 6060 33652 6112
rect 34336 6196 34388 6248
rect 34152 6128 34204 6180
rect 34796 6239 34848 6248
rect 34796 6205 34805 6239
rect 34805 6205 34839 6239
rect 34839 6205 34848 6239
rect 34796 6196 34848 6205
rect 34612 6060 34664 6112
rect 35716 6103 35768 6112
rect 35716 6069 35725 6103
rect 35725 6069 35759 6103
rect 35759 6069 35768 6103
rect 35716 6060 35768 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 6828 5856 6880 5908
rect 10876 5899 10928 5908
rect 10876 5865 10885 5899
rect 10885 5865 10919 5899
rect 10919 5865 10928 5899
rect 10876 5856 10928 5865
rect 18972 5856 19024 5908
rect 20260 5856 20312 5908
rect 20812 5856 20864 5908
rect 20996 5856 21048 5908
rect 21088 5899 21140 5908
rect 21088 5865 21097 5899
rect 21097 5865 21131 5899
rect 21131 5865 21140 5899
rect 21088 5856 21140 5865
rect 22008 5856 22060 5908
rect 22100 5856 22152 5908
rect 27804 5856 27856 5908
rect 33600 5856 33652 5908
rect 11152 5788 11204 5840
rect 15108 5788 15160 5840
rect 8116 5720 8168 5772
rect 9772 5720 9824 5772
rect 19340 5763 19392 5772
rect 19340 5729 19349 5763
rect 19349 5729 19383 5763
rect 19383 5729 19392 5763
rect 19340 5720 19392 5729
rect 27528 5788 27580 5840
rect 21824 5720 21876 5772
rect 21916 5720 21968 5772
rect 9404 5627 9456 5636
rect 9404 5593 9413 5627
rect 9413 5593 9447 5627
rect 9447 5593 9456 5627
rect 9404 5584 9456 5593
rect 9680 5584 9732 5636
rect 20720 5652 20772 5704
rect 22560 5652 22612 5704
rect 16304 5584 16356 5636
rect 16672 5584 16724 5636
rect 17868 5584 17920 5636
rect 18052 5584 18104 5636
rect 23204 5627 23256 5636
rect 23204 5593 23213 5627
rect 23213 5593 23247 5627
rect 23247 5593 23256 5627
rect 23204 5584 23256 5593
rect 27988 5652 28040 5704
rect 28172 5695 28224 5704
rect 28172 5661 28181 5695
rect 28181 5661 28215 5695
rect 28215 5661 28224 5695
rect 28172 5652 28224 5661
rect 28724 5695 28776 5704
rect 28724 5661 28733 5695
rect 28733 5661 28767 5695
rect 28767 5661 28776 5695
rect 28724 5652 28776 5661
rect 29368 5652 29420 5704
rect 30840 5720 30892 5772
rect 22468 5516 22520 5568
rect 26056 5516 26108 5568
rect 28264 5516 28316 5568
rect 30012 5584 30064 5636
rect 30748 5695 30800 5704
rect 30748 5661 30757 5695
rect 30757 5661 30791 5695
rect 30791 5661 30800 5695
rect 30748 5652 30800 5661
rect 34796 5720 34848 5772
rect 32588 5652 32640 5704
rect 33600 5652 33652 5704
rect 33692 5652 33744 5704
rect 34152 5695 34204 5704
rect 34152 5661 34161 5695
rect 34161 5661 34195 5695
rect 34195 5661 34204 5695
rect 36176 5856 36228 5908
rect 40960 5899 41012 5908
rect 40960 5865 40969 5899
rect 40969 5865 41003 5899
rect 41003 5865 41012 5899
rect 40960 5856 41012 5865
rect 34152 5652 34204 5661
rect 32772 5584 32824 5636
rect 35716 5652 35768 5704
rect 36912 5652 36964 5704
rect 29920 5516 29972 5568
rect 33232 5516 33284 5568
rect 34336 5559 34388 5568
rect 34336 5525 34345 5559
rect 34345 5525 34379 5559
rect 34379 5525 34388 5559
rect 34336 5516 34388 5525
rect 35348 5516 35400 5568
rect 41328 5516 41380 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 9404 5312 9456 5364
rect 10416 5312 10468 5364
rect 11980 5312 12032 5364
rect 12440 5312 12492 5364
rect 16304 5312 16356 5364
rect 13084 5244 13136 5296
rect 16672 5287 16724 5296
rect 16672 5253 16681 5287
rect 16681 5253 16715 5287
rect 16715 5253 16724 5287
rect 16672 5244 16724 5253
rect 16948 5176 17000 5228
rect 17132 5219 17184 5228
rect 17132 5185 17141 5219
rect 17141 5185 17175 5219
rect 17175 5185 17184 5219
rect 17132 5176 17184 5185
rect 18052 5176 18104 5228
rect 19340 5312 19392 5364
rect 20168 5312 20220 5364
rect 22468 5355 22520 5364
rect 22468 5321 22477 5355
rect 22477 5321 22511 5355
rect 22511 5321 22520 5355
rect 22468 5312 22520 5321
rect 18696 5244 18748 5296
rect 9956 5151 10008 5160
rect 9956 5117 9965 5151
rect 9965 5117 9999 5151
rect 9999 5117 10008 5151
rect 9956 5108 10008 5117
rect 9772 5040 9824 5092
rect 14372 4972 14424 5024
rect 17868 5108 17920 5160
rect 20628 5244 20680 5296
rect 29092 5244 29144 5296
rect 31576 5312 31628 5364
rect 31668 5312 31720 5364
rect 32680 5312 32732 5364
rect 32772 5312 32824 5364
rect 22284 5219 22336 5228
rect 22284 5185 22293 5219
rect 22293 5185 22327 5219
rect 22327 5185 22336 5219
rect 22284 5176 22336 5185
rect 23204 5108 23256 5160
rect 27252 5219 27304 5228
rect 27252 5185 27261 5219
rect 27261 5185 27295 5219
rect 27295 5185 27304 5219
rect 27252 5176 27304 5185
rect 27528 5219 27580 5228
rect 27528 5185 27537 5219
rect 27537 5185 27571 5219
rect 27571 5185 27580 5219
rect 27528 5176 27580 5185
rect 28172 5176 28224 5228
rect 28264 5176 28316 5228
rect 20076 4972 20128 5024
rect 20628 4972 20680 5024
rect 26976 5015 27028 5024
rect 26976 4981 26985 5015
rect 26985 4981 27019 5015
rect 27019 4981 27028 5015
rect 26976 4972 27028 4981
rect 27620 5040 27672 5092
rect 27712 5015 27764 5024
rect 27712 4981 27721 5015
rect 27721 4981 27755 5015
rect 27755 4981 27764 5015
rect 27712 4972 27764 4981
rect 29920 5176 29972 5228
rect 31024 5176 31076 5228
rect 31760 5176 31812 5228
rect 32588 5176 32640 5228
rect 33232 5176 33284 5228
rect 33508 5244 33560 5296
rect 34060 5244 34112 5296
rect 36912 5355 36964 5364
rect 36912 5321 36921 5355
rect 36921 5321 36955 5355
rect 36955 5321 36964 5355
rect 36912 5312 36964 5321
rect 35348 5244 35400 5296
rect 29000 4972 29052 5024
rect 29368 4972 29420 5024
rect 34796 5108 34848 5160
rect 36176 5108 36228 5160
rect 30932 5015 30984 5024
rect 30932 4981 30941 5015
rect 30941 4981 30975 5015
rect 30975 4981 30984 5015
rect 30932 4972 30984 4981
rect 31668 4972 31720 5024
rect 32956 5015 33008 5024
rect 32956 4981 32965 5015
rect 32965 4981 32999 5015
rect 32999 4981 33008 5015
rect 32956 4972 33008 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 9956 4768 10008 4820
rect 14372 4768 14424 4820
rect 17776 4811 17828 4820
rect 17776 4777 17785 4811
rect 17785 4777 17819 4811
rect 17819 4777 17828 4811
rect 17776 4768 17828 4777
rect 27528 4768 27580 4820
rect 28172 4768 28224 4820
rect 29092 4768 29144 4820
rect 31760 4811 31812 4820
rect 31760 4777 31769 4811
rect 31769 4777 31803 4811
rect 31803 4777 31812 4811
rect 31760 4768 31812 4777
rect 33600 4768 33652 4820
rect 1860 4675 1912 4684
rect 1860 4641 1869 4675
rect 1869 4641 1903 4675
rect 1903 4641 1912 4675
rect 1860 4632 1912 4641
rect 16304 4632 16356 4684
rect 26056 4632 26108 4684
rect 26976 4632 27028 4684
rect 6552 4564 6604 4616
rect 17868 4564 17920 4616
rect 27436 4564 27488 4616
rect 2136 4539 2188 4548
rect 2136 4505 2145 4539
rect 2145 4505 2179 4539
rect 2179 4505 2188 4539
rect 2136 4496 2188 4505
rect 29000 4632 29052 4684
rect 30012 4675 30064 4684
rect 30012 4641 30021 4675
rect 30021 4641 30055 4675
rect 30055 4641 30064 4675
rect 30012 4632 30064 4641
rect 31668 4632 31720 4684
rect 32956 4632 33008 4684
rect 29184 4564 29236 4616
rect 35992 4607 36044 4616
rect 35992 4573 36001 4607
rect 36001 4573 36035 4607
rect 36035 4573 36044 4607
rect 35992 4564 36044 4573
rect 30564 4496 30616 4548
rect 34060 4428 34112 4480
rect 36176 4471 36228 4480
rect 36176 4437 36185 4471
rect 36185 4437 36219 4471
rect 36219 4437 36228 4471
rect 36176 4428 36228 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 2136 4224 2188 4276
rect 30564 4267 30616 4276
rect 30564 4233 30573 4267
rect 30573 4233 30607 4267
rect 30607 4233 30616 4267
rect 30564 4224 30616 4233
rect 30932 4224 30984 4276
rect 940 4088 992 4140
rect 9772 4088 9824 4140
rect 10968 3927 11020 3936
rect 10968 3893 10977 3927
rect 10977 3893 11011 3927
rect 11011 3893 11020 3927
rect 10968 3884 11020 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 15016 3587 15068 3596
rect 15016 3553 15025 3587
rect 15025 3553 15059 3587
rect 15059 3553 15068 3587
rect 15016 3544 15068 3553
rect 20 3476 72 3528
rect 3608 3476 3660 3528
rect 14740 3519 14792 3528
rect 14740 3485 14749 3519
rect 14749 3485 14783 3519
rect 14783 3485 14792 3519
rect 14740 3476 14792 3485
rect 14188 3408 14240 3460
rect 23204 3408 23256 3460
rect 36728 3408 36780 3460
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 14740 3136 14792 3188
rect 3240 2796 3292 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 40776 2635 40828 2644
rect 40776 2601 40785 2635
rect 40785 2601 40819 2635
rect 40819 2601 40828 2635
rect 40776 2592 40828 2601
rect 20628 2456 20680 2508
rect 7288 2431 7340 2440
rect 7288 2397 7297 2431
rect 7297 2397 7331 2431
rect 7331 2397 7340 2431
rect 7288 2388 7340 2397
rect 22100 2431 22152 2440
rect 22100 2397 22109 2431
rect 22109 2397 22143 2431
rect 22143 2397 22152 2431
rect 22100 2388 22152 2397
rect 29000 2388 29052 2440
rect 29828 2499 29880 2508
rect 29828 2465 29837 2499
rect 29837 2465 29871 2499
rect 29871 2465 29880 2499
rect 29828 2456 29880 2465
rect 40684 2363 40736 2372
rect 40684 2329 40693 2363
rect 40693 2329 40727 2363
rect 40727 2329 40736 2363
rect 40684 2320 40736 2329
rect 7104 2252 7156 2304
rect 22008 2252 22060 2304
rect 33140 2295 33192 2304
rect 33140 2261 33149 2295
rect 33149 2261 33183 2295
rect 33183 2261 33192 2295
rect 33140 2252 33192 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 1306 43893 1362 44693
rect 5170 44010 5226 44693
rect 5170 43982 5396 44010
rect 5170 43893 5226 43982
rect 1320 42362 1348 43893
rect 3422 42936 3478 42945
rect 3422 42871 3478 42880
rect 1308 42356 1360 42362
rect 1308 42298 1360 42304
rect 1492 42220 1544 42226
rect 1492 42162 1544 42168
rect 1504 39506 1532 42162
rect 1676 41200 1728 41206
rect 1676 41142 1728 41148
rect 1688 40730 1716 41142
rect 3436 41070 3464 42871
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 3608 41132 3660 41138
rect 3608 41074 3660 41080
rect 2688 41064 2740 41070
rect 2688 41006 2740 41012
rect 2872 41064 2924 41070
rect 2872 41006 2924 41012
rect 3424 41064 3476 41070
rect 3424 41006 3476 41012
rect 1676 40724 1728 40730
rect 1676 40666 1728 40672
rect 2700 39982 2728 41006
rect 2884 40526 2912 41006
rect 3424 40588 3476 40594
rect 3424 40530 3476 40536
rect 2872 40520 2924 40526
rect 2872 40462 2924 40468
rect 2688 39976 2740 39982
rect 2688 39918 2740 39924
rect 1492 39500 1544 39506
rect 1492 39442 1544 39448
rect 1768 38888 1820 38894
rect 1768 38830 1820 38836
rect 1780 36786 1808 38830
rect 2700 38758 2728 39918
rect 3056 38888 3108 38894
rect 3056 38830 3108 38836
rect 2688 38752 2740 38758
rect 2688 38694 2740 38700
rect 3068 38554 3096 38830
rect 3056 38548 3108 38554
rect 3056 38490 3108 38496
rect 1768 36780 1820 36786
rect 1768 36722 1820 36728
rect 2044 36712 2096 36718
rect 2044 36654 2096 36660
rect 2056 36378 2084 36654
rect 2044 36372 2096 36378
rect 2044 36314 2096 36320
rect 3436 36242 3464 40530
rect 3620 39098 3648 41074
rect 5368 41070 5396 43982
rect 9034 43893 9090 44693
rect 12898 43893 12954 44693
rect 16118 43893 16174 44693
rect 19982 43893 20038 44693
rect 23846 43893 23902 44693
rect 27710 44010 27766 44693
rect 27632 43982 27766 44010
rect 9048 42294 9076 43893
rect 9036 42288 9088 42294
rect 9036 42230 9088 42236
rect 9312 42016 9364 42022
rect 9312 41958 9364 41964
rect 4068 41064 4120 41070
rect 4068 41006 4120 41012
rect 5356 41064 5408 41070
rect 5356 41006 5408 41012
rect 4080 40730 4108 41006
rect 5264 40928 5316 40934
rect 5264 40870 5316 40876
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4068 40724 4120 40730
rect 4068 40666 4120 40672
rect 4620 40520 4672 40526
rect 4620 40462 4672 40468
rect 4632 40390 4660 40462
rect 4620 40384 4672 40390
rect 4620 40326 4672 40332
rect 4804 40384 4856 40390
rect 4804 40326 4856 40332
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4068 39500 4120 39506
rect 4068 39442 4120 39448
rect 4080 39098 4108 39442
rect 4620 39296 4672 39302
rect 4620 39238 4672 39244
rect 3608 39092 3660 39098
rect 3608 39034 3660 39040
rect 4068 39092 4120 39098
rect 4068 39034 4120 39040
rect 3790 38856 3846 38865
rect 3790 38791 3846 38800
rect 3804 36854 3832 38791
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4632 38350 4660 39238
rect 4712 39024 4764 39030
rect 4712 38966 4764 38972
rect 4724 38554 4752 38966
rect 4712 38548 4764 38554
rect 4712 38490 4764 38496
rect 4620 38344 4672 38350
rect 4620 38286 4672 38292
rect 4620 38208 4672 38214
rect 4620 38150 4672 38156
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 3792 36848 3844 36854
rect 3792 36790 3844 36796
rect 3424 36236 3476 36242
rect 3424 36178 3476 36184
rect 1030 34776 1086 34785
rect 1030 34711 1032 34720
rect 1084 34711 1086 34720
rect 1032 34682 1084 34688
rect 1858 34640 1914 34649
rect 1858 34575 1860 34584
rect 1912 34575 1914 34584
rect 1860 34546 1912 34552
rect 2964 31816 3016 31822
rect 2964 31758 3016 31764
rect 2780 31680 2832 31686
rect 2780 31622 2832 31628
rect 2792 31414 2820 31622
rect 2780 31408 2832 31414
rect 2780 31350 2832 31356
rect 2044 31340 2096 31346
rect 2044 31282 2096 31288
rect 1768 31136 1820 31142
rect 1768 31078 1820 31084
rect 1780 30802 1808 31078
rect 1768 30796 1820 30802
rect 1768 30738 1820 30744
rect 1400 30728 1452 30734
rect 1400 30670 1452 30676
rect 1412 28558 1440 30670
rect 2056 30394 2084 31282
rect 2976 30938 3004 31758
rect 3056 31408 3108 31414
rect 3056 31350 3108 31356
rect 2964 30932 3016 30938
rect 2964 30874 3016 30880
rect 3068 30734 3096 31350
rect 3436 30818 3464 36178
rect 3804 36106 3832 36790
rect 4068 36576 4120 36582
rect 4068 36518 4120 36524
rect 4080 36378 4108 36518
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4068 36372 4120 36378
rect 4068 36314 4120 36320
rect 3792 36100 3844 36106
rect 3792 36042 3844 36048
rect 4160 36100 4212 36106
rect 4160 36042 4212 36048
rect 3976 36032 4028 36038
rect 4028 35980 4108 35986
rect 3976 35974 4108 35980
rect 3988 35958 4108 35974
rect 4080 35086 4108 35958
rect 4172 35834 4200 36042
rect 4160 35828 4212 35834
rect 4160 35770 4212 35776
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4068 35080 4120 35086
rect 4068 35022 4120 35028
rect 4080 34066 4108 35022
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4068 34060 4120 34066
rect 4068 34002 4120 34008
rect 4436 33992 4488 33998
rect 4436 33934 4488 33940
rect 4448 33522 4476 33934
rect 4528 33856 4580 33862
rect 4528 33798 4580 33804
rect 4436 33516 4488 33522
rect 4436 33458 4488 33464
rect 4540 33318 4568 33798
rect 4528 33312 4580 33318
rect 4528 33254 4580 33260
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 3700 31272 3752 31278
rect 3700 31214 3752 31220
rect 3344 30802 3464 30818
rect 3344 30796 3476 30802
rect 3344 30790 3424 30796
rect 3056 30728 3108 30734
rect 2778 30696 2834 30705
rect 3056 30670 3108 30676
rect 2964 30660 3016 30666
rect 2834 30640 2964 30648
rect 2778 30631 2964 30640
rect 2792 30620 2964 30631
rect 2792 30394 2820 30620
rect 2964 30602 3016 30608
rect 2044 30388 2096 30394
rect 2044 30330 2096 30336
rect 2780 30388 2832 30394
rect 2780 30330 2832 30336
rect 2872 30184 2924 30190
rect 2872 30126 2924 30132
rect 2884 29850 2912 30126
rect 2872 29844 2924 29850
rect 2872 29786 2924 29792
rect 2688 29640 2740 29646
rect 2688 29582 2740 29588
rect 2504 29504 2556 29510
rect 2504 29446 2556 29452
rect 1860 28960 1912 28966
rect 1860 28902 1912 28908
rect 1400 28552 1452 28558
rect 1400 28494 1452 28500
rect 1412 28082 1440 28494
rect 1872 28218 1900 28902
rect 2516 28626 2544 29446
rect 2700 29306 2728 29582
rect 2688 29300 2740 29306
rect 2688 29242 2740 29248
rect 3068 28626 3096 30670
rect 3344 30190 3372 30790
rect 3424 30738 3476 30744
rect 3712 30598 3740 31214
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4068 30660 4120 30666
rect 4068 30602 4120 30608
rect 3700 30592 3752 30598
rect 3700 30534 3752 30540
rect 3332 30184 3384 30190
rect 3332 30126 3384 30132
rect 3240 29164 3292 29170
rect 3240 29106 3292 29112
rect 3252 28914 3280 29106
rect 3344 29034 3372 30126
rect 3608 29232 3660 29238
rect 3422 29200 3478 29209
rect 3608 29174 3660 29180
rect 3422 29135 3424 29144
rect 3476 29135 3478 29144
rect 3424 29106 3476 29112
rect 3332 29028 3384 29034
rect 3332 28970 3384 28976
rect 3252 28886 3372 28914
rect 2504 28620 2556 28626
rect 2504 28562 2556 28568
rect 3056 28620 3108 28626
rect 3056 28562 3108 28568
rect 1860 28212 1912 28218
rect 1860 28154 1912 28160
rect 3068 28150 3096 28562
rect 3056 28144 3108 28150
rect 3056 28086 3108 28092
rect 1400 28076 1452 28082
rect 1400 28018 1452 28024
rect 1412 26926 1440 28018
rect 3068 27062 3096 28086
rect 3344 28014 3372 28886
rect 3620 28490 3648 29174
rect 3608 28484 3660 28490
rect 3608 28426 3660 28432
rect 3332 28008 3384 28014
rect 3332 27950 3384 27956
rect 3056 27056 3108 27062
rect 3056 26998 3108 27004
rect 1400 26920 1452 26926
rect 1400 26862 1452 26868
rect 1768 26920 1820 26926
rect 1768 26862 1820 26868
rect 1780 26586 1808 26862
rect 2872 26852 2924 26858
rect 2872 26794 2924 26800
rect 2412 26784 2464 26790
rect 2412 26726 2464 26732
rect 1768 26580 1820 26586
rect 1768 26522 1820 26528
rect 2424 25974 2452 26726
rect 2412 25968 2464 25974
rect 2412 25910 2464 25916
rect 2424 25362 2452 25910
rect 2412 25356 2464 25362
rect 2412 25298 2464 25304
rect 1676 25220 1728 25226
rect 1676 25162 1728 25168
rect 1688 24954 1716 25162
rect 1676 24948 1728 24954
rect 1676 24890 1728 24896
rect 2424 23662 2452 25298
rect 2884 24954 2912 26794
rect 2964 25900 3016 25906
rect 2964 25842 3016 25848
rect 2872 24948 2924 24954
rect 2872 24890 2924 24896
rect 2780 24064 2832 24070
rect 2780 24006 2832 24012
rect 2792 23866 2820 24006
rect 2780 23860 2832 23866
rect 2780 23802 2832 23808
rect 2412 23656 2464 23662
rect 2412 23598 2464 23604
rect 2424 23186 2452 23598
rect 2412 23180 2464 23186
rect 2412 23122 2464 23128
rect 1676 23044 1728 23050
rect 1676 22986 1728 22992
rect 1688 22778 1716 22986
rect 2884 22778 2912 24890
rect 1676 22772 1728 22778
rect 1676 22714 1728 22720
rect 2872 22772 2924 22778
rect 2872 22714 2924 22720
rect 2884 22094 2912 22714
rect 2792 22066 2912 22094
rect 2504 21888 2556 21894
rect 2504 21830 2556 21836
rect 2516 21690 2544 21830
rect 2504 21684 2556 21690
rect 2504 21626 2556 21632
rect 2688 21480 2740 21486
rect 2688 21422 2740 21428
rect 2700 21350 2728 21422
rect 1860 21344 1912 21350
rect 1860 21286 1912 21292
rect 2688 21344 2740 21350
rect 2688 21286 2740 21292
rect 1872 21146 1900 21286
rect 1860 21140 1912 21146
rect 1860 21082 1912 21088
rect 2700 21010 2728 21286
rect 1400 21004 1452 21010
rect 1400 20946 1452 20952
rect 2688 21004 2740 21010
rect 2688 20946 2740 20952
rect 1412 19922 1440 20946
rect 2596 20460 2648 20466
rect 2596 20402 2648 20408
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 1676 19780 1728 19786
rect 1676 19722 1728 19728
rect 1688 19514 1716 19722
rect 2608 19514 2636 20402
rect 2700 20398 2728 20946
rect 2688 20392 2740 20398
rect 2688 20334 2740 20340
rect 1676 19508 1728 19514
rect 1676 19450 1728 19456
rect 2596 19508 2648 19514
rect 2596 19450 2648 19456
rect 2792 19378 2820 22066
rect 2872 21888 2924 21894
rect 2872 21830 2924 21836
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 2504 18080 2556 18086
rect 2504 18022 2556 18028
rect 1676 17604 1728 17610
rect 1676 17546 1728 17552
rect 1688 17338 1716 17546
rect 2516 17338 2544 18022
rect 1676 17332 1728 17338
rect 1676 17274 1728 17280
rect 2504 17332 2556 17338
rect 2504 17274 2556 17280
rect 2136 16992 2188 16998
rect 2136 16934 2188 16940
rect 2148 16658 2176 16934
rect 2136 16652 2188 16658
rect 2136 16594 2188 16600
rect 2792 15366 2820 19314
rect 2884 19258 2912 21830
rect 2976 20534 3004 25842
rect 3068 25294 3096 26998
rect 3240 26784 3292 26790
rect 3240 26726 3292 26732
rect 3252 26382 3280 26726
rect 3240 26376 3292 26382
rect 3240 26318 3292 26324
rect 3056 25288 3108 25294
rect 3056 25230 3108 25236
rect 3068 23866 3096 25230
rect 3148 25152 3200 25158
rect 3148 25094 3200 25100
rect 3160 24954 3188 25094
rect 3148 24948 3200 24954
rect 3148 24890 3200 24896
rect 3056 23860 3108 23866
rect 3056 23802 3108 23808
rect 3068 23118 3096 23802
rect 3148 23248 3200 23254
rect 3148 23190 3200 23196
rect 3056 23112 3108 23118
rect 3056 23054 3108 23060
rect 3160 22778 3188 23190
rect 3148 22772 3200 22778
rect 3148 22714 3200 22720
rect 3148 22432 3200 22438
rect 3148 22374 3200 22380
rect 3160 22166 3188 22374
rect 3148 22160 3200 22166
rect 3148 22102 3200 22108
rect 3148 21888 3200 21894
rect 3148 21830 3200 21836
rect 3160 21010 3188 21830
rect 3240 21616 3292 21622
rect 3240 21558 3292 21564
rect 3252 21146 3280 21558
rect 3240 21140 3292 21146
rect 3240 21082 3292 21088
rect 3148 21004 3200 21010
rect 3148 20946 3200 20952
rect 3056 20868 3108 20874
rect 3056 20810 3108 20816
rect 2964 20528 3016 20534
rect 2964 20470 3016 20476
rect 3068 19786 3096 20810
rect 3056 19780 3108 19786
rect 3056 19722 3108 19728
rect 2884 19230 3004 19258
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 2884 18834 2912 19110
rect 2872 18828 2924 18834
rect 2872 18770 2924 18776
rect 2976 18222 3004 19230
rect 3344 19145 3372 27950
rect 3516 26784 3568 26790
rect 3516 26726 3568 26732
rect 3424 26444 3476 26450
rect 3424 26386 3476 26392
rect 3436 25770 3464 26386
rect 3528 26314 3556 26726
rect 3516 26308 3568 26314
rect 3516 26250 3568 26256
rect 3424 25764 3476 25770
rect 3424 25706 3476 25712
rect 3620 23225 3648 28426
rect 3606 23216 3662 23225
rect 3606 23151 3662 23160
rect 3424 20256 3476 20262
rect 3424 20198 3476 20204
rect 3608 20256 3660 20262
rect 3608 20198 3660 20204
rect 3436 19514 3464 20198
rect 3620 20058 3648 20198
rect 3608 20052 3660 20058
rect 3608 19994 3660 20000
rect 3608 19712 3660 19718
rect 3608 19654 3660 19660
rect 3424 19508 3476 19514
rect 3424 19450 3476 19456
rect 3620 19446 3648 19654
rect 3608 19440 3660 19446
rect 3608 19382 3660 19388
rect 3330 19136 3386 19145
rect 3330 19071 3386 19080
rect 2964 18216 3016 18222
rect 2964 18158 3016 18164
rect 3424 18216 3476 18222
rect 3424 18158 3476 18164
rect 2976 17270 3004 18158
rect 3436 17814 3464 18158
rect 3424 17808 3476 17814
rect 3424 17750 3476 17756
rect 3424 17604 3476 17610
rect 3424 17546 3476 17552
rect 2964 17264 3016 17270
rect 2964 17206 3016 17212
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 3344 15570 3372 16934
rect 3436 16522 3464 17546
rect 3712 17218 3740 30534
rect 4080 27305 4108 30602
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4526 29744 4582 29753
rect 4526 29679 4582 29688
rect 4160 29572 4212 29578
rect 4160 29514 4212 29520
rect 4172 29238 4200 29514
rect 4540 29306 4568 29679
rect 4528 29300 4580 29306
rect 4528 29242 4580 29248
rect 4160 29232 4212 29238
rect 4160 29174 4212 29180
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4632 27606 4660 38150
rect 4712 35148 4764 35154
rect 4712 35090 4764 35096
rect 4724 33998 4752 35090
rect 4712 33992 4764 33998
rect 4712 33934 4764 33940
rect 4816 32026 4844 40326
rect 5276 36922 5304 40870
rect 5368 40526 5396 41006
rect 5356 40520 5408 40526
rect 5356 40462 5408 40468
rect 8024 40452 8076 40458
rect 8024 40394 8076 40400
rect 7472 40112 7524 40118
rect 7472 40054 7524 40060
rect 7288 40044 7340 40050
rect 7288 39986 7340 39992
rect 7300 39506 7328 39986
rect 7380 39636 7432 39642
rect 7380 39578 7432 39584
rect 7288 39500 7340 39506
rect 7288 39442 7340 39448
rect 5724 39364 5776 39370
rect 5724 39306 5776 39312
rect 5736 38962 5764 39306
rect 7012 39296 7064 39302
rect 7012 39238 7064 39244
rect 7024 38962 7052 39238
rect 7300 39098 7328 39442
rect 7288 39092 7340 39098
rect 7288 39034 7340 39040
rect 5724 38956 5776 38962
rect 5724 38898 5776 38904
rect 7012 38956 7064 38962
rect 7012 38898 7064 38904
rect 5356 38412 5408 38418
rect 5356 38354 5408 38360
rect 5264 36916 5316 36922
rect 5264 36858 5316 36864
rect 5080 35692 5132 35698
rect 5080 35634 5132 35640
rect 4988 34468 5040 34474
rect 4988 34410 5040 34416
rect 5000 33998 5028 34410
rect 5092 34202 5120 35634
rect 5368 35630 5396 38354
rect 5540 38208 5592 38214
rect 5540 38150 5592 38156
rect 5552 37194 5580 38150
rect 5540 37188 5592 37194
rect 5540 37130 5592 37136
rect 5736 36786 5764 38898
rect 6460 38888 6512 38894
rect 6460 38830 6512 38836
rect 6472 38214 6500 38830
rect 6736 38752 6788 38758
rect 6736 38694 6788 38700
rect 6748 38554 6776 38694
rect 6552 38548 6604 38554
rect 6552 38490 6604 38496
rect 6736 38548 6788 38554
rect 6736 38490 6788 38496
rect 6460 38208 6512 38214
rect 6460 38150 6512 38156
rect 6472 37874 6500 38150
rect 6276 37868 6328 37874
rect 6276 37810 6328 37816
rect 6460 37868 6512 37874
rect 6460 37810 6512 37816
rect 5724 36780 5776 36786
rect 5724 36722 5776 36728
rect 5736 36310 5764 36722
rect 6092 36576 6144 36582
rect 6092 36518 6144 36524
rect 5724 36304 5776 36310
rect 5724 36246 5776 36252
rect 6104 36174 6132 36518
rect 6092 36168 6144 36174
rect 6092 36110 6144 36116
rect 5540 36032 5592 36038
rect 5540 35974 5592 35980
rect 5552 35698 5580 35974
rect 5540 35692 5592 35698
rect 5540 35634 5592 35640
rect 5356 35624 5408 35630
rect 5356 35566 5408 35572
rect 6184 34468 6236 34474
rect 6184 34410 6236 34416
rect 5080 34196 5132 34202
rect 5080 34138 5132 34144
rect 5264 34128 5316 34134
rect 5816 34128 5868 34134
rect 5316 34076 5764 34082
rect 5264 34070 5764 34076
rect 5816 34070 5868 34076
rect 5276 34054 5764 34070
rect 5736 33998 5764 34054
rect 4988 33992 5040 33998
rect 4988 33934 5040 33940
rect 5724 33992 5776 33998
rect 5724 33934 5776 33940
rect 4896 33924 4948 33930
rect 4896 33866 4948 33872
rect 5264 33924 5316 33930
rect 5264 33866 5316 33872
rect 4908 33522 4936 33866
rect 5276 33522 5304 33866
rect 4896 33516 4948 33522
rect 4896 33458 4948 33464
rect 5264 33516 5316 33522
rect 5264 33458 5316 33464
rect 4988 33312 5040 33318
rect 4988 33254 5040 33260
rect 5000 32502 5028 33254
rect 4988 32496 5040 32502
rect 4988 32438 5040 32444
rect 4896 32224 4948 32230
rect 4896 32166 4948 32172
rect 4908 32026 4936 32166
rect 4804 32020 4856 32026
rect 4804 31962 4856 31968
rect 4896 32020 4948 32026
rect 4896 31962 4948 31968
rect 4908 31346 4936 31962
rect 5000 31822 5028 32438
rect 5080 32360 5132 32366
rect 5080 32302 5132 32308
rect 4988 31816 5040 31822
rect 4988 31758 5040 31764
rect 5000 31346 5028 31758
rect 4896 31340 4948 31346
rect 4896 31282 4948 31288
rect 4988 31340 5040 31346
rect 4988 31282 5040 31288
rect 5092 31142 5120 32302
rect 5080 31136 5132 31142
rect 5080 31078 5132 31084
rect 5092 30802 5120 31078
rect 5080 30796 5132 30802
rect 5080 30738 5132 30744
rect 4804 30252 4856 30258
rect 4804 30194 4856 30200
rect 4816 29578 4844 30194
rect 4896 30116 4948 30122
rect 4896 30058 4948 30064
rect 4804 29572 4856 29578
rect 4804 29514 4856 29520
rect 4816 28626 4844 29514
rect 4908 29238 4936 30058
rect 5080 30048 5132 30054
rect 5080 29990 5132 29996
rect 4988 29776 5040 29782
rect 4988 29718 5040 29724
rect 4896 29232 4948 29238
rect 4896 29174 4948 29180
rect 4804 28620 4856 28626
rect 4804 28562 4856 28568
rect 5000 28082 5028 29718
rect 5092 29170 5120 29990
rect 5276 29850 5304 33458
rect 5828 33386 5856 34070
rect 5908 33924 5960 33930
rect 5908 33866 5960 33872
rect 5920 33590 5948 33866
rect 5908 33584 5960 33590
rect 5908 33526 5960 33532
rect 5816 33380 5868 33386
rect 5816 33322 5868 33328
rect 5724 32564 5776 32570
rect 5724 32506 5776 32512
rect 5356 31884 5408 31890
rect 5356 31826 5408 31832
rect 5368 31754 5396 31826
rect 5736 31822 5764 32506
rect 6092 32496 6144 32502
rect 6092 32438 6144 32444
rect 6000 32428 6052 32434
rect 6000 32370 6052 32376
rect 5908 32224 5960 32230
rect 5908 32166 5960 32172
rect 5920 31958 5948 32166
rect 6012 32026 6040 32370
rect 6104 32026 6132 32438
rect 6196 32434 6224 34410
rect 6288 33522 6316 37810
rect 6564 37466 6592 38490
rect 6748 38418 6776 38490
rect 6736 38412 6788 38418
rect 6736 38354 6788 38360
rect 6828 38412 6880 38418
rect 6828 38354 6880 38360
rect 6644 38344 6696 38350
rect 6644 38286 6696 38292
rect 6656 38010 6684 38286
rect 6644 38004 6696 38010
rect 6644 37946 6696 37952
rect 6748 37874 6776 38354
rect 6840 38214 6868 38354
rect 7288 38344 7340 38350
rect 7288 38286 7340 38292
rect 6828 38208 6880 38214
rect 6828 38150 6880 38156
rect 6736 37868 6788 37874
rect 6736 37810 6788 37816
rect 7012 37868 7064 37874
rect 7012 37810 7064 37816
rect 6736 37664 6788 37670
rect 6736 37606 6788 37612
rect 6748 37466 6776 37606
rect 6552 37460 6604 37466
rect 6552 37402 6604 37408
rect 6736 37460 6788 37466
rect 6736 37402 6788 37408
rect 6748 36786 6776 37402
rect 6920 37324 6972 37330
rect 6920 37266 6972 37272
rect 6932 36922 6960 37266
rect 6920 36916 6972 36922
rect 6920 36858 6972 36864
rect 6368 36780 6420 36786
rect 6368 36722 6420 36728
rect 6736 36780 6788 36786
rect 6736 36722 6788 36728
rect 6276 33516 6328 33522
rect 6276 33458 6328 33464
rect 6184 32428 6236 32434
rect 6184 32370 6236 32376
rect 6000 32020 6052 32026
rect 6000 31962 6052 31968
rect 6092 32020 6144 32026
rect 6092 31962 6144 31968
rect 5908 31952 5960 31958
rect 6196 31906 6224 32370
rect 6288 32366 6316 33458
rect 6276 32360 6328 32366
rect 6276 32302 6328 32308
rect 5908 31894 5960 31900
rect 6012 31878 6224 31906
rect 6012 31822 6040 31878
rect 5724 31816 5776 31822
rect 5724 31758 5776 31764
rect 6000 31816 6052 31822
rect 6000 31758 6052 31764
rect 6184 31816 6236 31822
rect 6184 31758 6236 31764
rect 5368 31726 5580 31754
rect 5264 29844 5316 29850
rect 5264 29786 5316 29792
rect 5356 29640 5408 29646
rect 5356 29582 5408 29588
rect 5368 29306 5396 29582
rect 5448 29504 5500 29510
rect 5448 29446 5500 29452
rect 5356 29300 5408 29306
rect 5356 29242 5408 29248
rect 5460 29186 5488 29446
rect 5552 29306 5580 31726
rect 6196 31210 6224 31758
rect 6184 31204 6236 31210
rect 6184 31146 6236 31152
rect 6184 30048 6236 30054
rect 6184 29990 6236 29996
rect 6196 29646 6224 29990
rect 5816 29640 5868 29646
rect 5816 29582 5868 29588
rect 6184 29640 6236 29646
rect 6184 29582 6236 29588
rect 5632 29572 5684 29578
rect 5632 29514 5684 29520
rect 5540 29300 5592 29306
rect 5540 29242 5592 29248
rect 5080 29164 5132 29170
rect 5080 29106 5132 29112
rect 5172 29164 5224 29170
rect 5172 29106 5224 29112
rect 5264 29164 5316 29170
rect 5264 29106 5316 29112
rect 5356 29164 5408 29170
rect 5460 29158 5580 29186
rect 5644 29170 5672 29514
rect 5828 29170 5856 29582
rect 5908 29232 5960 29238
rect 5908 29174 5960 29180
rect 5356 29106 5408 29112
rect 4988 28076 5040 28082
rect 4988 28018 5040 28024
rect 4712 27872 4764 27878
rect 4712 27814 4764 27820
rect 4620 27600 4672 27606
rect 4620 27542 4672 27548
rect 4066 27296 4122 27305
rect 4066 27231 4122 27240
rect 3884 27056 3936 27062
rect 3884 26998 3936 27004
rect 3792 26376 3844 26382
rect 3792 26318 3844 26324
rect 3804 25974 3832 26318
rect 3896 26246 3924 26998
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4620 26444 4672 26450
rect 4620 26386 4672 26392
rect 3976 26308 4028 26314
rect 3976 26250 4028 26256
rect 3884 26240 3936 26246
rect 3884 26182 3936 26188
rect 3792 25968 3844 25974
rect 3792 25910 3844 25916
rect 3884 25764 3936 25770
rect 3884 25706 3936 25712
rect 3896 24750 3924 25706
rect 3988 25498 4016 26250
rect 4068 25696 4120 25702
rect 4068 25638 4120 25644
rect 4080 25498 4108 25638
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 3976 25492 4028 25498
rect 3976 25434 4028 25440
rect 4068 25492 4120 25498
rect 4068 25434 4120 25440
rect 4068 25152 4120 25158
rect 4068 25094 4120 25100
rect 3976 24812 4028 24818
rect 3976 24754 4028 24760
rect 3884 24744 3936 24750
rect 3884 24686 3936 24692
rect 3896 24274 3924 24686
rect 3884 24268 3936 24274
rect 3884 24210 3936 24216
rect 3988 20058 4016 24754
rect 4080 23866 4108 25094
rect 4632 24682 4660 26386
rect 4620 24676 4672 24682
rect 4620 24618 4672 24624
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4724 24206 4752 27814
rect 5092 27402 5120 29106
rect 5184 28937 5212 29106
rect 5170 28928 5226 28937
rect 5170 28863 5226 28872
rect 5184 28558 5212 28863
rect 5172 28552 5224 28558
rect 5172 28494 5224 28500
rect 5276 28490 5304 29106
rect 5368 28762 5396 29106
rect 5552 29050 5580 29158
rect 5632 29164 5684 29170
rect 5632 29106 5684 29112
rect 5816 29164 5868 29170
rect 5816 29106 5868 29112
rect 5552 29022 5672 29050
rect 5356 28756 5408 28762
rect 5356 28698 5408 28704
rect 5540 28688 5592 28694
rect 5540 28630 5592 28636
rect 5264 28484 5316 28490
rect 5264 28426 5316 28432
rect 5448 28212 5500 28218
rect 5448 28154 5500 28160
rect 5356 28076 5408 28082
rect 5356 28018 5408 28024
rect 5368 27402 5396 28018
rect 4896 27396 4948 27402
rect 4896 27338 4948 27344
rect 5080 27396 5132 27402
rect 5080 27338 5132 27344
rect 5356 27396 5408 27402
rect 5356 27338 5408 27344
rect 4804 26784 4856 26790
rect 4804 26726 4856 26732
rect 4816 24290 4844 26726
rect 4908 24410 4936 27338
rect 5460 25906 5488 28154
rect 5552 27130 5580 28630
rect 5644 27962 5672 29022
rect 5724 29028 5776 29034
rect 5724 28970 5776 28976
rect 5816 29028 5868 29034
rect 5816 28970 5868 28976
rect 5736 28150 5764 28970
rect 5828 28762 5856 28970
rect 5816 28756 5868 28762
rect 5816 28698 5868 28704
rect 5920 28558 5948 29174
rect 6276 29164 6328 29170
rect 6276 29106 6328 29112
rect 6288 28937 6316 29106
rect 6380 28994 6408 36722
rect 6932 36582 6960 36858
rect 6460 36576 6512 36582
rect 6460 36518 6512 36524
rect 6920 36576 6972 36582
rect 6920 36518 6972 36524
rect 6472 35698 6500 36518
rect 6932 36378 6960 36518
rect 6920 36372 6972 36378
rect 6920 36314 6972 36320
rect 7024 36242 7052 37810
rect 7104 37664 7156 37670
rect 7104 37606 7156 37612
rect 7116 37262 7144 37606
rect 7300 37466 7328 38286
rect 7288 37460 7340 37466
rect 7288 37402 7340 37408
rect 7104 37256 7156 37262
rect 7104 37198 7156 37204
rect 7116 36786 7144 37198
rect 7196 37120 7248 37126
rect 7196 37062 7248 37068
rect 7104 36780 7156 36786
rect 7104 36722 7156 36728
rect 7208 36718 7236 37062
rect 7288 36916 7340 36922
rect 7288 36858 7340 36864
rect 7300 36786 7328 36858
rect 7288 36780 7340 36786
rect 7288 36722 7340 36728
rect 7392 36718 7420 39578
rect 7196 36712 7248 36718
rect 7196 36654 7248 36660
rect 7380 36712 7432 36718
rect 7380 36654 7432 36660
rect 7012 36236 7064 36242
rect 7012 36178 7064 36184
rect 7024 35698 7052 36178
rect 6460 35692 6512 35698
rect 6460 35634 6512 35640
rect 7012 35692 7064 35698
rect 7012 35634 7064 35640
rect 6552 35624 6604 35630
rect 6552 35566 6604 35572
rect 6564 34678 6592 35566
rect 6828 35488 6880 35494
rect 6828 35430 6880 35436
rect 6552 34672 6604 34678
rect 6552 34614 6604 34620
rect 6840 34490 6868 35430
rect 6920 34604 6972 34610
rect 7024 34592 7052 35634
rect 7392 35170 7420 36654
rect 6972 34564 7052 34592
rect 7116 35142 7420 35170
rect 6920 34546 6972 34552
rect 6748 34462 7052 34490
rect 6748 33590 6776 34462
rect 6920 34400 6972 34406
rect 6920 34342 6972 34348
rect 6932 34134 6960 34342
rect 6920 34128 6972 34134
rect 6920 34070 6972 34076
rect 6828 33992 6880 33998
rect 6932 33980 6960 34070
rect 7024 33998 7052 34462
rect 6880 33952 6960 33980
rect 7012 33992 7064 33998
rect 6828 33934 6880 33940
rect 7012 33934 7064 33940
rect 6840 33658 6868 33934
rect 6920 33856 6972 33862
rect 6920 33798 6972 33804
rect 6932 33658 6960 33798
rect 6828 33652 6880 33658
rect 6828 33594 6880 33600
rect 6920 33652 6972 33658
rect 6920 33594 6972 33600
rect 6736 33584 6788 33590
rect 6736 33526 6788 33532
rect 7116 33046 7144 35142
rect 7288 35080 7340 35086
rect 7288 35022 7340 35028
rect 7300 33946 7328 35022
rect 7380 34400 7432 34406
rect 7380 34342 7432 34348
rect 7392 34066 7420 34342
rect 7380 34060 7432 34066
rect 7380 34002 7432 34008
rect 7300 33918 7420 33946
rect 7196 33856 7248 33862
rect 7196 33798 7248 33804
rect 7104 33040 7156 33046
rect 7104 32982 7156 32988
rect 6828 32564 6880 32570
rect 6828 32506 6880 32512
rect 6920 32564 6972 32570
rect 6920 32506 6972 32512
rect 6840 32230 6868 32506
rect 6644 32224 6696 32230
rect 6644 32166 6696 32172
rect 6828 32224 6880 32230
rect 6828 32166 6880 32172
rect 6656 31890 6684 32166
rect 6644 31884 6696 31890
rect 6644 31826 6696 31832
rect 6932 31822 6960 32506
rect 7116 31822 7144 32982
rect 7208 32910 7236 33798
rect 7288 33108 7340 33114
rect 7288 33050 7340 33056
rect 7196 32904 7248 32910
rect 7196 32846 7248 32852
rect 7208 32026 7236 32846
rect 7300 32570 7328 33050
rect 7288 32564 7340 32570
rect 7288 32506 7340 32512
rect 7196 32020 7248 32026
rect 7196 31962 7248 31968
rect 6920 31816 6972 31822
rect 6920 31758 6972 31764
rect 7104 31816 7156 31822
rect 7104 31758 7156 31764
rect 7196 31408 7248 31414
rect 7196 31350 7248 31356
rect 7208 31226 7236 31350
rect 7208 31198 7328 31226
rect 7300 31142 7328 31198
rect 6736 31136 6788 31142
rect 6736 31078 6788 31084
rect 7288 31136 7340 31142
rect 7288 31078 7340 31084
rect 6552 30116 6604 30122
rect 6552 30058 6604 30064
rect 6460 30048 6512 30054
rect 6460 29990 6512 29996
rect 6472 29646 6500 29990
rect 6460 29640 6512 29646
rect 6460 29582 6512 29588
rect 6564 29510 6592 30058
rect 6748 29850 6776 31078
rect 6736 29844 6788 29850
rect 6736 29786 6788 29792
rect 7012 29776 7064 29782
rect 7012 29718 7064 29724
rect 6736 29708 6788 29714
rect 6736 29650 6788 29656
rect 6552 29504 6604 29510
rect 6552 29446 6604 29452
rect 6564 29170 6592 29446
rect 6748 29170 6776 29650
rect 7024 29578 7052 29718
rect 7104 29640 7156 29646
rect 7102 29608 7104 29617
rect 7196 29640 7248 29646
rect 7156 29608 7158 29617
rect 7012 29572 7064 29578
rect 7196 29582 7248 29588
rect 7102 29543 7158 29552
rect 7012 29514 7064 29520
rect 7116 29306 7144 29543
rect 7104 29300 7156 29306
rect 7104 29242 7156 29248
rect 6552 29164 6604 29170
rect 6552 29106 6604 29112
rect 6644 29164 6696 29170
rect 6644 29106 6696 29112
rect 6736 29164 6788 29170
rect 6736 29106 6788 29112
rect 6380 28966 6500 28994
rect 6274 28928 6330 28937
rect 6274 28863 6330 28872
rect 5908 28552 5960 28558
rect 5828 28500 5908 28506
rect 5828 28494 5960 28500
rect 5828 28478 5948 28494
rect 5724 28144 5776 28150
rect 5724 28086 5776 28092
rect 5644 27934 5764 27962
rect 5632 27464 5684 27470
rect 5632 27406 5684 27412
rect 5540 27124 5592 27130
rect 5540 27066 5592 27072
rect 5540 26580 5592 26586
rect 5540 26522 5592 26528
rect 5552 26042 5580 26522
rect 5540 26036 5592 26042
rect 5540 25978 5592 25984
rect 5448 25900 5500 25906
rect 5448 25842 5500 25848
rect 5080 24948 5132 24954
rect 5132 24908 5396 24936
rect 5080 24890 5132 24896
rect 5078 24848 5134 24857
rect 5078 24783 5080 24792
rect 5132 24783 5134 24792
rect 5172 24812 5224 24818
rect 5080 24754 5132 24760
rect 5172 24754 5224 24760
rect 4986 24712 5042 24721
rect 4986 24647 5042 24656
rect 5000 24410 5028 24647
rect 5092 24410 5120 24754
rect 5184 24682 5212 24754
rect 5264 24744 5316 24750
rect 5262 24712 5264 24721
rect 5316 24712 5318 24721
rect 5172 24676 5224 24682
rect 5262 24647 5318 24656
rect 5172 24618 5224 24624
rect 4896 24404 4948 24410
rect 4896 24346 4948 24352
rect 4988 24404 5040 24410
rect 4988 24346 5040 24352
rect 5080 24404 5132 24410
rect 5080 24346 5132 24352
rect 4816 24262 5212 24290
rect 4712 24200 4764 24206
rect 4712 24142 4764 24148
rect 4252 24064 4304 24070
rect 4252 24006 4304 24012
rect 4068 23860 4120 23866
rect 4068 23802 4120 23808
rect 4264 23798 4292 24006
rect 4252 23792 4304 23798
rect 4252 23734 4304 23740
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4160 22568 4212 22574
rect 4160 22510 4212 22516
rect 4528 22568 4580 22574
rect 4528 22510 4580 22516
rect 4172 22420 4200 22510
rect 4080 22392 4200 22420
rect 4540 22420 4568 22510
rect 4540 22392 4660 22420
rect 4080 22148 4108 22392
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 22234 4660 22392
rect 4620 22228 4672 22234
rect 4620 22170 4672 22176
rect 4080 22120 4200 22148
rect 4068 21412 4120 21418
rect 4068 21354 4120 21360
rect 4080 21010 4108 21354
rect 4172 21350 4200 22120
rect 4724 22094 4752 24142
rect 5080 23316 5132 23322
rect 5080 23258 5132 23264
rect 5092 23118 5120 23258
rect 5080 23112 5132 23118
rect 5080 23054 5132 23060
rect 4804 22976 4856 22982
rect 5092 22953 5120 23054
rect 4804 22918 4856 22924
rect 5078 22944 5134 22953
rect 4632 22066 4752 22094
rect 4632 21962 4660 22066
rect 4620 21956 4672 21962
rect 4620 21898 4672 21904
rect 4160 21344 4212 21350
rect 4160 21286 4212 21292
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 4816 20890 4844 22918
rect 5078 22879 5134 22888
rect 4988 21888 5040 21894
rect 4988 21830 5040 21836
rect 4632 20862 4844 20890
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3976 20052 4028 20058
rect 3976 19994 4028 20000
rect 3792 19984 3844 19990
rect 4632 19938 4660 20862
rect 4712 20800 4764 20806
rect 4712 20742 4764 20748
rect 3792 19926 3844 19932
rect 3620 17190 3740 17218
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3424 16516 3476 16522
rect 3424 16458 3476 16464
rect 3528 16114 3556 16730
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 3528 15570 3556 16050
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 3516 15564 3568 15570
rect 3516 15506 3568 15512
rect 3240 15428 3292 15434
rect 3240 15370 3292 15376
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 2044 15360 2096 15366
rect 2044 15302 2096 15308
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 1596 15201 1624 15302
rect 1582 15192 1638 15201
rect 2056 15162 2084 15302
rect 1582 15127 1638 15136
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 3148 15088 3200 15094
rect 3148 15030 3200 15036
rect 1584 14816 1636 14822
rect 1584 14758 1636 14764
rect 1596 14074 1624 14758
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1768 13864 1820 13870
rect 1768 13806 1820 13812
rect 1780 13530 1808 13806
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 2792 13326 2820 14214
rect 3160 14006 3188 15030
rect 3252 14482 3280 15370
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 3252 14006 3280 14418
rect 3528 14074 3556 15506
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3148 14000 3200 14006
rect 3148 13942 3200 13948
rect 3240 14000 3292 14006
rect 3240 13942 3292 13948
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 940 11756 992 11762
rect 940 11698 992 11704
rect 952 11665 980 11698
rect 1676 11688 1728 11694
rect 938 11656 994 11665
rect 1676 11630 1728 11636
rect 938 11591 994 11600
rect 1688 11354 1716 11630
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 940 7812 992 7818
rect 940 7754 992 7760
rect 952 7585 980 7754
rect 938 7576 994 7585
rect 938 7511 994 7520
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 1872 4690 1900 6734
rect 1860 4684 1912 4690
rect 1860 4626 1912 4632
rect 2136 4548 2188 4554
rect 2136 4490 2188 4496
rect 2148 4282 2176 4490
rect 2136 4276 2188 4282
rect 2136 4218 2188 4224
rect 940 4140 992 4146
rect 940 4082 992 4088
rect 20 3528 72 3534
rect 952 3505 980 4082
rect 3620 3534 3648 17190
rect 3804 16130 3832 19926
rect 4264 19910 4660 19938
rect 4264 19854 4292 19910
rect 3976 19848 4028 19854
rect 3976 19790 4028 19796
rect 4252 19848 4304 19854
rect 4252 19790 4304 19796
rect 3884 19168 3936 19174
rect 3884 19110 3936 19116
rect 3896 17134 3924 19110
rect 3988 18970 4016 19790
rect 4436 19780 4488 19786
rect 4436 19722 4488 19728
rect 4448 19378 4476 19722
rect 4620 19508 4672 19514
rect 4724 19496 4752 20742
rect 5000 20618 5028 21830
rect 5184 21706 5212 24262
rect 5368 24206 5396 24908
rect 5356 24200 5408 24206
rect 5356 24142 5408 24148
rect 5264 24132 5316 24138
rect 5264 24074 5316 24080
rect 5276 23798 5304 24074
rect 5460 24052 5488 25842
rect 5644 24954 5672 27406
rect 5736 26296 5764 27934
rect 5828 27470 5856 28478
rect 5908 28416 5960 28422
rect 5908 28358 5960 28364
rect 6184 28416 6236 28422
rect 6184 28358 6236 28364
rect 5816 27464 5868 27470
rect 5816 27406 5868 27412
rect 5920 27062 5948 28358
rect 6196 28218 6224 28358
rect 6184 28212 6236 28218
rect 6184 28154 6236 28160
rect 6092 28008 6144 28014
rect 6092 27950 6144 27956
rect 6000 27600 6052 27606
rect 6000 27542 6052 27548
rect 6012 27470 6040 27542
rect 6000 27464 6052 27470
rect 6000 27406 6052 27412
rect 6012 27130 6040 27406
rect 6000 27124 6052 27130
rect 6000 27066 6052 27072
rect 5908 27056 5960 27062
rect 5908 26998 5960 27004
rect 6104 26926 6132 27950
rect 6368 27396 6420 27402
rect 6368 27338 6420 27344
rect 6276 27328 6328 27334
rect 6276 27270 6328 27276
rect 6092 26920 6144 26926
rect 6092 26862 6144 26868
rect 5816 26308 5868 26314
rect 5736 26268 5816 26296
rect 5816 26250 5868 26256
rect 5724 25492 5776 25498
rect 5724 25434 5776 25440
rect 5632 24948 5684 24954
rect 5632 24890 5684 24896
rect 5538 24848 5594 24857
rect 5538 24783 5540 24792
rect 5592 24783 5594 24792
rect 5540 24754 5592 24760
rect 5632 24744 5684 24750
rect 5632 24686 5684 24692
rect 5644 24410 5672 24686
rect 5632 24404 5684 24410
rect 5632 24346 5684 24352
rect 5736 24138 5764 25434
rect 5828 24954 5856 26250
rect 5816 24948 5868 24954
rect 5816 24890 5868 24896
rect 5908 24744 5960 24750
rect 5906 24712 5908 24721
rect 5960 24712 5962 24721
rect 5906 24647 5962 24656
rect 5632 24132 5684 24138
rect 5632 24074 5684 24080
rect 5724 24132 5776 24138
rect 5724 24074 5776 24080
rect 5368 24024 5488 24052
rect 5264 23792 5316 23798
rect 5264 23734 5316 23740
rect 5264 23112 5316 23118
rect 5264 23054 5316 23060
rect 5092 21678 5212 21706
rect 5092 20806 5120 21678
rect 5172 21616 5224 21622
rect 5172 21558 5224 21564
rect 5184 20942 5212 21558
rect 5172 20936 5224 20942
rect 5276 20924 5304 23054
rect 5368 21962 5396 24024
rect 5540 23792 5592 23798
rect 5540 23734 5592 23740
rect 5448 22092 5500 22098
rect 5448 22034 5500 22040
rect 5356 21956 5408 21962
rect 5356 21898 5408 21904
rect 5460 21622 5488 22034
rect 5448 21616 5500 21622
rect 5448 21558 5500 21564
rect 5356 20936 5408 20942
rect 5276 20896 5356 20924
rect 5172 20878 5224 20884
rect 5356 20878 5408 20884
rect 5080 20800 5132 20806
rect 5080 20742 5132 20748
rect 5000 20590 5212 20618
rect 4988 20460 5040 20466
rect 4988 20402 5040 20408
rect 4724 19468 4844 19496
rect 4620 19450 4672 19456
rect 4436 19372 4488 19378
rect 4436 19314 4488 19320
rect 4068 19304 4120 19310
rect 4068 19246 4120 19252
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 4080 18290 4108 19246
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4436 18760 4488 18766
rect 4436 18702 4488 18708
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4448 18154 4476 18702
rect 4436 18148 4488 18154
rect 4436 18090 4488 18096
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17746 4660 19450
rect 4710 19408 4766 19417
rect 4710 19343 4712 19352
rect 4764 19343 4766 19352
rect 4712 19314 4764 19320
rect 4816 18630 4844 19468
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 4712 18080 4764 18086
rect 4712 18022 4764 18028
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4724 17542 4752 18022
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 3976 17264 4028 17270
rect 3976 17206 4028 17212
rect 3884 17128 3936 17134
rect 3884 17070 3936 17076
rect 3896 16794 3924 17070
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3712 16102 3832 16130
rect 3712 15502 3740 16102
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 3804 15706 3832 15982
rect 3792 15700 3844 15706
rect 3792 15642 3844 15648
rect 3700 15496 3752 15502
rect 3700 15438 3752 15444
rect 3712 15162 3740 15438
rect 3988 15162 4016 17206
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 4080 16794 4108 16934
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4816 16658 4844 18566
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4080 15586 4108 16390
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4080 15558 4200 15586
rect 4172 15502 4200 15558
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 3700 15156 3752 15162
rect 3700 15098 3752 15104
rect 3976 15156 4028 15162
rect 3976 15098 4028 15104
rect 4080 14618 4108 15302
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 3700 13864 3752 13870
rect 3700 13806 3752 13812
rect 3712 13530 3740 13806
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 3700 13524 3752 13530
rect 3700 13466 3752 13472
rect 4894 12744 4950 12753
rect 4620 12708 4672 12714
rect 4894 12679 4950 12688
rect 4620 12650 4672 12656
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4344 12232 4396 12238
rect 4632 12186 4660 12650
rect 4908 12374 4936 12679
rect 5000 12434 5028 20402
rect 5080 19848 5132 19854
rect 5080 19790 5132 19796
rect 5184 19802 5212 20590
rect 5368 20466 5396 20878
rect 5356 20460 5408 20466
rect 5356 20402 5408 20408
rect 5092 19514 5120 19790
rect 5184 19774 5304 19802
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 5080 19508 5132 19514
rect 5080 19450 5132 19456
rect 5092 18834 5120 19450
rect 5184 19378 5212 19654
rect 5172 19372 5224 19378
rect 5172 19314 5224 19320
rect 5080 18828 5132 18834
rect 5080 18770 5132 18776
rect 5276 18222 5304 19774
rect 5356 19780 5408 19786
rect 5356 19722 5408 19728
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 5092 16182 5120 16390
rect 5080 16176 5132 16182
rect 5080 16118 5132 16124
rect 5276 16046 5304 18158
rect 5368 16658 5396 19722
rect 5552 19514 5580 23734
rect 5644 22094 5672 24074
rect 5816 24064 5868 24070
rect 5816 24006 5868 24012
rect 5828 23866 5856 24006
rect 5816 23860 5868 23866
rect 5816 23802 5868 23808
rect 6000 23112 6052 23118
rect 6000 23054 6052 23060
rect 5908 22772 5960 22778
rect 5908 22714 5960 22720
rect 5816 22704 5868 22710
rect 5816 22646 5868 22652
rect 5828 22234 5856 22646
rect 5816 22228 5868 22234
rect 5816 22170 5868 22176
rect 5920 22098 5948 22714
rect 5644 22066 5764 22094
rect 5632 21888 5684 21894
rect 5632 21830 5684 21836
rect 5644 21690 5672 21830
rect 5632 21684 5684 21690
rect 5632 21626 5684 21632
rect 5632 20800 5684 20806
rect 5632 20742 5684 20748
rect 5540 19508 5592 19514
rect 5540 19450 5592 19456
rect 5644 19378 5672 20742
rect 5736 20058 5764 22066
rect 5908 22092 5960 22098
rect 5908 22034 5960 22040
rect 5816 21956 5868 21962
rect 5816 21898 5868 21904
rect 5828 20942 5856 21898
rect 5908 21344 5960 21350
rect 5908 21286 5960 21292
rect 5920 21010 5948 21286
rect 5908 21004 5960 21010
rect 5908 20946 5960 20952
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 6012 20806 6040 23054
rect 6092 22228 6144 22234
rect 6092 22170 6144 22176
rect 6000 20800 6052 20806
rect 6000 20742 6052 20748
rect 5816 20596 5868 20602
rect 5816 20538 5868 20544
rect 5828 20058 5856 20538
rect 5908 20528 5960 20534
rect 5908 20470 5960 20476
rect 5724 20052 5776 20058
rect 5724 19994 5776 20000
rect 5816 20052 5868 20058
rect 5816 19994 5868 20000
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 5736 19378 5764 19790
rect 5816 19780 5868 19786
rect 5816 19722 5868 19728
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 5724 19372 5776 19378
rect 5724 19314 5776 19320
rect 5632 19236 5684 19242
rect 5632 19178 5684 19184
rect 5644 18766 5672 19178
rect 5736 18970 5764 19314
rect 5828 19242 5856 19722
rect 5816 19236 5868 19242
rect 5816 19178 5868 19184
rect 5724 18964 5776 18970
rect 5724 18906 5776 18912
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5632 18760 5684 18766
rect 5632 18702 5684 18708
rect 5552 18306 5580 18702
rect 5552 18278 5672 18306
rect 5644 18222 5672 18278
rect 5632 18216 5684 18222
rect 5632 18158 5684 18164
rect 5644 17814 5672 18158
rect 5632 17808 5684 17814
rect 5632 17750 5684 17756
rect 5632 17672 5684 17678
rect 5632 17614 5684 17620
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5368 16250 5396 16594
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 5460 15706 5488 16390
rect 5644 16182 5672 17614
rect 5632 16176 5684 16182
rect 5632 16118 5684 16124
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5644 15434 5672 16118
rect 5632 15428 5684 15434
rect 5632 15370 5684 15376
rect 5354 15192 5410 15201
rect 5354 15127 5410 15136
rect 5368 13938 5396 15127
rect 5644 15094 5672 15370
rect 5632 15088 5684 15094
rect 5632 15030 5684 15036
rect 5644 14006 5672 15030
rect 5632 14000 5684 14006
rect 5632 13942 5684 13948
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5552 13326 5580 13738
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5000 12406 5120 12434
rect 4896 12368 4948 12374
rect 4896 12310 4948 12316
rect 4396 12180 4660 12186
rect 4344 12174 4660 12180
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 4356 12158 4660 12174
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 4344 12096 4396 12102
rect 4396 12056 4476 12084
rect 4344 12038 4396 12044
rect 3988 11898 4016 12038
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 4448 11694 4476 12056
rect 4632 11778 4660 12158
rect 4816 11898 4844 12174
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4908 11778 4936 12174
rect 4632 11750 4936 11778
rect 4436 11688 4488 11694
rect 4436 11630 4488 11636
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4816 10470 4844 11630
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4816 10266 4844 10406
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4908 9994 4936 11750
rect 5000 11354 5028 12174
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 4896 9988 4948 9994
rect 4896 9930 4948 9936
rect 5092 9586 5120 12406
rect 5276 12306 5304 13262
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 5368 12050 5396 12174
rect 5460 12102 5488 13262
rect 5920 12238 5948 20470
rect 6012 20466 6040 20742
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 6012 17882 6040 18702
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 6012 17202 6040 17818
rect 6104 17678 6132 22170
rect 6288 22094 6316 27270
rect 6380 26314 6408 27338
rect 6368 26308 6420 26314
rect 6368 26250 6420 26256
rect 6368 25832 6420 25838
rect 6368 25774 6420 25780
rect 6380 24818 6408 25774
rect 6368 24812 6420 24818
rect 6368 24754 6420 24760
rect 6380 22642 6408 24754
rect 6472 24206 6500 28966
rect 6656 28558 6684 29106
rect 7208 29073 7236 29582
rect 7194 29064 7250 29073
rect 6828 29028 6880 29034
rect 7194 28999 7250 29008
rect 6828 28970 6880 28976
rect 6644 28552 6696 28558
rect 6644 28494 6696 28500
rect 6840 27062 6868 28970
rect 7012 28960 7064 28966
rect 7012 28902 7064 28908
rect 7024 27402 7052 28902
rect 7012 27396 7064 27402
rect 7012 27338 7064 27344
rect 7024 27130 7052 27338
rect 7012 27124 7064 27130
rect 7012 27066 7064 27072
rect 6828 27056 6880 27062
rect 6828 26998 6880 27004
rect 6552 26512 6604 26518
rect 6552 26454 6604 26460
rect 6460 24200 6512 24206
rect 6458 24168 6460 24177
rect 6512 24168 6514 24177
rect 6458 24103 6514 24112
rect 6368 22636 6420 22642
rect 6368 22578 6420 22584
rect 6288 22066 6408 22094
rect 6276 21344 6328 21350
rect 6276 21286 6328 21292
rect 6288 21010 6316 21286
rect 6276 21004 6328 21010
rect 6276 20946 6328 20952
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6092 17672 6144 17678
rect 6092 17614 6144 17620
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 6104 16250 6132 16526
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 6196 16046 6224 18566
rect 6380 17882 6408 22066
rect 6368 17876 6420 17882
rect 6368 17818 6420 17824
rect 6564 17814 6592 26454
rect 7024 26314 7052 27066
rect 6828 26308 6880 26314
rect 6828 26250 6880 26256
rect 7012 26308 7064 26314
rect 7012 26250 7064 26256
rect 6644 25152 6696 25158
rect 6644 25094 6696 25100
rect 6656 24954 6684 25094
rect 6644 24948 6696 24954
rect 6644 24890 6696 24896
rect 6840 24410 6868 26250
rect 7104 26240 7156 26246
rect 7104 26182 7156 26188
rect 6920 25900 6972 25906
rect 6920 25842 6972 25848
rect 6828 24404 6880 24410
rect 6828 24346 6880 24352
rect 6932 24138 6960 25842
rect 7116 25838 7144 26182
rect 7104 25832 7156 25838
rect 7104 25774 7156 25780
rect 7116 24886 7144 25774
rect 7196 25696 7248 25702
rect 7196 25638 7248 25644
rect 7208 25362 7236 25638
rect 7196 25356 7248 25362
rect 7196 25298 7248 25304
rect 7300 25226 7328 31078
rect 7392 29850 7420 33918
rect 7484 33590 7512 40054
rect 7840 39432 7892 39438
rect 7840 39374 7892 39380
rect 7852 39302 7880 39374
rect 7840 39296 7892 39302
rect 7840 39238 7892 39244
rect 8036 38486 8064 40394
rect 8852 40384 8904 40390
rect 8852 40326 8904 40332
rect 8208 40112 8260 40118
rect 8208 40054 8260 40060
rect 8116 39840 8168 39846
rect 8116 39782 8168 39788
rect 8128 39370 8156 39782
rect 8220 39642 8248 40054
rect 8484 40044 8536 40050
rect 8484 39986 8536 39992
rect 8208 39636 8260 39642
rect 8208 39578 8260 39584
rect 8496 39522 8524 39986
rect 8576 39976 8628 39982
rect 8576 39918 8628 39924
rect 8588 39642 8616 39918
rect 8576 39636 8628 39642
rect 8576 39578 8628 39584
rect 8668 39636 8720 39642
rect 8668 39578 8720 39584
rect 8680 39522 8708 39578
rect 8496 39506 8708 39522
rect 8484 39500 8708 39506
rect 8536 39494 8708 39500
rect 8484 39442 8536 39448
rect 8116 39364 8168 39370
rect 8116 39306 8168 39312
rect 8392 39296 8444 39302
rect 8392 39238 8444 39244
rect 8484 39296 8536 39302
rect 8484 39238 8536 39244
rect 8404 39098 8432 39238
rect 8392 39092 8444 39098
rect 8392 39034 8444 39040
rect 8496 38962 8524 39238
rect 8864 38962 8892 40326
rect 9220 39500 9272 39506
rect 9220 39442 9272 39448
rect 9232 39098 9260 39442
rect 9220 39092 9272 39098
rect 9220 39034 9272 39040
rect 8484 38956 8536 38962
rect 8404 38916 8484 38944
rect 8208 38752 8260 38758
rect 8208 38694 8260 38700
rect 8024 38480 8076 38486
rect 8024 38422 8076 38428
rect 7748 38344 7800 38350
rect 7748 38286 7800 38292
rect 7760 37670 7788 38286
rect 7748 37664 7800 37670
rect 7748 37606 7800 37612
rect 7656 37460 7708 37466
rect 7656 37402 7708 37408
rect 7564 36712 7616 36718
rect 7564 36654 7616 36660
rect 7576 36378 7604 36654
rect 7564 36372 7616 36378
rect 7564 36314 7616 36320
rect 7564 35148 7616 35154
rect 7564 35090 7616 35096
rect 7576 34746 7604 35090
rect 7564 34740 7616 34746
rect 7564 34682 7616 34688
rect 7564 34536 7616 34542
rect 7564 34478 7616 34484
rect 7472 33584 7524 33590
rect 7472 33526 7524 33532
rect 7576 31754 7604 34478
rect 7668 34474 7696 37402
rect 7760 36786 7788 37606
rect 8036 37398 8064 38422
rect 8220 38350 8248 38694
rect 8208 38344 8260 38350
rect 8208 38286 8260 38292
rect 8116 38004 8168 38010
rect 8116 37946 8168 37952
rect 8128 37670 8156 37946
rect 8220 37942 8248 38286
rect 8208 37936 8260 37942
rect 8208 37878 8260 37884
rect 8116 37664 8168 37670
rect 8116 37606 8168 37612
rect 8024 37392 8076 37398
rect 8024 37334 8076 37340
rect 8300 37120 8352 37126
rect 8300 37062 8352 37068
rect 8312 36854 8340 37062
rect 8300 36848 8352 36854
rect 8300 36790 8352 36796
rect 7748 36780 7800 36786
rect 7748 36722 7800 36728
rect 7932 36304 7984 36310
rect 7932 36246 7984 36252
rect 7748 36100 7800 36106
rect 7748 36042 7800 36048
rect 7760 35290 7788 36042
rect 7748 35284 7800 35290
rect 7748 35226 7800 35232
rect 7656 34468 7708 34474
rect 7656 34410 7708 34416
rect 7656 32768 7708 32774
rect 7656 32710 7708 32716
rect 7668 32570 7696 32710
rect 7656 32564 7708 32570
rect 7656 32506 7708 32512
rect 7748 32224 7800 32230
rect 7748 32166 7800 32172
rect 7760 31890 7788 32166
rect 7944 32026 7972 36246
rect 8208 36168 8260 36174
rect 8208 36110 8260 36116
rect 8300 36168 8352 36174
rect 8404 36156 8432 38916
rect 8484 38898 8536 38904
rect 8668 38956 8720 38962
rect 8852 38956 8904 38962
rect 8720 38916 8800 38944
rect 8668 38898 8720 38904
rect 8484 38752 8536 38758
rect 8484 38694 8536 38700
rect 8352 36128 8432 36156
rect 8300 36110 8352 36116
rect 8116 36100 8168 36106
rect 8116 36042 8168 36048
rect 8128 35834 8156 36042
rect 8116 35828 8168 35834
rect 8116 35770 8168 35776
rect 8024 33040 8076 33046
rect 8024 32982 8076 32988
rect 8036 32570 8064 32982
rect 8024 32564 8076 32570
rect 8024 32506 8076 32512
rect 7932 32020 7984 32026
rect 7932 31962 7984 31968
rect 7748 31884 7800 31890
rect 7748 31826 7800 31832
rect 7576 31726 7880 31754
rect 7656 31680 7708 31686
rect 7656 31622 7708 31628
rect 7668 31278 7696 31622
rect 7656 31272 7708 31278
rect 7656 31214 7708 31220
rect 7852 30190 7880 31726
rect 7944 31142 7972 31962
rect 7932 31136 7984 31142
rect 7932 31078 7984 31084
rect 7932 30252 7984 30258
rect 7932 30194 7984 30200
rect 7840 30184 7892 30190
rect 7840 30126 7892 30132
rect 7380 29844 7432 29850
rect 7380 29786 7432 29792
rect 7852 29730 7880 30126
rect 7944 29850 7972 30194
rect 7932 29844 7984 29850
rect 7932 29786 7984 29792
rect 7852 29702 8064 29730
rect 7380 29640 7432 29646
rect 7748 29640 7800 29646
rect 7432 29600 7696 29628
rect 7380 29582 7432 29588
rect 7668 29170 7696 29600
rect 7746 29608 7748 29617
rect 7932 29640 7984 29646
rect 7800 29608 7802 29617
rect 7932 29582 7984 29588
rect 7746 29543 7802 29552
rect 7840 29504 7892 29510
rect 7840 29446 7892 29452
rect 7852 29306 7880 29446
rect 7840 29300 7892 29306
rect 7840 29242 7892 29248
rect 7944 29170 7972 29582
rect 7380 29164 7432 29170
rect 7380 29106 7432 29112
rect 7564 29164 7616 29170
rect 7564 29106 7616 29112
rect 7656 29164 7708 29170
rect 7656 29106 7708 29112
rect 7932 29164 7984 29170
rect 7932 29106 7984 29112
rect 7392 29034 7420 29106
rect 7380 29028 7432 29034
rect 7380 28970 7432 28976
rect 7576 28558 7604 29106
rect 7564 28552 7616 28558
rect 7564 28494 7616 28500
rect 7380 28484 7432 28490
rect 7380 28426 7432 28432
rect 7392 26926 7420 28426
rect 7380 26920 7432 26926
rect 7380 26862 7432 26868
rect 7392 25498 7420 26862
rect 7564 25832 7616 25838
rect 7564 25774 7616 25780
rect 7380 25492 7432 25498
rect 7380 25434 7432 25440
rect 7576 25430 7604 25774
rect 7564 25424 7616 25430
rect 7564 25366 7616 25372
rect 7472 25288 7524 25294
rect 7524 25248 7604 25276
rect 7472 25230 7524 25236
rect 7288 25220 7340 25226
rect 7288 25162 7340 25168
rect 7104 24880 7156 24886
rect 7104 24822 7156 24828
rect 7196 24268 7248 24274
rect 7300 24256 7328 25162
rect 7472 25152 7524 25158
rect 7472 25094 7524 25100
rect 7484 24954 7512 25094
rect 7472 24948 7524 24954
rect 7472 24890 7524 24896
rect 7248 24228 7328 24256
rect 7196 24210 7248 24216
rect 6920 24132 6972 24138
rect 6920 24074 6972 24080
rect 7196 24132 7248 24138
rect 7196 24074 7248 24080
rect 7208 23866 7236 24074
rect 7196 23860 7248 23866
rect 7196 23802 7248 23808
rect 7380 23724 7432 23730
rect 7380 23666 7432 23672
rect 7104 23520 7156 23526
rect 7104 23462 7156 23468
rect 7116 23322 7144 23462
rect 7104 23316 7156 23322
rect 7104 23258 7156 23264
rect 7104 23112 7156 23118
rect 7104 23054 7156 23060
rect 7116 22098 7144 23054
rect 7288 22704 7340 22710
rect 7288 22646 7340 22652
rect 7196 22568 7248 22574
rect 7196 22510 7248 22516
rect 7208 22234 7236 22510
rect 7196 22228 7248 22234
rect 7196 22170 7248 22176
rect 7104 22092 7156 22098
rect 7104 22034 7156 22040
rect 7300 21894 7328 22646
rect 7288 21888 7340 21894
rect 7288 21830 7340 21836
rect 6920 21412 6972 21418
rect 6920 21354 6972 21360
rect 6828 20528 6880 20534
rect 6828 20470 6880 20476
rect 6840 20233 6868 20470
rect 6932 20398 6960 21354
rect 7300 20942 7328 21830
rect 7288 20936 7340 20942
rect 7288 20878 7340 20884
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 6826 20224 6882 20233
rect 6826 20159 6882 20168
rect 7012 19780 7064 19786
rect 7012 19722 7064 19728
rect 6828 19712 6880 19718
rect 6828 19654 6880 19660
rect 6840 19242 6868 19654
rect 7024 19514 7052 19722
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 7300 19417 7328 20878
rect 7286 19408 7342 19417
rect 7286 19343 7342 19352
rect 6828 19236 6880 19242
rect 6828 19178 6880 19184
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 6932 18426 6960 19110
rect 7300 18630 7328 19343
rect 7392 18970 7420 23666
rect 7472 23588 7524 23594
rect 7472 23530 7524 23536
rect 7484 23322 7512 23530
rect 7472 23316 7524 23322
rect 7472 23258 7524 23264
rect 7472 23112 7524 23118
rect 7472 23054 7524 23060
rect 7484 22778 7512 23054
rect 7472 22772 7524 22778
rect 7472 22714 7524 22720
rect 7472 22092 7524 22098
rect 7472 22034 7524 22040
rect 7380 18964 7432 18970
rect 7380 18906 7432 18912
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 7288 18624 7340 18630
rect 7288 18566 7340 18572
rect 7116 18426 7144 18566
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 7104 18420 7156 18426
rect 7104 18362 7156 18368
rect 6552 17808 6604 17814
rect 6552 17750 6604 17756
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6656 16658 6684 16934
rect 6840 16810 6868 16934
rect 6748 16794 6868 16810
rect 6736 16788 6868 16794
rect 6788 16782 6868 16788
rect 6736 16730 6788 16736
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6644 16652 6696 16658
rect 6644 16594 6696 16600
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 6196 15706 6224 15982
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6288 15502 6316 16594
rect 6840 16046 6868 16782
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 6288 14958 6316 15438
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 6012 13326 6040 13670
rect 6092 13456 6144 13462
rect 6092 13398 6144 13404
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 5998 12744 6054 12753
rect 5998 12679 6054 12688
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 5276 12022 5396 12050
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5276 11558 5304 12022
rect 5644 11762 5672 12106
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5828 11898 5856 12038
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5368 11626 5580 11642
rect 5356 11620 5592 11626
rect 5408 11614 5540 11620
rect 5356 11562 5408 11568
rect 5540 11562 5592 11568
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 5276 11014 5304 11494
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 5276 9994 5304 10950
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5368 9994 5396 10406
rect 6012 10130 6040 12679
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 5356 9988 5408 9994
rect 5356 9930 5408 9936
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 5276 9450 5304 9930
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5736 9586 5764 9862
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 6000 9580 6052 9586
rect 6104 9568 6132 13398
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6196 11354 6224 11698
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 6052 9540 6132 9568
rect 6000 9522 6052 9528
rect 5264 9444 5316 9450
rect 5264 9386 5316 9392
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 5460 9110 5488 9522
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4080 6798 4108 8910
rect 6104 8294 6132 9540
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6196 9178 6224 9318
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5184 6322 5212 6734
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5552 6458 5580 6666
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 6288 6254 6316 14418
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6564 13530 6592 13874
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6472 12918 6500 13262
rect 6460 12912 6512 12918
rect 6460 12854 6512 12860
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6380 12306 6408 12786
rect 6472 12442 6500 12854
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6368 12096 6420 12102
rect 6368 12038 6420 12044
rect 6380 11354 6408 12038
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6472 11150 6500 12378
rect 6656 12170 6684 14758
rect 6748 14074 6776 14894
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6748 13462 6776 13874
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 6840 13530 6868 13670
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6736 13456 6788 13462
rect 6736 13398 6788 13404
rect 7024 13326 7052 13670
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 6748 12850 6776 13126
rect 7024 12986 7052 13262
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6644 12164 6696 12170
rect 6644 12106 6696 12112
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6472 10810 6500 11086
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6564 9178 6592 9522
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6656 9042 6684 12106
rect 6748 11898 6776 12582
rect 7024 12170 7052 12922
rect 7116 12782 7144 13806
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7208 12986 7236 13126
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7208 12850 7236 12922
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 7300 12306 7328 13738
rect 7380 13252 7432 13258
rect 7380 13194 7432 13200
rect 7392 13025 7420 13194
rect 7378 13016 7434 13025
rect 7378 12951 7434 12960
rect 7380 12708 7432 12714
rect 7380 12650 7432 12656
rect 7392 12374 7420 12650
rect 7380 12368 7432 12374
rect 7380 12310 7432 12316
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7012 12164 7064 12170
rect 7012 12106 7064 12112
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7300 11898 7328 12038
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 6748 11676 6776 11834
rect 6828 11688 6880 11694
rect 6748 11648 6828 11676
rect 6828 11630 6880 11636
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7116 10810 7144 10950
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7208 10674 7236 10950
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 6932 9586 6960 10610
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6932 9178 6960 9522
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 6552 8900 6604 8906
rect 6552 8842 6604 8848
rect 6564 6798 6592 8842
rect 7116 8838 7144 8910
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7208 7478 7236 9046
rect 7484 8022 7512 22034
rect 7576 21554 7604 25248
rect 7668 24138 7696 29106
rect 7840 28960 7892 28966
rect 7840 28902 7892 28908
rect 7852 28626 7880 28902
rect 7840 28620 7892 28626
rect 7840 28562 7892 28568
rect 7748 28416 7800 28422
rect 7748 28358 7800 28364
rect 7760 27554 7788 28358
rect 7760 27526 7880 27554
rect 7748 27464 7800 27470
rect 7748 27406 7800 27412
rect 7760 27130 7788 27406
rect 7748 27124 7800 27130
rect 7748 27066 7800 27072
rect 7852 26790 7880 27526
rect 7932 27396 7984 27402
rect 7932 27338 7984 27344
rect 7944 27130 7972 27338
rect 7932 27124 7984 27130
rect 7932 27066 7984 27072
rect 7932 26988 7984 26994
rect 7932 26930 7984 26936
rect 7944 26897 7972 26930
rect 7930 26888 7986 26897
rect 7930 26823 7986 26832
rect 7840 26784 7892 26790
rect 7840 26726 7892 26732
rect 7748 24336 7800 24342
rect 7748 24278 7800 24284
rect 7656 24132 7708 24138
rect 7656 24074 7708 24080
rect 7656 21684 7708 21690
rect 7656 21626 7708 21632
rect 7564 21548 7616 21554
rect 7564 21490 7616 21496
rect 7576 19378 7604 21490
rect 7668 21146 7696 21626
rect 7656 21140 7708 21146
rect 7656 21082 7708 21088
rect 7668 20602 7696 21082
rect 7760 20806 7788 24278
rect 7852 24138 7880 26726
rect 8036 26382 8064 29702
rect 8128 29646 8156 35770
rect 8220 32230 8248 36110
rect 8312 34202 8340 36110
rect 8300 34196 8352 34202
rect 8300 34138 8352 34144
rect 8300 32496 8352 32502
rect 8300 32438 8352 32444
rect 8312 32366 8340 32438
rect 8300 32360 8352 32366
rect 8352 32320 8432 32348
rect 8300 32302 8352 32308
rect 8208 32224 8260 32230
rect 8208 32166 8260 32172
rect 8220 31822 8248 32166
rect 8208 31816 8260 31822
rect 8208 31758 8260 31764
rect 8404 31142 8432 32320
rect 8392 31136 8444 31142
rect 8392 31078 8444 31084
rect 8208 30252 8260 30258
rect 8208 30194 8260 30200
rect 8220 29714 8248 30194
rect 8298 29880 8354 29889
rect 8298 29815 8354 29824
rect 8208 29708 8260 29714
rect 8208 29650 8260 29656
rect 8116 29640 8168 29646
rect 8116 29582 8168 29588
rect 8128 26994 8156 29582
rect 8208 29572 8260 29578
rect 8312 29560 8340 29815
rect 8260 29532 8340 29560
rect 8208 29514 8260 29520
rect 8220 29238 8248 29514
rect 8404 29306 8432 31078
rect 8392 29300 8444 29306
rect 8392 29242 8444 29248
rect 8208 29232 8260 29238
rect 8208 29174 8260 29180
rect 8300 29164 8352 29170
rect 8352 29124 8432 29152
rect 8300 29106 8352 29112
rect 8404 29034 8432 29124
rect 8300 29028 8352 29034
rect 8300 28970 8352 28976
rect 8392 29028 8444 29034
rect 8392 28970 8444 28976
rect 8208 28960 8260 28966
rect 8208 28902 8260 28908
rect 8116 26988 8168 26994
rect 8116 26930 8168 26936
rect 8024 26376 8076 26382
rect 8024 26318 8076 26324
rect 8116 25900 8168 25906
rect 8036 25860 8116 25888
rect 8036 24886 8064 25860
rect 8220 25888 8248 28902
rect 8312 28694 8340 28970
rect 8300 28688 8352 28694
rect 8300 28630 8352 28636
rect 8300 27872 8352 27878
rect 8300 27814 8352 27820
rect 8312 27674 8340 27814
rect 8300 27668 8352 27674
rect 8300 27610 8352 27616
rect 8390 27568 8446 27577
rect 8390 27503 8446 27512
rect 8300 27464 8352 27470
rect 8300 27406 8352 27412
rect 8312 27130 8340 27406
rect 8404 27334 8432 27503
rect 8496 27470 8524 38694
rect 8668 36644 8720 36650
rect 8668 36586 8720 36592
rect 8680 33522 8708 36586
rect 8772 35290 8800 38916
rect 8852 38898 8904 38904
rect 8864 36106 8892 38898
rect 8944 37868 8996 37874
rect 8944 37810 8996 37816
rect 8852 36100 8904 36106
rect 8852 36042 8904 36048
rect 8760 35284 8812 35290
rect 8760 35226 8812 35232
rect 8956 34474 8984 37810
rect 9036 37120 9088 37126
rect 9036 37062 9088 37068
rect 8944 34468 8996 34474
rect 8944 34410 8996 34416
rect 8668 33516 8720 33522
rect 8668 33458 8720 33464
rect 8576 32224 8628 32230
rect 8576 32166 8628 32172
rect 8588 31278 8616 32166
rect 9048 31754 9076 37062
rect 9128 33516 9180 33522
rect 9128 33458 9180 33464
rect 8772 31726 9076 31754
rect 8576 31272 8628 31278
rect 8576 31214 8628 31220
rect 8576 30252 8628 30258
rect 8576 30194 8628 30200
rect 8588 29646 8616 30194
rect 8668 29844 8720 29850
rect 8668 29786 8720 29792
rect 8576 29640 8628 29646
rect 8576 29582 8628 29588
rect 8588 29238 8616 29582
rect 8680 29238 8708 29786
rect 8576 29232 8628 29238
rect 8576 29174 8628 29180
rect 8668 29232 8720 29238
rect 8668 29174 8720 29180
rect 8668 27940 8720 27946
rect 8668 27882 8720 27888
rect 8484 27464 8536 27470
rect 8484 27406 8536 27412
rect 8576 27464 8628 27470
rect 8576 27406 8628 27412
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8300 27124 8352 27130
rect 8300 27066 8352 27072
rect 8300 26988 8352 26994
rect 8300 26930 8352 26936
rect 8312 26518 8340 26930
rect 8300 26512 8352 26518
rect 8300 26454 8352 26460
rect 8168 25860 8248 25888
rect 8116 25842 8168 25848
rect 8116 24948 8168 24954
rect 8116 24890 8168 24896
rect 8024 24880 8076 24886
rect 8024 24822 8076 24828
rect 7840 24132 7892 24138
rect 7840 24074 7892 24080
rect 7932 23112 7984 23118
rect 7932 23054 7984 23060
rect 7944 22012 7972 23054
rect 8036 22930 8064 24822
rect 8128 24206 8156 24890
rect 8206 24848 8262 24857
rect 8312 24818 8340 26454
rect 8206 24783 8208 24792
rect 8260 24783 8262 24792
rect 8300 24812 8352 24818
rect 8208 24754 8260 24760
rect 8300 24754 8352 24760
rect 8116 24200 8168 24206
rect 8116 24142 8168 24148
rect 8300 24132 8352 24138
rect 8300 24074 8352 24080
rect 8116 23316 8168 23322
rect 8116 23258 8168 23264
rect 8128 23050 8156 23258
rect 8116 23044 8168 23050
rect 8116 22986 8168 22992
rect 8036 22902 8156 22930
rect 7944 21984 8064 22012
rect 7932 21072 7984 21078
rect 7932 21014 7984 21020
rect 7748 20800 7800 20806
rect 7748 20742 7800 20748
rect 7656 20596 7708 20602
rect 7656 20538 7708 20544
rect 7656 20460 7708 20466
rect 7656 20402 7708 20408
rect 7748 20460 7800 20466
rect 7748 20402 7800 20408
rect 7668 19394 7696 20402
rect 7760 20330 7788 20402
rect 7748 20324 7800 20330
rect 7748 20266 7800 20272
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 7746 19408 7802 19417
rect 7564 19372 7616 19378
rect 7668 19366 7746 19394
rect 7746 19343 7802 19352
rect 7564 19314 7616 19320
rect 7576 17134 7604 19314
rect 7852 18970 7880 19790
rect 7840 18964 7892 18970
rect 7840 18906 7892 18912
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7576 11694 7604 17070
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 7852 15502 7880 15846
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7944 15178 7972 21014
rect 8036 20466 8064 21984
rect 8024 20460 8076 20466
rect 8024 20402 8076 20408
rect 8024 20324 8076 20330
rect 8024 20266 8076 20272
rect 8036 19990 8064 20266
rect 8024 19984 8076 19990
rect 8024 19926 8076 19932
rect 8128 19938 8156 22902
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 8220 21690 8248 22578
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 8220 20058 8248 20198
rect 8312 20058 8340 24074
rect 8404 23610 8432 27270
rect 8496 23730 8524 27406
rect 8588 27305 8616 27406
rect 8574 27296 8630 27305
rect 8574 27231 8630 27240
rect 8576 26988 8628 26994
rect 8576 26930 8628 26936
rect 8588 26382 8616 26930
rect 8680 26790 8708 27882
rect 8772 27577 8800 31726
rect 8944 31680 8996 31686
rect 9140 31634 9168 33458
rect 8996 31628 9168 31634
rect 8944 31622 9168 31628
rect 8956 31606 9168 31622
rect 8956 31482 8984 31606
rect 8944 31476 8996 31482
rect 8944 31418 8996 31424
rect 9324 30410 9352 41958
rect 11152 41676 11204 41682
rect 11152 41618 11204 41624
rect 10600 41540 10652 41546
rect 10600 41482 10652 41488
rect 10612 41414 10640 41482
rect 10968 41472 11020 41478
rect 10968 41414 11020 41420
rect 9692 41386 10640 41414
rect 10888 41386 11008 41414
rect 9588 39500 9640 39506
rect 9588 39442 9640 39448
rect 9600 38962 9628 39442
rect 9692 39370 9720 41386
rect 9772 40656 9824 40662
rect 9772 40598 9824 40604
rect 9680 39364 9732 39370
rect 9680 39306 9732 39312
rect 9588 38956 9640 38962
rect 9588 38898 9640 38904
rect 9404 38412 9456 38418
rect 9404 38354 9456 38360
rect 9416 38010 9444 38354
rect 9404 38004 9456 38010
rect 9404 37946 9456 37952
rect 9496 37868 9548 37874
rect 9496 37810 9548 37816
rect 9508 37466 9536 37810
rect 9496 37460 9548 37466
rect 9496 37402 9548 37408
rect 9404 32428 9456 32434
rect 9404 32370 9456 32376
rect 9416 31686 9444 32370
rect 9404 31680 9456 31686
rect 9404 31622 9456 31628
rect 9416 31328 9444 31622
rect 9496 31340 9548 31346
rect 9416 31300 9496 31328
rect 9496 31282 9548 31288
rect 8956 30394 9352 30410
rect 8944 30388 9352 30394
rect 8996 30382 9352 30388
rect 8944 30330 8996 30336
rect 8852 30184 8904 30190
rect 8852 30126 8904 30132
rect 8864 29889 8892 30126
rect 8850 29880 8906 29889
rect 8850 29815 8906 29824
rect 8852 28960 8904 28966
rect 8852 28902 8904 28908
rect 8864 28422 8892 28902
rect 8852 28416 8904 28422
rect 8852 28358 8904 28364
rect 8852 27600 8904 27606
rect 8758 27568 8814 27577
rect 8852 27542 8904 27548
rect 8758 27503 8814 27512
rect 8760 27464 8812 27470
rect 8864 27441 8892 27542
rect 8760 27406 8812 27412
rect 8850 27432 8906 27441
rect 8668 26784 8720 26790
rect 8668 26726 8720 26732
rect 8576 26376 8628 26382
rect 8576 26318 8628 26324
rect 8588 25838 8616 26318
rect 8576 25832 8628 25838
rect 8576 25774 8628 25780
rect 8680 24290 8708 26726
rect 8772 26518 8800 27406
rect 8850 27367 8906 27376
rect 8956 27130 8984 30330
rect 9508 30258 9536 31282
rect 9312 30252 9364 30258
rect 9312 30194 9364 30200
rect 9496 30252 9548 30258
rect 9496 30194 9548 30200
rect 9324 29714 9352 30194
rect 9312 29708 9364 29714
rect 9312 29650 9364 29656
rect 9404 29640 9456 29646
rect 9404 29582 9456 29588
rect 9220 29572 9272 29578
rect 9220 29514 9272 29520
rect 9128 29232 9180 29238
rect 9128 29174 9180 29180
rect 9036 29096 9088 29102
rect 9034 29064 9036 29073
rect 9088 29064 9090 29073
rect 9034 28999 9090 29008
rect 9140 27452 9168 29174
rect 9232 27577 9260 29514
rect 9312 29164 9364 29170
rect 9312 29106 9364 29112
rect 9324 28218 9352 29106
rect 9312 28212 9364 28218
rect 9312 28154 9364 28160
rect 9416 27614 9444 29582
rect 9508 27826 9536 30194
rect 9600 29646 9628 38898
rect 9784 38654 9812 40598
rect 10416 40520 10468 40526
rect 10416 40462 10468 40468
rect 9956 40384 10008 40390
rect 9956 40326 10008 40332
rect 9862 40216 9918 40225
rect 9862 40151 9864 40160
rect 9916 40151 9918 40160
rect 9864 40122 9916 40128
rect 9968 39302 9996 40326
rect 10428 40202 10456 40462
rect 10692 40452 10744 40458
rect 10692 40394 10744 40400
rect 10598 40216 10654 40225
rect 10428 40186 10548 40202
rect 10428 40180 10560 40186
rect 10428 40174 10508 40180
rect 10598 40151 10600 40160
rect 10508 40122 10560 40128
rect 10652 40151 10654 40160
rect 10600 40122 10652 40128
rect 10140 40112 10192 40118
rect 10046 40080 10102 40089
rect 10192 40072 10456 40100
rect 10140 40054 10192 40060
rect 10046 40015 10048 40024
rect 10100 40015 10102 40024
rect 10048 39986 10100 39992
rect 10428 39982 10456 40072
rect 10140 39976 10192 39982
rect 10140 39918 10192 39924
rect 10416 39976 10468 39982
rect 10416 39918 10468 39924
rect 10152 39302 10180 39918
rect 9956 39296 10008 39302
rect 9956 39238 10008 39244
rect 10140 39296 10192 39302
rect 10140 39238 10192 39244
rect 9784 38626 9996 38654
rect 9680 37800 9732 37806
rect 9680 37742 9732 37748
rect 9692 34746 9720 37742
rect 9968 37262 9996 38626
rect 10416 37664 10468 37670
rect 10416 37606 10468 37612
rect 10324 37324 10376 37330
rect 10324 37266 10376 37272
rect 9956 37256 10008 37262
rect 9956 37198 10008 37204
rect 9968 35630 9996 37198
rect 10232 36780 10284 36786
rect 10232 36722 10284 36728
rect 10244 36310 10272 36722
rect 10336 36378 10364 37266
rect 10324 36372 10376 36378
rect 10324 36314 10376 36320
rect 10232 36304 10284 36310
rect 10232 36246 10284 36252
rect 10048 36100 10100 36106
rect 10048 36042 10100 36048
rect 10060 35986 10088 36042
rect 10060 35958 10180 35986
rect 9956 35624 10008 35630
rect 9956 35566 10008 35572
rect 9864 35488 9916 35494
rect 9864 35430 9916 35436
rect 9876 35290 9904 35430
rect 9864 35284 9916 35290
rect 9864 35226 9916 35232
rect 9968 34950 9996 35566
rect 10152 35494 10180 35958
rect 10244 35630 10272 36246
rect 10428 35766 10456 37606
rect 10704 36922 10732 40394
rect 10782 40080 10838 40089
rect 10782 40015 10784 40024
rect 10836 40015 10838 40024
rect 10784 39986 10836 39992
rect 10796 39438 10824 39986
rect 10888 39914 10916 41386
rect 11060 40928 11112 40934
rect 11060 40870 11112 40876
rect 11072 40526 11100 40870
rect 11164 40730 11192 41618
rect 12072 41540 12124 41546
rect 12072 41482 12124 41488
rect 11520 41472 11572 41478
rect 11520 41414 11572 41420
rect 11532 41070 11560 41414
rect 12084 41274 12112 41482
rect 12912 41478 12940 43893
rect 16132 41614 16160 43893
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 17500 42220 17552 42226
rect 17500 42162 17552 42168
rect 19432 42220 19484 42226
rect 19432 42162 19484 42168
rect 17316 42016 17368 42022
rect 17316 41958 17368 41964
rect 17328 41818 17356 41958
rect 17316 41812 17368 41818
rect 17316 41754 17368 41760
rect 16120 41608 16172 41614
rect 16120 41550 16172 41556
rect 14004 41540 14056 41546
rect 14004 41482 14056 41488
rect 14372 41540 14424 41546
rect 14372 41482 14424 41488
rect 12900 41472 12952 41478
rect 12900 41414 12952 41420
rect 14016 41414 14044 41482
rect 12820 41386 12940 41414
rect 13924 41386 14044 41414
rect 12072 41268 12124 41274
rect 12072 41210 12124 41216
rect 12820 41138 12848 41386
rect 12532 41132 12584 41138
rect 12532 41074 12584 41080
rect 12808 41132 12860 41138
rect 12808 41074 12860 41080
rect 11520 41064 11572 41070
rect 11520 41006 11572 41012
rect 11152 40724 11204 40730
rect 11152 40666 11204 40672
rect 11532 40526 11560 41006
rect 11060 40520 11112 40526
rect 11060 40462 11112 40468
rect 11520 40520 11572 40526
rect 11520 40462 11572 40468
rect 11244 40384 11296 40390
rect 11244 40326 11296 40332
rect 11336 40384 11388 40390
rect 11336 40326 11388 40332
rect 11428 40384 11480 40390
rect 11428 40326 11480 40332
rect 11152 40180 11204 40186
rect 11152 40122 11204 40128
rect 11060 40112 11112 40118
rect 11060 40054 11112 40060
rect 10876 39908 10928 39914
rect 10876 39850 10928 39856
rect 10784 39432 10836 39438
rect 10784 39374 10836 39380
rect 11072 39370 11100 40054
rect 11060 39364 11112 39370
rect 11060 39306 11112 39312
rect 10784 38956 10836 38962
rect 10784 38898 10836 38904
rect 10796 37874 10824 38898
rect 11164 38350 11192 40122
rect 11256 39642 11284 40326
rect 11348 40186 11376 40326
rect 11336 40180 11388 40186
rect 11336 40122 11388 40128
rect 11440 40118 11468 40326
rect 11428 40112 11480 40118
rect 11428 40054 11480 40060
rect 11244 39636 11296 39642
rect 11244 39578 11296 39584
rect 11244 39432 11296 39438
rect 11244 39374 11296 39380
rect 11256 39098 11284 39374
rect 11244 39092 11296 39098
rect 11244 39034 11296 39040
rect 11440 39030 11468 40054
rect 11532 39982 11560 40462
rect 12348 40384 12400 40390
rect 12348 40326 12400 40332
rect 11520 39976 11572 39982
rect 11520 39918 11572 39924
rect 11888 39976 11940 39982
rect 11888 39918 11940 39924
rect 11428 39024 11480 39030
rect 11428 38966 11480 38972
rect 11336 38956 11388 38962
rect 11336 38898 11388 38904
rect 11348 38758 11376 38898
rect 11532 38842 11560 39918
rect 11796 39568 11848 39574
rect 11796 39510 11848 39516
rect 11612 39432 11664 39438
rect 11612 39374 11664 39380
rect 11440 38814 11560 38842
rect 11336 38752 11388 38758
rect 11256 38712 11336 38740
rect 11256 38350 11284 38712
rect 11336 38694 11388 38700
rect 11060 38344 11112 38350
rect 11060 38286 11112 38292
rect 11152 38344 11204 38350
rect 11152 38286 11204 38292
rect 11244 38344 11296 38350
rect 11244 38286 11296 38292
rect 11072 38010 11100 38286
rect 11060 38004 11112 38010
rect 11060 37946 11112 37952
rect 10784 37868 10836 37874
rect 10784 37810 10836 37816
rect 11060 37868 11112 37874
rect 11060 37810 11112 37816
rect 11072 37466 11100 37810
rect 11060 37460 11112 37466
rect 11060 37402 11112 37408
rect 11256 37262 11284 38286
rect 11336 37936 11388 37942
rect 11336 37878 11388 37884
rect 11060 37256 11112 37262
rect 11060 37198 11112 37204
rect 11244 37256 11296 37262
rect 11244 37198 11296 37204
rect 10692 36916 10744 36922
rect 10692 36858 10744 36864
rect 10784 36712 10836 36718
rect 10784 36654 10836 36660
rect 10796 36378 10824 36654
rect 10784 36372 10836 36378
rect 10784 36314 10836 36320
rect 10508 36168 10560 36174
rect 10508 36110 10560 36116
rect 10968 36168 11020 36174
rect 10968 36110 11020 36116
rect 10416 35760 10468 35766
rect 10416 35702 10468 35708
rect 10232 35624 10284 35630
rect 10232 35566 10284 35572
rect 10140 35488 10192 35494
rect 10140 35430 10192 35436
rect 10152 35086 10180 35430
rect 10048 35080 10100 35086
rect 10048 35022 10100 35028
rect 10140 35080 10192 35086
rect 10140 35022 10192 35028
rect 9772 34944 9824 34950
rect 9956 34944 10008 34950
rect 9772 34886 9824 34892
rect 9876 34904 9956 34932
rect 9680 34740 9732 34746
rect 9680 34682 9732 34688
rect 9784 34202 9812 34886
rect 9772 34196 9824 34202
rect 9772 34138 9824 34144
rect 9680 34128 9732 34134
rect 9732 34076 9812 34082
rect 9680 34070 9812 34076
rect 9692 34054 9812 34070
rect 9680 33992 9732 33998
rect 9680 33934 9732 33940
rect 9692 33658 9720 33934
rect 9680 33652 9732 33658
rect 9680 33594 9732 33600
rect 9680 33516 9732 33522
rect 9680 33458 9732 33464
rect 9692 32450 9720 33458
rect 9784 32570 9812 34054
rect 9876 33912 9904 34904
rect 9956 34886 10008 34892
rect 9876 33884 9996 33912
rect 9864 33448 9916 33454
rect 9864 33390 9916 33396
rect 9876 32774 9904 33390
rect 9968 33300 9996 33884
rect 10060 33674 10088 35022
rect 10244 33810 10272 35566
rect 10520 35018 10548 36110
rect 10692 36032 10744 36038
rect 10692 35974 10744 35980
rect 10600 35080 10652 35086
rect 10600 35022 10652 35028
rect 10508 35012 10560 35018
rect 10508 34954 10560 34960
rect 10324 34944 10376 34950
rect 10324 34886 10376 34892
rect 10336 34746 10364 34886
rect 10324 34740 10376 34746
rect 10324 34682 10376 34688
rect 10416 34604 10468 34610
rect 10416 34546 10468 34552
rect 10244 33782 10364 33810
rect 10060 33646 10272 33674
rect 10244 33318 10272 33646
rect 10336 33454 10364 33782
rect 10324 33448 10376 33454
rect 10324 33390 10376 33396
rect 10428 33318 10456 34546
rect 10048 33312 10100 33318
rect 9968 33272 10048 33300
rect 10048 33254 10100 33260
rect 10232 33312 10284 33318
rect 10232 33254 10284 33260
rect 10416 33312 10468 33318
rect 10416 33254 10468 33260
rect 9864 32768 9916 32774
rect 9864 32710 9916 32716
rect 9772 32564 9824 32570
rect 9772 32506 9824 32512
rect 9692 32422 9812 32450
rect 9680 32224 9732 32230
rect 9680 32166 9732 32172
rect 9692 31890 9720 32166
rect 9680 31884 9732 31890
rect 9680 31826 9732 31832
rect 9784 31124 9812 32422
rect 9864 32360 9916 32366
rect 9864 32302 9916 32308
rect 9876 31278 9904 32302
rect 10060 31482 10088 33254
rect 10244 31754 10272 33254
rect 10612 32434 10640 35022
rect 10704 33998 10732 35974
rect 10980 35834 11008 36110
rect 11072 36106 11100 37198
rect 11060 36100 11112 36106
rect 11060 36042 11112 36048
rect 10968 35828 11020 35834
rect 10968 35770 11020 35776
rect 10980 35698 11008 35770
rect 10968 35692 11020 35698
rect 10968 35634 11020 35640
rect 10980 34746 11008 35634
rect 11244 35080 11296 35086
rect 11244 35022 11296 35028
rect 11256 34746 11284 35022
rect 10968 34740 11020 34746
rect 11244 34740 11296 34746
rect 10968 34682 11020 34688
rect 11164 34700 11244 34728
rect 11164 34406 11192 34700
rect 11244 34682 11296 34688
rect 11348 34474 11376 37878
rect 11336 34468 11388 34474
rect 11256 34428 11336 34456
rect 11152 34400 11204 34406
rect 11152 34342 11204 34348
rect 11164 34066 11192 34342
rect 11152 34060 11204 34066
rect 11152 34002 11204 34008
rect 10692 33992 10744 33998
rect 10692 33934 10744 33940
rect 11060 33992 11112 33998
rect 11060 33934 11112 33940
rect 10876 33448 10928 33454
rect 10876 33390 10928 33396
rect 10784 32972 10836 32978
rect 10784 32914 10836 32920
rect 10600 32428 10652 32434
rect 10600 32370 10652 32376
rect 10244 31726 10364 31754
rect 10048 31476 10100 31482
rect 10048 31418 10100 31424
rect 9864 31272 9916 31278
rect 9864 31214 9916 31220
rect 9784 31096 9904 31124
rect 9772 30116 9824 30122
rect 9772 30058 9824 30064
rect 9680 29776 9732 29782
rect 9680 29718 9732 29724
rect 9588 29640 9640 29646
rect 9588 29582 9640 29588
rect 9692 29306 9720 29718
rect 9784 29578 9812 30058
rect 9876 29753 9904 31096
rect 10232 30660 10284 30666
rect 10232 30602 10284 30608
rect 9956 30252 10008 30258
rect 9956 30194 10008 30200
rect 9862 29744 9918 29753
rect 9862 29679 9918 29688
rect 9968 29646 9996 30194
rect 9956 29640 10008 29646
rect 9956 29582 10008 29588
rect 10138 29608 10194 29617
rect 9772 29572 9824 29578
rect 9772 29514 9824 29520
rect 9864 29572 9916 29578
rect 10138 29543 10194 29552
rect 9864 29514 9916 29520
rect 9876 29458 9904 29514
rect 10048 29504 10100 29510
rect 9954 29472 10010 29481
rect 9876 29430 9954 29458
rect 10048 29446 10100 29452
rect 9954 29407 10010 29416
rect 9680 29300 9732 29306
rect 9680 29242 9732 29248
rect 10060 29238 10088 29446
rect 10048 29232 10100 29238
rect 10048 29174 10100 29180
rect 9864 29164 9916 29170
rect 9864 29106 9916 29112
rect 9876 28422 9904 29106
rect 10060 28558 10088 29174
rect 10152 29170 10180 29543
rect 10140 29164 10192 29170
rect 10140 29106 10192 29112
rect 10244 28642 10272 30602
rect 10336 29209 10364 31726
rect 10322 29200 10378 29209
rect 10322 29135 10378 29144
rect 10336 28966 10364 29135
rect 10416 29096 10468 29102
rect 10416 29038 10468 29044
rect 10324 28960 10376 28966
rect 10324 28902 10376 28908
rect 10152 28614 10272 28642
rect 10048 28552 10100 28558
rect 10048 28494 10100 28500
rect 9864 28416 9916 28422
rect 9864 28358 9916 28364
rect 10048 27872 10100 27878
rect 9508 27798 9541 27826
rect 10048 27814 10100 27820
rect 9513 27614 9541 27798
rect 9324 27586 9444 27614
rect 9508 27586 9541 27614
rect 9218 27568 9274 27577
rect 9324 27554 9352 27586
rect 9324 27526 9398 27554
rect 9218 27503 9274 27512
rect 9370 27452 9398 27526
rect 9140 27424 9260 27452
rect 9370 27424 9444 27452
rect 8944 27124 8996 27130
rect 8944 27066 8996 27072
rect 9128 27124 9180 27130
rect 9128 27066 9180 27072
rect 8852 26988 8904 26994
rect 8852 26930 8904 26936
rect 8864 26586 8892 26930
rect 9036 26784 9088 26790
rect 9140 26761 9168 27066
rect 9036 26726 9088 26732
rect 9126 26752 9182 26761
rect 8852 26580 8904 26586
rect 8852 26522 8904 26528
rect 8760 26512 8812 26518
rect 8760 26454 8812 26460
rect 8944 26376 8996 26382
rect 8944 26318 8996 26324
rect 8956 26042 8984 26318
rect 8944 26036 8996 26042
rect 8944 25978 8996 25984
rect 9048 25906 9076 26726
rect 9126 26687 9182 26696
rect 9128 26376 9180 26382
rect 9128 26318 9180 26324
rect 9036 25900 9088 25906
rect 9036 25842 9088 25848
rect 9140 25809 9168 26318
rect 9232 26296 9260 27424
rect 9416 26994 9444 27424
rect 9508 27033 9536 27586
rect 9772 27464 9824 27470
rect 9600 27424 9772 27452
rect 9494 27024 9550 27033
rect 9404 26988 9456 26994
rect 9494 26959 9550 26968
rect 9404 26930 9456 26936
rect 9496 26852 9548 26858
rect 9496 26794 9548 26800
rect 9312 26308 9364 26314
rect 9232 26268 9312 26296
rect 9312 26250 9364 26256
rect 9404 26240 9456 26246
rect 9404 26182 9456 26188
rect 9312 25968 9364 25974
rect 9312 25910 9364 25916
rect 9126 25800 9182 25809
rect 9126 25735 9182 25744
rect 9220 25764 9272 25770
rect 9220 25706 9272 25712
rect 9232 25378 9260 25706
rect 9140 25350 9260 25378
rect 9036 25220 9088 25226
rect 9036 25162 9088 25168
rect 8760 24812 8812 24818
rect 8760 24754 8812 24760
rect 8588 24262 8708 24290
rect 8484 23724 8536 23730
rect 8484 23666 8536 23672
rect 8404 23582 8524 23610
rect 8392 22432 8444 22438
rect 8392 22374 8444 22380
rect 8404 22030 8432 22374
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8496 21622 8524 23582
rect 8588 23118 8616 24262
rect 8668 24200 8720 24206
rect 8668 24142 8720 24148
rect 8576 23112 8628 23118
rect 8576 23054 8628 23060
rect 8484 21616 8536 21622
rect 8484 21558 8536 21564
rect 8392 20800 8444 20806
rect 8392 20742 8444 20748
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 8128 19910 8248 19938
rect 8116 19780 8168 19786
rect 8116 19722 8168 19728
rect 8024 19236 8076 19242
rect 8024 19178 8076 19184
rect 8036 17746 8064 19178
rect 8024 17740 8076 17746
rect 8024 17682 8076 17688
rect 8036 17202 8064 17682
rect 8128 17678 8156 19722
rect 8116 17672 8168 17678
rect 8116 17614 8168 17620
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 8036 16114 8064 17138
rect 8128 16794 8156 17614
rect 8116 16788 8168 16794
rect 8116 16730 8168 16736
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 8024 16108 8076 16114
rect 8024 16050 8076 16056
rect 8128 15502 8156 16390
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 7944 15162 8064 15178
rect 7944 15156 8076 15162
rect 7944 15150 8024 15156
rect 7944 14482 7972 15150
rect 8024 15098 8076 15104
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 7840 14340 7892 14346
rect 7840 14282 7892 14288
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 7668 14074 7696 14214
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7852 13938 7880 14282
rect 7840 13932 7892 13938
rect 7760 13892 7840 13920
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7668 11354 7696 13262
rect 7760 12850 7788 13892
rect 7840 13874 7892 13880
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 7944 13462 7972 13874
rect 7932 13456 7984 13462
rect 7932 13398 7984 13404
rect 8116 13456 8168 13462
rect 8116 13398 8168 13404
rect 8128 13326 8156 13398
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 7838 13016 7894 13025
rect 7838 12951 7894 12960
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7656 11076 7708 11082
rect 7656 11018 7708 11024
rect 7668 9654 7696 11018
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7576 9450 7604 9522
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7576 9058 7604 9386
rect 7668 9178 7696 9590
rect 7760 9586 7788 10134
rect 7852 9654 7880 12951
rect 8036 12889 8064 13126
rect 8022 12880 8078 12889
rect 8022 12815 8078 12824
rect 8220 12442 8248 19910
rect 8300 19440 8352 19446
rect 8300 19382 8352 19388
rect 8312 18970 8340 19382
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8404 18290 8432 20742
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8484 20052 8536 20058
rect 8484 19994 8536 20000
rect 8496 19854 8524 19994
rect 8484 19848 8536 19854
rect 8484 19790 8536 19796
rect 8588 19514 8616 20198
rect 8576 19508 8628 19514
rect 8576 19450 8628 19456
rect 8680 18952 8708 24142
rect 8772 24138 8800 24754
rect 8852 24608 8904 24614
rect 8852 24550 8904 24556
rect 8760 24132 8812 24138
rect 8760 24074 8812 24080
rect 8864 23866 8892 24550
rect 9048 24206 9076 25162
rect 9036 24200 9088 24206
rect 9036 24142 9088 24148
rect 8852 23860 8904 23866
rect 8852 23802 8904 23808
rect 9036 23724 9088 23730
rect 9036 23666 9088 23672
rect 8852 23112 8904 23118
rect 9048 23100 9076 23666
rect 8904 23072 9076 23100
rect 8852 23054 8904 23060
rect 8864 22030 8892 23054
rect 9140 22710 9168 25350
rect 9220 25288 9272 25294
rect 9220 25230 9272 25236
rect 9232 24993 9260 25230
rect 9324 25140 9352 25910
rect 9416 25294 9444 26182
rect 9404 25288 9456 25294
rect 9404 25230 9456 25236
rect 9324 25112 9444 25140
rect 9218 24984 9274 24993
rect 9218 24919 9274 24928
rect 9312 24744 9364 24750
rect 9218 24712 9274 24721
rect 9312 24686 9364 24692
rect 9218 24647 9220 24656
rect 9272 24647 9274 24656
rect 9220 24618 9272 24624
rect 9324 24410 9352 24686
rect 9312 24404 9364 24410
rect 9312 24346 9364 24352
rect 9416 24290 9444 25112
rect 9508 24410 9536 26794
rect 9600 25974 9628 27424
rect 10060 27452 10088 27814
rect 9772 27406 9824 27412
rect 9876 27424 10088 27452
rect 9770 27160 9826 27169
rect 9876 27130 9904 27424
rect 10048 27328 10100 27334
rect 10048 27270 10100 27276
rect 10060 27130 10088 27270
rect 9770 27095 9772 27104
rect 9824 27095 9826 27104
rect 9864 27124 9916 27130
rect 9772 27066 9824 27072
rect 9864 27066 9916 27072
rect 10048 27124 10100 27130
rect 10048 27066 10100 27072
rect 10046 27024 10102 27033
rect 9956 26988 10008 26994
rect 10046 26959 10048 26968
rect 9956 26930 10008 26936
rect 10100 26959 10102 26968
rect 10048 26930 10100 26936
rect 9680 26852 9732 26858
rect 9680 26794 9732 26800
rect 9692 26586 9720 26794
rect 9680 26580 9732 26586
rect 9680 26522 9732 26528
rect 9588 25968 9640 25974
rect 9588 25910 9640 25916
rect 9588 25832 9640 25838
rect 9588 25774 9640 25780
rect 9600 25294 9628 25774
rect 9864 25696 9916 25702
rect 9864 25638 9916 25644
rect 9588 25288 9640 25294
rect 9588 25230 9640 25236
rect 9772 25288 9824 25294
rect 9772 25230 9824 25236
rect 9496 24404 9548 24410
rect 9496 24346 9548 24352
rect 9232 24262 9444 24290
rect 9128 22704 9180 22710
rect 9128 22646 9180 22652
rect 9140 22094 9168 22646
rect 9232 22234 9260 24262
rect 9600 24206 9628 25230
rect 9784 24954 9812 25230
rect 9680 24948 9732 24954
rect 9680 24890 9732 24896
rect 9772 24948 9824 24954
rect 9772 24890 9824 24896
rect 9588 24200 9640 24206
rect 9494 24168 9550 24177
rect 9588 24142 9640 24148
rect 9494 24103 9550 24112
rect 9508 23866 9536 24103
rect 9496 23860 9548 23866
rect 9496 23802 9548 23808
rect 9692 23730 9720 24890
rect 9404 23724 9456 23730
rect 9404 23666 9456 23672
rect 9588 23724 9640 23730
rect 9588 23666 9640 23672
rect 9680 23724 9732 23730
rect 9680 23666 9732 23672
rect 9416 23254 9444 23666
rect 9496 23588 9548 23594
rect 9496 23530 9548 23536
rect 9404 23248 9456 23254
rect 9404 23190 9456 23196
rect 9508 22982 9536 23530
rect 9600 22982 9628 23666
rect 9496 22976 9548 22982
rect 9496 22918 9548 22924
rect 9588 22976 9640 22982
rect 9588 22918 9640 22924
rect 9508 22658 9536 22918
rect 9324 22630 9536 22658
rect 9220 22228 9272 22234
rect 9220 22170 9272 22176
rect 9140 22066 9260 22094
rect 8852 22024 8904 22030
rect 8852 21966 8904 21972
rect 8864 21554 8892 21966
rect 9232 21842 9260 22066
rect 9324 22030 9352 22630
rect 9508 22574 9536 22630
rect 9404 22568 9456 22574
rect 9404 22510 9456 22516
rect 9496 22568 9548 22574
rect 9496 22510 9548 22516
rect 9312 22024 9364 22030
rect 9312 21966 9364 21972
rect 9140 21814 9260 21842
rect 8852 21548 8904 21554
rect 8852 21490 8904 21496
rect 8864 21350 8892 21490
rect 8852 21344 8904 21350
rect 8852 21286 8904 21292
rect 9140 20448 9168 21814
rect 9324 21690 9352 21966
rect 9220 21684 9272 21690
rect 9220 21626 9272 21632
rect 9312 21684 9364 21690
rect 9312 21626 9364 21632
rect 9232 21570 9260 21626
rect 9416 21570 9444 22510
rect 9600 22506 9628 22918
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 9588 22500 9640 22506
rect 9588 22442 9640 22448
rect 9600 22030 9628 22442
rect 9784 22166 9812 22578
rect 9772 22160 9824 22166
rect 9772 22102 9824 22108
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 9772 22024 9824 22030
rect 9772 21966 9824 21972
rect 9232 21542 9444 21570
rect 9600 21554 9628 21966
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 9692 21554 9720 21830
rect 9784 21690 9812 21966
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9416 21010 9444 21542
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 9404 21004 9456 21010
rect 9404 20946 9456 20952
rect 9876 20602 9904 25638
rect 9968 25498 9996 26930
rect 10048 26308 10100 26314
rect 10048 26250 10100 26256
rect 9956 25492 10008 25498
rect 9956 25434 10008 25440
rect 9956 24268 10008 24274
rect 9956 24210 10008 24216
rect 9968 23866 9996 24210
rect 9956 23860 10008 23866
rect 9956 23802 10008 23808
rect 10060 22642 10088 26250
rect 10048 22636 10100 22642
rect 10048 22578 10100 22584
rect 10152 22098 10180 28614
rect 10232 28552 10284 28558
rect 10232 28494 10284 28500
rect 10244 28422 10272 28494
rect 10232 28416 10284 28422
rect 10232 28358 10284 28364
rect 10244 25226 10272 28358
rect 10324 27872 10376 27878
rect 10324 27814 10376 27820
rect 10336 27538 10364 27814
rect 10428 27674 10456 29038
rect 10508 28416 10560 28422
rect 10508 28358 10560 28364
rect 10416 27668 10468 27674
rect 10416 27610 10468 27616
rect 10324 27532 10376 27538
rect 10324 27474 10376 27480
rect 10324 27396 10376 27402
rect 10324 27338 10376 27344
rect 10336 27305 10364 27338
rect 10416 27328 10468 27334
rect 10322 27296 10378 27305
rect 10416 27270 10468 27276
rect 10322 27231 10378 27240
rect 10324 26988 10376 26994
rect 10324 26930 10376 26936
rect 10336 26353 10364 26930
rect 10322 26344 10378 26353
rect 10428 26314 10456 27270
rect 10322 26279 10378 26288
rect 10416 26308 10468 26314
rect 10416 26250 10468 26256
rect 10416 25900 10468 25906
rect 10416 25842 10468 25848
rect 10232 25220 10284 25226
rect 10232 25162 10284 25168
rect 10232 24812 10284 24818
rect 10232 24754 10284 24760
rect 10244 24206 10272 24754
rect 10232 24200 10284 24206
rect 10232 24142 10284 24148
rect 10140 22092 10192 22098
rect 10140 22034 10192 22040
rect 10048 22024 10100 22030
rect 10046 21992 10048 22001
rect 10100 21992 10102 22001
rect 10046 21927 10102 21936
rect 9864 20596 9916 20602
rect 9864 20538 9916 20544
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 9220 20460 9272 20466
rect 9140 20420 9220 20448
rect 9220 20402 9272 20408
rect 8760 19848 8812 19854
rect 8760 19790 8812 19796
rect 9036 19848 9088 19854
rect 9126 19816 9182 19825
rect 9088 19796 9126 19802
rect 9036 19790 9126 19796
rect 8772 19514 8800 19790
rect 8944 19780 8996 19786
rect 9048 19774 9126 19790
rect 9126 19751 9182 19760
rect 8944 19722 8996 19728
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 8956 19310 8984 19722
rect 8944 19304 8996 19310
rect 8944 19246 8996 19252
rect 8760 18964 8812 18970
rect 8680 18924 8760 18952
rect 8760 18906 8812 18912
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 9232 18222 9260 20402
rect 9864 20392 9916 20398
rect 9864 20334 9916 20340
rect 9404 19848 9456 19854
rect 9404 19790 9456 19796
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 9416 19514 9444 19790
rect 9496 19712 9548 19718
rect 9496 19654 9548 19660
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 9508 19378 9536 19654
rect 9496 19372 9548 19378
rect 9496 19314 9548 19320
rect 9404 19168 9456 19174
rect 9404 19110 9456 19116
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8772 17678 8800 18022
rect 8760 17672 8812 17678
rect 8760 17614 8812 17620
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8496 17338 8524 17478
rect 8588 17338 8616 17478
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8576 17332 8628 17338
rect 8576 17274 8628 17280
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8312 15706 8340 15982
rect 8956 15706 8984 16390
rect 9048 16289 9076 16526
rect 9034 16280 9090 16289
rect 9034 16215 9090 16224
rect 9048 16182 9076 16215
rect 9036 16176 9088 16182
rect 9036 16118 9088 16124
rect 9036 16040 9088 16046
rect 9140 16028 9168 17614
rect 9232 16454 9260 18158
rect 9324 17270 9352 18566
rect 9416 18222 9444 19110
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9312 17264 9364 17270
rect 9312 17206 9364 17212
rect 9508 16590 9536 19314
rect 9600 17678 9628 19790
rect 9876 19310 9904 20334
rect 9968 19854 9996 20470
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 9968 19514 9996 19790
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 9956 19304 10008 19310
rect 9956 19246 10008 19252
rect 9772 18420 9824 18426
rect 9772 18362 9824 18368
rect 9680 17808 9732 17814
rect 9680 17750 9732 17756
rect 9588 17672 9640 17678
rect 9588 17614 9640 17620
rect 9692 17202 9720 17750
rect 9784 17338 9812 18362
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9876 17218 9904 19246
rect 9968 18766 9996 19246
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9968 17746 9996 18702
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9784 17190 9904 17218
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9692 16794 9720 16934
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9220 16448 9272 16454
rect 9220 16390 9272 16396
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9088 16000 9168 16028
rect 9036 15982 9088 15988
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 8404 15026 8432 15438
rect 8760 15428 8812 15434
rect 8760 15370 8812 15376
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8496 14618 8524 14962
rect 8576 14816 8628 14822
rect 8576 14758 8628 14764
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8588 13870 8616 14758
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8668 13796 8720 13802
rect 8668 13738 8720 13744
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8312 12866 8340 13466
rect 8496 13258 8524 13670
rect 8680 13326 8708 13738
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 8404 12986 8432 13194
rect 8680 13138 8708 13262
rect 8772 13240 8800 15370
rect 9128 14884 9180 14890
rect 9128 14826 9180 14832
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 9048 14006 9076 14214
rect 8852 14000 8904 14006
rect 8852 13942 8904 13948
rect 9036 14000 9088 14006
rect 9036 13942 9088 13948
rect 8864 13394 8892 13942
rect 9140 13938 9168 14826
rect 9232 14482 9260 16390
rect 9324 16130 9352 16390
rect 9586 16280 9642 16289
rect 9586 16215 9588 16224
rect 9640 16215 9642 16224
rect 9680 16244 9732 16250
rect 9588 16186 9640 16192
rect 9680 16186 9732 16192
rect 9692 16130 9720 16186
rect 9324 16102 9720 16130
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9416 13938 9444 14758
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 9220 13864 9272 13870
rect 9496 13864 9548 13870
rect 9272 13824 9352 13852
rect 9220 13806 9272 13812
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 8772 13212 8892 13240
rect 8680 13110 8800 13138
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8496 12940 8708 12968
rect 8496 12866 8524 12940
rect 8312 12850 8524 12866
rect 8300 12844 8524 12850
rect 8352 12838 8524 12844
rect 8576 12844 8628 12850
rect 8300 12786 8352 12792
rect 8576 12786 8628 12792
rect 8208 12436 8260 12442
rect 8036 12406 8208 12434
rect 7932 11280 7984 11286
rect 8036 11268 8064 12406
rect 8208 12378 8260 12384
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8128 11354 8156 11834
rect 8300 11824 8352 11830
rect 8300 11766 8352 11772
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 7984 11240 8064 11268
rect 7932 11222 7984 11228
rect 7932 11144 7984 11150
rect 8220 11098 8248 11698
rect 8312 11354 8340 11766
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8588 11150 8616 12786
rect 7932 11086 7984 11092
rect 7944 10810 7972 11086
rect 8036 11070 8248 11098
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 8036 10690 8064 11070
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 7944 10662 8064 10690
rect 7840 9648 7892 9654
rect 7840 9590 7892 9596
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7576 9030 7788 9058
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7576 8090 7604 8298
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7472 8016 7524 8022
rect 7472 7958 7524 7964
rect 7196 7472 7248 7478
rect 7196 7414 7248 7420
rect 7668 7426 7696 8774
rect 7760 8090 7788 9030
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7852 7546 7880 9590
rect 7944 9450 7972 10662
rect 8128 10062 8156 10950
rect 8680 10674 8708 12940
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 7932 9444 7984 9450
rect 7932 9386 7984 9392
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 8036 9178 8064 9318
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8220 8974 8248 10542
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8404 10266 8432 10406
rect 8496 10266 8524 10610
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8680 9722 8708 10610
rect 8772 10198 8800 13110
rect 8760 10192 8812 10198
rect 8760 10134 8812 10140
rect 8864 10062 8892 13212
rect 8956 10674 8984 13262
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 9048 12850 9076 13126
rect 9218 13016 9274 13025
rect 9128 12980 9180 12986
rect 9218 12951 9274 12960
rect 9128 12922 9180 12928
rect 9140 12889 9168 12922
rect 9232 12918 9260 12951
rect 9220 12912 9272 12918
rect 9126 12880 9182 12889
rect 9036 12844 9088 12850
rect 9220 12854 9272 12860
rect 9126 12815 9182 12824
rect 9036 12786 9088 12792
rect 9048 12238 9076 12786
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9140 11898 9168 12174
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9324 10674 9352 13824
rect 9496 13806 9548 13812
rect 9404 13388 9456 13394
rect 9508 13376 9536 13806
rect 9456 13348 9536 13376
rect 9404 13330 9456 13336
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 9416 10674 9444 13194
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9508 10674 9536 13126
rect 9692 12850 9720 13126
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9784 12434 9812 17190
rect 9968 16658 9996 17682
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 10060 16114 10088 21927
rect 10138 20224 10194 20233
rect 10138 20159 10194 20168
rect 10152 19446 10180 20159
rect 10244 19990 10272 24142
rect 10428 22094 10456 25842
rect 10520 25294 10548 28358
rect 10690 27568 10746 27577
rect 10612 27526 10690 27554
rect 10508 25288 10560 25294
rect 10508 25230 10560 25236
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 10520 23118 10548 23666
rect 10612 23186 10640 27526
rect 10690 27503 10746 27512
rect 10796 27334 10824 32914
rect 10888 30734 10916 33390
rect 11072 31754 11100 33934
rect 11152 33380 11204 33386
rect 11152 33322 11204 33328
rect 11164 33114 11192 33322
rect 11152 33108 11204 33114
rect 11152 33050 11204 33056
rect 11072 31726 11192 31754
rect 10876 30728 10928 30734
rect 10876 30670 10928 30676
rect 11164 30666 11192 31726
rect 11152 30660 11204 30666
rect 11152 30602 11204 30608
rect 10876 30320 10928 30326
rect 10876 30262 10928 30268
rect 10784 27328 10836 27334
rect 10784 27270 10836 27276
rect 10692 27056 10744 27062
rect 10692 26998 10744 27004
rect 10704 26586 10732 26998
rect 10784 26784 10836 26790
rect 10784 26726 10836 26732
rect 10692 26580 10744 26586
rect 10692 26522 10744 26528
rect 10692 26240 10744 26246
rect 10692 26182 10744 26188
rect 10704 25378 10732 26182
rect 10796 25906 10824 26726
rect 10784 25900 10836 25906
rect 10784 25842 10836 25848
rect 10704 25362 10824 25378
rect 10704 25356 10836 25362
rect 10704 25350 10784 25356
rect 10784 25298 10836 25304
rect 10690 25256 10746 25265
rect 10690 25191 10746 25200
rect 10600 23180 10652 23186
rect 10600 23122 10652 23128
rect 10508 23112 10560 23118
rect 10508 23054 10560 23060
rect 10704 22098 10732 25191
rect 10784 22432 10836 22438
rect 10784 22374 10836 22380
rect 10336 22066 10456 22094
rect 10692 22092 10744 22098
rect 10336 20602 10364 22066
rect 10692 22034 10744 22040
rect 10600 22024 10652 22030
rect 10796 22012 10824 22374
rect 10888 22094 10916 30262
rect 11060 29164 11112 29170
rect 11060 29106 11112 29112
rect 11072 28762 11100 29106
rect 11060 28756 11112 28762
rect 11060 28698 11112 28704
rect 10968 28688 11020 28694
rect 10968 28630 11020 28636
rect 10980 28529 11008 28630
rect 11164 28608 11192 30602
rect 11256 30054 11284 34428
rect 11336 34410 11388 34416
rect 11336 33516 11388 33522
rect 11336 33458 11388 33464
rect 11348 32570 11376 33458
rect 11336 32564 11388 32570
rect 11336 32506 11388 32512
rect 11440 32450 11468 38814
rect 11624 38486 11652 39374
rect 11808 39098 11836 39510
rect 11900 39506 11928 39918
rect 11888 39500 11940 39506
rect 11888 39442 11940 39448
rect 11796 39092 11848 39098
rect 11796 39034 11848 39040
rect 11704 38956 11756 38962
rect 11704 38898 11756 38904
rect 11716 38554 11744 38898
rect 12256 38820 12308 38826
rect 12256 38762 12308 38768
rect 11704 38548 11756 38554
rect 11704 38490 11756 38496
rect 11612 38480 11664 38486
rect 11612 38422 11664 38428
rect 11520 38344 11572 38350
rect 11520 38286 11572 38292
rect 11980 38344 12032 38350
rect 11980 38286 12032 38292
rect 11532 37466 11560 38286
rect 11992 38010 12020 38286
rect 12268 38282 12296 38762
rect 12256 38276 12308 38282
rect 12256 38218 12308 38224
rect 11980 38004 12032 38010
rect 11980 37946 12032 37952
rect 11520 37460 11572 37466
rect 11520 37402 11572 37408
rect 12360 35170 12388 40326
rect 12440 37120 12492 37126
rect 12440 37062 12492 37068
rect 12452 36854 12480 37062
rect 12440 36848 12492 36854
rect 12440 36790 12492 36796
rect 12544 36174 12572 41074
rect 13268 40588 13320 40594
rect 13268 40530 13320 40536
rect 13176 39976 13228 39982
rect 13176 39918 13228 39924
rect 12624 39840 12676 39846
rect 12624 39782 12676 39788
rect 12716 39840 12768 39846
rect 12716 39782 12768 39788
rect 12636 38962 12664 39782
rect 12728 39574 12756 39782
rect 13188 39642 13216 39918
rect 12900 39636 12952 39642
rect 12900 39578 12952 39584
rect 13176 39636 13228 39642
rect 13176 39578 13228 39584
rect 12716 39568 12768 39574
rect 12716 39510 12768 39516
rect 12912 39438 12940 39578
rect 13280 39438 13308 40530
rect 13924 40118 13952 41386
rect 14384 41274 14412 41482
rect 14372 41268 14424 41274
rect 14372 41210 14424 41216
rect 16132 41138 16160 41550
rect 17408 41540 17460 41546
rect 17408 41482 17460 41488
rect 14280 41132 14332 41138
rect 14280 41074 14332 41080
rect 16120 41132 16172 41138
rect 16120 41074 16172 41080
rect 17224 41132 17276 41138
rect 17224 41074 17276 41080
rect 14188 40520 14240 40526
rect 14188 40462 14240 40468
rect 14200 40186 14228 40462
rect 14292 40390 14320 41074
rect 15384 40996 15436 41002
rect 15384 40938 15436 40944
rect 15396 40730 15424 40938
rect 16028 40928 16080 40934
rect 16028 40870 16080 40876
rect 15384 40724 15436 40730
rect 15384 40666 15436 40672
rect 15476 40724 15528 40730
rect 15476 40666 15528 40672
rect 14740 40520 14792 40526
rect 15016 40520 15068 40526
rect 14792 40480 15016 40508
rect 14740 40462 14792 40468
rect 15016 40462 15068 40468
rect 15384 40520 15436 40526
rect 15384 40462 15436 40468
rect 14280 40384 14332 40390
rect 14280 40326 14332 40332
rect 14740 40384 14792 40390
rect 14740 40326 14792 40332
rect 14188 40180 14240 40186
rect 14188 40122 14240 40128
rect 13912 40112 13964 40118
rect 13912 40054 13964 40060
rect 12900 39432 12952 39438
rect 12900 39374 12952 39380
rect 13268 39432 13320 39438
rect 13268 39374 13320 39380
rect 12912 39098 12940 39374
rect 13084 39364 13136 39370
rect 13084 39306 13136 39312
rect 12992 39296 13044 39302
rect 12992 39238 13044 39244
rect 12900 39092 12952 39098
rect 12900 39034 12952 39040
rect 13004 39030 13032 39238
rect 12992 39024 13044 39030
rect 12992 38966 13044 38972
rect 12624 38956 12676 38962
rect 12624 38898 12676 38904
rect 12900 38888 12952 38894
rect 12900 38830 12952 38836
rect 12912 38554 12940 38830
rect 12900 38548 12952 38554
rect 12900 38490 12952 38496
rect 12992 37732 13044 37738
rect 12992 37674 13044 37680
rect 12808 37120 12860 37126
rect 12808 37062 12860 37068
rect 12820 36378 12848 37062
rect 12808 36372 12860 36378
rect 12808 36314 12860 36320
rect 12716 36236 12768 36242
rect 12716 36178 12768 36184
rect 12532 36168 12584 36174
rect 12532 36110 12584 36116
rect 12268 35154 12388 35170
rect 11520 35148 11572 35154
rect 11520 35090 11572 35096
rect 12256 35148 12388 35154
rect 12308 35142 12388 35148
rect 12256 35090 12308 35096
rect 11532 34678 11560 35090
rect 11704 35080 11756 35086
rect 11610 35048 11666 35057
rect 11704 35022 11756 35028
rect 11610 34983 11666 34992
rect 11624 34950 11652 34983
rect 11612 34944 11664 34950
rect 11612 34886 11664 34892
rect 11520 34672 11572 34678
rect 11520 34614 11572 34620
rect 11532 33590 11560 34614
rect 11624 34610 11652 34886
rect 11612 34604 11664 34610
rect 11612 34546 11664 34552
rect 11520 33584 11572 33590
rect 11520 33526 11572 33532
rect 11348 32422 11468 32450
rect 11532 32450 11560 33526
rect 11624 32910 11652 34546
rect 11716 34542 11744 35022
rect 11888 34944 11940 34950
rect 11888 34886 11940 34892
rect 11900 34610 11928 34886
rect 12072 34672 12124 34678
rect 12072 34614 12124 34620
rect 11888 34604 11940 34610
rect 11888 34546 11940 34552
rect 11704 34536 11756 34542
rect 11704 34478 11756 34484
rect 11716 34202 11744 34478
rect 11704 34196 11756 34202
rect 11704 34138 11756 34144
rect 11888 33992 11940 33998
rect 11888 33934 11940 33940
rect 11900 33658 11928 33934
rect 12084 33658 12112 34614
rect 12360 34610 12388 35142
rect 12348 34604 12400 34610
rect 12348 34546 12400 34552
rect 12348 34400 12400 34406
rect 12544 34388 12572 36110
rect 12624 34604 12676 34610
rect 12624 34546 12676 34552
rect 12400 34360 12572 34388
rect 12348 34342 12400 34348
rect 11888 33652 11940 33658
rect 11888 33594 11940 33600
rect 12072 33652 12124 33658
rect 12072 33594 12124 33600
rect 12360 33318 12388 34342
rect 12636 33930 12664 34546
rect 12728 34202 12756 36178
rect 12808 34604 12860 34610
rect 12808 34546 12860 34552
rect 12716 34196 12768 34202
rect 12716 34138 12768 34144
rect 12820 33998 12848 34546
rect 12808 33992 12860 33998
rect 12808 33934 12860 33940
rect 12624 33924 12676 33930
rect 12624 33866 12676 33872
rect 12636 33658 12664 33866
rect 12624 33652 12676 33658
rect 12624 33594 12676 33600
rect 12624 33516 12676 33522
rect 12624 33458 12676 33464
rect 12348 33312 12400 33318
rect 12348 33254 12400 33260
rect 11612 32904 11664 32910
rect 11610 32872 11612 32881
rect 12072 32904 12124 32910
rect 11664 32872 11666 32881
rect 12072 32846 12124 32852
rect 11610 32807 11666 32816
rect 11980 32836 12032 32842
rect 11980 32778 12032 32784
rect 11532 32434 11928 32450
rect 11532 32428 11940 32434
rect 11532 32422 11888 32428
rect 11244 30048 11296 30054
rect 11244 29990 11296 29996
rect 11072 28580 11192 28608
rect 10966 28520 11022 28529
rect 10966 28455 11022 28464
rect 10968 28416 11020 28422
rect 10968 28358 11020 28364
rect 10980 28121 11008 28358
rect 10966 28112 11022 28121
rect 10966 28047 11022 28056
rect 10968 27668 11020 27674
rect 10968 27610 11020 27616
rect 10980 26450 11008 27610
rect 10968 26444 11020 26450
rect 10968 26386 11020 26392
rect 11072 23866 11100 28580
rect 11348 28558 11376 32422
rect 11532 31754 11560 32422
rect 11888 32370 11940 32376
rect 11612 31884 11664 31890
rect 11612 31826 11664 31832
rect 11440 31726 11560 31754
rect 11440 30666 11468 31726
rect 11624 30954 11652 31826
rect 11796 31272 11848 31278
rect 11796 31214 11848 31220
rect 11532 30926 11652 30954
rect 11808 30938 11836 31214
rect 11796 30932 11848 30938
rect 11532 30666 11560 30926
rect 11796 30874 11848 30880
rect 11612 30864 11664 30870
rect 11612 30806 11664 30812
rect 11428 30660 11480 30666
rect 11428 30602 11480 30608
rect 11520 30660 11572 30666
rect 11520 30602 11572 30608
rect 11336 28552 11388 28558
rect 11336 28494 11388 28500
rect 11152 28416 11204 28422
rect 11152 28358 11204 28364
rect 11244 28416 11296 28422
rect 11244 28358 11296 28364
rect 11164 25362 11192 28358
rect 11256 28218 11284 28358
rect 11244 28212 11296 28218
rect 11244 28154 11296 28160
rect 11348 26586 11376 28494
rect 11336 26580 11388 26586
rect 11336 26522 11388 26528
rect 11440 26466 11468 30602
rect 11532 30308 11560 30602
rect 11624 30433 11652 30806
rect 11992 30598 12020 32778
rect 12084 32570 12112 32846
rect 12072 32564 12124 32570
rect 12072 32506 12124 32512
rect 12360 32366 12388 33254
rect 12348 32360 12400 32366
rect 12348 32302 12400 32308
rect 12360 30870 12388 32302
rect 12532 32292 12584 32298
rect 12532 32234 12584 32240
rect 12440 32224 12492 32230
rect 12440 32166 12492 32172
rect 12452 31822 12480 32166
rect 12544 31822 12572 32234
rect 12636 32026 12664 33458
rect 12624 32020 12676 32026
rect 12624 31962 12676 31968
rect 12440 31816 12492 31822
rect 12440 31758 12492 31764
rect 12532 31816 12584 31822
rect 12532 31758 12584 31764
rect 12440 31680 12492 31686
rect 12440 31622 12492 31628
rect 12348 30864 12400 30870
rect 12348 30806 12400 30812
rect 12452 30734 12480 31622
rect 12072 30728 12124 30734
rect 12072 30670 12124 30676
rect 12440 30728 12492 30734
rect 12440 30670 12492 30676
rect 12532 30728 12584 30734
rect 12532 30670 12584 30676
rect 11980 30592 12032 30598
rect 11978 30560 11980 30569
rect 12032 30560 12034 30569
rect 11978 30495 12034 30504
rect 11610 30424 11666 30433
rect 11610 30359 11666 30368
rect 11532 30280 11836 30308
rect 11520 29708 11572 29714
rect 11520 29650 11572 29656
rect 11532 29238 11560 29650
rect 11704 29572 11756 29578
rect 11704 29514 11756 29520
rect 11716 29306 11744 29514
rect 11704 29300 11756 29306
rect 11704 29242 11756 29248
rect 11520 29232 11572 29238
rect 11520 29174 11572 29180
rect 11612 28960 11664 28966
rect 11612 28902 11664 28908
rect 11624 28490 11652 28902
rect 11716 28558 11744 29242
rect 11704 28552 11756 28558
rect 11704 28494 11756 28500
rect 11612 28484 11664 28490
rect 11612 28426 11664 28432
rect 11520 28416 11572 28422
rect 11808 28370 11836 30280
rect 11980 29640 12032 29646
rect 11980 29582 12032 29588
rect 11888 29572 11940 29578
rect 11888 29514 11940 29520
rect 11520 28358 11572 28364
rect 11532 28098 11560 28358
rect 11716 28342 11836 28370
rect 11532 28070 11652 28098
rect 11348 26438 11468 26466
rect 11244 26376 11296 26382
rect 11244 26318 11296 26324
rect 11256 26042 11284 26318
rect 11244 26036 11296 26042
rect 11244 25978 11296 25984
rect 11152 25356 11204 25362
rect 11152 25298 11204 25304
rect 11152 24812 11204 24818
rect 11152 24754 11204 24760
rect 11164 24342 11192 24754
rect 11152 24336 11204 24342
rect 11152 24278 11204 24284
rect 11060 23860 11112 23866
rect 11060 23802 11112 23808
rect 11244 23656 11296 23662
rect 11244 23598 11296 23604
rect 11256 22982 11284 23598
rect 11152 22976 11204 22982
rect 11152 22918 11204 22924
rect 11244 22976 11296 22982
rect 11244 22918 11296 22924
rect 10888 22066 11008 22094
rect 10876 22024 10928 22030
rect 10796 21984 10876 22012
rect 10600 21966 10652 21972
rect 10876 21966 10928 21972
rect 10416 21888 10468 21894
rect 10416 21830 10468 21836
rect 10428 21554 10456 21830
rect 10416 21548 10468 21554
rect 10416 21490 10468 21496
rect 10508 21548 10560 21554
rect 10508 21490 10560 21496
rect 10520 21146 10548 21490
rect 10508 21140 10560 21146
rect 10508 21082 10560 21088
rect 10612 20618 10640 21966
rect 10692 21956 10744 21962
rect 10692 21898 10744 21904
rect 10704 21554 10732 21898
rect 10980 21876 11008 22066
rect 11164 21962 11192 22918
rect 11256 22098 11284 22918
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 11152 21956 11204 21962
rect 11152 21898 11204 21904
rect 11244 21956 11296 21962
rect 11244 21898 11296 21904
rect 10888 21848 11008 21876
rect 10888 21622 10916 21848
rect 10876 21616 10928 21622
rect 10876 21558 10928 21564
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10876 20936 10928 20942
rect 10876 20878 10928 20884
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10428 20590 10640 20618
rect 10428 20262 10456 20590
rect 10508 20460 10560 20466
rect 10508 20402 10560 20408
rect 10416 20256 10468 20262
rect 10416 20198 10468 20204
rect 10232 19984 10284 19990
rect 10232 19926 10284 19932
rect 10416 19916 10468 19922
rect 10416 19858 10468 19864
rect 10140 19440 10192 19446
rect 10140 19382 10192 19388
rect 10230 19408 10286 19417
rect 10230 19343 10286 19352
rect 10244 19292 10272 19343
rect 10152 19264 10272 19292
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 9864 14340 9916 14346
rect 9864 14282 9916 14288
rect 9876 14074 9904 14282
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9876 13326 9904 14010
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 9876 12646 9904 12922
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9692 12406 9812 12434
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8956 9674 8984 10610
rect 9416 10554 9444 10610
rect 9232 10526 9444 10554
rect 8956 9654 9076 9674
rect 8944 9648 9076 9654
rect 8996 9646 9076 9648
rect 8944 9590 8996 9596
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 8036 7954 8064 8842
rect 8944 8832 8996 8838
rect 8944 8774 8996 8780
rect 8956 8634 8984 8774
rect 9048 8634 9076 9646
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 9140 8498 9168 9590
rect 9232 9382 9260 10526
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9324 8974 9352 10066
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9416 8922 9444 9658
rect 9508 9586 9536 10610
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9600 9654 9628 9862
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9588 9444 9640 9450
rect 9588 9386 9640 9392
rect 9600 9178 9628 9386
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9416 8906 9536 8922
rect 9416 8900 9548 8906
rect 9416 8894 9496 8900
rect 9496 8842 9548 8848
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 8116 8084 8168 8090
rect 8116 8026 8168 8032
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 8128 7886 8156 8026
rect 8208 8016 8260 8022
rect 8208 7958 8260 7964
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8128 7546 8156 7686
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 7668 7410 7788 7426
rect 7852 7410 7880 7482
rect 7668 7404 7800 7410
rect 7668 7398 7748 7404
rect 7748 7346 7800 7352
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 6564 4622 6592 6734
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6840 5914 6868 6190
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3608 3528 3660 3534
rect 20 3470 72 3476
rect 938 3496 994 3505
rect 32 800 60 3470
rect 3608 3470 3660 3476
rect 938 3431 994 3440
rect 3240 2848 3292 2854
rect 3240 2790 3292 2796
rect 3252 800 3280 2790
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 7300 2446 7328 6734
rect 7392 6730 7420 7142
rect 7484 6798 7512 7142
rect 7576 7002 7604 7278
rect 7760 7206 7788 7346
rect 8220 7342 8248 7958
rect 8312 7410 8340 8230
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8668 7812 8720 7818
rect 8668 7754 8720 7760
rect 8404 7410 8432 7754
rect 8680 7546 8708 7754
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 8220 6934 8248 7278
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7380 6724 7432 6730
rect 7380 6666 7432 6672
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7668 6458 7696 6598
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7944 6390 7972 6598
rect 7932 6384 7984 6390
rect 7932 6326 7984 6332
rect 8116 6248 8168 6254
rect 8312 6236 8340 7346
rect 8496 7206 8524 7346
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8496 6798 8524 7142
rect 8680 6798 8708 7482
rect 9140 7478 9168 8230
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8864 6798 8892 7278
rect 9692 6798 9720 12406
rect 9968 11150 9996 15302
rect 10046 12880 10102 12889
rect 10046 12815 10048 12824
rect 10100 12815 10102 12824
rect 10048 12786 10100 12792
rect 10152 12434 10180 19264
rect 10428 18426 10456 19858
rect 10520 19417 10548 20402
rect 10600 20256 10652 20262
rect 10600 20198 10652 20204
rect 10506 19408 10562 19417
rect 10506 19343 10562 19352
rect 10612 18834 10640 20198
rect 10784 19848 10836 19854
rect 10784 19790 10836 19796
rect 10796 19310 10824 19790
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10416 18420 10468 18426
rect 10416 18362 10468 18368
rect 10232 17604 10284 17610
rect 10232 17546 10284 17552
rect 10244 17338 10272 17546
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10692 17060 10744 17066
rect 10692 17002 10744 17008
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10612 14414 10640 14758
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 10244 12850 10272 13670
rect 10416 13456 10468 13462
rect 10416 13398 10468 13404
rect 10428 12986 10456 13398
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10612 13297 10640 13330
rect 10598 13288 10654 13297
rect 10598 13223 10654 13232
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10520 12986 10548 13126
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10428 12866 10456 12922
rect 10232 12844 10284 12850
rect 10428 12838 10548 12866
rect 10232 12786 10284 12792
rect 10520 12782 10548 12838
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 10232 12640 10284 12646
rect 10612 12628 10640 13126
rect 10284 12600 10640 12628
rect 10232 12582 10284 12588
rect 10704 12434 10732 17002
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10796 16658 10824 16934
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 10796 15162 10824 15302
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10796 14090 10824 14894
rect 10888 14346 10916 20878
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10980 20602 11008 20742
rect 10968 20596 11020 20602
rect 10968 20538 11020 20544
rect 11060 19984 11112 19990
rect 11060 19926 11112 19932
rect 11072 19446 11100 19926
rect 11150 19544 11206 19553
rect 11256 19530 11284 21898
rect 11348 20942 11376 26438
rect 11428 26376 11480 26382
rect 11426 26344 11428 26353
rect 11520 26376 11572 26382
rect 11480 26344 11482 26353
rect 11520 26318 11572 26324
rect 11426 26279 11482 26288
rect 11532 26042 11560 26318
rect 11520 26036 11572 26042
rect 11520 25978 11572 25984
rect 11624 25906 11652 28070
rect 11612 25900 11664 25906
rect 11612 25842 11664 25848
rect 11520 25152 11572 25158
rect 11520 25094 11572 25100
rect 11428 22228 11480 22234
rect 11428 22170 11480 22176
rect 11440 21690 11468 22170
rect 11532 22094 11560 25094
rect 11624 24993 11652 25842
rect 11610 24984 11666 24993
rect 11610 24919 11666 24928
rect 11716 24868 11744 28342
rect 11900 28150 11928 29514
rect 11992 28937 12020 29582
rect 12084 29322 12112 30670
rect 12256 29640 12308 29646
rect 12256 29582 12308 29588
rect 12084 29294 12168 29322
rect 12140 29220 12168 29294
rect 12085 29192 12168 29220
rect 12085 29186 12113 29192
rect 12084 29158 12113 29186
rect 11978 28928 12034 28937
rect 11978 28863 12034 28872
rect 11992 28558 12020 28863
rect 11980 28552 12032 28558
rect 11980 28494 12032 28500
rect 11980 28416 12032 28422
rect 11980 28358 12032 28364
rect 11888 28144 11940 28150
rect 11888 28086 11940 28092
rect 11796 27056 11848 27062
rect 11796 26998 11848 27004
rect 11808 26382 11836 26998
rect 11888 26920 11940 26926
rect 11888 26862 11940 26868
rect 11900 26586 11928 26862
rect 11888 26580 11940 26586
rect 11888 26522 11940 26528
rect 11796 26376 11848 26382
rect 11796 26318 11848 26324
rect 11796 25696 11848 25702
rect 11796 25638 11848 25644
rect 11808 25430 11836 25638
rect 11888 25492 11940 25498
rect 11888 25434 11940 25440
rect 11796 25424 11848 25430
rect 11796 25366 11848 25372
rect 11900 25294 11928 25434
rect 11888 25288 11940 25294
rect 11888 25230 11940 25236
rect 11624 24840 11744 24868
rect 11624 23050 11652 24840
rect 11992 24614 12020 28358
rect 12084 27962 12112 29158
rect 12268 28762 12296 29582
rect 12348 29504 12400 29510
rect 12348 29446 12400 29452
rect 12360 29238 12388 29446
rect 12348 29232 12400 29238
rect 12348 29174 12400 29180
rect 12256 28756 12308 28762
rect 12256 28698 12308 28704
rect 12164 28552 12216 28558
rect 12162 28520 12164 28529
rect 12216 28520 12218 28529
rect 12162 28455 12218 28464
rect 12176 28082 12204 28455
rect 12268 28082 12296 28698
rect 12164 28076 12216 28082
rect 12164 28018 12216 28024
rect 12256 28076 12308 28082
rect 12256 28018 12308 28024
rect 12084 27934 12296 27962
rect 12164 27872 12216 27878
rect 12164 27814 12216 27820
rect 12072 27056 12124 27062
rect 12070 27024 12072 27033
rect 12124 27024 12126 27033
rect 12070 26959 12126 26968
rect 12176 25294 12204 27814
rect 12072 25288 12124 25294
rect 12072 25230 12124 25236
rect 12164 25288 12216 25294
rect 12164 25230 12216 25236
rect 12084 24954 12112 25230
rect 12268 24954 12296 27934
rect 12348 27668 12400 27674
rect 12348 27610 12400 27616
rect 12360 27130 12388 27610
rect 12452 27554 12480 30670
rect 12544 30410 12572 30670
rect 12716 30592 12768 30598
rect 12716 30534 12768 30540
rect 12728 30433 12756 30534
rect 12714 30424 12770 30433
rect 12544 30382 12714 30410
rect 12714 30359 12770 30368
rect 12808 29776 12860 29782
rect 12530 29744 12586 29753
rect 12808 29718 12860 29724
rect 12530 29679 12586 29688
rect 12544 29306 12572 29679
rect 12716 29504 12768 29510
rect 12716 29446 12768 29452
rect 12532 29300 12584 29306
rect 12532 29242 12584 29248
rect 12728 29170 12756 29446
rect 12820 29170 12848 29718
rect 13004 29170 13032 37674
rect 13096 34746 13124 39306
rect 13280 38350 13308 39374
rect 13924 38962 13952 40054
rect 14200 39302 14228 40122
rect 14752 39982 14780 40326
rect 15028 40050 15056 40462
rect 15292 40384 15344 40390
rect 15292 40326 15344 40332
rect 15304 40050 15332 40326
rect 15396 40118 15424 40462
rect 15384 40112 15436 40118
rect 15384 40054 15436 40060
rect 15488 40050 15516 40666
rect 15660 40656 15712 40662
rect 15660 40598 15712 40604
rect 15568 40112 15620 40118
rect 15568 40054 15620 40060
rect 15016 40044 15068 40050
rect 15016 39986 15068 39992
rect 15292 40044 15344 40050
rect 15292 39986 15344 39992
rect 15476 40044 15528 40050
rect 15476 39986 15528 39992
rect 14740 39976 14792 39982
rect 14740 39918 14792 39924
rect 14752 39438 14780 39918
rect 15028 39642 15056 39986
rect 15016 39636 15068 39642
rect 15016 39578 15068 39584
rect 15200 39568 15252 39574
rect 15120 39516 15200 39522
rect 15120 39510 15252 39516
rect 15120 39494 15240 39510
rect 14740 39432 14792 39438
rect 14740 39374 14792 39380
rect 14188 39296 14240 39302
rect 14188 39238 14240 39244
rect 13912 38956 13964 38962
rect 13912 38898 13964 38904
rect 13268 38344 13320 38350
rect 13268 38286 13320 38292
rect 13728 37868 13780 37874
rect 13728 37810 13780 37816
rect 13740 36242 13768 37810
rect 13924 36718 13952 38898
rect 14372 38888 14424 38894
rect 14372 38830 14424 38836
rect 14280 38208 14332 38214
rect 14280 38150 14332 38156
rect 14292 37398 14320 38150
rect 14280 37392 14332 37398
rect 14280 37334 14332 37340
rect 14096 37256 14148 37262
rect 14096 37198 14148 37204
rect 14108 36854 14136 37198
rect 14280 37188 14332 37194
rect 14280 37130 14332 37136
rect 14096 36848 14148 36854
rect 14096 36790 14148 36796
rect 13912 36712 13964 36718
rect 13912 36654 13964 36660
rect 14292 36650 14320 37130
rect 14280 36644 14332 36650
rect 14280 36586 14332 36592
rect 13728 36236 13780 36242
rect 13728 36178 13780 36184
rect 13636 35624 13688 35630
rect 13636 35566 13688 35572
rect 13544 35284 13596 35290
rect 13544 35226 13596 35232
rect 13084 34740 13136 34746
rect 13084 34682 13136 34688
rect 13556 34610 13584 35226
rect 13544 34604 13596 34610
rect 13544 34546 13596 34552
rect 13556 33998 13584 34546
rect 13176 33992 13228 33998
rect 13176 33934 13228 33940
rect 13544 33992 13596 33998
rect 13544 33934 13596 33940
rect 13188 33590 13216 33934
rect 13452 33924 13504 33930
rect 13452 33866 13504 33872
rect 13464 33658 13492 33866
rect 13452 33652 13504 33658
rect 13452 33594 13504 33600
rect 13176 33584 13228 33590
rect 13176 33526 13228 33532
rect 13084 33516 13136 33522
rect 13084 33458 13136 33464
rect 13096 32026 13124 33458
rect 13084 32020 13136 32026
rect 13084 31962 13136 31968
rect 13544 31272 13596 31278
rect 13544 31214 13596 31220
rect 13556 30938 13584 31214
rect 13544 30932 13596 30938
rect 13544 30874 13596 30880
rect 13188 29702 13584 29730
rect 13188 29646 13216 29702
rect 13176 29640 13228 29646
rect 13176 29582 13228 29588
rect 13268 29640 13320 29646
rect 13268 29582 13320 29588
rect 13280 29481 13308 29582
rect 13360 29572 13412 29578
rect 13360 29514 13412 29520
rect 13266 29472 13322 29481
rect 13266 29407 13322 29416
rect 13372 29306 13400 29514
rect 13556 29306 13584 29702
rect 13360 29300 13412 29306
rect 13280 29260 13360 29288
rect 12716 29164 12768 29170
rect 12716 29106 12768 29112
rect 12808 29164 12860 29170
rect 12808 29106 12860 29112
rect 12992 29164 13044 29170
rect 12992 29106 13044 29112
rect 13176 29164 13228 29170
rect 13176 29106 13228 29112
rect 12532 28960 12584 28966
rect 12532 28902 12584 28908
rect 12544 28218 12572 28902
rect 12728 28762 12756 29106
rect 12808 29028 12860 29034
rect 13188 28994 13216 29106
rect 12808 28970 12860 28976
rect 12716 28756 12768 28762
rect 12716 28698 12768 28704
rect 12716 28552 12768 28558
rect 12622 28520 12678 28529
rect 12716 28494 12768 28500
rect 12622 28455 12678 28464
rect 12636 28422 12664 28455
rect 12624 28416 12676 28422
rect 12624 28358 12676 28364
rect 12728 28218 12756 28494
rect 12532 28212 12584 28218
rect 12532 28154 12584 28160
rect 12716 28212 12768 28218
rect 12716 28154 12768 28160
rect 12624 28076 12676 28082
rect 12624 28018 12676 28024
rect 12636 27674 12664 28018
rect 12624 27668 12676 27674
rect 12624 27610 12676 27616
rect 12820 27614 12848 28970
rect 12912 28966 13216 28994
rect 12912 28370 12940 28966
rect 13280 28676 13308 29260
rect 13360 29242 13412 29248
rect 13544 29300 13596 29306
rect 13544 29242 13596 29248
rect 13452 29164 13504 29170
rect 13452 29106 13504 29112
rect 13464 29073 13492 29106
rect 13450 29064 13506 29073
rect 13360 29028 13412 29034
rect 13450 28999 13506 29008
rect 13360 28970 13412 28976
rect 13096 28648 13308 28676
rect 13096 28558 13124 28648
rect 13084 28552 13136 28558
rect 13084 28494 13136 28500
rect 13268 28416 13320 28422
rect 12912 28342 13032 28370
rect 13268 28358 13320 28364
rect 12820 27586 12940 27614
rect 12452 27526 12664 27554
rect 12440 27464 12492 27470
rect 12440 27406 12492 27412
rect 12348 27124 12400 27130
rect 12348 27066 12400 27072
rect 12452 26976 12480 27406
rect 12530 27160 12586 27169
rect 12530 27095 12532 27104
rect 12584 27095 12586 27104
rect 12532 27066 12584 27072
rect 12532 26988 12584 26994
rect 12452 26948 12532 26976
rect 12532 26930 12584 26936
rect 12440 26852 12492 26858
rect 12440 26794 12492 26800
rect 12452 26586 12480 26794
rect 12440 26580 12492 26586
rect 12440 26522 12492 26528
rect 12544 26518 12572 26930
rect 12532 26512 12584 26518
rect 12532 26454 12584 26460
rect 12636 26466 12664 27526
rect 12808 27328 12860 27334
rect 12808 27270 12860 27276
rect 12820 27130 12848 27270
rect 12808 27124 12860 27130
rect 12808 27066 12860 27072
rect 12636 26438 12756 26466
rect 12624 26376 12676 26382
rect 12624 26318 12676 26324
rect 12532 26308 12584 26314
rect 12532 26250 12584 26256
rect 12348 26240 12400 26246
rect 12348 26182 12400 26188
rect 12360 25294 12388 26182
rect 12544 25294 12572 26250
rect 12348 25288 12400 25294
rect 12348 25230 12400 25236
rect 12532 25288 12584 25294
rect 12532 25230 12584 25236
rect 12072 24948 12124 24954
rect 12072 24890 12124 24896
rect 12256 24948 12308 24954
rect 12256 24890 12308 24896
rect 12348 24880 12400 24886
rect 12348 24822 12400 24828
rect 11980 24608 12032 24614
rect 11980 24550 12032 24556
rect 12256 24404 12308 24410
rect 12256 24346 12308 24352
rect 11796 24268 11848 24274
rect 11796 24210 11848 24216
rect 11702 23488 11758 23497
rect 11702 23423 11758 23432
rect 11612 23044 11664 23050
rect 11612 22986 11664 22992
rect 11716 22506 11744 23423
rect 11704 22500 11756 22506
rect 11704 22442 11756 22448
rect 11532 22066 11652 22094
rect 11520 21888 11572 21894
rect 11520 21830 11572 21836
rect 11532 21690 11560 21830
rect 11428 21684 11480 21690
rect 11428 21626 11480 21632
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 11624 21486 11652 22066
rect 11612 21480 11664 21486
rect 11612 21422 11664 21428
rect 11716 21298 11744 22442
rect 11440 21270 11744 21298
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 11206 19502 11284 19530
rect 11150 19479 11206 19488
rect 11060 19440 11112 19446
rect 11060 19382 11112 19388
rect 11244 17604 11296 17610
rect 11244 17546 11296 17552
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11164 16561 11192 16934
rect 11150 16552 11206 16561
rect 11256 16522 11284 17546
rect 11150 16487 11206 16496
rect 11244 16516 11296 16522
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 10980 15162 11008 15370
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 11072 15026 11100 15302
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 11164 14958 11192 16487
rect 11244 16458 11296 16464
rect 11256 16182 11284 16458
rect 11244 16176 11296 16182
rect 11244 16118 11296 16124
rect 11440 15162 11468 21270
rect 11520 21140 11572 21146
rect 11520 21082 11572 21088
rect 11532 19854 11560 21082
rect 11808 20641 11836 24210
rect 11980 24200 12032 24206
rect 11980 24142 12032 24148
rect 11992 23322 12020 24142
rect 12164 23588 12216 23594
rect 12164 23530 12216 23536
rect 11980 23316 12032 23322
rect 11980 23258 12032 23264
rect 11980 23112 12032 23118
rect 11900 23060 11980 23066
rect 11900 23054 12032 23060
rect 11900 23038 12020 23054
rect 11900 22778 11928 23038
rect 12176 22794 12204 23530
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 11992 22766 12204 22794
rect 11992 22030 12020 22766
rect 12070 22672 12126 22681
rect 12070 22607 12072 22616
rect 12124 22607 12126 22616
rect 12164 22636 12216 22642
rect 12072 22578 12124 22584
rect 12164 22578 12216 22584
rect 12176 22234 12204 22578
rect 12164 22228 12216 22234
rect 12164 22170 12216 22176
rect 12268 22094 12296 24346
rect 12360 24206 12388 24822
rect 12532 24336 12584 24342
rect 12530 24304 12532 24313
rect 12584 24304 12586 24313
rect 12530 24239 12586 24248
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12530 23488 12586 23497
rect 12530 23423 12586 23432
rect 12348 23044 12400 23050
rect 12348 22986 12400 22992
rect 12176 22066 12296 22094
rect 12176 22030 12204 22066
rect 11980 22024 12032 22030
rect 11980 21966 12032 21972
rect 12164 22024 12216 22030
rect 12164 21966 12216 21972
rect 11888 21956 11940 21962
rect 11888 21898 11940 21904
rect 11900 20806 11928 21898
rect 11992 21418 12020 21966
rect 12072 21480 12124 21486
rect 12072 21422 12124 21428
rect 11980 21412 12032 21418
rect 11980 21354 12032 21360
rect 11888 20800 11940 20806
rect 11888 20742 11940 20748
rect 11794 20632 11850 20641
rect 11794 20567 11850 20576
rect 11808 20466 11836 20567
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11704 20392 11756 20398
rect 11704 20334 11756 20340
rect 11612 20256 11664 20262
rect 11612 20198 11664 20204
rect 11520 19848 11572 19854
rect 11520 19790 11572 19796
rect 11624 18766 11652 20198
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 11612 17604 11664 17610
rect 11612 17546 11664 17552
rect 11624 15570 11652 17546
rect 11612 15564 11664 15570
rect 11612 15506 11664 15512
rect 11520 15428 11572 15434
rect 11520 15370 11572 15376
rect 11428 15156 11480 15162
rect 11428 15098 11480 15104
rect 11440 15042 11468 15098
rect 11256 15014 11468 15042
rect 11152 14952 11204 14958
rect 11152 14894 11204 14900
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 10876 14340 10928 14346
rect 10876 14282 10928 14288
rect 10980 14090 11008 14418
rect 11072 14346 11100 14758
rect 11060 14340 11112 14346
rect 11060 14282 11112 14288
rect 10796 14062 11008 14090
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10796 12918 10824 13466
rect 10784 12912 10836 12918
rect 10784 12854 10836 12860
rect 10784 12776 10836 12782
rect 10784 12718 10836 12724
rect 10060 12406 10180 12434
rect 10612 12406 10732 12434
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9784 9654 9812 10066
rect 9876 10062 9904 10950
rect 9968 10674 9996 11086
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9876 9654 9904 9862
rect 9772 9648 9824 9654
rect 9772 9590 9824 9596
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 9968 9586 9996 10610
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 9876 8974 9904 9386
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9784 8362 9812 8910
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8404 6458 8432 6598
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 9692 6322 9720 6734
rect 10060 6458 10088 12406
rect 10612 12050 10640 12406
rect 10796 12322 10824 12718
rect 10704 12294 10824 12322
rect 10704 12238 10732 12294
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10612 12022 10732 12050
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10244 11558 10272 11834
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10152 10674 10180 11154
rect 10336 11150 10364 11494
rect 10704 11218 10732 12022
rect 10888 11762 10916 14062
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 11072 12442 11100 13262
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 11164 12306 11192 13262
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 11152 12164 11204 12170
rect 11152 12106 11204 12112
rect 11058 12064 11114 12073
rect 11058 11999 11114 12008
rect 11072 11762 11100 11999
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10336 10606 10364 11086
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10428 10538 10456 10950
rect 10888 10742 10916 11698
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 10876 10736 10928 10742
rect 10876 10678 10928 10684
rect 10416 10532 10468 10538
rect 10416 10474 10468 10480
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10244 10130 10272 10406
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10324 6928 10376 6934
rect 10324 6870 10376 6876
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10336 6390 10364 6870
rect 10980 6730 11008 11154
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 11072 8974 11100 9454
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11164 8294 11192 12106
rect 11256 11370 11284 15014
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11348 11898 11376 12718
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11440 11506 11468 14758
rect 11532 12594 11560 15370
rect 11610 12744 11666 12753
rect 11610 12679 11612 12688
rect 11664 12679 11666 12688
rect 11612 12650 11664 12656
rect 11532 12566 11652 12594
rect 11440 11478 11560 11506
rect 11256 11342 11468 11370
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11256 10810 11284 10950
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11440 10266 11468 11342
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 11532 9674 11560 11478
rect 11624 11082 11652 12566
rect 11612 11076 11664 11082
rect 11612 11018 11664 11024
rect 11256 9646 11560 9674
rect 11256 9518 11284 9646
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 11610 9480 11666 9489
rect 11256 9081 11284 9454
rect 11242 9072 11298 9081
rect 11242 9007 11244 9016
rect 11296 9007 11298 9016
rect 11244 8978 11296 8984
rect 11348 8906 11376 9454
rect 11610 9415 11666 9424
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11440 8974 11468 9318
rect 11624 9178 11652 9415
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11532 8974 11560 9046
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11336 8900 11388 8906
rect 11336 8842 11388 8848
rect 11348 8634 11376 8842
rect 11532 8809 11560 8910
rect 11518 8800 11574 8809
rect 11518 8735 11574 8744
rect 11336 8628 11388 8634
rect 11716 8616 11744 20334
rect 11796 20256 11848 20262
rect 11796 20198 11848 20204
rect 11808 19718 11836 20198
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 12084 19174 12112 21422
rect 12164 20800 12216 20806
rect 12164 20742 12216 20748
rect 12176 20466 12204 20742
rect 12360 20602 12388 22986
rect 12544 22642 12572 23423
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12440 22568 12492 22574
rect 12440 22510 12492 22516
rect 12452 22030 12480 22510
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12440 20936 12492 20942
rect 12636 20924 12664 26318
rect 12728 24154 12756 26438
rect 12808 26036 12860 26042
rect 12808 25978 12860 25984
rect 12820 24886 12848 25978
rect 12808 24880 12860 24886
rect 12808 24822 12860 24828
rect 12808 24608 12860 24614
rect 12808 24550 12860 24556
rect 12820 24449 12848 24550
rect 12806 24440 12862 24449
rect 12806 24375 12862 24384
rect 12820 24274 12848 24375
rect 12912 24342 12940 27586
rect 13004 27130 13032 28342
rect 12992 27124 13044 27130
rect 12992 27066 13044 27072
rect 13004 24585 13032 27066
rect 13174 27024 13230 27033
rect 13174 26959 13176 26968
rect 13228 26959 13230 26968
rect 13176 26930 13228 26936
rect 13176 26852 13228 26858
rect 13176 26794 13228 26800
rect 13188 26058 13216 26794
rect 13280 26382 13308 28358
rect 13372 26858 13400 28970
rect 13544 28960 13596 28966
rect 13544 28902 13596 28908
rect 13452 28688 13504 28694
rect 13452 28630 13504 28636
rect 13464 28218 13492 28630
rect 13452 28212 13504 28218
rect 13452 28154 13504 28160
rect 13360 26852 13412 26858
rect 13360 26794 13412 26800
rect 13464 26382 13492 28154
rect 13556 28014 13584 28902
rect 13544 28008 13596 28014
rect 13544 27950 13596 27956
rect 13648 27946 13676 35566
rect 14280 35556 14332 35562
rect 14280 35498 14332 35504
rect 14096 34944 14148 34950
rect 14096 34886 14148 34892
rect 14108 34542 14136 34886
rect 14292 34746 14320 35498
rect 14280 34740 14332 34746
rect 14280 34682 14332 34688
rect 14096 34536 14148 34542
rect 14096 34478 14148 34484
rect 13912 33992 13964 33998
rect 13912 33934 13964 33940
rect 13924 32570 13952 33934
rect 14004 33584 14056 33590
rect 14004 33526 14056 33532
rect 14016 32842 14044 33526
rect 14004 32836 14056 32842
rect 14004 32778 14056 32784
rect 13912 32564 13964 32570
rect 13912 32506 13964 32512
rect 14016 32434 14044 32778
rect 14004 32428 14056 32434
rect 14004 32370 14056 32376
rect 14280 32360 14332 32366
rect 14280 32302 14332 32308
rect 14188 32224 14240 32230
rect 14188 32166 14240 32172
rect 14200 31822 14228 32166
rect 14188 31816 14240 31822
rect 14188 31758 14240 31764
rect 14200 31278 14228 31758
rect 14292 31346 14320 32302
rect 14384 31754 14412 38830
rect 14832 38480 14884 38486
rect 14832 38422 14884 38428
rect 14464 38344 14516 38350
rect 14464 38286 14516 38292
rect 14476 35834 14504 38286
rect 14556 37868 14608 37874
rect 14556 37810 14608 37816
rect 14740 37868 14792 37874
rect 14740 37810 14792 37816
rect 14568 37466 14596 37810
rect 14648 37664 14700 37670
rect 14648 37606 14700 37612
rect 14556 37460 14608 37466
rect 14556 37402 14608 37408
rect 14660 36718 14688 37606
rect 14752 37126 14780 37810
rect 14740 37120 14792 37126
rect 14740 37062 14792 37068
rect 14648 36712 14700 36718
rect 14844 36666 14872 38422
rect 15016 36780 15068 36786
rect 15016 36722 15068 36728
rect 14648 36654 14700 36660
rect 14752 36638 14872 36666
rect 14464 35828 14516 35834
rect 14464 35770 14516 35776
rect 14476 35306 14504 35770
rect 14476 35278 14688 35306
rect 14556 35012 14608 35018
rect 14556 34954 14608 34960
rect 14464 34672 14516 34678
rect 14464 34614 14516 34620
rect 14476 34202 14504 34614
rect 14568 34542 14596 34954
rect 14660 34610 14688 35278
rect 14648 34604 14700 34610
rect 14648 34546 14700 34552
rect 14556 34536 14608 34542
rect 14556 34478 14608 34484
rect 14464 34196 14516 34202
rect 14464 34138 14516 34144
rect 14464 33992 14516 33998
rect 14464 33934 14516 33940
rect 14556 33992 14608 33998
rect 14556 33934 14608 33940
rect 14476 33658 14504 33934
rect 14464 33652 14516 33658
rect 14464 33594 14516 33600
rect 14568 33386 14596 33934
rect 14648 33516 14700 33522
rect 14752 33504 14780 36638
rect 14832 36576 14884 36582
rect 14832 36518 14884 36524
rect 14924 36576 14976 36582
rect 14924 36518 14976 36524
rect 14844 36378 14872 36518
rect 14832 36372 14884 36378
rect 14832 36314 14884 36320
rect 14936 35698 14964 36518
rect 15028 36378 15056 36722
rect 15016 36372 15068 36378
rect 15016 36314 15068 36320
rect 14924 35692 14976 35698
rect 14924 35634 14976 35640
rect 14700 33476 14780 33504
rect 14832 33516 14884 33522
rect 14648 33458 14700 33464
rect 14832 33458 14884 33464
rect 14556 33380 14608 33386
rect 14556 33322 14608 33328
rect 14556 33108 14608 33114
rect 14556 33050 14608 33056
rect 14568 32570 14596 33050
rect 14844 32570 14872 33458
rect 14556 32564 14608 32570
rect 14556 32506 14608 32512
rect 14832 32564 14884 32570
rect 14832 32506 14884 32512
rect 14568 31890 14596 32506
rect 14936 32026 14964 35634
rect 15120 35601 15148 39494
rect 15304 39370 15332 39986
rect 15488 39438 15516 39986
rect 15476 39432 15528 39438
rect 15476 39374 15528 39380
rect 15580 39370 15608 40054
rect 15672 39914 15700 40598
rect 15844 40384 15896 40390
rect 15844 40326 15896 40332
rect 15856 40186 15884 40326
rect 15844 40180 15896 40186
rect 15844 40122 15896 40128
rect 15844 40044 15896 40050
rect 15844 39986 15896 39992
rect 15660 39908 15712 39914
rect 15660 39850 15712 39856
rect 15856 39370 15884 39986
rect 15936 39840 15988 39846
rect 15936 39782 15988 39788
rect 15292 39364 15344 39370
rect 15292 39306 15344 39312
rect 15568 39364 15620 39370
rect 15568 39306 15620 39312
rect 15844 39364 15896 39370
rect 15844 39306 15896 39312
rect 15304 37398 15332 39306
rect 15476 38888 15528 38894
rect 15476 38830 15528 38836
rect 15384 38752 15436 38758
rect 15384 38694 15436 38700
rect 15396 38282 15424 38694
rect 15384 38276 15436 38282
rect 15384 38218 15436 38224
rect 15292 37392 15344 37398
rect 15292 37334 15344 37340
rect 15200 36576 15252 36582
rect 15200 36518 15252 36524
rect 15384 36576 15436 36582
rect 15384 36518 15436 36524
rect 15106 35592 15162 35601
rect 15106 35527 15162 35536
rect 15108 35488 15160 35494
rect 15108 35430 15160 35436
rect 15120 34678 15148 35430
rect 15108 34672 15160 34678
rect 15108 34614 15160 34620
rect 15212 33930 15240 36518
rect 15396 35562 15424 36518
rect 15384 35556 15436 35562
rect 15384 35498 15436 35504
rect 15200 33924 15252 33930
rect 15200 33866 15252 33872
rect 15200 32224 15252 32230
rect 15200 32166 15252 32172
rect 15212 32026 15240 32166
rect 14924 32020 14976 32026
rect 14924 31962 14976 31968
rect 15200 32020 15252 32026
rect 15200 31962 15252 31968
rect 14936 31890 14964 31962
rect 14556 31884 14608 31890
rect 14556 31826 14608 31832
rect 14924 31884 14976 31890
rect 14924 31826 14976 31832
rect 14648 31816 14700 31822
rect 14648 31758 14700 31764
rect 14384 31726 14596 31754
rect 14464 31680 14516 31686
rect 14464 31622 14516 31628
rect 14372 31476 14424 31482
rect 14372 31418 14424 31424
rect 14280 31340 14332 31346
rect 14280 31282 14332 31288
rect 14188 31272 14240 31278
rect 14188 31214 14240 31220
rect 13820 30048 13872 30054
rect 13820 29990 13872 29996
rect 13912 30048 13964 30054
rect 13912 29990 13964 29996
rect 13832 29850 13860 29990
rect 13820 29844 13872 29850
rect 13820 29786 13872 29792
rect 13924 29646 13952 29990
rect 14384 29850 14412 31418
rect 14476 31278 14504 31622
rect 14464 31272 14516 31278
rect 14464 31214 14516 31220
rect 14372 29844 14424 29850
rect 14372 29786 14424 29792
rect 14372 29708 14424 29714
rect 14372 29650 14424 29656
rect 13912 29640 13964 29646
rect 13912 29582 13964 29588
rect 14096 29640 14148 29646
rect 14096 29582 14148 29588
rect 14002 29472 14058 29481
rect 14002 29407 14058 29416
rect 13728 29164 13780 29170
rect 13728 29106 13780 29112
rect 13636 27940 13688 27946
rect 13636 27882 13688 27888
rect 13544 27532 13596 27538
rect 13544 27474 13596 27480
rect 13556 26994 13584 27474
rect 13740 27402 13768 29106
rect 14016 28540 14044 29407
rect 14108 29306 14136 29582
rect 14384 29306 14412 29650
rect 14096 29300 14148 29306
rect 14096 29242 14148 29248
rect 14372 29300 14424 29306
rect 14372 29242 14424 29248
rect 14280 29164 14332 29170
rect 14280 29106 14332 29112
rect 14188 28960 14240 28966
rect 14188 28902 14240 28908
rect 14096 28552 14148 28558
rect 14016 28512 14096 28540
rect 14096 28494 14148 28500
rect 13820 27668 13872 27674
rect 13820 27610 13872 27616
rect 13728 27396 13780 27402
rect 13728 27338 13780 27344
rect 13740 27062 13768 27338
rect 13728 27056 13780 27062
rect 13728 26998 13780 27004
rect 13832 26994 13860 27610
rect 13912 27396 13964 27402
rect 13912 27338 13964 27344
rect 13544 26988 13596 26994
rect 13544 26930 13596 26936
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 13832 26874 13860 26930
rect 13648 26846 13860 26874
rect 13648 26586 13676 26846
rect 13924 26790 13952 27338
rect 14004 27124 14056 27130
rect 14004 27066 14056 27072
rect 13728 26784 13780 26790
rect 13726 26752 13728 26761
rect 13912 26784 13964 26790
rect 13780 26752 13782 26761
rect 13912 26726 13964 26732
rect 13726 26687 13782 26696
rect 13636 26580 13688 26586
rect 13636 26522 13688 26528
rect 13268 26376 13320 26382
rect 13268 26318 13320 26324
rect 13452 26376 13504 26382
rect 13452 26318 13504 26324
rect 13544 26376 13596 26382
rect 13544 26318 13596 26324
rect 13188 26030 13308 26058
rect 13176 25968 13228 25974
rect 13176 25910 13228 25916
rect 13188 25242 13216 25910
rect 13096 25214 13216 25242
rect 12990 24576 13046 24585
rect 12990 24511 13046 24520
rect 12900 24336 12952 24342
rect 12900 24278 12952 24284
rect 12808 24268 12860 24274
rect 12808 24210 12860 24216
rect 12728 24126 12940 24154
rect 12716 23520 12768 23526
rect 12716 23462 12768 23468
rect 12728 22642 12756 23462
rect 12716 22636 12768 22642
rect 12716 22578 12768 22584
rect 12728 22234 12756 22578
rect 12716 22228 12768 22234
rect 12716 22170 12768 22176
rect 12808 22160 12860 22166
rect 12808 22102 12860 22108
rect 12492 20896 12664 20924
rect 12440 20878 12492 20884
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 12360 20466 12388 20538
rect 12164 20460 12216 20466
rect 12164 20402 12216 20408
rect 12348 20460 12400 20466
rect 12348 20402 12400 20408
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 12176 18970 12204 20402
rect 12452 19802 12480 20878
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12624 20324 12676 20330
rect 12624 20266 12676 20272
rect 12532 20256 12584 20262
rect 12532 20198 12584 20204
rect 12544 19922 12572 20198
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12452 19774 12572 19802
rect 12348 19440 12400 19446
rect 12348 19382 12400 19388
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12360 18766 12388 19382
rect 12544 19378 12572 19774
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12348 18760 12400 18766
rect 12348 18702 12400 18708
rect 12176 17814 12204 18702
rect 12256 18624 12308 18630
rect 12256 18566 12308 18572
rect 12164 17808 12216 17814
rect 12164 17750 12216 17756
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11808 17338 11836 17478
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 12268 17134 12296 18566
rect 12440 18148 12492 18154
rect 12440 18090 12492 18096
rect 12452 17746 12480 18090
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 12544 17678 12572 19314
rect 12636 18850 12664 20266
rect 12728 19514 12756 20402
rect 12716 19508 12768 19514
rect 12716 19450 12768 19456
rect 12714 19408 12770 19417
rect 12714 19343 12770 19352
rect 12728 19310 12756 19343
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12820 18970 12848 22102
rect 12912 22094 12940 24126
rect 12992 24064 13044 24070
rect 12992 24006 13044 24012
rect 13004 23730 13032 24006
rect 13096 23866 13124 25214
rect 13280 24936 13308 26030
rect 13464 25498 13492 26318
rect 13452 25492 13504 25498
rect 13452 25434 13504 25440
rect 13556 25362 13584 26318
rect 13924 26314 13952 26726
rect 13912 26308 13964 26314
rect 13912 26250 13964 26256
rect 13636 25900 13688 25906
rect 13636 25842 13688 25848
rect 13544 25356 13596 25362
rect 13544 25298 13596 25304
rect 13544 25152 13596 25158
rect 13544 25094 13596 25100
rect 13188 24908 13308 24936
rect 13188 24682 13216 24908
rect 13268 24812 13320 24818
rect 13320 24772 13492 24800
rect 13268 24754 13320 24760
rect 13176 24676 13228 24682
rect 13176 24618 13228 24624
rect 13268 24608 13320 24614
rect 13268 24550 13320 24556
rect 13176 24336 13228 24342
rect 13176 24278 13228 24284
rect 13084 23860 13136 23866
rect 13084 23802 13136 23808
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 13096 22166 13124 23666
rect 13084 22160 13136 22166
rect 13084 22102 13136 22108
rect 12912 22080 12996 22094
rect 12912 22066 13032 22080
rect 12968 22052 13032 22066
rect 12898 21992 12954 22001
rect 12898 21927 12954 21936
rect 12912 21894 12940 21927
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 13004 21418 13032 22052
rect 13084 21956 13136 21962
rect 13084 21898 13136 21904
rect 12992 21412 13044 21418
rect 12992 21354 13044 21360
rect 13096 20534 13124 21898
rect 13084 20528 13136 20534
rect 13084 20470 13136 20476
rect 13084 20392 13136 20398
rect 13084 20334 13136 20340
rect 13096 20058 13124 20334
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 12900 19236 12952 19242
rect 12900 19178 12952 19184
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12636 18834 12756 18850
rect 12636 18828 12768 18834
rect 12636 18822 12716 18828
rect 12716 18770 12768 18776
rect 12912 18766 12940 19178
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 13188 17954 13216 24278
rect 13096 17926 13216 17954
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12544 17338 12572 17614
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 12256 17128 12308 17134
rect 12256 17070 12308 17076
rect 12084 16726 12112 17070
rect 12268 16794 12296 17070
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 12072 16720 12124 16726
rect 12072 16662 12124 16668
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12452 14482 12480 14894
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12544 14362 12572 17274
rect 13096 16182 13124 17926
rect 13188 17882 13216 17926
rect 13280 17898 13308 24550
rect 13360 24200 13412 24206
rect 13464 24188 13492 24772
rect 13412 24160 13492 24188
rect 13360 24142 13412 24148
rect 13360 22976 13412 22982
rect 13360 22918 13412 22924
rect 13372 21962 13400 22918
rect 13360 21956 13412 21962
rect 13360 21898 13412 21904
rect 13360 20392 13412 20398
rect 13360 20334 13412 20340
rect 13372 20058 13400 20334
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13360 19712 13412 19718
rect 13464 19700 13492 24160
rect 13412 19672 13492 19700
rect 13360 19654 13412 19660
rect 13372 19378 13400 19654
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 13176 17876 13228 17882
rect 13280 17870 13492 17898
rect 13176 17818 13228 17824
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 13188 16726 13216 17070
rect 13176 16720 13228 16726
rect 13176 16662 13228 16668
rect 13084 16176 13136 16182
rect 13084 16118 13136 16124
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12728 15706 12756 15846
rect 12912 15706 12940 15846
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 13268 15632 13320 15638
rect 13268 15574 13320 15580
rect 12900 15428 12952 15434
rect 12900 15370 12952 15376
rect 12912 15162 12940 15370
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12256 14340 12308 14346
rect 12256 14282 12308 14288
rect 12452 14334 12572 14362
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11992 13326 12020 14214
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12072 13796 12124 13802
rect 12072 13738 12124 13744
rect 12084 13569 12112 13738
rect 12070 13560 12126 13569
rect 12070 13495 12126 13504
rect 12176 13326 12204 13874
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 11794 13016 11850 13025
rect 11794 12951 11850 12960
rect 11808 12850 11836 12951
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11900 11082 11928 13262
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 11992 12866 12020 13126
rect 11992 12838 12112 12866
rect 12176 12850 12204 13126
rect 12084 12782 12112 12838
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 12268 11354 12296 14282
rect 12348 14000 12400 14006
rect 12348 13942 12400 13948
rect 12360 12850 12388 13942
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12268 11218 12296 11290
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 11888 11076 11940 11082
rect 11888 11018 11940 11024
rect 11900 9654 11928 11018
rect 11978 10976 12034 10985
rect 11978 10911 12034 10920
rect 11992 10810 12020 10911
rect 12176 10810 12204 11154
rect 12452 11150 12480 14334
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12544 12345 12572 13262
rect 12820 13258 12848 13874
rect 12808 13252 12860 13258
rect 12808 13194 12860 13200
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12636 12986 12664 13126
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 12636 12889 12664 12922
rect 12622 12880 12678 12889
rect 12622 12815 12678 12824
rect 12530 12336 12586 12345
rect 12530 12271 12586 12280
rect 12716 12164 12768 12170
rect 12716 12106 12768 12112
rect 12728 11898 12756 12106
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12544 11150 12572 11766
rect 12912 11286 12940 14758
rect 13176 14000 13228 14006
rect 13176 13942 13228 13948
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 13004 13462 13032 13874
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 12992 13456 13044 13462
rect 12992 13398 13044 13404
rect 13096 13394 13124 13806
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 13188 13326 13216 13942
rect 13176 13320 13228 13326
rect 13176 13262 13228 13268
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 12900 11280 12952 11286
rect 12900 11222 12952 11228
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12636 10606 12664 10950
rect 13004 10674 13032 12582
rect 13084 12164 13136 12170
rect 13280 12152 13308 15574
rect 13372 14822 13400 16050
rect 13464 15552 13492 17870
rect 13556 17678 13584 25094
rect 13648 24886 13676 25842
rect 13924 25430 13952 26250
rect 13912 25424 13964 25430
rect 13912 25366 13964 25372
rect 13912 24948 13964 24954
rect 13912 24890 13964 24896
rect 13636 24880 13688 24886
rect 13636 24822 13688 24828
rect 13648 24682 13676 24822
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 13636 24676 13688 24682
rect 13636 24618 13688 24624
rect 13636 24336 13688 24342
rect 13636 24278 13688 24284
rect 13648 23866 13676 24278
rect 13636 23860 13688 23866
rect 13636 23802 13688 23808
rect 13832 23594 13860 24754
rect 13820 23588 13872 23594
rect 13820 23530 13872 23536
rect 13818 22672 13874 22681
rect 13728 22636 13780 22642
rect 13924 22624 13952 24890
rect 14016 24410 14044 27066
rect 14108 26858 14136 28494
rect 14200 28218 14228 28902
rect 14292 28762 14320 29106
rect 14280 28756 14332 28762
rect 14280 28698 14332 28704
rect 14384 28558 14412 29242
rect 14372 28552 14424 28558
rect 14372 28494 14424 28500
rect 14188 28212 14240 28218
rect 14188 28154 14240 28160
rect 14464 28144 14516 28150
rect 14186 28112 14242 28121
rect 14464 28086 14516 28092
rect 14186 28047 14188 28056
rect 14240 28047 14242 28056
rect 14188 28018 14240 28024
rect 14200 26994 14228 28018
rect 14280 27940 14332 27946
rect 14280 27882 14332 27888
rect 14188 26988 14240 26994
rect 14188 26930 14240 26936
rect 14096 26852 14148 26858
rect 14096 26794 14148 26800
rect 14108 25974 14136 26794
rect 14096 25968 14148 25974
rect 14096 25910 14148 25916
rect 14096 25424 14148 25430
rect 14096 25366 14148 25372
rect 14004 24404 14056 24410
rect 14004 24346 14056 24352
rect 14004 24132 14056 24138
rect 14004 24074 14056 24080
rect 14016 23186 14044 24074
rect 14004 23180 14056 23186
rect 14004 23122 14056 23128
rect 14108 22642 14136 25366
rect 14200 24313 14228 26930
rect 14292 26450 14320 27882
rect 14372 27328 14424 27334
rect 14372 27270 14424 27276
rect 14384 26994 14412 27270
rect 14372 26988 14424 26994
rect 14372 26930 14424 26936
rect 14476 26874 14504 28086
rect 14568 27130 14596 31726
rect 14660 31686 14688 31758
rect 15488 31754 15516 38830
rect 15856 38010 15884 39306
rect 15948 38418 15976 39782
rect 15936 38412 15988 38418
rect 15936 38354 15988 38360
rect 15844 38004 15896 38010
rect 15844 37946 15896 37952
rect 15856 37466 15884 37946
rect 15844 37460 15896 37466
rect 15844 37402 15896 37408
rect 15752 36780 15804 36786
rect 15752 36722 15804 36728
rect 15568 35556 15620 35562
rect 15568 35498 15620 35504
rect 15580 35290 15608 35498
rect 15568 35284 15620 35290
rect 15568 35226 15620 35232
rect 15764 35086 15792 36722
rect 15844 36304 15896 36310
rect 15844 36246 15896 36252
rect 15856 35222 15884 36246
rect 15948 36174 15976 38354
rect 16040 37942 16068 40870
rect 17236 40730 17264 41074
rect 17316 41064 17368 41070
rect 17420 41052 17448 41482
rect 17512 41274 17540 42162
rect 19340 41676 19392 41682
rect 19340 41618 19392 41624
rect 18788 41608 18840 41614
rect 18788 41550 18840 41556
rect 17500 41268 17552 41274
rect 17500 41210 17552 41216
rect 17368 41024 17448 41052
rect 17316 41006 17368 41012
rect 17224 40724 17276 40730
rect 17224 40666 17276 40672
rect 16580 40588 16632 40594
rect 16580 40530 16632 40536
rect 16212 40112 16264 40118
rect 16212 40054 16264 40060
rect 16224 39642 16252 40054
rect 16396 39840 16448 39846
rect 16396 39782 16448 39788
rect 16212 39636 16264 39642
rect 16212 39578 16264 39584
rect 16408 39506 16436 39782
rect 16396 39500 16448 39506
rect 16396 39442 16448 39448
rect 16592 39098 16620 40530
rect 16948 40520 17000 40526
rect 16948 40462 17000 40468
rect 16672 39976 16724 39982
rect 16672 39918 16724 39924
rect 16684 39438 16712 39918
rect 16672 39432 16724 39438
rect 16672 39374 16724 39380
rect 16580 39092 16632 39098
rect 16580 39034 16632 39040
rect 16592 38418 16620 39034
rect 16580 38412 16632 38418
rect 16580 38354 16632 38360
rect 16028 37936 16080 37942
rect 16028 37878 16080 37884
rect 16488 37868 16540 37874
rect 16488 37810 16540 37816
rect 16500 37262 16528 37810
rect 16580 37664 16632 37670
rect 16580 37606 16632 37612
rect 16212 37256 16264 37262
rect 16212 37198 16264 37204
rect 16304 37256 16356 37262
rect 16304 37198 16356 37204
rect 16488 37256 16540 37262
rect 16488 37198 16540 37204
rect 16224 36786 16252 37198
rect 16212 36780 16264 36786
rect 16212 36722 16264 36728
rect 15936 36168 15988 36174
rect 15936 36110 15988 36116
rect 16224 36106 16252 36722
rect 16316 36378 16344 37198
rect 16500 36718 16528 37198
rect 16488 36712 16540 36718
rect 16488 36654 16540 36660
rect 16304 36372 16356 36378
rect 16304 36314 16356 36320
rect 16488 36168 16540 36174
rect 16488 36110 16540 36116
rect 16212 36100 16264 36106
rect 16212 36042 16264 36048
rect 16224 35834 16252 36042
rect 16212 35828 16264 35834
rect 16212 35770 16264 35776
rect 15936 35692 15988 35698
rect 15936 35634 15988 35640
rect 15844 35216 15896 35222
rect 15844 35158 15896 35164
rect 15752 35080 15804 35086
rect 15752 35022 15804 35028
rect 15752 33992 15804 33998
rect 15752 33934 15804 33940
rect 15660 33312 15712 33318
rect 15660 33254 15712 33260
rect 15672 32910 15700 33254
rect 15660 32904 15712 32910
rect 15660 32846 15712 32852
rect 15660 32768 15712 32774
rect 15660 32710 15712 32716
rect 15568 32496 15620 32502
rect 15568 32438 15620 32444
rect 15580 31822 15608 32438
rect 15672 32026 15700 32710
rect 15660 32020 15712 32026
rect 15660 31962 15712 31968
rect 15764 31822 15792 33934
rect 15856 33114 15884 35158
rect 15844 33108 15896 33114
rect 15844 33050 15896 33056
rect 15856 32774 15884 33050
rect 15948 32978 15976 35634
rect 16500 35494 16528 36110
rect 16488 35488 16540 35494
rect 16488 35430 16540 35436
rect 16304 35148 16356 35154
rect 16304 35090 16356 35096
rect 16212 35080 16264 35086
rect 16212 35022 16264 35028
rect 16120 34400 16172 34406
rect 16120 34342 16172 34348
rect 16132 33930 16160 34342
rect 16224 34202 16252 35022
rect 16212 34196 16264 34202
rect 16212 34138 16264 34144
rect 16316 34066 16344 35090
rect 16488 35080 16540 35086
rect 16486 35048 16488 35057
rect 16540 35048 16542 35057
rect 16486 34983 16542 34992
rect 16304 34060 16356 34066
rect 16304 34002 16356 34008
rect 16120 33924 16172 33930
rect 16120 33866 16172 33872
rect 16212 33856 16264 33862
rect 16212 33798 16264 33804
rect 16224 33522 16252 33798
rect 16120 33516 16172 33522
rect 16120 33458 16172 33464
rect 16212 33516 16264 33522
rect 16212 33458 16264 33464
rect 16028 33448 16080 33454
rect 16028 33390 16080 33396
rect 15936 32972 15988 32978
rect 15936 32914 15988 32920
rect 15936 32836 15988 32842
rect 15936 32778 15988 32784
rect 15844 32768 15896 32774
rect 15844 32710 15896 32716
rect 15948 32230 15976 32778
rect 16040 32570 16068 33390
rect 16132 33114 16160 33458
rect 16120 33108 16172 33114
rect 16120 33050 16172 33056
rect 16028 32564 16080 32570
rect 16028 32506 16080 32512
rect 16212 32360 16264 32366
rect 16212 32302 16264 32308
rect 15936 32224 15988 32230
rect 15936 32166 15988 32172
rect 15568 31816 15620 31822
rect 15568 31758 15620 31764
rect 15752 31816 15804 31822
rect 15752 31758 15804 31764
rect 15396 31726 15516 31754
rect 15660 31748 15712 31754
rect 14648 31680 14700 31686
rect 14648 31622 14700 31628
rect 14660 30802 14688 31622
rect 15108 31408 15160 31414
rect 15108 31350 15160 31356
rect 14740 31272 14792 31278
rect 14740 31214 14792 31220
rect 14648 30796 14700 30802
rect 14648 30738 14700 30744
rect 14648 29504 14700 29510
rect 14648 29446 14700 29452
rect 14556 27124 14608 27130
rect 14556 27066 14608 27072
rect 14556 26988 14608 26994
rect 14660 26976 14688 29446
rect 14608 26948 14688 26976
rect 14556 26930 14608 26936
rect 14384 26846 14504 26874
rect 14280 26444 14332 26450
rect 14280 26386 14332 26392
rect 14384 26330 14412 26846
rect 14464 26784 14516 26790
rect 14464 26726 14516 26732
rect 14476 26586 14504 26726
rect 14464 26580 14516 26586
rect 14464 26522 14516 26528
rect 14292 26302 14412 26330
rect 14292 24886 14320 26302
rect 14280 24880 14332 24886
rect 14280 24822 14332 24828
rect 14372 24880 14424 24886
rect 14372 24822 14424 24828
rect 14384 24426 14412 24822
rect 14464 24812 14516 24818
rect 14464 24754 14516 24760
rect 14476 24721 14504 24754
rect 14462 24712 14518 24721
rect 14462 24647 14518 24656
rect 14292 24398 14412 24426
rect 14462 24440 14518 24449
rect 14186 24304 14242 24313
rect 14186 24239 14242 24248
rect 13874 22616 13952 22624
rect 13818 22607 13952 22616
rect 13728 22578 13780 22584
rect 13832 22596 13952 22607
rect 14096 22636 14148 22642
rect 13740 22166 13768 22578
rect 13832 22234 13860 22596
rect 14096 22578 14148 22584
rect 13912 22500 13964 22506
rect 13912 22442 13964 22448
rect 13820 22228 13872 22234
rect 13820 22170 13872 22176
rect 13728 22160 13780 22166
rect 13728 22102 13780 22108
rect 13924 22012 13952 22442
rect 14200 22438 14228 24239
rect 14188 22432 14240 22438
rect 14188 22374 14240 22380
rect 14096 22024 14148 22030
rect 13924 21984 14096 22012
rect 14096 21966 14148 21972
rect 13912 21888 13964 21894
rect 13912 21830 13964 21836
rect 13924 21622 13952 21830
rect 13912 21616 13964 21622
rect 13912 21558 13964 21564
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 13636 21412 13688 21418
rect 13636 21354 13688 21360
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13556 16114 13584 17614
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13464 15524 13584 15552
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 13556 13734 13584 15524
rect 13648 15094 13676 21354
rect 13820 21344 13872 21350
rect 13820 21286 13872 21292
rect 13832 19825 13860 21286
rect 13912 20528 13964 20534
rect 13912 20470 13964 20476
rect 13818 19816 13874 19825
rect 13924 19786 13952 20470
rect 13818 19751 13874 19760
rect 13912 19780 13964 19786
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 13740 19242 13768 19450
rect 13728 19236 13780 19242
rect 13728 19178 13780 19184
rect 13728 17264 13780 17270
rect 13728 17206 13780 17212
rect 13740 15638 13768 17206
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13636 15088 13688 15094
rect 13636 15030 13688 15036
rect 13544 13728 13596 13734
rect 13542 13696 13544 13705
rect 13596 13696 13598 13705
rect 13542 13631 13598 13640
rect 13636 13252 13688 13258
rect 13636 13194 13688 13200
rect 13136 12124 13308 12152
rect 13084 12106 13136 12112
rect 13096 10713 13124 12106
rect 13450 10840 13506 10849
rect 13450 10775 13506 10784
rect 13082 10704 13138 10713
rect 12992 10668 13044 10674
rect 13082 10639 13138 10648
rect 12992 10610 13044 10616
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12636 10062 12664 10542
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 11888 9648 11940 9654
rect 11888 9590 11940 9596
rect 12176 9382 12204 9862
rect 12912 9722 12940 10406
rect 12900 9716 12952 9722
rect 12900 9658 12952 9664
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12544 9489 12572 9522
rect 12530 9480 12586 9489
rect 12530 9415 12586 9424
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 11978 9072 12034 9081
rect 11978 9007 12034 9016
rect 11992 8974 12020 9007
rect 12176 8974 12204 9318
rect 12268 9178 12296 9318
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 11796 8968 11848 8974
rect 11980 8968 12032 8974
rect 11848 8928 11928 8956
rect 11796 8910 11848 8916
rect 11336 8570 11388 8576
rect 11440 8588 11744 8616
rect 11440 8514 11468 8588
rect 11256 8486 11468 8514
rect 11518 8528 11574 8537
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 10968 6724 11020 6730
rect 10968 6666 11020 6672
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 10324 6384 10376 6390
rect 10324 6326 10376 6332
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 8668 6248 8720 6254
rect 8312 6208 8668 6236
rect 8116 6190 8168 6196
rect 8668 6190 8720 6196
rect 8128 5778 8156 6190
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 9692 5642 9720 6258
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9416 5370 9444 5578
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9784 5098 9812 5714
rect 10428 5370 10456 6054
rect 10888 5914 10916 6394
rect 11072 6322 11100 7958
rect 11164 7886 11192 8230
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11256 6798 11284 8486
rect 11518 8463 11520 8472
rect 11572 8463 11574 8472
rect 11612 8492 11664 8498
rect 11520 8434 11572 8440
rect 11900 8480 11928 8928
rect 11980 8910 12032 8916
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 11978 8800 12034 8809
rect 11978 8735 12034 8744
rect 11992 8634 12020 8735
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 11980 8492 12032 8498
rect 11900 8452 11980 8480
rect 11612 8434 11664 8440
rect 11980 8434 12032 8440
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11348 6798 11376 8298
rect 11428 7744 11480 7750
rect 11428 7686 11480 7692
rect 11520 7744 11572 7750
rect 11624 7732 11652 8434
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11808 7886 11836 8230
rect 12084 7886 12112 8910
rect 12728 8634 12756 9522
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12176 8378 12204 8434
rect 12176 8362 12388 8378
rect 12164 8356 12388 8362
rect 12216 8350 12388 8356
rect 12164 8298 12216 8304
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 11704 7744 11756 7750
rect 11624 7704 11704 7732
rect 11520 7686 11572 7692
rect 11704 7686 11756 7692
rect 11440 7002 11468 7686
rect 11532 7478 11560 7686
rect 11520 7472 11572 7478
rect 11520 7414 11572 7420
rect 11716 7410 11744 7686
rect 11808 7546 11836 7822
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11612 7268 11664 7274
rect 11612 7210 11664 7216
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11164 6390 11192 6598
rect 11532 6458 11560 6734
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11152 6384 11204 6390
rect 11152 6326 11204 6332
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 11164 5846 11192 6326
rect 11624 6254 11652 7210
rect 11704 6724 11756 6730
rect 11704 6666 11756 6672
rect 11716 6458 11744 6666
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11808 6322 11836 7482
rect 11900 7342 11928 7822
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 12268 7410 12296 7754
rect 12256 7404 12308 7410
rect 12360 7392 12388 8350
rect 12728 8022 12756 8570
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12728 7478 12756 7822
rect 12716 7472 12768 7478
rect 12716 7414 12768 7420
rect 12532 7404 12584 7410
rect 12360 7364 12532 7392
rect 12256 7346 12308 7352
rect 12532 7346 12584 7352
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 12268 6882 12296 7346
rect 12728 7313 12756 7414
rect 12808 7336 12860 7342
rect 12714 7304 12770 7313
rect 12808 7278 12860 7284
rect 12714 7239 12770 7248
rect 12820 7002 12848 7278
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12636 6905 12664 6938
rect 12176 6854 12296 6882
rect 12622 6896 12678 6905
rect 12072 6724 12124 6730
rect 12072 6666 12124 6672
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 11992 5370 12020 6598
rect 12084 6458 12112 6666
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 12176 6118 12204 6854
rect 12622 6831 12678 6840
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 12268 6254 12296 6666
rect 12820 6458 12848 6938
rect 12992 6724 13044 6730
rect 12992 6666 13044 6672
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12360 6066 12388 6326
rect 12820 6118 12848 6394
rect 13004 6322 13032 6666
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 12808 6112 12860 6118
rect 12360 6038 12480 6066
rect 12808 6054 12860 6060
rect 12452 5370 12480 6038
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 13096 5302 13124 10639
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 13188 9178 13216 9318
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13464 6186 13492 10775
rect 13648 10198 13676 13194
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13740 11626 13768 12106
rect 13832 12102 13860 19751
rect 13912 19722 13964 19728
rect 13924 17882 13952 19722
rect 13912 17876 13964 17882
rect 13912 17818 13964 17824
rect 13924 17270 13952 17818
rect 13912 17264 13964 17270
rect 13912 17206 13964 17212
rect 13912 16584 13964 16590
rect 13912 16526 13964 16532
rect 13924 16250 13952 16526
rect 13912 16244 13964 16250
rect 13912 16186 13964 16192
rect 14016 16130 14044 21490
rect 14096 18080 14148 18086
rect 14096 18022 14148 18028
rect 14108 17678 14136 18022
rect 14200 17746 14228 22374
rect 14292 22094 14320 24398
rect 14462 24375 14464 24384
rect 14516 24375 14518 24384
rect 14464 24346 14516 24352
rect 14372 24200 14424 24206
rect 14372 24142 14424 24148
rect 14384 23730 14412 24142
rect 14568 23798 14596 26930
rect 14648 26308 14700 26314
rect 14648 26250 14700 26256
rect 14660 24818 14688 26250
rect 14752 25362 14780 31214
rect 15120 30938 15148 31350
rect 15200 31340 15252 31346
rect 15200 31282 15252 31288
rect 15108 30932 15160 30938
rect 15108 30874 15160 30880
rect 14832 30048 14884 30054
rect 14832 29990 14884 29996
rect 14844 29646 14872 29990
rect 15016 29844 15068 29850
rect 15016 29786 15068 29792
rect 15028 29646 15056 29786
rect 14832 29640 14884 29646
rect 15016 29640 15068 29646
rect 14884 29600 14964 29628
rect 14832 29582 14884 29588
rect 14832 29164 14884 29170
rect 14832 29106 14884 29112
rect 14844 28694 14872 29106
rect 14832 28688 14884 28694
rect 14832 28630 14884 28636
rect 14844 28529 14872 28630
rect 14830 28520 14886 28529
rect 14830 28455 14886 28464
rect 14936 28422 14964 29600
rect 15016 29582 15068 29588
rect 15028 29186 15056 29582
rect 15108 29572 15160 29578
rect 15108 29514 15160 29520
rect 15120 29306 15148 29514
rect 15108 29300 15160 29306
rect 15108 29242 15160 29248
rect 15028 29170 15148 29186
rect 15028 29164 15160 29170
rect 15028 29158 15108 29164
rect 15108 29106 15160 29112
rect 15016 29096 15068 29102
rect 15016 29038 15068 29044
rect 15028 28762 15056 29038
rect 15108 29028 15160 29034
rect 15108 28970 15160 28976
rect 15016 28756 15068 28762
rect 15016 28698 15068 28704
rect 15120 28558 15148 28970
rect 15016 28552 15068 28558
rect 15016 28494 15068 28500
rect 15108 28552 15160 28558
rect 15108 28494 15160 28500
rect 14832 28416 14884 28422
rect 14832 28358 14884 28364
rect 14924 28416 14976 28422
rect 14924 28358 14976 28364
rect 14740 25356 14792 25362
rect 14740 25298 14792 25304
rect 14844 24954 14872 28358
rect 15028 27946 15056 28494
rect 15016 27940 15068 27946
rect 15016 27882 15068 27888
rect 15120 27606 15148 28494
rect 15108 27600 15160 27606
rect 15108 27542 15160 27548
rect 14922 27160 14978 27169
rect 15120 27112 15148 27542
rect 14922 27095 14924 27104
rect 14976 27095 14978 27104
rect 14924 27066 14976 27072
rect 15028 27084 15148 27112
rect 15028 26858 15056 27084
rect 15108 26988 15160 26994
rect 15108 26930 15160 26936
rect 15016 26852 15068 26858
rect 15016 26794 15068 26800
rect 14924 26240 14976 26246
rect 14924 26182 14976 26188
rect 14832 24948 14884 24954
rect 14832 24890 14884 24896
rect 14648 24812 14700 24818
rect 14648 24754 14700 24760
rect 14740 24812 14792 24818
rect 14740 24754 14792 24760
rect 14752 24698 14780 24754
rect 14752 24670 14872 24698
rect 14648 24132 14700 24138
rect 14648 24074 14700 24080
rect 14556 23792 14608 23798
rect 14556 23734 14608 23740
rect 14372 23724 14424 23730
rect 14372 23666 14424 23672
rect 14464 23724 14516 23730
rect 14464 23666 14516 23672
rect 14476 23322 14504 23666
rect 14464 23316 14516 23322
rect 14464 23258 14516 23264
rect 14660 23118 14688 24074
rect 14648 23112 14700 23118
rect 14648 23054 14700 23060
rect 14844 23050 14872 24670
rect 14832 23044 14884 23050
rect 14832 22986 14884 22992
rect 14556 22976 14608 22982
rect 14556 22918 14608 22924
rect 14292 22066 14412 22094
rect 14278 21992 14334 22001
rect 14278 21927 14280 21936
rect 14332 21927 14334 21936
rect 14280 21898 14332 21904
rect 14292 21554 14320 21898
rect 14280 21548 14332 21554
rect 14280 21490 14332 21496
rect 14384 19718 14412 22066
rect 14464 21956 14516 21962
rect 14464 21898 14516 21904
rect 14476 21350 14504 21898
rect 14464 21344 14516 21350
rect 14464 21286 14516 21292
rect 14568 21146 14596 22918
rect 14740 22636 14792 22642
rect 14740 22578 14792 22584
rect 14752 22234 14780 22578
rect 14740 22228 14792 22234
rect 14740 22170 14792 22176
rect 14556 21140 14608 21146
rect 14556 21082 14608 21088
rect 14844 20602 14872 22986
rect 14936 22506 14964 26182
rect 15016 25696 15068 25702
rect 15016 25638 15068 25644
rect 15028 25362 15056 25638
rect 15016 25356 15068 25362
rect 15016 25298 15068 25304
rect 15120 24614 15148 26930
rect 15212 26246 15240 31282
rect 15396 29170 15424 31726
rect 15660 31690 15712 31696
rect 15476 31476 15528 31482
rect 15476 31418 15528 31424
rect 15488 31362 15516 31418
rect 15672 31362 15700 31690
rect 15948 31414 15976 32166
rect 16224 31754 16252 32302
rect 16304 32292 16356 32298
rect 16304 32234 16356 32240
rect 16316 31822 16344 32234
rect 16488 32224 16540 32230
rect 16488 32166 16540 32172
rect 16304 31816 16356 31822
rect 16304 31758 16356 31764
rect 16212 31748 16264 31754
rect 16212 31690 16264 31696
rect 16120 31680 16172 31686
rect 16120 31622 16172 31628
rect 15488 31334 15700 31362
rect 15936 31408 15988 31414
rect 15936 31350 15988 31356
rect 16132 31346 16160 31622
rect 16224 31482 16252 31690
rect 16316 31482 16344 31758
rect 16212 31476 16264 31482
rect 16212 31418 16264 31424
rect 16304 31476 16356 31482
rect 16304 31418 16356 31424
rect 16500 31346 16528 32166
rect 16120 31340 16172 31346
rect 16120 31282 16172 31288
rect 16488 31340 16540 31346
rect 16488 31282 16540 31288
rect 15568 29572 15620 29578
rect 15568 29514 15620 29520
rect 15476 29504 15528 29510
rect 15476 29446 15528 29452
rect 15384 29164 15436 29170
rect 15304 29124 15384 29152
rect 15304 26994 15332 29124
rect 15384 29106 15436 29112
rect 15488 28558 15516 29446
rect 15580 29034 15608 29514
rect 15844 29232 15896 29238
rect 15750 29200 15806 29209
rect 15660 29164 15712 29170
rect 15844 29174 15896 29180
rect 15750 29135 15806 29144
rect 15660 29106 15712 29112
rect 15568 29028 15620 29034
rect 15568 28970 15620 28976
rect 15580 28762 15608 28970
rect 15568 28756 15620 28762
rect 15568 28698 15620 28704
rect 15384 28552 15436 28558
rect 15384 28494 15436 28500
rect 15476 28552 15528 28558
rect 15476 28494 15528 28500
rect 15396 28082 15424 28494
rect 15568 28484 15620 28490
rect 15568 28426 15620 28432
rect 15580 28150 15608 28426
rect 15568 28144 15620 28150
rect 15568 28086 15620 28092
rect 15384 28076 15436 28082
rect 15384 28018 15436 28024
rect 15672 27614 15700 29106
rect 15764 29034 15792 29135
rect 15752 29028 15804 29034
rect 15752 28970 15804 28976
rect 15764 28762 15792 28970
rect 15752 28756 15804 28762
rect 15752 28698 15804 28704
rect 15856 28490 15884 29174
rect 15936 29096 15988 29102
rect 15934 29064 15936 29073
rect 15988 29064 15990 29073
rect 15934 28999 15990 29008
rect 15948 28558 15976 28999
rect 16132 28994 16160 31282
rect 16592 31210 16620 37606
rect 16856 36780 16908 36786
rect 16856 36722 16908 36728
rect 16868 36378 16896 36722
rect 16856 36372 16908 36378
rect 16856 36314 16908 36320
rect 16764 34400 16816 34406
rect 16764 34342 16816 34348
rect 16776 33998 16804 34342
rect 16764 33992 16816 33998
rect 16764 33934 16816 33940
rect 16856 33992 16908 33998
rect 16856 33934 16908 33940
rect 16868 33658 16896 33934
rect 16856 33652 16908 33658
rect 16856 33594 16908 33600
rect 16764 33516 16816 33522
rect 16764 33458 16816 33464
rect 16776 33114 16804 33458
rect 16960 33318 16988 40462
rect 17420 39982 17448 41024
rect 17592 41064 17644 41070
rect 17592 41006 17644 41012
rect 17500 40384 17552 40390
rect 17500 40326 17552 40332
rect 17408 39976 17460 39982
rect 17408 39918 17460 39924
rect 17224 39432 17276 39438
rect 17224 39374 17276 39380
rect 17236 39098 17264 39374
rect 17224 39092 17276 39098
rect 17224 39034 17276 39040
rect 17316 38888 17368 38894
rect 17316 38830 17368 38836
rect 17040 38344 17092 38350
rect 17040 38286 17092 38292
rect 17052 37942 17080 38286
rect 17328 38214 17356 38830
rect 17316 38208 17368 38214
rect 17316 38150 17368 38156
rect 17040 37936 17092 37942
rect 17040 37878 17092 37884
rect 17316 37120 17368 37126
rect 17316 37062 17368 37068
rect 17328 36582 17356 37062
rect 17040 36576 17092 36582
rect 17040 36518 17092 36524
rect 17316 36576 17368 36582
rect 17316 36518 17368 36524
rect 17052 33862 17080 36518
rect 17328 36378 17356 36518
rect 17316 36372 17368 36378
rect 17316 36314 17368 36320
rect 17316 35760 17368 35766
rect 17316 35702 17368 35708
rect 17224 35488 17276 35494
rect 17224 35430 17276 35436
rect 17236 34610 17264 35430
rect 17224 34604 17276 34610
rect 17224 34546 17276 34552
rect 17040 33856 17092 33862
rect 17040 33798 17092 33804
rect 17132 33856 17184 33862
rect 17132 33798 17184 33804
rect 17144 33658 17172 33798
rect 17132 33652 17184 33658
rect 17132 33594 17184 33600
rect 17236 33454 17264 34546
rect 17328 34474 17356 35702
rect 17408 35624 17460 35630
rect 17408 35566 17460 35572
rect 17316 34468 17368 34474
rect 17316 34410 17368 34416
rect 17316 33516 17368 33522
rect 17316 33458 17368 33464
rect 17224 33448 17276 33454
rect 17224 33390 17276 33396
rect 16948 33312 17000 33318
rect 16948 33254 17000 33260
rect 16764 33108 16816 33114
rect 16764 33050 16816 33056
rect 17328 32910 17356 33458
rect 17316 32904 17368 32910
rect 17316 32846 17368 32852
rect 17420 31958 17448 35566
rect 17512 35290 17540 40326
rect 17604 38894 17632 41006
rect 18328 40384 18380 40390
rect 18328 40326 18380 40332
rect 18340 39982 18368 40326
rect 18052 39976 18104 39982
rect 18052 39918 18104 39924
rect 18328 39976 18380 39982
rect 18328 39918 18380 39924
rect 17960 39092 18012 39098
rect 17960 39034 18012 39040
rect 17592 38888 17644 38894
rect 17592 38830 17644 38836
rect 17972 38554 18000 39034
rect 17960 38548 18012 38554
rect 17960 38490 18012 38496
rect 17592 38344 17644 38350
rect 17592 38286 17644 38292
rect 17604 36582 17632 38286
rect 17684 38276 17736 38282
rect 17684 38218 17736 38224
rect 17776 38276 17828 38282
rect 17776 38218 17828 38224
rect 17696 37670 17724 38218
rect 17788 38010 17816 38218
rect 17776 38004 17828 38010
rect 17776 37946 17828 37952
rect 17868 37936 17920 37942
rect 17868 37878 17920 37884
rect 18064 37890 18092 39918
rect 18800 39302 18828 41550
rect 19352 40610 19380 41618
rect 19444 41274 19472 42162
rect 19616 42016 19668 42022
rect 19616 41958 19668 41964
rect 19628 41682 19656 41958
rect 19996 41682 20024 43893
rect 19616 41676 19668 41682
rect 19616 41618 19668 41624
rect 19984 41676 20036 41682
rect 19984 41618 20036 41624
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19996 41274 20024 41618
rect 22100 41608 22152 41614
rect 22100 41550 22152 41556
rect 20904 41540 20956 41546
rect 20904 41482 20956 41488
rect 20916 41414 20944 41482
rect 20916 41386 21220 41414
rect 19432 41268 19484 41274
rect 19432 41210 19484 41216
rect 19984 41268 20036 41274
rect 19984 41210 20036 41216
rect 21088 41064 21140 41070
rect 21088 41006 21140 41012
rect 19352 40594 19472 40610
rect 19352 40588 19484 40594
rect 19352 40582 19432 40588
rect 19432 40530 19484 40536
rect 20720 40520 20772 40526
rect 20720 40462 20772 40468
rect 19432 40452 19484 40458
rect 19432 40394 19484 40400
rect 19444 40186 19472 40394
rect 20076 40384 20128 40390
rect 20076 40326 20128 40332
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19432 40180 19484 40186
rect 19432 40122 19484 40128
rect 19340 40112 19392 40118
rect 19340 40054 19392 40060
rect 18880 40044 18932 40050
rect 18880 39986 18932 39992
rect 18236 39296 18288 39302
rect 18236 39238 18288 39244
rect 18788 39296 18840 39302
rect 18788 39238 18840 39244
rect 18248 39030 18276 39238
rect 18800 39030 18828 39238
rect 18236 39024 18288 39030
rect 18236 38966 18288 38972
rect 18788 39024 18840 39030
rect 18788 38966 18840 38972
rect 18144 38344 18196 38350
rect 18144 38286 18196 38292
rect 18156 38010 18184 38286
rect 18604 38208 18656 38214
rect 18892 38196 18920 39986
rect 18656 38168 18920 38196
rect 18604 38150 18656 38156
rect 18144 38004 18196 38010
rect 18144 37946 18196 37952
rect 17684 37664 17736 37670
rect 17684 37606 17736 37612
rect 17684 37460 17736 37466
rect 17684 37402 17736 37408
rect 17696 36854 17724 37402
rect 17684 36848 17736 36854
rect 17684 36790 17736 36796
rect 17592 36576 17644 36582
rect 17592 36518 17644 36524
rect 17880 36106 17908 37878
rect 18064 37862 18184 37890
rect 18052 37120 18104 37126
rect 18052 37062 18104 37068
rect 18064 36786 18092 37062
rect 18052 36780 18104 36786
rect 18052 36722 18104 36728
rect 18052 36168 18104 36174
rect 18052 36110 18104 36116
rect 17868 36100 17920 36106
rect 17868 36042 17920 36048
rect 17880 35894 17908 36042
rect 17880 35866 18000 35894
rect 17972 35494 18000 35866
rect 18064 35698 18092 36110
rect 18052 35692 18104 35698
rect 18052 35634 18104 35640
rect 17960 35488 18012 35494
rect 17960 35430 18012 35436
rect 17500 35284 17552 35290
rect 17500 35226 17552 35232
rect 17684 34740 17736 34746
rect 17684 34682 17736 34688
rect 17592 34536 17644 34542
rect 17592 34478 17644 34484
rect 17408 31952 17460 31958
rect 17408 31894 17460 31900
rect 16856 31680 16908 31686
rect 16856 31622 16908 31628
rect 16580 31204 16632 31210
rect 16580 31146 16632 31152
rect 16396 31136 16448 31142
rect 16396 31078 16448 31084
rect 16408 30977 16436 31078
rect 16394 30968 16450 30977
rect 16394 30903 16450 30912
rect 16408 30802 16436 30903
rect 16396 30796 16448 30802
rect 16396 30738 16448 30744
rect 16580 30796 16632 30802
rect 16580 30738 16632 30744
rect 16396 29776 16448 29782
rect 16396 29718 16448 29724
rect 16408 29288 16436 29718
rect 16316 29260 16436 29288
rect 16212 29164 16264 29170
rect 16212 29106 16264 29112
rect 16040 28966 16160 28994
rect 15936 28552 15988 28558
rect 15936 28494 15988 28500
rect 15844 28484 15896 28490
rect 15844 28426 15896 28432
rect 15844 28076 15896 28082
rect 15844 28018 15896 28024
rect 15856 27674 15884 28018
rect 15488 27586 15700 27614
rect 15844 27668 15896 27674
rect 15844 27610 15896 27616
rect 15936 27668 15988 27674
rect 15936 27610 15988 27616
rect 15382 27024 15438 27033
rect 15292 26988 15344 26994
rect 15488 26994 15516 27586
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 15568 27396 15620 27402
rect 15568 27338 15620 27344
rect 15580 26994 15608 27338
rect 15764 27130 15792 27406
rect 15948 27402 15976 27610
rect 15936 27396 15988 27402
rect 15936 27338 15988 27344
rect 15934 27160 15990 27169
rect 15752 27124 15804 27130
rect 15934 27095 15936 27104
rect 15752 27066 15804 27072
rect 15988 27095 15990 27104
rect 15936 27066 15988 27072
rect 15382 26959 15384 26968
rect 15292 26930 15344 26936
rect 15436 26959 15438 26968
rect 15476 26988 15528 26994
rect 15384 26930 15436 26936
rect 15476 26930 15528 26936
rect 15568 26988 15620 26994
rect 15568 26930 15620 26936
rect 15396 26858 15424 26930
rect 15384 26852 15436 26858
rect 15384 26794 15436 26800
rect 15200 26240 15252 26246
rect 15200 26182 15252 26188
rect 15200 25900 15252 25906
rect 15200 25842 15252 25848
rect 15212 24954 15240 25842
rect 15200 24948 15252 24954
rect 15200 24890 15252 24896
rect 15488 24614 15516 26930
rect 15752 25696 15804 25702
rect 15752 25638 15804 25644
rect 15660 25152 15712 25158
rect 15660 25094 15712 25100
rect 15672 24886 15700 25094
rect 15660 24880 15712 24886
rect 15660 24822 15712 24828
rect 15568 24744 15620 24750
rect 15568 24686 15620 24692
rect 15108 24608 15160 24614
rect 15108 24550 15160 24556
rect 15476 24608 15528 24614
rect 15476 24550 15528 24556
rect 15200 24336 15252 24342
rect 15200 24278 15252 24284
rect 15016 23860 15068 23866
rect 15016 23802 15068 23808
rect 15028 22642 15056 23802
rect 15108 23724 15160 23730
rect 15108 23666 15160 23672
rect 15016 22636 15068 22642
rect 15016 22578 15068 22584
rect 14924 22500 14976 22506
rect 14924 22442 14976 22448
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 14738 20088 14794 20097
rect 14738 20023 14794 20032
rect 14752 19922 14780 20023
rect 14844 19922 14872 20538
rect 14740 19916 14792 19922
rect 14740 19858 14792 19864
rect 14832 19916 14884 19922
rect 14832 19858 14884 19864
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 14384 18290 14412 19654
rect 14568 19446 14596 19654
rect 14556 19440 14608 19446
rect 14556 19382 14608 19388
rect 14752 19378 14780 19858
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14476 18426 14504 19246
rect 14648 19236 14700 19242
rect 14648 19178 14700 19184
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14188 17740 14240 17746
rect 14188 17682 14240 17688
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 14108 17338 14136 17478
rect 14096 17332 14148 17338
rect 14096 17274 14148 17280
rect 13924 16102 14044 16130
rect 14200 16114 14228 17682
rect 14384 17082 14412 18226
rect 14476 17338 14504 18362
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 14384 17054 14596 17082
rect 14188 16108 14240 16114
rect 13924 12209 13952 16102
rect 14188 16050 14240 16056
rect 14568 16046 14596 17054
rect 14660 16522 14688 19178
rect 14832 18896 14884 18902
rect 14832 18838 14884 18844
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14752 18222 14780 18566
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 14648 16516 14700 16522
rect 14648 16458 14700 16464
rect 14660 16250 14688 16458
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 14752 16046 14780 16730
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14464 15360 14516 15366
rect 14464 15302 14516 15308
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 14016 13258 14044 14894
rect 14292 14414 14320 15302
rect 14476 15026 14504 15302
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14004 13252 14056 13258
rect 14004 13194 14056 13200
rect 14096 13252 14148 13258
rect 14096 13194 14148 13200
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 13910 12200 13966 12209
rect 13910 12135 13966 12144
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13832 11762 13860 12038
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 14016 11676 14044 12922
rect 14108 12850 14136 13194
rect 14200 12850 14228 13194
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14292 12850 14320 13126
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14384 12322 14412 12582
rect 14292 12294 14412 12322
rect 14462 12336 14518 12345
rect 14292 12238 14320 12294
rect 14462 12271 14518 12280
rect 14476 12238 14504 12271
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14096 12164 14148 12170
rect 14096 12106 14148 12112
rect 14108 11830 14136 12106
rect 14096 11824 14148 11830
rect 14096 11766 14148 11772
rect 14016 11648 14136 11676
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13636 10192 13688 10198
rect 13636 10134 13688 10140
rect 13740 9568 13768 11562
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13832 9994 13860 10950
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13832 9586 13860 9930
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 14004 9920 14056 9926
rect 14004 9862 14056 9868
rect 13924 9586 13952 9862
rect 13648 9540 13768 9568
rect 13820 9580 13872 9586
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13556 8498 13584 9046
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13556 8022 13584 8434
rect 13648 8378 13676 9540
rect 13820 9522 13872 9528
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13740 8634 13768 9386
rect 13832 9178 13860 9522
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 14016 8974 14044 9862
rect 14108 9466 14136 11648
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14200 9586 14228 9998
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14108 9438 14320 9466
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13740 8498 13768 8570
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13648 8350 13768 8378
rect 13544 8016 13596 8022
rect 13544 7958 13596 7964
rect 13740 6882 13768 8350
rect 14016 7886 14044 8910
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 14108 7546 14136 8774
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14004 7472 14056 7478
rect 14004 7414 14056 7420
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13556 6854 13768 6882
rect 13556 6730 13584 6854
rect 13740 6798 13768 6854
rect 13636 6792 13688 6798
rect 13634 6760 13636 6769
rect 13728 6792 13780 6798
rect 13688 6760 13690 6769
rect 13544 6724 13596 6730
rect 13728 6734 13780 6740
rect 13634 6695 13690 6704
rect 13544 6666 13596 6672
rect 13648 6458 13676 6695
rect 13832 6662 13860 7210
rect 14016 6798 14044 7414
rect 14292 6866 14320 9438
rect 14372 8560 14424 8566
rect 14372 8502 14424 8508
rect 14384 7410 14412 8502
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13452 6180 13504 6186
rect 13452 6122 13504 6128
rect 14108 6118 14136 6598
rect 14384 6322 14412 7346
rect 14476 7313 14504 12174
rect 14568 11354 14596 15982
rect 14648 14544 14700 14550
rect 14648 14486 14700 14492
rect 14660 13530 14688 14486
rect 14844 13734 14872 18838
rect 14936 14618 14964 22442
rect 15016 20324 15068 20330
rect 15016 20266 15068 20272
rect 15028 15026 15056 20266
rect 15120 19242 15148 23666
rect 15212 23050 15240 24278
rect 15384 24064 15436 24070
rect 15384 24006 15436 24012
rect 15396 23798 15424 24006
rect 15384 23792 15436 23798
rect 15384 23734 15436 23740
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 15200 23044 15252 23050
rect 15200 22986 15252 22992
rect 15488 22710 15516 23666
rect 15476 22704 15528 22710
rect 15476 22646 15528 22652
rect 15384 21480 15436 21486
rect 15384 21422 15436 21428
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15396 21010 15424 21422
rect 15488 21078 15516 21422
rect 15580 21146 15608 24686
rect 15672 23798 15700 24822
rect 15764 24750 15792 25638
rect 15752 24744 15804 24750
rect 15752 24686 15804 24692
rect 15844 24064 15896 24070
rect 15842 24032 15844 24041
rect 15896 24032 15898 24041
rect 15842 23967 15898 23976
rect 15660 23792 15712 23798
rect 15660 23734 15712 23740
rect 15672 22642 15700 23734
rect 15844 23724 15896 23730
rect 15844 23666 15896 23672
rect 15856 23322 15884 23666
rect 15844 23316 15896 23322
rect 15844 23258 15896 23264
rect 15752 23112 15804 23118
rect 15752 23054 15804 23060
rect 15936 23112 15988 23118
rect 15936 23054 15988 23060
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 15764 22506 15792 23054
rect 15948 22794 15976 23054
rect 16040 22953 16068 28966
rect 16224 28762 16252 29106
rect 16212 28756 16264 28762
rect 16212 28698 16264 28704
rect 16212 27464 16264 27470
rect 16212 27406 16264 27412
rect 16224 27044 16252 27406
rect 16316 27169 16344 29260
rect 16486 29200 16542 29209
rect 16486 29135 16488 29144
rect 16540 29135 16542 29144
rect 16488 29106 16540 29112
rect 16592 28994 16620 30738
rect 16868 30598 16896 31622
rect 16948 31408 17000 31414
rect 16948 31350 17000 31356
rect 17500 31408 17552 31414
rect 17500 31350 17552 31356
rect 16960 30705 16988 31350
rect 17224 31272 17276 31278
rect 17224 31214 17276 31220
rect 17236 30938 17264 31214
rect 17224 30932 17276 30938
rect 17224 30874 17276 30880
rect 17512 30870 17540 31350
rect 17132 30864 17184 30870
rect 17132 30806 17184 30812
rect 17500 30864 17552 30870
rect 17500 30806 17552 30812
rect 16946 30696 17002 30705
rect 16946 30631 17002 30640
rect 16856 30592 16908 30598
rect 16856 30534 16908 30540
rect 16948 29572 17000 29578
rect 16948 29514 17000 29520
rect 16960 29306 16988 29514
rect 16948 29300 17000 29306
rect 16948 29242 17000 29248
rect 16948 29164 17000 29170
rect 16948 29106 17000 29112
rect 16960 29034 16988 29106
rect 16408 28966 16620 28994
rect 16948 29028 17000 29034
rect 16948 28970 17000 28976
rect 17040 29028 17092 29034
rect 17040 28970 17092 28976
rect 16302 27160 16358 27169
rect 16302 27095 16358 27104
rect 16408 27044 16436 28966
rect 17052 28762 17080 28970
rect 17040 28756 17092 28762
rect 17040 28698 17092 28704
rect 16946 28112 17002 28121
rect 16946 28047 17002 28056
rect 16486 27568 16542 27577
rect 16486 27503 16542 27512
rect 16224 27016 16436 27044
rect 16304 26852 16356 26858
rect 16304 26794 16356 26800
rect 16212 26376 16264 26382
rect 16316 26353 16344 26794
rect 16408 26466 16436 27016
rect 16500 26586 16528 27503
rect 16580 27464 16632 27470
rect 16580 27406 16632 27412
rect 16764 27464 16816 27470
rect 16764 27406 16816 27412
rect 16592 27130 16620 27406
rect 16580 27124 16632 27130
rect 16580 27066 16632 27072
rect 16592 26790 16620 27066
rect 16670 26888 16726 26897
rect 16670 26823 16726 26832
rect 16580 26784 16632 26790
rect 16580 26726 16632 26732
rect 16684 26586 16712 26823
rect 16776 26586 16804 27406
rect 16488 26580 16540 26586
rect 16488 26522 16540 26528
rect 16672 26580 16724 26586
rect 16672 26522 16724 26528
rect 16764 26580 16816 26586
rect 16764 26522 16816 26528
rect 16408 26438 16620 26466
rect 16212 26318 16264 26324
rect 16302 26344 16358 26353
rect 16224 26234 16252 26318
rect 16302 26279 16358 26288
rect 16224 26206 16344 26234
rect 16212 24200 16264 24206
rect 16212 24142 16264 24148
rect 16120 23180 16172 23186
rect 16120 23122 16172 23128
rect 16026 22944 16082 22953
rect 16026 22879 16082 22888
rect 15948 22766 16068 22794
rect 16040 22710 16068 22766
rect 16028 22704 16080 22710
rect 16028 22646 16080 22652
rect 15844 22636 15896 22642
rect 15844 22578 15896 22584
rect 15936 22636 15988 22642
rect 15936 22578 15988 22584
rect 15752 22500 15804 22506
rect 15752 22442 15804 22448
rect 15764 21690 15792 22442
rect 15752 21684 15804 21690
rect 15752 21626 15804 21632
rect 15660 21616 15712 21622
rect 15660 21558 15712 21564
rect 15568 21140 15620 21146
rect 15568 21082 15620 21088
rect 15476 21072 15528 21078
rect 15476 21014 15528 21020
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 15396 20466 15424 20946
rect 15488 20466 15516 21014
rect 15672 20874 15700 21558
rect 15752 21480 15804 21486
rect 15752 21422 15804 21428
rect 15764 21350 15792 21422
rect 15752 21344 15804 21350
rect 15752 21286 15804 21292
rect 15764 21078 15792 21286
rect 15752 21072 15804 21078
rect 15752 21014 15804 21020
rect 15660 20868 15712 20874
rect 15660 20810 15712 20816
rect 15672 20534 15700 20810
rect 15764 20806 15792 21014
rect 15752 20800 15804 20806
rect 15752 20742 15804 20748
rect 15764 20534 15792 20742
rect 15660 20528 15712 20534
rect 15660 20470 15712 20476
rect 15752 20528 15804 20534
rect 15752 20470 15804 20476
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 15856 20398 15884 22578
rect 15948 20602 15976 22578
rect 16132 22420 16160 23122
rect 16224 22982 16252 24142
rect 16316 23186 16344 26206
rect 16486 24712 16542 24721
rect 16408 24670 16486 24698
rect 16408 23848 16436 24670
rect 16486 24647 16542 24656
rect 16488 24200 16540 24206
rect 16486 24168 16488 24177
rect 16540 24168 16542 24177
rect 16486 24103 16542 24112
rect 16408 23820 16528 23848
rect 16304 23180 16356 23186
rect 16500 23168 16528 23820
rect 16592 23730 16620 26438
rect 16960 25906 16988 28047
rect 17040 26512 17092 26518
rect 17040 26454 17092 26460
rect 16948 25900 17000 25906
rect 16948 25842 17000 25848
rect 16672 25220 16724 25226
rect 16672 25162 16724 25168
rect 16580 23724 16632 23730
rect 16580 23666 16632 23672
rect 16684 23474 16712 25162
rect 17052 24818 17080 26454
rect 17144 25294 17172 30806
rect 17604 30802 17632 34478
rect 17696 33658 17724 34682
rect 17868 34604 17920 34610
rect 17868 34546 17920 34552
rect 17776 34536 17828 34542
rect 17776 34478 17828 34484
rect 17788 33658 17816 34478
rect 17880 33658 17908 34546
rect 17684 33652 17736 33658
rect 17684 33594 17736 33600
rect 17776 33652 17828 33658
rect 17776 33594 17828 33600
rect 17868 33652 17920 33658
rect 17868 33594 17920 33600
rect 17880 33538 17908 33594
rect 17696 33510 17908 33538
rect 17592 30796 17644 30802
rect 17592 30738 17644 30744
rect 17696 30569 17724 33510
rect 17868 33380 17920 33386
rect 17868 33322 17920 33328
rect 17682 30560 17738 30569
rect 17682 30495 17738 30504
rect 17684 29504 17736 29510
rect 17684 29446 17736 29452
rect 17696 29306 17724 29446
rect 17684 29300 17736 29306
rect 17684 29242 17736 29248
rect 17500 29232 17552 29238
rect 17500 29174 17552 29180
rect 17224 29164 17276 29170
rect 17224 29106 17276 29112
rect 17408 29164 17460 29170
rect 17408 29106 17460 29112
rect 17236 27946 17264 29106
rect 17420 28558 17448 29106
rect 17408 28552 17460 28558
rect 17408 28494 17460 28500
rect 17512 28490 17540 29174
rect 17592 29028 17644 29034
rect 17592 28970 17644 28976
rect 17500 28484 17552 28490
rect 17500 28426 17552 28432
rect 17408 28416 17460 28422
rect 17604 28370 17632 28970
rect 17684 28756 17736 28762
rect 17684 28698 17736 28704
rect 17696 28490 17724 28698
rect 17684 28484 17736 28490
rect 17684 28426 17736 28432
rect 17460 28364 17632 28370
rect 17408 28358 17632 28364
rect 17420 28342 17632 28358
rect 17224 27940 17276 27946
rect 17224 27882 17276 27888
rect 17132 25288 17184 25294
rect 17132 25230 17184 25236
rect 17040 24812 17092 24818
rect 17040 24754 17092 24760
rect 17040 24608 17092 24614
rect 17040 24550 17092 24556
rect 17316 24608 17368 24614
rect 17316 24550 17368 24556
rect 16684 23446 16896 23474
rect 16500 23140 16620 23168
rect 16304 23122 16356 23128
rect 16488 23044 16540 23050
rect 16488 22986 16540 22992
rect 16212 22976 16264 22982
rect 16212 22918 16264 22924
rect 16394 22944 16450 22953
rect 16394 22879 16450 22888
rect 16304 22568 16356 22574
rect 16304 22510 16356 22516
rect 16212 22432 16264 22438
rect 16132 22392 16212 22420
rect 16212 22374 16264 22380
rect 16120 21344 16172 21350
rect 16120 21286 16172 21292
rect 16028 21072 16080 21078
rect 16028 21014 16080 21020
rect 15936 20596 15988 20602
rect 15936 20538 15988 20544
rect 15844 20392 15896 20398
rect 15844 20334 15896 20340
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 15212 19854 15240 20198
rect 16040 19854 16068 21014
rect 16132 20466 16160 21286
rect 16224 21078 16252 22374
rect 16212 21072 16264 21078
rect 16212 21014 16264 21020
rect 16210 20904 16266 20913
rect 16210 20839 16212 20848
rect 16264 20839 16266 20848
rect 16212 20810 16264 20816
rect 16210 20768 16266 20777
rect 16210 20703 16266 20712
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 15764 19378 15792 19654
rect 16040 19446 16068 19790
rect 16028 19440 16080 19446
rect 16028 19382 16080 19388
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 16118 19272 16174 19281
rect 15108 19236 15160 19242
rect 16118 19207 16174 19216
rect 15108 19178 15160 19184
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 15488 17882 15516 18226
rect 15580 18222 15608 19110
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 15948 18290 15976 18906
rect 16028 18420 16080 18426
rect 16028 18362 16080 18368
rect 16040 18290 16068 18362
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 15568 18216 15620 18222
rect 15568 18158 15620 18164
rect 15750 18184 15806 18193
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15476 17876 15528 17882
rect 15476 17818 15528 17824
rect 15304 17678 15332 17818
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15292 17536 15344 17542
rect 15292 17478 15344 17484
rect 15304 17202 15332 17478
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 15200 15632 15252 15638
rect 15200 15574 15252 15580
rect 15108 15088 15160 15094
rect 15212 15076 15240 15574
rect 15292 15496 15344 15502
rect 15290 15464 15292 15473
rect 15344 15464 15346 15473
rect 15290 15399 15346 15408
rect 15304 15162 15332 15399
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15160 15048 15240 15076
rect 15108 15030 15160 15036
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14924 14408 14976 14414
rect 15212 14396 15240 15048
rect 15580 14958 15608 18158
rect 15750 18119 15806 18128
rect 15764 18086 15792 18119
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 15764 15434 15792 18022
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 15752 15428 15804 15434
rect 15752 15370 15804 15376
rect 15856 15162 15884 16934
rect 15844 15156 15896 15162
rect 15844 15098 15896 15104
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15580 14550 15608 14894
rect 15658 14784 15714 14793
rect 15658 14719 15714 14728
rect 15568 14544 15620 14550
rect 15568 14486 15620 14492
rect 14976 14368 15608 14396
rect 14924 14350 14976 14356
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 14648 13524 14700 13530
rect 14648 13466 14700 13472
rect 14660 12850 14688 13466
rect 15304 13462 15332 14214
rect 15292 13456 15344 13462
rect 15292 13398 15344 13404
rect 15304 12918 15332 13398
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15292 12912 15344 12918
rect 15292 12854 15344 12860
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 14740 12368 14792 12374
rect 14740 12310 14792 12316
rect 14832 12368 14884 12374
rect 14832 12310 14884 12316
rect 15028 12322 15056 12786
rect 15108 12708 15160 12714
rect 15108 12650 15160 12656
rect 15120 12442 15148 12650
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 14646 12200 14702 12209
rect 14646 12135 14702 12144
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14660 8537 14688 12135
rect 14752 11830 14780 12310
rect 14740 11824 14792 11830
rect 14740 11766 14792 11772
rect 14844 11694 14872 12310
rect 15028 12294 15148 12322
rect 15120 12238 15148 12294
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 15106 11792 15162 11801
rect 15106 11727 15108 11736
rect 15160 11727 15162 11736
rect 15108 11698 15160 11704
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14646 8528 14702 8537
rect 14646 8463 14702 8472
rect 14844 7410 14872 8774
rect 15120 8498 15148 11698
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15212 9110 15240 9318
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 15304 8974 15332 12582
rect 15396 12442 15424 13126
rect 15474 13016 15530 13025
rect 15474 12951 15530 12960
rect 15580 12968 15608 14368
rect 15672 13326 15700 14719
rect 16040 14618 16068 18226
rect 16132 17785 16160 19207
rect 16118 17776 16174 17785
rect 16118 17711 16174 17720
rect 16224 17082 16252 20703
rect 16316 20262 16344 22510
rect 16408 21690 16436 22879
rect 16500 22778 16528 22986
rect 16488 22772 16540 22778
rect 16488 22714 16540 22720
rect 16488 22568 16540 22574
rect 16488 22510 16540 22516
rect 16500 21962 16528 22510
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 16396 21684 16448 21690
rect 16396 21626 16448 21632
rect 16408 20330 16436 21626
rect 16396 20324 16448 20330
rect 16396 20266 16448 20272
rect 16304 20256 16356 20262
rect 16304 20198 16356 20204
rect 16396 19440 16448 19446
rect 16396 19382 16448 19388
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16316 17338 16344 18226
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 16408 17202 16436 19382
rect 16592 19174 16620 23140
rect 16672 23044 16724 23050
rect 16672 22986 16724 22992
rect 16684 22642 16712 22986
rect 16764 22704 16816 22710
rect 16764 22646 16816 22652
rect 16672 22636 16724 22642
rect 16672 22578 16724 22584
rect 16776 22438 16804 22646
rect 16764 22432 16816 22438
rect 16764 22374 16816 22380
rect 16672 20868 16724 20874
rect 16672 20810 16724 20816
rect 16684 20534 16712 20810
rect 16672 20528 16724 20534
rect 16672 20470 16724 20476
rect 16580 19168 16632 19174
rect 16580 19110 16632 19116
rect 16488 18148 16540 18154
rect 16488 18090 16540 18096
rect 16500 17270 16528 18090
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16672 18080 16724 18086
rect 16672 18022 16724 18028
rect 16592 17338 16620 18022
rect 16684 17882 16712 18022
rect 16672 17876 16724 17882
rect 16672 17818 16724 17824
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16684 17270 16712 17478
rect 16488 17264 16540 17270
rect 16488 17206 16540 17212
rect 16672 17264 16724 17270
rect 16672 17206 16724 17212
rect 16396 17196 16448 17202
rect 16396 17138 16448 17144
rect 16224 17054 16436 17082
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 16132 15094 16160 15982
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16120 15088 16172 15094
rect 16120 15030 16172 15036
rect 16028 14612 16080 14618
rect 16028 14554 16080 14560
rect 15750 13560 15806 13569
rect 15750 13495 15806 13504
rect 16028 13524 16080 13530
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15304 8498 15332 8910
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 15016 7336 15068 7342
rect 14462 7304 14518 7313
rect 15016 7278 15068 7284
rect 14462 7239 14518 7248
rect 15028 6905 15056 7278
rect 15014 6896 15070 6905
rect 15014 6831 15016 6840
rect 15068 6831 15070 6840
rect 15016 6802 15068 6808
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14568 6458 14596 6598
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 15120 5846 15148 8434
rect 15488 7750 15516 12951
rect 15580 12940 15700 12968
rect 15566 12880 15622 12889
rect 15566 12815 15568 12824
rect 15620 12815 15622 12824
rect 15568 12786 15620 12792
rect 15568 11620 15620 11626
rect 15568 11562 15620 11568
rect 15580 11218 15608 11562
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15672 10538 15700 12940
rect 15764 12238 15792 13495
rect 16028 13466 16080 13472
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15856 12782 15884 13126
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15948 11354 15976 12786
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15948 9994 15976 11290
rect 16040 10554 16068 13466
rect 16118 13152 16174 13161
rect 16118 13087 16174 13096
rect 16132 12850 16160 13087
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16132 11354 16160 12786
rect 16224 12434 16252 15846
rect 16304 14952 16356 14958
rect 16304 14894 16356 14900
rect 16316 13410 16344 14894
rect 16408 14804 16436 17054
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16592 15026 16620 16594
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16488 14816 16540 14822
rect 16408 14776 16488 14804
rect 16488 14758 16540 14764
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 16394 13560 16450 13569
rect 16394 13495 16396 13504
rect 16448 13495 16450 13504
rect 16396 13466 16448 13472
rect 16316 13382 16436 13410
rect 16224 12406 16344 12434
rect 16316 11626 16344 12406
rect 16304 11620 16356 11626
rect 16304 11562 16356 11568
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16316 11150 16344 11562
rect 16408 11558 16436 13382
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 16304 11008 16356 11014
rect 16304 10950 16356 10956
rect 16040 10526 16252 10554
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 15936 9988 15988 9994
rect 15936 9930 15988 9936
rect 15844 9920 15896 9926
rect 15844 9862 15896 9868
rect 15856 9586 15884 9862
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 16040 9042 16068 10134
rect 16132 10062 16160 10406
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16132 9722 16160 9998
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 16120 9580 16172 9586
rect 16224 9568 16252 10526
rect 16316 10130 16344 10950
rect 16500 10810 16528 14554
rect 16592 14006 16620 14962
rect 16776 14090 16804 22374
rect 16868 21298 16896 23446
rect 17052 22778 17080 24550
rect 17328 24410 17356 24550
rect 17316 24404 17368 24410
rect 17316 24346 17368 24352
rect 17328 23866 17356 24346
rect 17420 24041 17448 28342
rect 17696 28014 17724 28426
rect 17684 28008 17736 28014
rect 17684 27950 17736 27956
rect 17592 27464 17644 27470
rect 17592 27406 17644 27412
rect 17604 26994 17632 27406
rect 17592 26988 17644 26994
rect 17592 26930 17644 26936
rect 17604 26314 17632 26930
rect 17592 26308 17644 26314
rect 17592 26250 17644 26256
rect 17592 25900 17644 25906
rect 17592 25842 17644 25848
rect 17500 24064 17552 24070
rect 17406 24032 17462 24041
rect 17500 24006 17552 24012
rect 17406 23967 17462 23976
rect 17316 23860 17368 23866
rect 17316 23802 17368 23808
rect 17512 23594 17540 24006
rect 17500 23588 17552 23594
rect 17500 23530 17552 23536
rect 17224 23520 17276 23526
rect 17224 23462 17276 23468
rect 17236 23050 17264 23462
rect 17500 23248 17552 23254
rect 17406 23216 17462 23225
rect 17500 23190 17552 23196
rect 17406 23151 17462 23160
rect 17420 23118 17448 23151
rect 17316 23112 17368 23118
rect 17316 23054 17368 23060
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 17224 23044 17276 23050
rect 17224 22986 17276 22992
rect 17328 22778 17356 23054
rect 17408 22976 17460 22982
rect 17408 22918 17460 22924
rect 17040 22772 17092 22778
rect 17040 22714 17092 22720
rect 17316 22772 17368 22778
rect 17316 22714 17368 22720
rect 16868 21270 16988 21298
rect 16856 21140 16908 21146
rect 16856 21082 16908 21088
rect 16868 20942 16896 21082
rect 16856 20936 16908 20942
rect 16856 20878 16908 20884
rect 16854 20632 16910 20641
rect 16960 20618 16988 21270
rect 16910 20590 16988 20618
rect 16854 20567 16910 20576
rect 16856 20256 16908 20262
rect 16856 20198 16908 20204
rect 16868 19514 16896 20198
rect 16960 19786 16988 20590
rect 16948 19780 17000 19786
rect 16948 19722 17000 19728
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16856 18828 16908 18834
rect 16856 18770 16908 18776
rect 16868 15450 16896 18770
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 16960 16114 16988 18362
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16868 15422 16988 15450
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16868 15094 16896 15302
rect 16856 15088 16908 15094
rect 16856 15030 16908 15036
rect 16960 14958 16988 15422
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16960 14618 16988 14894
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 16776 14062 16896 14090
rect 16580 14000 16632 14006
rect 16580 13942 16632 13948
rect 16592 12306 16620 13942
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16776 13841 16804 13874
rect 16762 13832 16818 13841
rect 16762 13767 16818 13776
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16684 13297 16712 13330
rect 16670 13288 16726 13297
rect 16670 13223 16726 13232
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 16592 11762 16620 12242
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16172 9540 16252 9568
rect 16120 9522 16172 9528
rect 16132 9110 16160 9522
rect 16580 9512 16632 9518
rect 16684 9466 16712 13223
rect 16868 12832 16896 14062
rect 16632 9460 16712 9466
rect 16580 9454 16712 9460
rect 16592 9438 16712 9454
rect 16776 12804 16896 12832
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 16488 9376 16540 9382
rect 16488 9318 16540 9324
rect 16120 9104 16172 9110
rect 16120 9046 16172 9052
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 16040 8498 16068 8978
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 16224 8498 16252 8910
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 16408 8430 16436 9318
rect 16500 9178 16528 9318
rect 16592 9178 16620 9438
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16776 8566 16804 12804
rect 17052 12730 17080 22714
rect 17420 22642 17448 22918
rect 17224 22636 17276 22642
rect 17408 22636 17460 22642
rect 17224 22578 17276 22584
rect 17328 22596 17408 22624
rect 17236 22438 17264 22578
rect 17224 22432 17276 22438
rect 17224 22374 17276 22380
rect 17328 22030 17356 22596
rect 17408 22578 17460 22584
rect 17408 22432 17460 22438
rect 17408 22374 17460 22380
rect 17420 22098 17448 22374
rect 17408 22092 17460 22098
rect 17408 22034 17460 22040
rect 17316 22024 17368 22030
rect 17316 21966 17368 21972
rect 17406 21992 17462 22001
rect 17406 21927 17408 21936
rect 17460 21927 17462 21936
rect 17408 21898 17460 21904
rect 17314 21176 17370 21185
rect 17314 21111 17370 21120
rect 17130 20904 17186 20913
rect 17130 20839 17186 20848
rect 17144 20806 17172 20839
rect 17132 20800 17184 20806
rect 17132 20742 17184 20748
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 17236 20058 17264 20198
rect 17328 20058 17356 21111
rect 17408 20460 17460 20466
rect 17408 20402 17460 20408
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 17316 20052 17368 20058
rect 17316 19994 17368 20000
rect 17328 19378 17356 19994
rect 17420 19514 17448 20402
rect 17512 20233 17540 23190
rect 17498 20224 17554 20233
rect 17498 20159 17554 20168
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17512 19417 17540 20159
rect 17604 19446 17632 25842
rect 17776 24676 17828 24682
rect 17776 24618 17828 24624
rect 17788 24410 17816 24618
rect 17776 24404 17828 24410
rect 17776 24346 17828 24352
rect 17684 24064 17736 24070
rect 17684 24006 17736 24012
rect 17696 23730 17724 24006
rect 17684 23724 17736 23730
rect 17684 23666 17736 23672
rect 17788 23594 17816 24346
rect 17776 23588 17828 23594
rect 17776 23530 17828 23536
rect 17684 23316 17736 23322
rect 17684 23258 17736 23264
rect 17696 21146 17724 23258
rect 17776 22024 17828 22030
rect 17776 21966 17828 21972
rect 17788 21690 17816 21966
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 17684 21140 17736 21146
rect 17684 21082 17736 21088
rect 17880 21026 17908 33322
rect 17972 32570 18000 35430
rect 18052 32768 18104 32774
rect 18052 32710 18104 32716
rect 17960 32564 18012 32570
rect 17960 32506 18012 32512
rect 18064 32502 18092 32710
rect 18052 32496 18104 32502
rect 18052 32438 18104 32444
rect 17960 30728 18012 30734
rect 17960 30670 18012 30676
rect 17972 30258 18000 30670
rect 18156 30666 18184 37862
rect 18512 37868 18564 37874
rect 18512 37810 18564 37816
rect 18328 37732 18380 37738
rect 18328 37674 18380 37680
rect 18236 37256 18288 37262
rect 18236 37198 18288 37204
rect 18248 36650 18276 37198
rect 18340 36786 18368 37674
rect 18524 37330 18552 37810
rect 18512 37324 18564 37330
rect 18512 37266 18564 37272
rect 18328 36780 18380 36786
rect 18328 36722 18380 36728
rect 18420 36780 18472 36786
rect 18420 36722 18472 36728
rect 18236 36644 18288 36650
rect 18236 36586 18288 36592
rect 18248 36106 18276 36586
rect 18432 36378 18460 36722
rect 18420 36372 18472 36378
rect 18420 36314 18472 36320
rect 18524 36310 18552 37266
rect 18616 36718 18644 38150
rect 19064 37936 19116 37942
rect 19064 37878 19116 37884
rect 19076 37262 19104 37878
rect 19248 37732 19300 37738
rect 19248 37674 19300 37680
rect 19260 37466 19288 37674
rect 19248 37460 19300 37466
rect 19248 37402 19300 37408
rect 19260 37330 19288 37402
rect 19248 37324 19300 37330
rect 19248 37266 19300 37272
rect 19064 37256 19116 37262
rect 19064 37198 19116 37204
rect 18972 37120 19024 37126
rect 18972 37062 19024 37068
rect 18604 36712 18656 36718
rect 18604 36654 18656 36660
rect 18512 36304 18564 36310
rect 18512 36246 18564 36252
rect 18236 36100 18288 36106
rect 18236 36042 18288 36048
rect 18236 34128 18288 34134
rect 18236 34070 18288 34076
rect 18248 33930 18276 34070
rect 18236 33924 18288 33930
rect 18236 33866 18288 33872
rect 18248 33590 18276 33866
rect 18616 33862 18644 36654
rect 18984 36650 19012 37062
rect 19156 36780 19208 36786
rect 19156 36722 19208 36728
rect 18972 36644 19024 36650
rect 18972 36586 19024 36592
rect 18880 36576 18932 36582
rect 18880 36518 18932 36524
rect 18892 36242 18920 36518
rect 18880 36236 18932 36242
rect 18880 36178 18932 36184
rect 18984 36174 19012 36586
rect 18972 36168 19024 36174
rect 18972 36110 19024 36116
rect 19168 35698 19196 36722
rect 19248 36168 19300 36174
rect 19248 36110 19300 36116
rect 19156 35692 19208 35698
rect 19156 35634 19208 35640
rect 19260 35630 19288 36110
rect 19248 35624 19300 35630
rect 19248 35566 19300 35572
rect 18786 35184 18842 35193
rect 18786 35119 18842 35128
rect 18696 34060 18748 34066
rect 18696 34002 18748 34008
rect 18604 33856 18656 33862
rect 18604 33798 18656 33804
rect 18236 33584 18288 33590
rect 18236 33526 18288 33532
rect 18616 33454 18644 33798
rect 18604 33448 18656 33454
rect 18604 33390 18656 33396
rect 18708 31890 18736 34002
rect 18696 31884 18748 31890
rect 18696 31826 18748 31832
rect 18708 31278 18736 31826
rect 18696 31272 18748 31278
rect 18696 31214 18748 31220
rect 18800 30682 18828 35119
rect 19064 34468 19116 34474
rect 19064 34410 19116 34416
rect 18972 34400 19024 34406
rect 18972 34342 19024 34348
rect 18984 33930 19012 34342
rect 19076 34066 19104 34410
rect 19064 34060 19116 34066
rect 19064 34002 19116 34008
rect 18972 33924 19024 33930
rect 18972 33866 19024 33872
rect 19064 33924 19116 33930
rect 19064 33866 19116 33872
rect 19076 31754 19104 33866
rect 19156 32360 19208 32366
rect 19156 32302 19208 32308
rect 18052 30660 18104 30666
rect 18052 30602 18104 30608
rect 18144 30660 18196 30666
rect 18144 30602 18196 30608
rect 18236 30660 18288 30666
rect 18236 30602 18288 30608
rect 18432 30654 18828 30682
rect 18984 31726 19104 31754
rect 18064 30394 18092 30602
rect 18052 30388 18104 30394
rect 18052 30330 18104 30336
rect 17960 30252 18012 30258
rect 17960 30194 18012 30200
rect 17972 29753 18000 30194
rect 18052 30048 18104 30054
rect 18156 30036 18184 30602
rect 18248 30258 18276 30602
rect 18236 30252 18288 30258
rect 18236 30194 18288 30200
rect 18104 30008 18184 30036
rect 18052 29990 18104 29996
rect 17958 29744 18014 29753
rect 17958 29679 18014 29688
rect 18064 28082 18092 29990
rect 18144 29640 18196 29646
rect 18144 29582 18196 29588
rect 18156 28558 18184 29582
rect 18236 29572 18288 29578
rect 18236 29514 18288 29520
rect 18248 28558 18276 29514
rect 18328 29164 18380 29170
rect 18328 29106 18380 29112
rect 18340 28665 18368 29106
rect 18432 29034 18460 30654
rect 18604 30592 18656 30598
rect 18604 30534 18656 30540
rect 18696 30592 18748 30598
rect 18984 30580 19012 31726
rect 19064 31272 19116 31278
rect 19064 31214 19116 31220
rect 19076 30938 19104 31214
rect 19168 30954 19196 32302
rect 19352 31958 19380 40054
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19432 38820 19484 38826
rect 19432 38762 19484 38768
rect 19444 37806 19472 38762
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19524 37868 19576 37874
rect 19524 37810 19576 37816
rect 19432 37800 19484 37806
rect 19432 37742 19484 37748
rect 19444 37330 19472 37742
rect 19432 37324 19484 37330
rect 19432 37266 19484 37272
rect 19536 37210 19564 37810
rect 19444 37194 19564 37210
rect 19444 37188 19576 37194
rect 19444 37182 19524 37188
rect 19444 36718 19472 37182
rect 19524 37130 19576 37136
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19432 36712 19484 36718
rect 19432 36654 19484 36660
rect 19892 36712 19944 36718
rect 19892 36654 19944 36660
rect 19444 36310 19472 36654
rect 19616 36644 19668 36650
rect 19616 36586 19668 36592
rect 19628 36310 19656 36586
rect 19904 36378 19932 36654
rect 19892 36372 19944 36378
rect 19892 36314 19944 36320
rect 19432 36304 19484 36310
rect 19432 36246 19484 36252
rect 19616 36304 19668 36310
rect 19616 36246 19668 36252
rect 19444 35834 19472 36246
rect 19984 36168 20036 36174
rect 19984 36110 20036 36116
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19432 35828 19484 35834
rect 19432 35770 19484 35776
rect 19432 35080 19484 35086
rect 19432 35022 19484 35028
rect 19444 34474 19472 35022
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19996 34746 20024 36110
rect 20088 34746 20116 40326
rect 20732 39982 20760 40462
rect 20720 39976 20772 39982
rect 20720 39918 20772 39924
rect 20732 39438 20760 39918
rect 20168 39432 20220 39438
rect 20168 39374 20220 39380
rect 20720 39432 20772 39438
rect 20720 39374 20772 39380
rect 20180 39098 20208 39374
rect 20628 39296 20680 39302
rect 20628 39238 20680 39244
rect 20168 39092 20220 39098
rect 20168 39034 20220 39040
rect 20180 38350 20208 39034
rect 20168 38344 20220 38350
rect 20168 38286 20220 38292
rect 20180 37330 20208 38286
rect 20640 38282 20668 39238
rect 20904 38752 20956 38758
rect 20904 38694 20956 38700
rect 20628 38276 20680 38282
rect 20628 38218 20680 38224
rect 20352 38208 20404 38214
rect 20352 38150 20404 38156
rect 20364 37670 20392 38150
rect 20916 37806 20944 38694
rect 20996 38276 21048 38282
rect 20996 38218 21048 38224
rect 20904 37800 20956 37806
rect 20904 37742 20956 37748
rect 20352 37664 20404 37670
rect 20352 37606 20404 37612
rect 20168 37324 20220 37330
rect 20168 37266 20220 37272
rect 20180 36854 20208 37266
rect 20168 36848 20220 36854
rect 20168 36790 20220 36796
rect 20168 36304 20220 36310
rect 20168 36246 20220 36252
rect 19984 34740 20036 34746
rect 19984 34682 20036 34688
rect 20076 34740 20128 34746
rect 20076 34682 20128 34688
rect 19892 34604 19944 34610
rect 19892 34546 19944 34552
rect 19432 34468 19484 34474
rect 19432 34410 19484 34416
rect 19444 33522 19472 34410
rect 19904 34202 19932 34546
rect 19984 34400 20036 34406
rect 19984 34342 20036 34348
rect 19892 34196 19944 34202
rect 19892 34138 19944 34144
rect 19614 34096 19670 34105
rect 19614 34031 19670 34040
rect 19628 33998 19656 34031
rect 19996 33998 20024 34342
rect 19616 33992 19668 33998
rect 19616 33934 19668 33940
rect 19984 33992 20036 33998
rect 19984 33934 20036 33940
rect 20074 33960 20130 33969
rect 19996 33833 20024 33934
rect 20074 33895 20130 33904
rect 20088 33862 20116 33895
rect 20076 33856 20128 33862
rect 19982 33824 20038 33833
rect 20076 33798 20128 33804
rect 19574 33756 19882 33765
rect 19982 33759 20038 33768
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19432 33516 19484 33522
rect 19432 33458 19484 33464
rect 19524 33516 19576 33522
rect 19524 33458 19576 33464
rect 19536 33114 19564 33458
rect 19524 33108 19576 33114
rect 19524 33050 19576 33056
rect 20180 32978 20208 36246
rect 20364 35018 20392 37606
rect 20536 36576 20588 36582
rect 20536 36518 20588 36524
rect 20352 35012 20404 35018
rect 20352 34954 20404 34960
rect 20260 34944 20312 34950
rect 20260 34886 20312 34892
rect 20272 34649 20300 34886
rect 20258 34640 20314 34649
rect 20258 34575 20314 34584
rect 20260 34468 20312 34474
rect 20260 34410 20312 34416
rect 20272 33998 20300 34410
rect 20260 33992 20312 33998
rect 20260 33934 20312 33940
rect 20272 33454 20300 33934
rect 20260 33448 20312 33454
rect 20260 33390 20312 33396
rect 20260 33312 20312 33318
rect 20260 33254 20312 33260
rect 20168 32972 20220 32978
rect 20168 32914 20220 32920
rect 20180 32881 20208 32914
rect 20166 32872 20222 32881
rect 20166 32807 20222 32816
rect 19984 32768 20036 32774
rect 19984 32710 20036 32716
rect 20076 32768 20128 32774
rect 20076 32710 20128 32716
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19996 32337 20024 32710
rect 19982 32328 20038 32337
rect 19982 32263 20038 32272
rect 19340 31952 19392 31958
rect 19340 31894 19392 31900
rect 19352 31822 19380 31894
rect 19340 31816 19392 31822
rect 19340 31758 19392 31764
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19248 31136 19300 31142
rect 19300 31096 19380 31124
rect 19248 31078 19300 31084
rect 19064 30932 19116 30938
rect 19168 30926 19288 30954
rect 19064 30874 19116 30880
rect 19156 30864 19208 30870
rect 19156 30806 19208 30812
rect 18748 30552 19012 30580
rect 19064 30592 19116 30598
rect 18696 30534 18748 30540
rect 18616 30190 18644 30534
rect 18800 30258 18828 30552
rect 19064 30534 19116 30540
rect 19076 30394 19104 30534
rect 19064 30388 19116 30394
rect 19064 30330 19116 30336
rect 18972 30320 19024 30326
rect 18892 30280 18972 30308
rect 18788 30252 18840 30258
rect 18788 30194 18840 30200
rect 18604 30184 18656 30190
rect 18604 30126 18656 30132
rect 18512 29844 18564 29850
rect 18512 29786 18564 29792
rect 18524 29170 18552 29786
rect 18694 29200 18750 29209
rect 18512 29164 18564 29170
rect 18564 29124 18644 29152
rect 18694 29135 18750 29144
rect 18512 29106 18564 29112
rect 18420 29028 18472 29034
rect 18420 28970 18472 28976
rect 18326 28656 18382 28665
rect 18326 28591 18382 28600
rect 18144 28552 18196 28558
rect 18144 28494 18196 28500
rect 18236 28552 18288 28558
rect 18236 28494 18288 28500
rect 18052 28076 18104 28082
rect 18052 28018 18104 28024
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 17972 27130 18000 27406
rect 18144 27396 18196 27402
rect 18144 27338 18196 27344
rect 18328 27396 18380 27402
rect 18328 27338 18380 27344
rect 17960 27124 18012 27130
rect 17960 27066 18012 27072
rect 18156 26382 18184 27338
rect 18340 26926 18368 27338
rect 18328 26920 18380 26926
rect 18328 26862 18380 26868
rect 18340 26382 18368 26862
rect 18144 26376 18196 26382
rect 18144 26318 18196 26324
rect 18328 26376 18380 26382
rect 18328 26318 18380 26324
rect 18236 26308 18288 26314
rect 18236 26250 18288 26256
rect 18248 25974 18276 26250
rect 18236 25968 18288 25974
rect 18236 25910 18288 25916
rect 18052 25288 18104 25294
rect 18052 25230 18104 25236
rect 18064 24886 18092 25230
rect 18144 25152 18196 25158
rect 18144 25094 18196 25100
rect 18052 24880 18104 24886
rect 18052 24822 18104 24828
rect 18156 24206 18184 25094
rect 18144 24200 18196 24206
rect 18144 24142 18196 24148
rect 18328 24200 18380 24206
rect 18328 24142 18380 24148
rect 18052 24132 18104 24138
rect 18052 24074 18104 24080
rect 17960 23588 18012 23594
rect 17960 23530 18012 23536
rect 17972 23225 18000 23530
rect 17958 23216 18014 23225
rect 17958 23151 18014 23160
rect 18064 23118 18092 24074
rect 18340 23866 18368 24142
rect 18432 24120 18460 28970
rect 18512 28960 18564 28966
rect 18512 28902 18564 28908
rect 18524 28558 18552 28902
rect 18512 28552 18564 28558
rect 18512 28494 18564 28500
rect 18512 28416 18564 28422
rect 18512 28358 18564 28364
rect 18524 25226 18552 28358
rect 18512 25220 18564 25226
rect 18512 25162 18564 25168
rect 18524 24614 18552 25162
rect 18616 24698 18644 29124
rect 18708 29034 18736 29135
rect 18696 29028 18748 29034
rect 18696 28970 18748 28976
rect 18696 26988 18748 26994
rect 18696 26930 18748 26936
rect 18708 26382 18736 26930
rect 18696 26376 18748 26382
rect 18696 26318 18748 26324
rect 18616 24670 18736 24698
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18604 24608 18656 24614
rect 18604 24550 18656 24556
rect 18432 24092 18552 24120
rect 18418 24032 18474 24041
rect 18418 23967 18474 23976
rect 18328 23860 18380 23866
rect 18328 23802 18380 23808
rect 18144 23520 18196 23526
rect 18144 23462 18196 23468
rect 18052 23112 18104 23118
rect 18052 23054 18104 23060
rect 18052 22976 18104 22982
rect 18052 22918 18104 22924
rect 18064 22710 18092 22918
rect 18156 22710 18184 23462
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 18052 22704 18104 22710
rect 18052 22646 18104 22652
rect 18144 22704 18196 22710
rect 18144 22646 18196 22652
rect 18156 22094 18184 22646
rect 18064 22066 18184 22094
rect 18064 22030 18092 22066
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 17972 21554 18000 21966
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 17696 20998 17908 21026
rect 17592 19440 17644 19446
rect 17498 19408 17554 19417
rect 17316 19372 17368 19378
rect 17592 19382 17644 19388
rect 17498 19343 17554 19352
rect 17316 19314 17368 19320
rect 17224 19168 17276 19174
rect 17224 19110 17276 19116
rect 17236 18290 17264 19110
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17132 18216 17184 18222
rect 17132 18158 17184 18164
rect 17144 16998 17172 18158
rect 17236 17678 17264 18226
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17604 17513 17632 17546
rect 17590 17504 17646 17513
rect 17590 17439 17646 17448
rect 17222 17232 17278 17241
rect 17222 17167 17278 17176
rect 17236 17134 17264 17167
rect 17224 17128 17276 17134
rect 17276 17088 17632 17116
rect 17224 17070 17276 17076
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 17604 16266 17632 17088
rect 17696 16454 17724 20998
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 17880 19514 17908 19858
rect 18234 19816 18290 19825
rect 18234 19751 18290 19760
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 17868 19508 17920 19514
rect 17868 19450 17920 19456
rect 17776 18284 17828 18290
rect 17776 18226 17828 18232
rect 17788 18086 17816 18226
rect 17776 18080 17828 18086
rect 17776 18022 17828 18028
rect 17774 17912 17830 17921
rect 17774 17847 17830 17856
rect 17788 17678 17816 17847
rect 17880 17746 17908 19450
rect 17972 19122 18000 19654
rect 18156 19446 18184 19654
rect 18248 19446 18276 19751
rect 18144 19440 18196 19446
rect 18144 19382 18196 19388
rect 18236 19440 18288 19446
rect 18236 19382 18288 19388
rect 18156 19334 18184 19382
rect 18156 19306 18276 19334
rect 18144 19168 18196 19174
rect 17972 19116 18144 19122
rect 17972 19110 18196 19116
rect 17972 19094 18184 19110
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 17972 18766 18000 18906
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 17776 17672 17828 17678
rect 17776 17614 17828 17620
rect 17880 17270 17908 17682
rect 17972 17542 18000 18702
rect 18052 17808 18104 17814
rect 18052 17750 18104 17756
rect 18064 17678 18092 17750
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 17868 16992 17920 16998
rect 18064 16980 18092 17614
rect 17920 16952 18092 16980
rect 17868 16934 17920 16940
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 17604 16238 17816 16266
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17500 15904 17552 15910
rect 17500 15846 17552 15852
rect 17224 15700 17276 15706
rect 17224 15642 17276 15648
rect 17130 15464 17186 15473
rect 17130 15399 17186 15408
rect 16868 12702 17080 12730
rect 16868 11626 16896 12702
rect 17144 12238 17172 15399
rect 17236 15094 17264 15642
rect 17420 15434 17448 15846
rect 17408 15428 17460 15434
rect 17408 15370 17460 15376
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 17328 14822 17356 14894
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17512 14634 17540 15846
rect 17592 14816 17644 14822
rect 17592 14758 17644 14764
rect 17420 14606 17540 14634
rect 17420 14414 17448 14606
rect 17500 14544 17552 14550
rect 17500 14486 17552 14492
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17316 13796 17368 13802
rect 17316 13738 17368 13744
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 17236 12442 17264 13466
rect 17328 12782 17356 13738
rect 17420 13394 17448 14214
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17316 12776 17368 12782
rect 17316 12718 17368 12724
rect 17224 12436 17276 12442
rect 17224 12378 17276 12384
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 16854 10840 16910 10849
rect 16854 10775 16910 10784
rect 16868 10742 16896 10775
rect 17052 10742 17080 10950
rect 16856 10736 16908 10742
rect 16856 10678 16908 10684
rect 17040 10736 17092 10742
rect 17040 10678 17092 10684
rect 16868 10130 16896 10678
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16960 9586 16988 9862
rect 17144 9586 17172 11018
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 16868 9178 16896 9522
rect 16946 9480 17002 9489
rect 17236 9466 17264 12378
rect 17420 12322 17448 13330
rect 17512 12986 17540 14486
rect 17604 14346 17632 14758
rect 17684 14612 17736 14618
rect 17684 14554 17736 14560
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 17604 13705 17632 14282
rect 17696 13938 17724 14554
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 17590 13696 17646 13705
rect 17590 13631 17646 13640
rect 17604 13326 17632 13631
rect 17696 13326 17724 13874
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17684 13184 17736 13190
rect 17684 13126 17736 13132
rect 17696 13025 17724 13126
rect 17682 13016 17738 13025
rect 17500 12980 17552 12986
rect 17682 12951 17738 12960
rect 17500 12922 17552 12928
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17512 12434 17540 12786
rect 17512 12406 17724 12434
rect 17420 12294 17540 12322
rect 17512 12238 17540 12294
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17328 11014 17356 12174
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17420 11218 17448 11698
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17512 11218 17540 11494
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 17420 10674 17448 11154
rect 17696 10742 17724 12406
rect 17788 11218 17816 16238
rect 17880 16114 17908 16934
rect 18156 16590 18184 19094
rect 18248 18290 18276 19306
rect 18340 18766 18368 23054
rect 18432 22574 18460 23967
rect 18420 22568 18472 22574
rect 18420 22510 18472 22516
rect 18432 22030 18460 22510
rect 18524 22030 18552 24092
rect 18616 23866 18644 24550
rect 18604 23860 18656 23866
rect 18604 23802 18656 23808
rect 18708 23050 18736 24670
rect 18696 23044 18748 23050
rect 18696 22986 18748 22992
rect 18708 22574 18736 22986
rect 18696 22568 18748 22574
rect 18696 22510 18748 22516
rect 18708 22030 18736 22510
rect 18420 22024 18472 22030
rect 18420 21966 18472 21972
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 18696 22024 18748 22030
rect 18696 21966 18748 21972
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 18248 17649 18276 18226
rect 18328 17876 18380 17882
rect 18328 17818 18380 17824
rect 18340 17746 18368 17818
rect 18328 17740 18380 17746
rect 18328 17682 18380 17688
rect 18234 17640 18290 17649
rect 18234 17575 18290 17584
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18248 17134 18276 17478
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 17880 15434 17908 16050
rect 17972 15706 18000 16186
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 18064 15706 18092 16050
rect 17960 15700 18012 15706
rect 17960 15642 18012 15648
rect 18052 15700 18104 15706
rect 18052 15642 18104 15648
rect 18144 15496 18196 15502
rect 18248 15484 18276 16050
rect 18196 15456 18276 15484
rect 18144 15438 18196 15444
rect 17868 15428 17920 15434
rect 17868 15370 17920 15376
rect 17880 12850 17908 15370
rect 18340 15094 18368 17682
rect 18432 16522 18460 21966
rect 18512 21480 18564 21486
rect 18512 21422 18564 21428
rect 18524 18426 18552 21422
rect 18800 18970 18828 30194
rect 18892 29170 18920 30280
rect 18972 30262 19024 30268
rect 18880 29164 18932 29170
rect 19168 29152 19196 30806
rect 19260 30394 19288 30926
rect 19352 30734 19380 31096
rect 19340 30728 19392 30734
rect 19340 30670 19392 30676
rect 19248 30388 19300 30394
rect 19248 30330 19300 30336
rect 19352 30258 19380 30670
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19340 30252 19392 30258
rect 19340 30194 19392 30200
rect 19248 30184 19300 30190
rect 19248 30126 19300 30132
rect 18880 29106 18932 29112
rect 18984 29124 19196 29152
rect 18880 27328 18932 27334
rect 18880 27270 18932 27276
rect 18892 26790 18920 27270
rect 18880 26784 18932 26790
rect 18880 26726 18932 26732
rect 18892 26586 18920 26726
rect 18880 26580 18932 26586
rect 18880 26522 18932 26528
rect 18892 26382 18920 26522
rect 18880 26376 18932 26382
rect 18880 26318 18932 26324
rect 18880 26240 18932 26246
rect 18880 26182 18932 26188
rect 18892 25702 18920 26182
rect 18880 25696 18932 25702
rect 18880 25638 18932 25644
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 18892 22030 18920 22578
rect 18984 22094 19012 29124
rect 19260 29050 19288 30126
rect 19890 29744 19946 29753
rect 19946 29702 20024 29730
rect 19890 29679 19946 29688
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19432 29164 19484 29170
rect 19432 29106 19484 29112
rect 19168 29022 19288 29050
rect 19168 28490 19196 29022
rect 19248 28960 19300 28966
rect 19248 28902 19300 28908
rect 19260 28490 19288 28902
rect 19444 28762 19472 29106
rect 19524 29096 19576 29102
rect 19524 29038 19576 29044
rect 19432 28756 19484 28762
rect 19432 28698 19484 28704
rect 19156 28484 19208 28490
rect 19156 28426 19208 28432
rect 19248 28484 19300 28490
rect 19248 28426 19300 28432
rect 19064 28144 19116 28150
rect 19064 28086 19116 28092
rect 19076 26246 19104 28086
rect 19168 26518 19196 28426
rect 19260 28150 19288 28426
rect 19248 28144 19300 28150
rect 19248 28086 19300 28092
rect 19340 28008 19392 28014
rect 19340 27950 19392 27956
rect 19248 27396 19300 27402
rect 19248 27338 19300 27344
rect 19260 27130 19288 27338
rect 19248 27124 19300 27130
rect 19248 27066 19300 27072
rect 19352 26994 19380 27950
rect 19340 26988 19392 26994
rect 19340 26930 19392 26936
rect 19248 26852 19300 26858
rect 19248 26794 19300 26800
rect 19156 26512 19208 26518
rect 19156 26454 19208 26460
rect 19064 26240 19116 26246
rect 19064 26182 19116 26188
rect 19260 26058 19288 26794
rect 19444 26586 19472 28698
rect 19536 28490 19564 29038
rect 19892 29028 19944 29034
rect 19892 28970 19944 28976
rect 19798 28792 19854 28801
rect 19798 28727 19800 28736
rect 19852 28727 19854 28736
rect 19800 28698 19852 28704
rect 19904 28694 19932 28970
rect 19892 28688 19944 28694
rect 19892 28630 19944 28636
rect 19798 28520 19854 28529
rect 19524 28484 19576 28490
rect 19798 28455 19800 28464
rect 19524 28426 19576 28432
rect 19852 28455 19854 28464
rect 19800 28426 19852 28432
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19524 27872 19576 27878
rect 19524 27814 19576 27820
rect 19536 27674 19564 27814
rect 19996 27713 20024 29702
rect 19982 27704 20038 27713
rect 19524 27668 19576 27674
rect 19982 27639 20038 27648
rect 19524 27610 19576 27616
rect 19616 27600 19668 27606
rect 19616 27542 19668 27548
rect 19628 27334 19656 27542
rect 19984 27464 20036 27470
rect 19984 27406 20036 27412
rect 19616 27328 19668 27334
rect 19616 27270 19668 27276
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19996 27062 20024 27406
rect 19984 27056 20036 27062
rect 19984 26998 20036 27004
rect 19616 26920 19668 26926
rect 19616 26862 19668 26868
rect 19340 26580 19392 26586
rect 19340 26522 19392 26528
rect 19432 26580 19484 26586
rect 19432 26522 19484 26528
rect 19076 26030 19288 26058
rect 19076 25362 19104 26030
rect 19156 25968 19208 25974
rect 19156 25910 19208 25916
rect 19064 25356 19116 25362
rect 19064 25298 19116 25304
rect 19076 24954 19104 25298
rect 19064 24948 19116 24954
rect 19064 24890 19116 24896
rect 19168 24800 19196 25910
rect 19352 25838 19380 26522
rect 19628 26518 19656 26862
rect 20088 26586 20116 32710
rect 20168 31748 20220 31754
rect 20168 31690 20220 31696
rect 20180 26874 20208 31690
rect 20272 26976 20300 33254
rect 20364 31754 20392 34954
rect 20444 34672 20496 34678
rect 20444 34614 20496 34620
rect 20456 34202 20484 34614
rect 20548 34490 20576 36518
rect 20628 35692 20680 35698
rect 20628 35634 20680 35640
rect 20640 34746 20668 35634
rect 20628 34740 20680 34746
rect 20628 34682 20680 34688
rect 20548 34462 20668 34490
rect 20536 34400 20588 34406
rect 20536 34342 20588 34348
rect 20548 34202 20576 34342
rect 20444 34196 20496 34202
rect 20444 34138 20496 34144
rect 20536 34196 20588 34202
rect 20536 34138 20588 34144
rect 20456 33114 20484 34138
rect 20534 34096 20590 34105
rect 20534 34031 20536 34040
rect 20588 34031 20590 34040
rect 20536 34002 20588 34008
rect 20536 33924 20588 33930
rect 20536 33866 20588 33872
rect 20548 33833 20576 33866
rect 20534 33824 20590 33833
rect 20534 33759 20590 33768
rect 20444 33108 20496 33114
rect 20444 33050 20496 33056
rect 20640 31754 20668 34462
rect 20916 33318 20944 37742
rect 21008 36786 21036 38218
rect 20996 36780 21048 36786
rect 20996 36722 21048 36728
rect 21008 33640 21036 36722
rect 21100 35290 21128 41006
rect 21192 40458 21220 41386
rect 22112 41206 22140 41550
rect 22468 41540 22520 41546
rect 22468 41482 22520 41488
rect 22100 41200 22152 41206
rect 22100 41142 22152 41148
rect 21364 41132 21416 41138
rect 21364 41074 21416 41080
rect 21640 41132 21692 41138
rect 21640 41074 21692 41080
rect 21376 40730 21404 41074
rect 21364 40724 21416 40730
rect 21364 40666 21416 40672
rect 21652 40594 21680 41074
rect 21824 41064 21876 41070
rect 21824 41006 21876 41012
rect 21640 40588 21692 40594
rect 21640 40530 21692 40536
rect 21180 40452 21232 40458
rect 21180 40394 21232 40400
rect 21088 35284 21140 35290
rect 21088 35226 21140 35232
rect 21008 33612 21128 33640
rect 20904 33312 20956 33318
rect 20904 33254 20956 33260
rect 21100 32994 21128 33612
rect 21192 33522 21220 40394
rect 21836 39982 21864 41006
rect 22480 40730 22508 41482
rect 23860 41274 23888 43893
rect 23940 41540 23992 41546
rect 23940 41482 23992 41488
rect 24216 41540 24268 41546
rect 24216 41482 24268 41488
rect 23848 41268 23900 41274
rect 23848 41210 23900 41216
rect 23388 41132 23440 41138
rect 23388 41074 23440 41080
rect 22468 40724 22520 40730
rect 22468 40666 22520 40672
rect 22284 40588 22336 40594
rect 22284 40530 22336 40536
rect 22008 40044 22060 40050
rect 22008 39986 22060 39992
rect 21824 39976 21876 39982
rect 21824 39918 21876 39924
rect 21824 39840 21876 39846
rect 21824 39782 21876 39788
rect 21836 39506 21864 39782
rect 21824 39500 21876 39506
rect 21824 39442 21876 39448
rect 22020 39098 22048 39986
rect 22008 39092 22060 39098
rect 22008 39034 22060 39040
rect 22008 38956 22060 38962
rect 22008 38898 22060 38904
rect 22020 38554 22048 38898
rect 22008 38548 22060 38554
rect 22008 38490 22060 38496
rect 22008 37868 22060 37874
rect 22008 37810 22060 37816
rect 22020 37369 22048 37810
rect 22100 37732 22152 37738
rect 22100 37674 22152 37680
rect 22006 37360 22062 37369
rect 22006 37295 22062 37304
rect 22112 35894 22140 37674
rect 21928 35866 22140 35894
rect 21928 35698 21956 35866
rect 21916 35692 21968 35698
rect 21916 35634 21968 35640
rect 21824 35488 21876 35494
rect 21824 35430 21876 35436
rect 21836 35154 21864 35430
rect 21824 35148 21876 35154
rect 21824 35090 21876 35096
rect 21732 34944 21784 34950
rect 21732 34886 21784 34892
rect 21548 34604 21600 34610
rect 21548 34546 21600 34552
rect 21454 34096 21510 34105
rect 21454 34031 21456 34040
rect 21508 34031 21510 34040
rect 21456 34002 21508 34008
rect 21364 33992 21416 33998
rect 21362 33960 21364 33969
rect 21416 33960 21418 33969
rect 21362 33895 21418 33904
rect 21180 33516 21232 33522
rect 21180 33458 21232 33464
rect 21008 32966 21128 32994
rect 21008 32910 21036 32966
rect 21192 32910 21220 33458
rect 21364 33312 21416 33318
rect 21364 33254 21416 33260
rect 21376 32978 21404 33254
rect 21364 32972 21416 32978
rect 21364 32914 21416 32920
rect 20996 32904 21048 32910
rect 20996 32846 21048 32852
rect 21180 32904 21232 32910
rect 21180 32846 21232 32852
rect 20904 31816 20956 31822
rect 20904 31758 20956 31764
rect 20352 31748 20404 31754
rect 20352 31690 20404 31696
rect 20456 31726 20668 31754
rect 20456 31226 20484 31726
rect 20916 31362 20944 31758
rect 21008 31482 21036 32846
rect 21376 32473 21404 32914
rect 21362 32464 21418 32473
rect 21180 32428 21232 32434
rect 21362 32399 21418 32408
rect 21180 32370 21232 32376
rect 21088 31680 21140 31686
rect 21088 31622 21140 31628
rect 21100 31482 21128 31622
rect 20996 31476 21048 31482
rect 20996 31418 21048 31424
rect 21088 31476 21140 31482
rect 21088 31418 21140 31424
rect 20916 31334 21036 31362
rect 20364 31198 20484 31226
rect 20364 28642 20392 31198
rect 20444 31136 20496 31142
rect 20444 31078 20496 31084
rect 20628 31136 20680 31142
rect 20628 31078 20680 31084
rect 20456 30734 20484 31078
rect 20444 30728 20496 30734
rect 20444 30670 20496 30676
rect 20456 30326 20484 30670
rect 20536 30660 20588 30666
rect 20536 30602 20588 30608
rect 20444 30320 20496 30326
rect 20444 30262 20496 30268
rect 20442 30152 20498 30161
rect 20442 30087 20444 30096
rect 20496 30087 20498 30096
rect 20444 30058 20496 30064
rect 20548 29170 20576 30602
rect 20640 30190 20668 31078
rect 20904 30592 20956 30598
rect 20904 30534 20956 30540
rect 20628 30184 20680 30190
rect 20628 30126 20680 30132
rect 20812 30048 20864 30054
rect 20732 30008 20812 30036
rect 20628 29232 20680 29238
rect 20628 29174 20680 29180
rect 20536 29164 20588 29170
rect 20536 29106 20588 29112
rect 20364 28614 20484 28642
rect 20352 28552 20404 28558
rect 20352 28494 20404 28500
rect 20364 28014 20392 28494
rect 20352 28008 20404 28014
rect 20352 27950 20404 27956
rect 20456 27044 20484 28614
rect 20548 27470 20576 29106
rect 20536 27464 20588 27470
rect 20536 27406 20588 27412
rect 20456 27016 20576 27044
rect 20272 26948 20484 26976
rect 20180 26846 20300 26874
rect 20168 26784 20220 26790
rect 20168 26726 20220 26732
rect 20076 26580 20128 26586
rect 20076 26522 20128 26528
rect 19616 26512 19668 26518
rect 19616 26454 19668 26460
rect 19432 26376 19484 26382
rect 19432 26318 19484 26324
rect 19444 25906 19472 26318
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19432 25900 19484 25906
rect 19432 25842 19484 25848
rect 20076 25900 20128 25906
rect 20076 25842 20128 25848
rect 19340 25832 19392 25838
rect 19340 25774 19392 25780
rect 19340 25696 19392 25702
rect 19340 25638 19392 25644
rect 19248 25288 19300 25294
rect 19248 25230 19300 25236
rect 19260 24954 19288 25230
rect 19248 24948 19300 24954
rect 19248 24890 19300 24896
rect 19248 24812 19300 24818
rect 19168 24772 19248 24800
rect 19248 24754 19300 24760
rect 19352 24410 19380 25638
rect 19340 24404 19392 24410
rect 19340 24346 19392 24352
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19352 22166 19380 23122
rect 19340 22160 19392 22166
rect 19340 22102 19392 22108
rect 18984 22066 19104 22094
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 19076 21842 19104 22066
rect 19156 21956 19208 21962
rect 19156 21898 19208 21904
rect 18892 21814 19104 21842
rect 18788 18964 18840 18970
rect 18788 18906 18840 18912
rect 18604 18692 18656 18698
rect 18604 18634 18656 18640
rect 18616 18426 18644 18634
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 18512 18420 18564 18426
rect 18512 18362 18564 18368
rect 18604 18420 18656 18426
rect 18604 18362 18656 18368
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18512 17672 18564 17678
rect 18510 17640 18512 17649
rect 18564 17640 18566 17649
rect 18510 17575 18566 17584
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 18420 16516 18472 16522
rect 18420 16458 18472 16464
rect 18432 16182 18460 16458
rect 18420 16176 18472 16182
rect 18420 16118 18472 16124
rect 18524 16046 18552 17070
rect 18512 16040 18564 16046
rect 18512 15982 18564 15988
rect 18524 15910 18552 15982
rect 18512 15904 18564 15910
rect 18432 15864 18512 15892
rect 18328 15088 18380 15094
rect 18328 15030 18380 15036
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 17972 14414 18000 14554
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17960 14272 18012 14278
rect 17960 14214 18012 14220
rect 17972 12850 18000 14214
rect 18156 13938 18184 14554
rect 18144 13932 18196 13938
rect 18144 13874 18196 13880
rect 18340 13870 18368 14758
rect 18432 14414 18460 15864
rect 18512 15846 18564 15852
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18052 13728 18104 13734
rect 18052 13670 18104 13676
rect 18064 12850 18092 13670
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 18156 12442 18184 13262
rect 18432 13161 18460 14214
rect 18418 13152 18474 13161
rect 18418 13087 18474 13096
rect 18616 12850 18644 18022
rect 18708 17814 18736 18566
rect 18696 17808 18748 17814
rect 18696 17750 18748 17756
rect 18696 17536 18748 17542
rect 18696 17478 18748 17484
rect 18708 17338 18736 17478
rect 18696 17332 18748 17338
rect 18696 17274 18748 17280
rect 18800 16250 18828 18906
rect 18892 17882 18920 21814
rect 19064 21684 19116 21690
rect 19064 21626 19116 21632
rect 18972 21548 19024 21554
rect 18972 21490 19024 21496
rect 18984 21146 19012 21490
rect 19076 21418 19104 21626
rect 19064 21412 19116 21418
rect 19064 21354 19116 21360
rect 18972 21140 19024 21146
rect 19168 21128 19196 21898
rect 19340 21616 19392 21622
rect 19340 21558 19392 21564
rect 19248 21344 19300 21350
rect 19248 21286 19300 21292
rect 18972 21082 19024 21088
rect 19076 21100 19196 21128
rect 19076 20398 19104 21100
rect 19260 21026 19288 21286
rect 19168 21010 19288 21026
rect 19156 21004 19288 21010
rect 19208 20998 19288 21004
rect 19156 20946 19208 20952
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 19064 20392 19116 20398
rect 19064 20334 19116 20340
rect 19064 19984 19116 19990
rect 19064 19926 19116 19932
rect 19076 19310 19104 19926
rect 19064 19304 19116 19310
rect 19064 19246 19116 19252
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 19076 18290 19104 19110
rect 19168 18902 19196 19246
rect 19260 19009 19288 20878
rect 19352 20330 19380 21558
rect 19444 21554 19472 25842
rect 19984 25288 20036 25294
rect 19984 25230 20036 25236
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19616 24880 19668 24886
rect 19668 24840 19748 24868
rect 19616 24822 19668 24828
rect 19720 24449 19748 24840
rect 19800 24608 19852 24614
rect 19800 24550 19852 24556
rect 19706 24440 19762 24449
rect 19706 24375 19708 24384
rect 19760 24375 19762 24384
rect 19708 24346 19760 24352
rect 19812 24138 19840 24550
rect 19996 24206 20024 25230
rect 20088 25158 20116 25842
rect 20076 25152 20128 25158
rect 20076 25094 20128 25100
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 19800 24132 19852 24138
rect 19800 24074 19852 24080
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19892 22704 19944 22710
rect 19892 22646 19944 22652
rect 19904 22098 19932 22646
rect 19892 22092 19944 22098
rect 19892 22034 19944 22040
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19524 21684 19576 21690
rect 19524 21626 19576 21632
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19444 21010 19472 21490
rect 19536 21457 19564 21626
rect 19522 21448 19578 21457
rect 19522 21383 19578 21392
rect 19432 21004 19484 21010
rect 19432 20946 19484 20952
rect 19536 20788 19564 21383
rect 19444 20760 19564 20788
rect 19444 20534 19472 20760
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19996 20602 20024 21830
rect 20088 21350 20116 25094
rect 20180 23866 20208 26726
rect 20272 25974 20300 26846
rect 20352 26580 20404 26586
rect 20352 26522 20404 26528
rect 20260 25968 20312 25974
rect 20260 25910 20312 25916
rect 20260 25492 20312 25498
rect 20260 25434 20312 25440
rect 20272 24818 20300 25434
rect 20260 24812 20312 24818
rect 20260 24754 20312 24760
rect 20260 24064 20312 24070
rect 20260 24006 20312 24012
rect 20168 23860 20220 23866
rect 20168 23802 20220 23808
rect 20272 23633 20300 24006
rect 20258 23624 20314 23633
rect 20168 23588 20220 23594
rect 20258 23559 20314 23568
rect 20168 23530 20220 23536
rect 20180 22778 20208 23530
rect 20260 23520 20312 23526
rect 20260 23462 20312 23468
rect 20168 22772 20220 22778
rect 20168 22714 20220 22720
rect 20168 21956 20220 21962
rect 20168 21898 20220 21904
rect 20180 21622 20208 21898
rect 20168 21616 20220 21622
rect 20168 21558 20220 21564
rect 20076 21344 20128 21350
rect 20076 21286 20128 21292
rect 20088 21146 20116 21286
rect 20076 21140 20128 21146
rect 20076 21082 20128 21088
rect 20272 21010 20300 23462
rect 20260 21004 20312 21010
rect 20260 20946 20312 20952
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 19432 20528 19484 20534
rect 19432 20470 19484 20476
rect 20076 20528 20128 20534
rect 20076 20470 20128 20476
rect 19706 20360 19762 20369
rect 19340 20324 19392 20330
rect 19706 20295 19762 20304
rect 19984 20324 20036 20330
rect 19340 20266 19392 20272
rect 19614 20088 19670 20097
rect 19614 20023 19670 20032
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19246 19000 19302 19009
rect 19246 18935 19302 18944
rect 19156 18896 19208 18902
rect 19156 18838 19208 18844
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 18972 18216 19024 18222
rect 19168 18170 19196 18838
rect 19352 18408 19380 19858
rect 19628 19854 19656 20023
rect 19720 19990 19748 20295
rect 19984 20266 20036 20272
rect 19708 19984 19760 19990
rect 19708 19926 19760 19932
rect 19616 19848 19668 19854
rect 19616 19790 19668 19796
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19444 19310 19472 19654
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 19304 19484 19310
rect 19432 19246 19484 19252
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19352 18380 19472 18408
rect 19340 18284 19392 18290
rect 19340 18226 19392 18232
rect 19024 18164 19196 18170
rect 18972 18158 19196 18164
rect 18984 18142 19196 18158
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18984 17921 19012 18022
rect 18970 17912 19026 17921
rect 18880 17876 18932 17882
rect 18970 17847 19026 17856
rect 18880 17818 18932 17824
rect 19168 17678 19196 18142
rect 19352 17882 19380 18226
rect 19444 18222 19472 18380
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19338 17776 19394 17785
rect 19248 17740 19300 17746
rect 19338 17711 19394 17720
rect 19248 17682 19300 17688
rect 18880 17672 18932 17678
rect 19156 17672 19208 17678
rect 18880 17614 18932 17620
rect 19062 17640 19118 17649
rect 18892 17513 18920 17614
rect 19156 17614 19208 17620
rect 19062 17575 19118 17584
rect 18878 17504 18934 17513
rect 18878 17439 18934 17448
rect 18972 16516 19024 16522
rect 18972 16458 19024 16464
rect 18788 16244 18840 16250
rect 18788 16186 18840 16192
rect 18800 15638 18828 16186
rect 18984 16114 19012 16458
rect 18972 16108 19024 16114
rect 18892 16068 18972 16096
rect 18788 15632 18840 15638
rect 18788 15574 18840 15580
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18708 14890 18736 15438
rect 18788 15088 18840 15094
rect 18788 15030 18840 15036
rect 18696 14884 18748 14890
rect 18696 14826 18748 14832
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18708 13802 18736 14214
rect 18696 13796 18748 13802
rect 18696 13738 18748 13744
rect 18800 12918 18828 15030
rect 18892 14414 18920 16068
rect 18972 16050 19024 16056
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 19076 14278 19104 17575
rect 19260 16590 19288 17682
rect 19352 17270 19380 17711
rect 19340 17264 19392 17270
rect 19340 17206 19392 17212
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 19246 16144 19302 16153
rect 19246 16079 19248 16088
rect 19300 16079 19302 16088
rect 19248 16050 19300 16056
rect 19156 15972 19208 15978
rect 19156 15914 19208 15920
rect 19168 15473 19196 15914
rect 19154 15464 19210 15473
rect 19154 15399 19210 15408
rect 19156 15360 19208 15366
rect 19156 15302 19208 15308
rect 19064 14272 19116 14278
rect 19064 14214 19116 14220
rect 19168 14226 19196 15302
rect 19352 14906 19380 16934
rect 19444 15366 19472 18158
rect 19616 18080 19668 18086
rect 19616 18022 19668 18028
rect 19628 17746 19656 18022
rect 19616 17740 19668 17746
rect 19616 17682 19668 17688
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19890 16824 19946 16833
rect 19890 16759 19946 16768
rect 19904 16726 19932 16759
rect 19892 16720 19944 16726
rect 19892 16662 19944 16668
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19616 15156 19668 15162
rect 19616 15098 19668 15104
rect 19432 15088 19484 15094
rect 19432 15030 19484 15036
rect 19444 14929 19472 15030
rect 19524 15020 19576 15026
rect 19524 14962 19576 14968
rect 19260 14890 19380 14906
rect 19248 14884 19380 14890
rect 19300 14878 19380 14884
rect 19430 14920 19486 14929
rect 19430 14855 19486 14864
rect 19248 14826 19300 14832
rect 19260 14414 19288 14826
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19248 14408 19300 14414
rect 19248 14350 19300 14356
rect 19168 14198 19288 14226
rect 19260 13954 19288 14198
rect 19352 14074 19380 14758
rect 19444 14550 19472 14758
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 19536 14498 19564 14962
rect 19628 14618 19656 15098
rect 19996 14770 20024 20266
rect 20088 19145 20116 20470
rect 20168 20392 20220 20398
rect 20168 20334 20220 20340
rect 20180 19922 20208 20334
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 20168 19440 20220 19446
rect 20168 19382 20220 19388
rect 20074 19136 20130 19145
rect 20074 19071 20130 19080
rect 20180 18465 20208 19382
rect 20166 18456 20222 18465
rect 20166 18391 20222 18400
rect 20180 16998 20208 18391
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20076 16652 20128 16658
rect 20076 16594 20128 16600
rect 19904 14742 20024 14770
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19800 14544 19852 14550
rect 19720 14504 19800 14532
rect 19720 14498 19748 14504
rect 19536 14470 19748 14498
rect 19800 14486 19852 14492
rect 19904 14385 19932 14742
rect 20088 14634 20116 16594
rect 20166 15192 20222 15201
rect 20166 15127 20168 15136
rect 20220 15127 20222 15136
rect 20168 15098 20220 15104
rect 19996 14606 20116 14634
rect 19996 14550 20024 14606
rect 19984 14544 20036 14550
rect 19984 14486 20036 14492
rect 19890 14376 19946 14385
rect 19432 14340 19484 14346
rect 19890 14311 19946 14320
rect 19432 14282 19484 14288
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19260 13926 19380 13954
rect 19064 13728 19116 13734
rect 19064 13670 19116 13676
rect 19076 13138 19104 13670
rect 18892 13110 19104 13138
rect 18788 12912 18840 12918
rect 18788 12854 18840 12860
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18616 11898 18644 12038
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18328 11620 18380 11626
rect 18328 11562 18380 11568
rect 17776 11212 17828 11218
rect 17776 11154 17828 11160
rect 17960 10804 18012 10810
rect 17960 10746 18012 10752
rect 17684 10736 17736 10742
rect 17684 10678 17736 10684
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17002 9438 17264 9466
rect 16946 9415 16948 9424
rect 17000 9415 17002 9424
rect 16948 9386 17000 9392
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16764 8560 16816 8566
rect 16764 8502 16816 8508
rect 17316 8560 17368 8566
rect 17316 8502 17368 8508
rect 16304 8424 16356 8430
rect 16304 8366 16356 8372
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 15488 7410 15516 7686
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 16040 7410 16068 7482
rect 16224 7410 16252 7686
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 15384 7336 15436 7342
rect 15844 7336 15896 7342
rect 15842 7304 15844 7313
rect 15896 7304 15898 7313
rect 15436 7284 15608 7290
rect 15384 7278 15608 7284
rect 15396 7262 15608 7278
rect 15396 6769 15424 7262
rect 15580 7206 15608 7262
rect 15842 7239 15898 7248
rect 16316 7206 16344 8366
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16684 7410 16712 8230
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 15488 7002 15516 7142
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 17328 6866 17356 8502
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 15382 6760 15438 6769
rect 15382 6695 15438 6704
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15304 6458 15332 6598
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15108 5840 15160 5846
rect 15108 5782 15160 5788
rect 16316 5642 16344 6802
rect 17512 6798 17540 10202
rect 17592 8900 17644 8906
rect 17592 8842 17644 8848
rect 17604 8634 17632 8842
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17130 5672 17186 5681
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 16672 5636 16724 5642
rect 17130 5607 17186 5616
rect 16672 5578 16724 5584
rect 16316 5370 16344 5578
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 13084 5296 13136 5302
rect 13084 5238 13136 5244
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9772 5092 9824 5098
rect 9772 5034 9824 5040
rect 9784 4146 9812 5034
rect 9968 4826 9996 5102
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14384 4826 14412 4966
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 16316 4690 16344 5306
rect 16684 5302 16712 5578
rect 16946 5536 17002 5545
rect 16946 5471 17002 5480
rect 16672 5296 16724 5302
rect 16672 5238 16724 5244
rect 16960 5234 16988 5471
rect 17144 5234 17172 5607
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 17132 5228 17184 5234
rect 17132 5170 17184 5176
rect 17788 4826 17816 7822
rect 17868 6724 17920 6730
rect 17868 6666 17920 6672
rect 17880 5642 17908 6666
rect 17972 6390 18000 10746
rect 18340 8430 18368 11562
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18418 9208 18474 9217
rect 18418 9143 18474 9152
rect 18432 8537 18460 9143
rect 18418 8528 18474 8537
rect 18418 8463 18474 8472
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 18432 6866 18460 8463
rect 18616 8294 18644 11154
rect 18708 10674 18736 12786
rect 18800 12753 18828 12854
rect 18786 12744 18842 12753
rect 18786 12679 18842 12688
rect 18892 12434 18920 13110
rect 18972 12708 19024 12714
rect 18972 12650 19024 12656
rect 18984 12442 19012 12650
rect 19064 12640 19116 12646
rect 19064 12582 19116 12588
rect 18800 12406 18920 12434
rect 18972 12436 19024 12442
rect 18800 12238 18828 12406
rect 18972 12378 19024 12384
rect 19076 12238 19104 12582
rect 19352 12442 19380 13926
rect 19444 13734 19472 14282
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19522 13968 19578 13977
rect 19522 13903 19578 13912
rect 19798 13968 19854 13977
rect 19996 13938 20024 14486
rect 19798 13903 19800 13912
rect 19432 13728 19484 13734
rect 19432 13670 19484 13676
rect 19536 13240 19564 13903
rect 19852 13903 19854 13912
rect 19984 13932 20036 13938
rect 19800 13874 19852 13880
rect 19984 13874 20036 13880
rect 19708 13864 19760 13870
rect 19708 13806 19760 13812
rect 19720 13326 19748 13806
rect 19996 13394 20024 13874
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19444 13212 19564 13240
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 19064 12232 19116 12238
rect 19064 12174 19116 12180
rect 19340 11824 19392 11830
rect 19340 11766 19392 11772
rect 19352 10810 19380 11766
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 18972 10736 19024 10742
rect 19064 10736 19116 10742
rect 18972 10678 19024 10684
rect 19062 10704 19064 10713
rect 19116 10704 19118 10713
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18984 8974 19012 10678
rect 19062 10639 19118 10648
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19340 10600 19392 10606
rect 19340 10542 19392 10548
rect 19168 10062 19196 10542
rect 19352 10266 19380 10542
rect 19340 10260 19392 10266
rect 19340 10202 19392 10208
rect 19156 10056 19208 10062
rect 19444 10033 19472 13212
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19628 12442 19656 12718
rect 19616 12436 19668 12442
rect 19616 12378 19668 12384
rect 20076 12436 20128 12442
rect 20076 12378 20128 12384
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19996 10674 20024 12038
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 19156 9998 19208 10004
rect 19430 10024 19486 10033
rect 19430 9959 19486 9968
rect 19444 9654 19472 9959
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19996 9654 20024 10406
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19800 9648 19852 9654
rect 19800 9590 19852 9596
rect 19984 9648 20036 9654
rect 19984 9590 20036 9596
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 19168 9178 19196 9522
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19156 9172 19208 9178
rect 19156 9114 19208 9120
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 18972 8968 19024 8974
rect 18892 8928 18972 8956
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18892 7886 18920 8928
rect 18972 8910 19024 8916
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 18972 8832 19024 8838
rect 19076 8786 19104 8910
rect 19024 8780 19104 8786
rect 18972 8774 19104 8780
rect 19248 8832 19300 8838
rect 19248 8774 19300 8780
rect 18984 8758 19104 8774
rect 18984 8090 19012 8758
rect 19260 8634 19288 8774
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 19062 8120 19118 8129
rect 18972 8084 19024 8090
rect 19062 8055 19118 8064
rect 18972 8026 19024 8032
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18696 7812 18748 7818
rect 18696 7754 18748 7760
rect 18708 7478 18736 7754
rect 18892 7478 18920 7822
rect 18696 7472 18748 7478
rect 18696 7414 18748 7420
rect 18880 7472 18932 7478
rect 18880 7414 18932 7420
rect 19076 6866 19104 8055
rect 19352 7546 19380 8978
rect 19444 8634 19472 9318
rect 19720 9042 19748 9318
rect 19708 9036 19760 9042
rect 19812 9024 19840 9590
rect 19812 8996 20024 9024
rect 19708 8978 19760 8984
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19996 8566 20024 8996
rect 19984 8560 20036 8566
rect 19984 8502 20036 8508
rect 20088 8498 20116 12378
rect 20180 11830 20208 15098
rect 20272 12238 20300 20198
rect 20364 15094 20392 26522
rect 20456 26450 20484 26948
rect 20444 26444 20496 26450
rect 20444 26386 20496 26392
rect 20444 26036 20496 26042
rect 20444 25978 20496 25984
rect 20456 25362 20484 25978
rect 20444 25356 20496 25362
rect 20444 25298 20496 25304
rect 20456 23866 20484 25298
rect 20444 23860 20496 23866
rect 20444 23802 20496 23808
rect 20548 23118 20576 27016
rect 20640 26586 20668 29174
rect 20732 28966 20760 30008
rect 20812 29990 20864 29996
rect 20812 29708 20864 29714
rect 20812 29650 20864 29656
rect 20720 28960 20772 28966
rect 20720 28902 20772 28908
rect 20718 28792 20774 28801
rect 20718 28727 20774 28736
rect 20732 28422 20760 28727
rect 20720 28416 20772 28422
rect 20720 28358 20772 28364
rect 20824 28200 20852 29650
rect 20732 28172 20852 28200
rect 20628 26580 20680 26586
rect 20628 26522 20680 26528
rect 20628 26444 20680 26450
rect 20628 26386 20680 26392
rect 20640 24274 20668 26386
rect 20732 25786 20760 28172
rect 20812 28076 20864 28082
rect 20916 28064 20944 30534
rect 21008 28665 21036 31334
rect 21086 30832 21142 30841
rect 21192 30818 21220 32370
rect 21364 32292 21416 32298
rect 21364 32234 21416 32240
rect 21272 31136 21324 31142
rect 21272 31078 21324 31084
rect 21284 30938 21312 31078
rect 21272 30932 21324 30938
rect 21272 30874 21324 30880
rect 21192 30790 21312 30818
rect 21086 30767 21142 30776
rect 21100 29714 21128 30767
rect 21180 30728 21232 30734
rect 21180 30670 21232 30676
rect 21192 30326 21220 30670
rect 21180 30320 21232 30326
rect 21180 30262 21232 30268
rect 21180 30184 21232 30190
rect 21178 30152 21180 30161
rect 21232 30152 21234 30161
rect 21178 30087 21234 30096
rect 21088 29708 21140 29714
rect 21088 29650 21140 29656
rect 21088 29504 21140 29510
rect 21088 29446 21140 29452
rect 20994 28656 21050 28665
rect 20994 28591 21050 28600
rect 21100 28558 21128 29446
rect 21284 29102 21312 30790
rect 21272 29096 21324 29102
rect 21272 29038 21324 29044
rect 21284 28762 21312 29038
rect 21272 28756 21324 28762
rect 21272 28698 21324 28704
rect 21180 28620 21232 28626
rect 21180 28562 21232 28568
rect 20996 28552 21048 28558
rect 20994 28520 20996 28529
rect 21088 28552 21140 28558
rect 21048 28520 21050 28529
rect 21088 28494 21140 28500
rect 20994 28455 21050 28464
rect 20996 28212 21048 28218
rect 20996 28154 21048 28160
rect 20864 28036 20944 28064
rect 20812 28018 20864 28024
rect 20824 27713 20852 28018
rect 20810 27704 20866 27713
rect 20810 27639 20866 27648
rect 21008 27614 21036 28154
rect 21100 27690 21128 28494
rect 21192 28218 21220 28562
rect 21272 28484 21324 28490
rect 21272 28426 21324 28432
rect 21180 28212 21232 28218
rect 21180 28154 21232 28160
rect 21284 28150 21312 28426
rect 21272 28144 21324 28150
rect 21272 28086 21324 28092
rect 21272 27872 21324 27878
rect 21272 27814 21324 27820
rect 21100 27662 21220 27690
rect 20916 27586 21036 27614
rect 20916 26246 20944 27586
rect 20996 27056 21048 27062
rect 20996 26998 21048 27004
rect 20904 26240 20956 26246
rect 20904 26182 20956 26188
rect 21008 25945 21036 26998
rect 21088 26920 21140 26926
rect 21088 26862 21140 26868
rect 20994 25936 21050 25945
rect 20904 25900 20956 25906
rect 20994 25871 21050 25880
rect 20904 25842 20956 25848
rect 20732 25758 20852 25786
rect 20720 25696 20772 25702
rect 20720 25638 20772 25644
rect 20628 24268 20680 24274
rect 20628 24210 20680 24216
rect 20536 23112 20588 23118
rect 20536 23054 20588 23060
rect 20640 22094 20668 24210
rect 20732 23866 20760 25638
rect 20824 25498 20852 25758
rect 20916 25498 20944 25842
rect 20996 25696 21048 25702
rect 20996 25638 21048 25644
rect 20812 25492 20864 25498
rect 20812 25434 20864 25440
rect 20904 25492 20956 25498
rect 20904 25434 20956 25440
rect 20916 25362 20944 25434
rect 20904 25356 20956 25362
rect 20904 25298 20956 25304
rect 21008 25294 21036 25638
rect 20996 25288 21048 25294
rect 20996 25230 21048 25236
rect 20812 24812 20864 24818
rect 20812 24754 20864 24760
rect 20720 23860 20772 23866
rect 20720 23802 20772 23808
rect 20720 23656 20772 23662
rect 20718 23624 20720 23633
rect 20772 23624 20774 23633
rect 20718 23559 20774 23568
rect 20720 22976 20772 22982
rect 20720 22918 20772 22924
rect 20732 22574 20760 22918
rect 20720 22568 20772 22574
rect 20720 22510 20772 22516
rect 20548 22066 20668 22094
rect 20444 21888 20496 21894
rect 20444 21830 20496 21836
rect 20456 21418 20484 21830
rect 20444 21412 20496 21418
rect 20444 21354 20496 21360
rect 20444 20460 20496 20466
rect 20444 20402 20496 20408
rect 20456 19718 20484 20402
rect 20548 19718 20576 22066
rect 20628 22024 20680 22030
rect 20626 21992 20628 22001
rect 20680 21992 20682 22001
rect 20626 21927 20682 21936
rect 20732 21876 20760 22510
rect 20824 22438 20852 24754
rect 20904 24336 20956 24342
rect 20904 24278 20956 24284
rect 20812 22432 20864 22438
rect 20812 22374 20864 22380
rect 20640 21848 20760 21876
rect 20640 20942 20668 21848
rect 20720 21616 20772 21622
rect 20824 21604 20852 22374
rect 20772 21576 20852 21604
rect 20720 21558 20772 21564
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20732 21185 20760 21422
rect 20718 21176 20774 21185
rect 20718 21111 20774 21120
rect 20628 20936 20680 20942
rect 20628 20878 20680 20884
rect 20916 20754 20944 24278
rect 21008 23594 21036 25230
rect 20996 23588 21048 23594
rect 20996 23530 21048 23536
rect 20994 22944 21050 22953
rect 20994 22879 21050 22888
rect 21008 22030 21036 22879
rect 21100 22273 21128 26862
rect 21192 25129 21220 27662
rect 21178 25120 21234 25129
rect 21178 25055 21234 25064
rect 21284 24682 21312 27814
rect 21272 24676 21324 24682
rect 21272 24618 21324 24624
rect 21272 24404 21324 24410
rect 21272 24346 21324 24352
rect 21284 23866 21312 24346
rect 21376 24342 21404 32234
rect 21456 32224 21508 32230
rect 21456 32166 21508 32172
rect 21468 31822 21496 32166
rect 21560 31822 21588 34546
rect 21640 33856 21692 33862
rect 21640 33798 21692 33804
rect 21652 32434 21680 33798
rect 21640 32428 21692 32434
rect 21640 32370 21692 32376
rect 21456 31816 21508 31822
rect 21456 31758 21508 31764
rect 21548 31816 21600 31822
rect 21548 31758 21600 31764
rect 21744 31686 21772 34886
rect 21824 32768 21876 32774
rect 21928 32756 21956 35634
rect 22296 34898 22324 40530
rect 22468 40520 22520 40526
rect 22468 40462 22520 40468
rect 22480 38418 22508 40462
rect 23400 40066 23428 41074
rect 23860 41070 23888 41210
rect 23952 41138 23980 41482
rect 24228 41274 24256 41482
rect 24216 41268 24268 41274
rect 24216 41210 24268 41216
rect 23940 41132 23992 41138
rect 23940 41074 23992 41080
rect 23848 41064 23900 41070
rect 23848 41006 23900 41012
rect 24228 40526 24256 41210
rect 24216 40520 24268 40526
rect 24216 40462 24268 40468
rect 24952 40180 25004 40186
rect 24952 40122 25004 40128
rect 23572 40112 23624 40118
rect 23400 40060 23572 40066
rect 23400 40054 23624 40060
rect 23112 40044 23164 40050
rect 23112 39986 23164 39992
rect 23400 40038 23612 40054
rect 23124 39642 23152 39986
rect 23112 39636 23164 39642
rect 23112 39578 23164 39584
rect 22836 39568 22888 39574
rect 22836 39510 22888 39516
rect 22468 38412 22520 38418
rect 22468 38354 22520 38360
rect 22652 37868 22704 37874
rect 22652 37810 22704 37816
rect 22376 37664 22428 37670
rect 22376 37606 22428 37612
rect 22388 37330 22416 37606
rect 22376 37324 22428 37330
rect 22376 37266 22428 37272
rect 22664 36922 22692 37810
rect 22652 36916 22704 36922
rect 22652 36858 22704 36864
rect 22848 36718 22876 39510
rect 23400 39302 23428 40038
rect 24964 39438 24992 40122
rect 26148 39500 26200 39506
rect 26148 39442 26200 39448
rect 24952 39432 25004 39438
rect 24952 39374 25004 39380
rect 26056 39364 26108 39370
rect 26056 39306 26108 39312
rect 22928 39296 22980 39302
rect 22928 39238 22980 39244
rect 23388 39296 23440 39302
rect 23388 39238 23440 39244
rect 22940 39098 22968 39238
rect 22928 39092 22980 39098
rect 22928 39034 22980 39040
rect 23204 38548 23256 38554
rect 23204 38490 23256 38496
rect 23216 37874 23244 38490
rect 23400 38214 23428 39238
rect 26068 39098 26096 39306
rect 26056 39092 26108 39098
rect 26056 39034 26108 39040
rect 25596 38956 25648 38962
rect 25596 38898 25648 38904
rect 25780 38956 25832 38962
rect 25780 38898 25832 38904
rect 26056 38956 26108 38962
rect 26056 38898 26108 38904
rect 24952 38412 25004 38418
rect 24952 38354 25004 38360
rect 23388 38208 23440 38214
rect 23388 38150 23440 38156
rect 23112 37868 23164 37874
rect 23112 37810 23164 37816
rect 23204 37868 23256 37874
rect 23204 37810 23256 37816
rect 22836 36712 22888 36718
rect 22836 36654 22888 36660
rect 22848 36310 22876 36654
rect 22836 36304 22888 36310
rect 22836 36246 22888 36252
rect 22376 36236 22428 36242
rect 22376 36178 22428 36184
rect 22388 35698 22416 36178
rect 22376 35692 22428 35698
rect 22428 35652 22508 35680
rect 22376 35634 22428 35640
rect 22204 34870 22324 34898
rect 22100 34060 22152 34066
rect 22100 34002 22152 34008
rect 22008 33516 22060 33522
rect 22008 33458 22060 33464
rect 21876 32728 21956 32756
rect 21824 32710 21876 32716
rect 22020 32586 22048 33458
rect 22112 33386 22140 34002
rect 22100 33380 22152 33386
rect 22100 33322 22152 33328
rect 21928 32558 22048 32586
rect 21824 32496 21876 32502
rect 21824 32438 21876 32444
rect 21732 31680 21784 31686
rect 21560 31640 21732 31668
rect 21560 30258 21588 31640
rect 21732 31622 21784 31628
rect 21732 31136 21784 31142
rect 21730 31104 21732 31113
rect 21784 31104 21786 31113
rect 21730 31039 21786 31048
rect 21836 30938 21864 32438
rect 21824 30932 21876 30938
rect 21824 30874 21876 30880
rect 21640 30728 21692 30734
rect 21640 30670 21692 30676
rect 21548 30252 21600 30258
rect 21548 30194 21600 30200
rect 21456 30116 21508 30122
rect 21508 30076 21588 30104
rect 21456 30058 21508 30064
rect 21456 29164 21508 29170
rect 21456 29106 21508 29112
rect 21468 28558 21496 29106
rect 21560 28994 21588 30076
rect 21652 30054 21680 30670
rect 21928 30190 21956 32558
rect 22112 31793 22140 33322
rect 22204 32026 22232 34870
rect 22284 33992 22336 33998
rect 22284 33934 22336 33940
rect 22296 33658 22324 33934
rect 22284 33652 22336 33658
rect 22284 33594 22336 33600
rect 22376 33380 22428 33386
rect 22376 33322 22428 33328
rect 22284 32768 22336 32774
rect 22284 32710 22336 32716
rect 22296 32502 22324 32710
rect 22284 32496 22336 32502
rect 22284 32438 22336 32444
rect 22192 32020 22244 32026
rect 22192 31962 22244 31968
rect 22098 31784 22154 31793
rect 22098 31719 22154 31728
rect 22100 31680 22152 31686
rect 22100 31622 22152 31628
rect 22008 31272 22060 31278
rect 22008 31214 22060 31220
rect 22020 30870 22048 31214
rect 22112 31142 22140 31622
rect 22204 31482 22232 31962
rect 22388 31754 22416 33322
rect 22480 32502 22508 35652
rect 23124 35630 23152 37810
rect 23400 37262 23428 38150
rect 24964 38010 24992 38354
rect 25044 38276 25096 38282
rect 25044 38218 25096 38224
rect 24952 38004 25004 38010
rect 24952 37946 25004 37952
rect 23480 37868 23532 37874
rect 23480 37810 23532 37816
rect 23572 37868 23624 37874
rect 23572 37810 23624 37816
rect 23492 37466 23520 37810
rect 23480 37460 23532 37466
rect 23480 37402 23532 37408
rect 23584 37262 23612 37810
rect 24584 37664 24636 37670
rect 24584 37606 24636 37612
rect 24768 37664 24820 37670
rect 24768 37606 24820 37612
rect 23388 37256 23440 37262
rect 23388 37198 23440 37204
rect 23572 37256 23624 37262
rect 23572 37198 23624 37204
rect 24492 37256 24544 37262
rect 24492 37198 24544 37204
rect 22560 35624 22612 35630
rect 22560 35566 22612 35572
rect 23112 35624 23164 35630
rect 23112 35566 23164 35572
rect 22572 34950 22600 35566
rect 23296 35556 23348 35562
rect 23296 35498 23348 35504
rect 22652 35488 22704 35494
rect 22652 35430 22704 35436
rect 22560 34944 22612 34950
rect 22560 34886 22612 34892
rect 22572 34785 22600 34886
rect 22558 34776 22614 34785
rect 22558 34711 22614 34720
rect 22664 34660 22692 35430
rect 23020 35284 23072 35290
rect 23020 35226 23072 35232
rect 22834 35048 22890 35057
rect 22834 34983 22890 34992
rect 22928 35012 22980 35018
rect 22572 34632 22692 34660
rect 22572 34202 22600 34632
rect 22848 34610 22876 34983
rect 22928 34954 22980 34960
rect 22940 34746 22968 34954
rect 22928 34740 22980 34746
rect 22928 34682 22980 34688
rect 23032 34626 23060 35226
rect 23112 35080 23164 35086
rect 23112 35022 23164 35028
rect 23204 35080 23256 35086
rect 23204 35022 23256 35028
rect 23124 34746 23152 35022
rect 23112 34740 23164 34746
rect 23112 34682 23164 34688
rect 22836 34604 22888 34610
rect 23032 34598 23152 34626
rect 22836 34546 22888 34552
rect 22652 34400 22704 34406
rect 22652 34342 22704 34348
rect 22560 34196 22612 34202
rect 22560 34138 22612 34144
rect 22468 32496 22520 32502
rect 22468 32438 22520 32444
rect 22572 32178 22600 34138
rect 22664 33998 22692 34342
rect 22836 34128 22888 34134
rect 22836 34070 22888 34076
rect 22652 33992 22704 33998
rect 22848 33969 22876 34070
rect 22652 33934 22704 33940
rect 22834 33960 22890 33969
rect 22664 32366 22692 33934
rect 22834 33895 22890 33904
rect 22928 33856 22980 33862
rect 22928 33798 22980 33804
rect 22744 32836 22796 32842
rect 22744 32778 22796 32784
rect 22756 32570 22784 32778
rect 22744 32564 22796 32570
rect 22744 32506 22796 32512
rect 22836 32496 22888 32502
rect 22836 32438 22888 32444
rect 22652 32360 22704 32366
rect 22652 32302 22704 32308
rect 22572 32150 22784 32178
rect 22558 31784 22614 31793
rect 22376 31748 22428 31754
rect 22376 31690 22428 31696
rect 22480 31728 22558 31754
rect 22480 31726 22614 31728
rect 22192 31476 22244 31482
rect 22192 31418 22244 31424
rect 22192 31272 22244 31278
rect 22244 31249 22324 31260
rect 22244 31240 22338 31249
rect 22244 31232 22282 31240
rect 22192 31214 22244 31220
rect 22282 31175 22338 31184
rect 22100 31136 22152 31142
rect 22100 31078 22152 31084
rect 22192 31136 22244 31142
rect 22192 31078 22244 31084
rect 22284 31136 22336 31142
rect 22284 31078 22336 31084
rect 22008 30864 22060 30870
rect 22204 30841 22232 31078
rect 22296 30938 22324 31078
rect 22284 30932 22336 30938
rect 22284 30874 22336 30880
rect 22008 30806 22060 30812
rect 22190 30832 22246 30841
rect 22190 30767 22246 30776
rect 22008 30728 22060 30734
rect 22008 30670 22060 30676
rect 22020 30308 22048 30670
rect 22192 30388 22244 30394
rect 22192 30330 22244 30336
rect 22020 30280 22140 30308
rect 21916 30184 21968 30190
rect 21916 30126 21968 30132
rect 21824 30116 21876 30122
rect 21824 30058 21876 30064
rect 21640 30048 21692 30054
rect 21640 29990 21692 29996
rect 21640 29776 21692 29782
rect 21640 29718 21692 29724
rect 21652 29306 21680 29718
rect 21732 29708 21784 29714
rect 21732 29650 21784 29656
rect 21640 29300 21692 29306
rect 21640 29242 21692 29248
rect 21560 28966 21680 28994
rect 21548 28756 21600 28762
rect 21548 28698 21600 28704
rect 21560 28558 21588 28698
rect 21456 28552 21508 28558
rect 21456 28494 21508 28500
rect 21548 28552 21600 28558
rect 21548 28494 21600 28500
rect 21560 28393 21588 28494
rect 21546 28384 21602 28393
rect 21546 28319 21602 28328
rect 21454 28248 21510 28257
rect 21454 28183 21510 28192
rect 21468 27713 21496 28183
rect 21454 27704 21510 27713
rect 21454 27639 21510 27648
rect 21364 24336 21416 24342
rect 21364 24278 21416 24284
rect 21468 23866 21496 27639
rect 21548 26376 21600 26382
rect 21546 26344 21548 26353
rect 21600 26344 21602 26353
rect 21546 26279 21602 26288
rect 21548 25696 21600 25702
rect 21546 25664 21548 25673
rect 21600 25664 21602 25673
rect 21546 25599 21602 25608
rect 21546 25528 21602 25537
rect 21546 25463 21602 25472
rect 21560 25226 21588 25463
rect 21548 25220 21600 25226
rect 21548 25162 21600 25168
rect 21560 24818 21588 25162
rect 21548 24812 21600 24818
rect 21548 24754 21600 24760
rect 21272 23860 21324 23866
rect 21272 23802 21324 23808
rect 21456 23860 21508 23866
rect 21456 23802 21508 23808
rect 21180 23724 21232 23730
rect 21180 23666 21232 23672
rect 21364 23724 21416 23730
rect 21364 23666 21416 23672
rect 21192 23186 21220 23666
rect 21180 23180 21232 23186
rect 21180 23122 21232 23128
rect 21086 22264 21142 22273
rect 21086 22199 21142 22208
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 21086 21992 21142 22001
rect 21086 21927 21142 21936
rect 20996 21888 21048 21894
rect 20996 21830 21048 21836
rect 21008 21690 21036 21830
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 20916 20726 21036 20754
rect 21008 20398 21036 20726
rect 21100 20398 21128 21927
rect 21192 21690 21220 23122
rect 21270 23080 21326 23089
rect 21270 23015 21272 23024
rect 21324 23015 21326 23024
rect 21272 22986 21324 22992
rect 21270 22672 21326 22681
rect 21270 22607 21272 22616
rect 21324 22607 21326 22616
rect 21272 22578 21324 22584
rect 21376 22574 21404 23666
rect 21560 23526 21588 24754
rect 21652 24018 21680 28966
rect 21744 28762 21772 29650
rect 21836 29510 21864 30058
rect 21824 29504 21876 29510
rect 21824 29446 21876 29452
rect 21928 29322 21956 30126
rect 22006 29336 22062 29345
rect 21928 29294 22006 29322
rect 21928 29170 21956 29294
rect 22006 29271 22062 29280
rect 22008 29232 22060 29238
rect 22006 29200 22008 29209
rect 22060 29200 22062 29209
rect 21916 29164 21968 29170
rect 22006 29135 22062 29144
rect 21916 29106 21968 29112
rect 21822 28928 21878 28937
rect 21822 28863 21878 28872
rect 21836 28762 21864 28863
rect 21732 28756 21784 28762
rect 21732 28698 21784 28704
rect 21824 28756 21876 28762
rect 21824 28698 21876 28704
rect 21744 28257 21772 28698
rect 21730 28248 21786 28257
rect 21730 28183 21786 28192
rect 21824 28076 21876 28082
rect 21824 28018 21876 28024
rect 21730 26752 21786 26761
rect 21730 26687 21786 26696
rect 21744 26382 21772 26687
rect 21732 26376 21784 26382
rect 21732 26318 21784 26324
rect 21732 26240 21784 26246
rect 21732 26182 21784 26188
rect 21744 24274 21772 26182
rect 21836 25537 21864 28018
rect 21928 27305 21956 29106
rect 21914 27296 21970 27305
rect 21914 27231 21970 27240
rect 22020 27112 22048 29135
rect 22112 28762 22140 30280
rect 22204 29850 22232 30330
rect 22192 29844 22244 29850
rect 22192 29786 22244 29792
rect 22388 29714 22416 31690
rect 22480 29850 22508 31726
rect 22558 31719 22614 31726
rect 22560 31476 22612 31482
rect 22560 31418 22612 31424
rect 22468 29844 22520 29850
rect 22468 29786 22520 29792
rect 22376 29708 22428 29714
rect 22376 29650 22428 29656
rect 22192 29572 22244 29578
rect 22192 29514 22244 29520
rect 22204 29034 22232 29514
rect 22468 29504 22520 29510
rect 22466 29472 22468 29481
rect 22520 29472 22522 29481
rect 22466 29407 22522 29416
rect 22468 29164 22520 29170
rect 22468 29106 22520 29112
rect 22192 29028 22244 29034
rect 22192 28970 22244 28976
rect 22100 28756 22152 28762
rect 22100 28698 22152 28704
rect 22098 28656 22154 28665
rect 22098 28591 22100 28600
rect 22152 28591 22154 28600
rect 22100 28562 22152 28568
rect 22204 28490 22232 28970
rect 22480 28744 22508 29106
rect 22572 29102 22600 31418
rect 22756 30394 22784 32150
rect 22848 31822 22876 32438
rect 22836 31816 22888 31822
rect 22836 31758 22888 31764
rect 22848 30938 22876 31758
rect 22940 31482 22968 33798
rect 23020 33584 23072 33590
rect 23020 33526 23072 33532
rect 22928 31476 22980 31482
rect 22928 31418 22980 31424
rect 22928 31340 22980 31346
rect 22928 31282 22980 31288
rect 22836 30932 22888 30938
rect 22836 30874 22888 30880
rect 22836 30728 22888 30734
rect 22836 30670 22888 30676
rect 22744 30388 22796 30394
rect 22744 30330 22796 30336
rect 22744 29572 22796 29578
rect 22744 29514 22796 29520
rect 22652 29504 22704 29510
rect 22652 29446 22704 29452
rect 22560 29096 22612 29102
rect 22560 29038 22612 29044
rect 22296 28716 22508 28744
rect 22558 28792 22614 28801
rect 22558 28727 22614 28736
rect 22192 28484 22244 28490
rect 22192 28426 22244 28432
rect 22296 28218 22324 28716
rect 22572 28694 22600 28727
rect 22560 28688 22612 28694
rect 22560 28630 22612 28636
rect 22468 28620 22520 28626
rect 22468 28562 22520 28568
rect 22284 28212 22336 28218
rect 22284 28154 22336 28160
rect 22190 27976 22246 27985
rect 22190 27911 22246 27920
rect 22100 27328 22152 27334
rect 22100 27270 22152 27276
rect 22112 27130 22140 27270
rect 21928 27084 22048 27112
rect 22100 27124 22152 27130
rect 21822 25528 21878 25537
rect 21822 25463 21878 25472
rect 21824 25356 21876 25362
rect 21824 25298 21876 25304
rect 21836 24886 21864 25298
rect 21824 24880 21876 24886
rect 21824 24822 21876 24828
rect 21928 24614 21956 27084
rect 22100 27066 22152 27072
rect 22008 26988 22060 26994
rect 22008 26930 22060 26936
rect 22020 26364 22048 26930
rect 22204 26897 22232 27911
rect 22284 27872 22336 27878
rect 22284 27814 22336 27820
rect 22190 26888 22246 26897
rect 22190 26823 22246 26832
rect 22100 26784 22152 26790
rect 22100 26726 22152 26732
rect 22112 26518 22140 26726
rect 22100 26512 22152 26518
rect 22100 26454 22152 26460
rect 22192 26376 22244 26382
rect 22020 26336 22192 26364
rect 22020 26042 22048 26336
rect 22192 26318 22244 26324
rect 22100 26240 22152 26246
rect 22100 26182 22152 26188
rect 22112 26042 22140 26182
rect 22008 26036 22060 26042
rect 22008 25978 22060 25984
rect 22100 26036 22152 26042
rect 22100 25978 22152 25984
rect 22296 25974 22324 27814
rect 22376 27532 22428 27538
rect 22376 27474 22428 27480
rect 22388 26246 22416 27474
rect 22376 26240 22428 26246
rect 22376 26182 22428 26188
rect 22284 25968 22336 25974
rect 22284 25910 22336 25916
rect 22008 25832 22060 25838
rect 22008 25774 22060 25780
rect 22020 25226 22048 25774
rect 22100 25288 22152 25294
rect 22480 25242 22508 28562
rect 22560 28552 22612 28558
rect 22560 28494 22612 28500
rect 22572 28082 22600 28494
rect 22560 28076 22612 28082
rect 22560 28018 22612 28024
rect 22560 27396 22612 27402
rect 22560 27338 22612 27344
rect 22572 25430 22600 27338
rect 22560 25424 22612 25430
rect 22560 25366 22612 25372
rect 22100 25230 22152 25236
rect 22008 25220 22060 25226
rect 22008 25162 22060 25168
rect 22006 25120 22062 25129
rect 22006 25055 22062 25064
rect 22020 24954 22048 25055
rect 22008 24948 22060 24954
rect 22008 24890 22060 24896
rect 22112 24886 22140 25230
rect 22296 25214 22508 25242
rect 22192 25152 22244 25158
rect 22192 25094 22244 25100
rect 22204 24886 22232 25094
rect 22100 24880 22152 24886
rect 22100 24822 22152 24828
rect 22192 24880 22244 24886
rect 22192 24822 22244 24828
rect 21916 24608 21968 24614
rect 21916 24550 21968 24556
rect 21928 24410 21956 24550
rect 21916 24404 21968 24410
rect 21916 24346 21968 24352
rect 21732 24268 21784 24274
rect 21732 24210 21784 24216
rect 21928 24188 21956 24346
rect 21928 24160 22048 24188
rect 21652 23990 21956 24018
rect 21732 23860 21784 23866
rect 21732 23802 21784 23808
rect 21548 23520 21600 23526
rect 21548 23462 21600 23468
rect 21456 23112 21508 23118
rect 21456 23054 21508 23060
rect 21548 23112 21600 23118
rect 21548 23054 21600 23060
rect 21468 22778 21496 23054
rect 21456 22772 21508 22778
rect 21456 22714 21508 22720
rect 21560 22710 21588 23054
rect 21548 22704 21600 22710
rect 21548 22646 21600 22652
rect 21364 22568 21416 22574
rect 21364 22510 21416 22516
rect 21272 22432 21324 22438
rect 21272 22374 21324 22380
rect 21180 21684 21232 21690
rect 21180 21626 21232 21632
rect 21284 21554 21312 22374
rect 21362 22264 21418 22273
rect 21362 22199 21418 22208
rect 21638 22264 21694 22273
rect 21638 22199 21640 22208
rect 21272 21548 21324 21554
rect 21272 21490 21324 21496
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 21088 20392 21140 20398
rect 21088 20334 21140 20340
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 20640 19922 20852 19938
rect 20628 19916 20864 19922
rect 20680 19910 20812 19916
rect 20628 19858 20680 19864
rect 20812 19858 20864 19864
rect 20444 19712 20496 19718
rect 20444 19654 20496 19660
rect 20536 19712 20588 19718
rect 20536 19654 20588 19660
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 20352 15088 20404 15094
rect 20352 15030 20404 15036
rect 20350 14512 20406 14521
rect 20350 14447 20406 14456
rect 20364 14414 20392 14447
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 20272 11218 20300 11494
rect 20260 11212 20312 11218
rect 20260 11154 20312 11160
rect 20260 10600 20312 10606
rect 20260 10542 20312 10548
rect 20168 10124 20220 10130
rect 20168 10066 20220 10072
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 19432 7948 19484 7954
rect 19536 7936 19564 8434
rect 19484 7908 19564 7936
rect 19432 7890 19484 7896
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 17960 6384 18012 6390
rect 17960 6326 18012 6332
rect 18064 6186 18092 6734
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18052 6180 18104 6186
rect 18052 6122 18104 6128
rect 17868 5636 17920 5642
rect 17868 5578 17920 5584
rect 18052 5636 18104 5642
rect 18052 5578 18104 5584
rect 17880 5166 17908 5578
rect 18064 5234 18092 5578
rect 18708 5302 18736 6598
rect 19076 6390 19104 6802
rect 19352 6390 19380 7482
rect 19444 7342 19472 7890
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19444 6458 19472 6734
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19064 6384 19116 6390
rect 19064 6326 19116 6332
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 18972 6248 19024 6254
rect 18972 6190 19024 6196
rect 18984 6118 19012 6190
rect 18972 6112 19024 6118
rect 18972 6054 19024 6060
rect 18984 5914 19012 6054
rect 18972 5908 19024 5914
rect 18972 5850 19024 5856
rect 19352 5778 19380 6326
rect 20076 6316 20128 6322
rect 20076 6258 20128 6264
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19352 5370 19380 5714
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 18696 5296 18748 5302
rect 18696 5238 18748 5244
rect 18052 5228 18104 5234
rect 18052 5170 18104 5176
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 17880 4622 17908 5102
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 15014 4040 15070 4049
rect 15014 3975 15070 3984
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7116 800 7144 2246
rect 10980 800 11008 3878
rect 14738 3632 14794 3641
rect 15028 3602 15056 3975
rect 14738 3567 14794 3576
rect 15016 3596 15068 3602
rect 14752 3534 14780 3567
rect 15016 3538 15068 3544
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14188 3460 14240 3466
rect 14188 3402 14240 3408
rect 14200 800 14228 3402
rect 14752 3194 14780 3470
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 18064 800 18092 5170
rect 20088 5030 20116 6258
rect 20180 5370 20208 10066
rect 20272 8090 20300 10542
rect 20456 10266 20484 19654
rect 20548 19446 20576 19654
rect 20536 19440 20588 19446
rect 20536 19382 20588 19388
rect 20732 19378 20760 19654
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 20628 19236 20680 19242
rect 20628 19178 20680 19184
rect 20640 18834 20668 19178
rect 20916 18834 20944 20198
rect 21008 19854 21036 20334
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 20904 18828 20956 18834
rect 20904 18770 20956 18776
rect 20996 18828 21048 18834
rect 20996 18770 21048 18776
rect 20536 18624 20588 18630
rect 20536 18566 20588 18572
rect 20548 14822 20576 18566
rect 20640 18426 20668 18770
rect 20628 18420 20680 18426
rect 20628 18362 20680 18368
rect 20916 18154 20944 18770
rect 21008 18737 21036 18770
rect 21100 18766 21128 20334
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 21192 18834 21220 19110
rect 21180 18828 21232 18834
rect 21180 18770 21232 18776
rect 21088 18760 21140 18766
rect 20994 18728 21050 18737
rect 21284 18714 21312 21490
rect 21088 18702 21140 18708
rect 20994 18663 21050 18672
rect 21192 18686 21312 18714
rect 21086 18320 21142 18329
rect 21086 18255 21142 18264
rect 20904 18148 20956 18154
rect 20904 18090 20956 18096
rect 20718 18048 20774 18057
rect 20774 18006 20852 18034
rect 20718 17983 20774 17992
rect 20628 17808 20680 17814
rect 20628 17750 20680 17756
rect 20640 17270 20668 17750
rect 20628 17264 20680 17270
rect 20628 17206 20680 17212
rect 20824 17202 20852 18006
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20718 16960 20774 16969
rect 20640 16590 20668 16934
rect 20718 16895 20774 16904
rect 20732 16794 20760 16895
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20824 16726 20852 17138
rect 20812 16720 20864 16726
rect 20812 16662 20864 16668
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20548 14414 20576 14758
rect 20640 14618 20668 16050
rect 20732 15706 20760 16390
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20536 14408 20588 14414
rect 20536 14350 20588 14356
rect 20732 14346 20760 15370
rect 20824 15026 20852 16662
rect 20904 15088 20956 15094
rect 20902 15056 20904 15065
rect 20956 15056 20958 15065
rect 20812 15020 20864 15026
rect 20902 14991 20958 15000
rect 20812 14962 20864 14968
rect 20720 14340 20772 14346
rect 20720 14282 20772 14288
rect 20732 14074 20760 14282
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20812 13796 20864 13802
rect 20812 13738 20864 13744
rect 20824 13462 20852 13738
rect 20812 13456 20864 13462
rect 20812 13398 20864 13404
rect 20812 13252 20864 13258
rect 20812 13194 20864 13200
rect 20824 12434 20852 13194
rect 20824 12406 21036 12434
rect 20904 12096 20956 12102
rect 20904 12038 20956 12044
rect 20916 11898 20944 12038
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 20720 10736 20772 10742
rect 20720 10678 20772 10684
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 20732 9722 20760 10678
rect 20812 10260 20864 10266
rect 20812 10202 20864 10208
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20824 9178 20852 10202
rect 20916 9994 20944 10746
rect 21008 10248 21036 12406
rect 21100 12306 21128 18255
rect 21192 17610 21220 18686
rect 21180 17604 21232 17610
rect 21180 17546 21232 17552
rect 21192 15502 21220 17546
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 21284 17202 21312 17478
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 21376 17134 21404 22199
rect 21692 22199 21694 22208
rect 21640 22170 21692 22176
rect 21744 22001 21772 23802
rect 21824 23792 21876 23798
rect 21824 23734 21876 23740
rect 21836 22030 21864 23734
rect 21824 22024 21876 22030
rect 21730 21992 21786 22001
rect 21824 21966 21876 21972
rect 21730 21927 21786 21936
rect 21548 21888 21600 21894
rect 21548 21830 21600 21836
rect 21640 21888 21692 21894
rect 21640 21830 21692 21836
rect 21732 21888 21784 21894
rect 21732 21830 21784 21836
rect 21454 21720 21510 21729
rect 21454 21655 21510 21664
rect 21468 20534 21496 21655
rect 21456 20528 21508 20534
rect 21456 20470 21508 20476
rect 21456 20052 21508 20058
rect 21456 19994 21508 20000
rect 21468 18970 21496 19994
rect 21560 19310 21588 21830
rect 21652 21350 21680 21830
rect 21640 21344 21692 21350
rect 21640 21286 21692 21292
rect 21744 21146 21772 21830
rect 21824 21548 21876 21554
rect 21824 21490 21876 21496
rect 21732 21140 21784 21146
rect 21732 21082 21784 21088
rect 21640 20800 21692 20806
rect 21640 20742 21692 20748
rect 21548 19304 21600 19310
rect 21548 19246 21600 19252
rect 21456 18964 21508 18970
rect 21456 18906 21508 18912
rect 21560 18714 21588 19246
rect 21468 18686 21588 18714
rect 21468 17882 21496 18686
rect 21548 18624 21600 18630
rect 21548 18566 21600 18572
rect 21560 18426 21588 18566
rect 21548 18420 21600 18426
rect 21548 18362 21600 18368
rect 21548 18148 21600 18154
rect 21548 18090 21600 18096
rect 21456 17876 21508 17882
rect 21456 17818 21508 17824
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21468 17134 21496 17614
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 21456 17128 21508 17134
rect 21456 17070 21508 17076
rect 21468 16522 21496 17070
rect 21560 16590 21588 18090
rect 21652 17202 21680 20742
rect 21744 19446 21772 21082
rect 21836 21010 21864 21490
rect 21928 21146 21956 23990
rect 22020 22234 22048 24160
rect 22190 23352 22246 23361
rect 22190 23287 22192 23296
rect 22244 23287 22246 23296
rect 22192 23258 22244 23264
rect 22190 22808 22246 22817
rect 22112 22766 22190 22794
rect 22112 22710 22140 22766
rect 22190 22743 22246 22752
rect 22100 22704 22152 22710
rect 22100 22646 22152 22652
rect 22190 22672 22246 22681
rect 22296 22658 22324 25214
rect 22560 24812 22612 24818
rect 22560 24754 22612 24760
rect 22468 24744 22520 24750
rect 22468 24686 22520 24692
rect 22480 24290 22508 24686
rect 22572 24410 22600 24754
rect 22560 24404 22612 24410
rect 22560 24346 22612 24352
rect 22480 24262 22600 24290
rect 22468 24200 22520 24206
rect 22468 24142 22520 24148
rect 22480 23769 22508 24142
rect 22466 23760 22522 23769
rect 22466 23695 22522 23704
rect 22468 23656 22520 23662
rect 22468 23598 22520 23604
rect 22376 23520 22428 23526
rect 22376 23462 22428 23468
rect 22246 22630 22324 22658
rect 22190 22607 22246 22616
rect 22100 22432 22152 22438
rect 22100 22374 22152 22380
rect 22192 22432 22244 22438
rect 22192 22374 22244 22380
rect 22008 22228 22060 22234
rect 22008 22170 22060 22176
rect 22112 22166 22140 22374
rect 22100 22160 22152 22166
rect 22100 22102 22152 22108
rect 22204 21978 22232 22374
rect 22282 22264 22338 22273
rect 22282 22199 22284 22208
rect 22336 22199 22338 22208
rect 22284 22170 22336 22176
rect 22112 21950 22232 21978
rect 22008 21888 22060 21894
rect 22008 21830 22060 21836
rect 21916 21140 21968 21146
rect 21916 21082 21968 21088
rect 22020 21026 22048 21830
rect 21824 21004 21876 21010
rect 21824 20946 21876 20952
rect 21928 20998 22048 21026
rect 22112 21010 22140 21950
rect 22388 21865 22416 23462
rect 22480 22409 22508 23598
rect 22466 22400 22522 22409
rect 22466 22335 22522 22344
rect 22572 22273 22600 24262
rect 22558 22264 22614 22273
rect 22558 22199 22614 22208
rect 22468 22024 22520 22030
rect 22466 21992 22468 22001
rect 22520 21992 22522 22001
rect 22466 21927 22522 21936
rect 22468 21888 22520 21894
rect 22374 21856 22430 21865
rect 22468 21830 22520 21836
rect 22374 21791 22430 21800
rect 22192 21548 22244 21554
rect 22244 21508 22324 21536
rect 22192 21490 22244 21496
rect 22190 21312 22246 21321
rect 22190 21247 22246 21256
rect 22100 21004 22152 21010
rect 21732 19440 21784 19446
rect 21732 19382 21784 19388
rect 21732 18624 21784 18630
rect 21732 18566 21784 18572
rect 21640 17196 21692 17202
rect 21640 17138 21692 17144
rect 21640 16652 21692 16658
rect 21744 16640 21772 18566
rect 21928 17105 21956 20998
rect 22100 20946 22152 20952
rect 22008 20936 22060 20942
rect 22008 20878 22060 20884
rect 22020 20777 22048 20878
rect 22006 20768 22062 20777
rect 22006 20703 22062 20712
rect 22204 20058 22232 21247
rect 22296 21010 22324 21508
rect 22284 21004 22336 21010
rect 22284 20946 22336 20952
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 22296 19854 22324 20946
rect 22480 20890 22508 21830
rect 22388 20874 22508 20890
rect 22376 20868 22508 20874
rect 22428 20862 22508 20868
rect 22376 20810 22428 20816
rect 22468 20800 22520 20806
rect 22468 20742 22520 20748
rect 22374 20360 22430 20369
rect 22374 20295 22430 20304
rect 22388 20262 22416 20295
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 22296 19428 22324 19790
rect 22376 19440 22428 19446
rect 22296 19400 22376 19428
rect 22376 19382 22428 19388
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22006 18864 22062 18873
rect 22006 18799 22008 18808
rect 22060 18799 22062 18808
rect 22008 18770 22060 18776
rect 22204 18698 22232 19314
rect 22376 19304 22428 19310
rect 22376 19246 22428 19252
rect 22192 18692 22244 18698
rect 22192 18634 22244 18640
rect 22008 17672 22060 17678
rect 22008 17614 22060 17620
rect 21914 17096 21970 17105
rect 22020 17082 22048 17614
rect 22020 17054 22140 17082
rect 21914 17031 21970 17040
rect 21928 16980 21956 17031
rect 21928 16952 22048 16980
rect 21824 16788 21876 16794
rect 21824 16730 21876 16736
rect 21692 16612 21772 16640
rect 21640 16594 21692 16600
rect 21548 16584 21600 16590
rect 21548 16526 21600 16532
rect 21456 16516 21508 16522
rect 21456 16458 21508 16464
rect 21456 16176 21508 16182
rect 21376 16124 21456 16130
rect 21376 16118 21508 16124
rect 21376 16102 21496 16118
rect 21180 15496 21232 15502
rect 21180 15438 21232 15444
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 21192 13190 21220 15302
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 21284 15065 21312 15098
rect 21270 15056 21326 15065
rect 21270 14991 21326 15000
rect 21272 14544 21324 14550
rect 21272 14486 21324 14492
rect 21284 13326 21312 14486
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21180 13184 21232 13190
rect 21180 13126 21232 13132
rect 21376 13002 21404 16102
rect 21638 16008 21694 16017
rect 21638 15943 21694 15952
rect 21456 15632 21508 15638
rect 21456 15574 21508 15580
rect 21284 12974 21404 13002
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 21284 12186 21312 12974
rect 21364 12844 21416 12850
rect 21364 12786 21416 12792
rect 21376 12306 21404 12786
rect 21364 12300 21416 12306
rect 21364 12242 21416 12248
rect 21284 12158 21404 12186
rect 21376 12102 21404 12158
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21376 11354 21404 12038
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21468 11014 21496 15574
rect 21652 15502 21680 15943
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21744 15366 21772 16612
rect 21548 15360 21600 15366
rect 21548 15302 21600 15308
rect 21732 15360 21784 15366
rect 21732 15302 21784 15308
rect 21560 12306 21588 15302
rect 21836 15094 21864 16730
rect 21916 16652 21968 16658
rect 21916 16594 21968 16600
rect 21928 16250 21956 16594
rect 22020 16454 22048 16952
rect 22112 16454 22140 17054
rect 22192 16992 22244 16998
rect 22244 16940 22324 16946
rect 22192 16934 22324 16940
rect 22204 16918 22324 16934
rect 22296 16726 22324 16918
rect 22284 16720 22336 16726
rect 22284 16662 22336 16668
rect 22008 16448 22060 16454
rect 22008 16390 22060 16396
rect 22100 16448 22152 16454
rect 22100 16390 22152 16396
rect 21916 16244 21968 16250
rect 21916 16186 21968 16192
rect 22008 15972 22060 15978
rect 22008 15914 22060 15920
rect 22020 15162 22048 15914
rect 22190 15736 22246 15745
rect 22100 15700 22152 15706
rect 22190 15671 22246 15680
rect 22100 15642 22152 15648
rect 22008 15156 22060 15162
rect 22008 15098 22060 15104
rect 21824 15088 21876 15094
rect 21824 15030 21876 15036
rect 21914 15056 21970 15065
rect 21970 15026 22048 15042
rect 21970 15020 22060 15026
rect 21970 15014 22008 15020
rect 21914 14991 21970 15000
rect 22008 14962 22060 14968
rect 21638 14920 21694 14929
rect 21638 14855 21640 14864
rect 21692 14855 21694 14864
rect 21640 14826 21692 14832
rect 22008 14816 22060 14822
rect 22008 14758 22060 14764
rect 22020 14074 22048 14758
rect 22008 14068 22060 14074
rect 22008 14010 22060 14016
rect 21916 12640 21968 12646
rect 21916 12582 21968 12588
rect 21928 12434 21956 12582
rect 21836 12406 21956 12434
rect 21548 12300 21600 12306
rect 21548 12242 21600 12248
rect 21836 11626 21864 12406
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 21824 11620 21876 11626
rect 21824 11562 21876 11568
rect 21456 11008 21508 11014
rect 21456 10950 21508 10956
rect 21638 10976 21694 10985
rect 21638 10911 21694 10920
rect 21456 10532 21508 10538
rect 21456 10474 21508 10480
rect 21468 10266 21496 10474
rect 21652 10470 21680 10911
rect 21640 10464 21692 10470
rect 21640 10406 21692 10412
rect 21456 10260 21508 10266
rect 21008 10220 21128 10248
rect 20996 10124 21048 10130
rect 20996 10066 21048 10072
rect 20904 9988 20956 9994
rect 20904 9930 20956 9936
rect 20812 9172 20864 9178
rect 20812 9114 20864 9120
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20260 8084 20312 8090
rect 20260 8026 20312 8032
rect 20272 7970 20300 8026
rect 20272 7942 20392 7970
rect 20260 7812 20312 7818
rect 20260 7754 20312 7760
rect 20272 7546 20300 7754
rect 20260 7540 20312 7546
rect 20260 7482 20312 7488
rect 20364 7478 20392 7942
rect 20352 7472 20404 7478
rect 20352 7414 20404 7420
rect 20444 6656 20496 6662
rect 20444 6598 20496 6604
rect 20456 6458 20484 6598
rect 20640 6458 20668 8230
rect 20824 8090 20852 9114
rect 21008 9042 21036 10066
rect 20996 9036 21048 9042
rect 20996 8978 21048 8984
rect 21100 8838 21128 10220
rect 21456 10202 21508 10208
rect 21652 10062 21680 10406
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 21640 10056 21692 10062
rect 21640 9998 21692 10004
rect 21192 9654 21220 9998
rect 21272 9988 21324 9994
rect 21272 9930 21324 9936
rect 21180 9648 21232 9654
rect 21180 9590 21232 9596
rect 21284 9110 21312 9930
rect 21824 9512 21876 9518
rect 21824 9454 21876 9460
rect 21836 9178 21864 9454
rect 21824 9172 21876 9178
rect 21824 9114 21876 9120
rect 21272 9104 21324 9110
rect 21272 9046 21324 9052
rect 21928 8906 21956 12242
rect 22112 11286 22140 15642
rect 22204 15502 22232 15671
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 22192 15156 22244 15162
rect 22192 15098 22244 15104
rect 22204 13462 22232 15098
rect 22296 14822 22324 16662
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22192 13456 22244 13462
rect 22192 13398 22244 13404
rect 22388 13258 22416 19246
rect 22192 13252 22244 13258
rect 22376 13252 22428 13258
rect 22192 13194 22244 13200
rect 22296 13212 22376 13240
rect 22204 12850 22232 13194
rect 22296 12986 22324 13212
rect 22376 13194 22428 13200
rect 22284 12980 22336 12986
rect 22284 12922 22336 12928
rect 22480 12918 22508 20742
rect 22572 19174 22600 22199
rect 22560 19168 22612 19174
rect 22560 19110 22612 19116
rect 22664 17954 22692 29446
rect 22756 29238 22784 29514
rect 22744 29232 22796 29238
rect 22744 29174 22796 29180
rect 22744 28416 22796 28422
rect 22744 28358 22796 28364
rect 22756 28014 22784 28358
rect 22848 28150 22876 30670
rect 22836 28144 22888 28150
rect 22836 28086 22888 28092
rect 22744 28008 22796 28014
rect 22744 27950 22796 27956
rect 22744 27328 22796 27334
rect 22744 27270 22796 27276
rect 22756 26790 22784 27270
rect 22940 27130 22968 31282
rect 23032 30666 23060 33526
rect 23124 30938 23152 34598
rect 23216 33930 23244 35022
rect 23204 33924 23256 33930
rect 23204 33866 23256 33872
rect 23112 30932 23164 30938
rect 23112 30874 23164 30880
rect 23216 30818 23244 33866
rect 23308 31754 23336 35498
rect 23400 35222 23428 37198
rect 23756 37120 23808 37126
rect 23756 37062 23808 37068
rect 24504 37074 24532 37198
rect 24596 37194 24624 37606
rect 24780 37482 24808 37606
rect 24688 37454 24900 37482
rect 24688 37262 24716 37454
rect 24676 37256 24728 37262
rect 24676 37198 24728 37204
rect 24584 37188 24636 37194
rect 24584 37130 24636 37136
rect 23768 36786 23796 37062
rect 24504 37046 24808 37074
rect 24780 36922 24808 37046
rect 24768 36916 24820 36922
rect 24768 36858 24820 36864
rect 23756 36780 23808 36786
rect 23756 36722 23808 36728
rect 23940 36780 23992 36786
rect 23940 36722 23992 36728
rect 23768 36378 23796 36722
rect 23756 36372 23808 36378
rect 23756 36314 23808 36320
rect 23480 35828 23532 35834
rect 23480 35770 23532 35776
rect 23388 35216 23440 35222
rect 23388 35158 23440 35164
rect 23492 34746 23520 35770
rect 23952 35766 23980 36722
rect 24216 36304 24268 36310
rect 24216 36246 24268 36252
rect 24124 36032 24176 36038
rect 24124 35974 24176 35980
rect 23940 35760 23992 35766
rect 23940 35702 23992 35708
rect 24136 35698 24164 35974
rect 24124 35692 24176 35698
rect 24124 35634 24176 35640
rect 24122 35320 24178 35329
rect 24122 35255 24178 35264
rect 23572 35216 23624 35222
rect 23572 35158 23624 35164
rect 23938 35184 23994 35193
rect 23480 34740 23532 34746
rect 23480 34682 23532 34688
rect 23584 33998 23612 35158
rect 23938 35119 23994 35128
rect 23664 34944 23716 34950
rect 23664 34886 23716 34892
rect 23572 33992 23624 33998
rect 23572 33934 23624 33940
rect 23388 33040 23440 33046
rect 23388 32982 23440 32988
rect 23296 31748 23348 31754
rect 23296 31690 23348 31696
rect 23308 31657 23336 31690
rect 23294 31648 23350 31657
rect 23294 31583 23350 31592
rect 23124 30790 23244 30818
rect 23020 30660 23072 30666
rect 23020 30602 23072 30608
rect 23020 29708 23072 29714
rect 23020 29650 23072 29656
rect 23032 28762 23060 29650
rect 23020 28756 23072 28762
rect 23020 28698 23072 28704
rect 23020 28552 23072 28558
rect 23018 28520 23020 28529
rect 23072 28520 23074 28529
rect 23018 28455 23074 28464
rect 23020 28144 23072 28150
rect 23020 28086 23072 28092
rect 23032 27452 23060 28086
rect 23124 27606 23152 30790
rect 23400 30682 23428 32982
rect 23480 32768 23532 32774
rect 23480 32710 23532 32716
rect 23492 31906 23520 32710
rect 23676 32026 23704 34886
rect 23952 34678 23980 35119
rect 24136 35086 24164 35255
rect 24228 35154 24256 36246
rect 24676 35828 24728 35834
rect 24676 35770 24728 35776
rect 24688 35698 24716 35770
rect 24584 35692 24636 35698
rect 24584 35634 24636 35640
rect 24676 35692 24728 35698
rect 24676 35634 24728 35640
rect 24596 35494 24624 35634
rect 24400 35488 24452 35494
rect 24584 35488 24636 35494
rect 24452 35448 24532 35476
rect 24400 35430 24452 35436
rect 24216 35148 24268 35154
rect 24216 35090 24268 35096
rect 24124 35080 24176 35086
rect 24124 35022 24176 35028
rect 24400 35080 24452 35086
rect 24400 35022 24452 35028
rect 24308 34944 24360 34950
rect 24308 34886 24360 34892
rect 23940 34672 23992 34678
rect 23940 34614 23992 34620
rect 24320 34542 24348 34886
rect 24308 34536 24360 34542
rect 24308 34478 24360 34484
rect 24412 34406 24440 35022
rect 23848 34400 23900 34406
rect 23848 34342 23900 34348
rect 24400 34400 24452 34406
rect 24400 34342 24452 34348
rect 23756 32292 23808 32298
rect 23756 32234 23808 32240
rect 23664 32020 23716 32026
rect 23664 31962 23716 31968
rect 23492 31878 23704 31906
rect 23480 31816 23532 31822
rect 23480 31758 23532 31764
rect 23216 30654 23428 30682
rect 23216 29646 23244 30654
rect 23296 30592 23348 30598
rect 23296 30534 23348 30540
rect 23204 29640 23256 29646
rect 23204 29582 23256 29588
rect 23204 29504 23256 29510
rect 23204 29446 23256 29452
rect 23216 27606 23244 29446
rect 23112 27600 23164 27606
rect 23112 27542 23164 27548
rect 23204 27600 23256 27606
rect 23204 27542 23256 27548
rect 23032 27424 23244 27452
rect 23020 27328 23072 27334
rect 23020 27270 23072 27276
rect 22928 27124 22980 27130
rect 22848 27084 22928 27112
rect 22848 26994 22876 27084
rect 22928 27066 22980 27072
rect 22836 26988 22888 26994
rect 22836 26930 22888 26936
rect 22744 26784 22796 26790
rect 22744 26726 22796 26732
rect 22756 26586 22784 26726
rect 22744 26580 22796 26586
rect 22744 26522 22796 26528
rect 22744 26376 22796 26382
rect 22744 26318 22796 26324
rect 22756 25294 22784 26318
rect 23032 25770 23060 27270
rect 23110 26888 23166 26897
rect 23110 26823 23166 26832
rect 23020 25764 23072 25770
rect 23020 25706 23072 25712
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 22928 24812 22980 24818
rect 22928 24754 22980 24760
rect 23020 24812 23072 24818
rect 23020 24754 23072 24760
rect 22744 24200 22796 24206
rect 22742 24168 22744 24177
rect 22796 24168 22798 24177
rect 22742 24103 22798 24112
rect 22756 23322 22784 24103
rect 22940 23866 22968 24754
rect 23032 24614 23060 24754
rect 23020 24608 23072 24614
rect 23020 24550 23072 24556
rect 23020 24200 23072 24206
rect 23020 24142 23072 24148
rect 22928 23860 22980 23866
rect 22928 23802 22980 23808
rect 22834 23760 22890 23769
rect 22834 23695 22890 23704
rect 22744 23316 22796 23322
rect 22744 23258 22796 23264
rect 22756 22438 22784 23258
rect 22848 22982 22876 23695
rect 22928 23180 22980 23186
rect 22928 23122 22980 23128
rect 22836 22976 22888 22982
rect 22940 22953 22968 23122
rect 22836 22918 22888 22924
rect 22926 22944 22982 22953
rect 22848 22642 22876 22918
rect 22926 22879 22982 22888
rect 22926 22808 22982 22817
rect 22926 22743 22928 22752
rect 22980 22743 22982 22752
rect 22928 22714 22980 22720
rect 22836 22636 22888 22642
rect 22836 22578 22888 22584
rect 22744 22432 22796 22438
rect 22744 22374 22796 22380
rect 22848 22250 22876 22578
rect 22756 22222 22876 22250
rect 22756 21554 22784 22222
rect 22836 22024 22888 22030
rect 22836 21966 22888 21972
rect 22744 21548 22796 21554
rect 22744 21490 22796 21496
rect 22744 21412 22796 21418
rect 22744 21354 22796 21360
rect 22756 21060 22784 21354
rect 22848 21128 22876 21966
rect 22940 21690 22968 22714
rect 23032 22710 23060 24142
rect 23020 22704 23072 22710
rect 23020 22646 23072 22652
rect 23032 22506 23060 22646
rect 23020 22500 23072 22506
rect 23020 22442 23072 22448
rect 23020 22160 23072 22166
rect 23020 22102 23072 22108
rect 23032 21894 23060 22102
rect 23020 21888 23072 21894
rect 23020 21830 23072 21836
rect 22928 21684 22980 21690
rect 22928 21626 22980 21632
rect 23032 21418 23060 21830
rect 23020 21412 23072 21418
rect 23020 21354 23072 21360
rect 22848 21100 23060 21128
rect 22756 21032 22876 21060
rect 22848 18834 22876 21032
rect 22928 20936 22980 20942
rect 22928 20878 22980 20884
rect 22940 20602 22968 20878
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 23032 20346 23060 21100
rect 23124 20942 23152 26823
rect 23216 26790 23244 27424
rect 23204 26784 23256 26790
rect 23204 26726 23256 26732
rect 23216 24154 23244 26726
rect 23308 24410 23336 30534
rect 23388 29640 23440 29646
rect 23388 29582 23440 29588
rect 23400 29034 23428 29582
rect 23492 29306 23520 31758
rect 23572 31680 23624 31686
rect 23572 31622 23624 31628
rect 23584 31346 23612 31622
rect 23572 31340 23624 31346
rect 23572 31282 23624 31288
rect 23676 30104 23704 31878
rect 23768 31482 23796 32234
rect 23860 31929 23888 34342
rect 24124 33992 24176 33998
rect 24044 33952 24124 33980
rect 24044 33454 24072 33952
rect 24124 33934 24176 33940
rect 24216 33856 24268 33862
rect 24216 33798 24268 33804
rect 24032 33448 24084 33454
rect 24032 33390 24084 33396
rect 24228 32502 24256 33798
rect 24216 32496 24268 32502
rect 24216 32438 24268 32444
rect 24400 32360 24452 32366
rect 24400 32302 24452 32308
rect 24216 32292 24268 32298
rect 24216 32234 24268 32240
rect 24228 32026 24256 32234
rect 24308 32224 24360 32230
rect 24308 32166 24360 32172
rect 24124 32020 24176 32026
rect 24124 31962 24176 31968
rect 24216 32020 24268 32026
rect 24216 31962 24268 31968
rect 23846 31920 23902 31929
rect 23846 31855 23902 31864
rect 23756 31476 23808 31482
rect 23756 31418 23808 31424
rect 23860 31346 23888 31855
rect 24136 31482 24164 31962
rect 24320 31521 24348 32166
rect 24306 31512 24362 31521
rect 24032 31476 24084 31482
rect 24032 31418 24084 31424
rect 24124 31476 24176 31482
rect 24306 31447 24362 31456
rect 24124 31418 24176 31424
rect 24044 31385 24072 31418
rect 24030 31376 24086 31385
rect 23848 31340 23900 31346
rect 24320 31362 24348 31447
rect 24030 31311 24086 31320
rect 24129 31340 24181 31346
rect 23848 31282 23900 31288
rect 24228 31334 24348 31362
rect 24228 31328 24256 31334
rect 24181 31300 24256 31328
rect 24129 31282 24181 31288
rect 23940 31272 23992 31278
rect 23940 31214 23992 31220
rect 23756 30728 23808 30734
rect 23756 30670 23808 30676
rect 23768 30394 23796 30670
rect 23756 30388 23808 30394
rect 23756 30330 23808 30336
rect 23584 30076 23704 30104
rect 23480 29300 23532 29306
rect 23480 29242 23532 29248
rect 23480 29164 23532 29170
rect 23480 29106 23532 29112
rect 23388 29028 23440 29034
rect 23388 28970 23440 28976
rect 23492 28558 23520 29106
rect 23584 28694 23612 30076
rect 23848 29708 23900 29714
rect 23848 29650 23900 29656
rect 23664 29504 23716 29510
rect 23664 29446 23716 29452
rect 23572 28688 23624 28694
rect 23572 28630 23624 28636
rect 23676 28558 23704 29446
rect 23388 28552 23440 28558
rect 23388 28494 23440 28500
rect 23480 28552 23532 28558
rect 23664 28552 23716 28558
rect 23480 28494 23532 28500
rect 23570 28520 23626 28529
rect 23400 28218 23428 28494
rect 23756 28552 23808 28558
rect 23664 28494 23716 28500
rect 23754 28520 23756 28529
rect 23808 28520 23810 28529
rect 23570 28455 23626 28464
rect 23754 28455 23810 28464
rect 23388 28212 23440 28218
rect 23388 28154 23440 28160
rect 23480 28008 23532 28014
rect 23480 27950 23532 27956
rect 23388 27600 23440 27606
rect 23388 27542 23440 27548
rect 23400 27130 23428 27542
rect 23388 27124 23440 27130
rect 23388 27066 23440 27072
rect 23388 26444 23440 26450
rect 23388 26386 23440 26392
rect 23400 26353 23428 26386
rect 23386 26344 23442 26353
rect 23386 26279 23442 26288
rect 23388 25220 23440 25226
rect 23388 25162 23440 25168
rect 23296 24404 23348 24410
rect 23296 24346 23348 24352
rect 23294 24304 23350 24313
rect 23294 24239 23296 24248
rect 23348 24239 23350 24248
rect 23296 24210 23348 24216
rect 23216 24138 23336 24154
rect 23216 24132 23348 24138
rect 23216 24126 23296 24132
rect 23296 24074 23348 24080
rect 23202 22944 23258 22953
rect 23202 22879 23258 22888
rect 23216 22166 23244 22879
rect 23204 22160 23256 22166
rect 23202 22128 23204 22137
rect 23256 22128 23258 22137
rect 23202 22063 23258 22072
rect 23308 22030 23336 24074
rect 23400 23118 23428 25162
rect 23492 23798 23520 27950
rect 23584 27130 23612 28455
rect 23860 28218 23888 29650
rect 23952 29209 23980 31214
rect 23938 29200 23994 29209
rect 23938 29135 23994 29144
rect 24032 28756 24084 28762
rect 24032 28698 24084 28704
rect 24044 28422 24072 28698
rect 24032 28416 24084 28422
rect 24032 28358 24084 28364
rect 23848 28212 23900 28218
rect 24044 28200 24072 28358
rect 23848 28154 23900 28160
rect 23952 28172 24072 28200
rect 23756 28144 23808 28150
rect 23756 28086 23808 28092
rect 23664 28008 23716 28014
rect 23664 27950 23716 27956
rect 23572 27124 23624 27130
rect 23572 27066 23624 27072
rect 23572 26920 23624 26926
rect 23572 26862 23624 26868
rect 23584 26234 23612 26862
rect 23676 26586 23704 27950
rect 23768 26586 23796 28086
rect 23848 27532 23900 27538
rect 23848 27474 23900 27480
rect 23664 26580 23716 26586
rect 23664 26522 23716 26528
rect 23756 26580 23808 26586
rect 23756 26522 23808 26528
rect 23664 26376 23716 26382
rect 23662 26344 23664 26353
rect 23756 26376 23808 26382
rect 23716 26344 23718 26353
rect 23756 26318 23808 26324
rect 23662 26279 23718 26288
rect 23584 26206 23704 26234
rect 23572 26036 23624 26042
rect 23572 25978 23624 25984
rect 23480 23792 23532 23798
rect 23480 23734 23532 23740
rect 23478 23624 23534 23633
rect 23478 23559 23480 23568
rect 23532 23559 23534 23568
rect 23480 23530 23532 23536
rect 23584 23497 23612 25978
rect 23676 24954 23704 26206
rect 23768 26042 23796 26318
rect 23756 26036 23808 26042
rect 23756 25978 23808 25984
rect 23664 24948 23716 24954
rect 23664 24890 23716 24896
rect 23860 24698 23888 27474
rect 23952 26246 23980 28172
rect 24032 28076 24084 28082
rect 24032 28018 24084 28024
rect 24044 27985 24072 28018
rect 24030 27976 24086 27985
rect 24030 27911 24086 27920
rect 24044 26926 24072 27911
rect 24032 26920 24084 26926
rect 24032 26862 24084 26868
rect 24032 26784 24084 26790
rect 24032 26726 24084 26732
rect 24044 26586 24072 26726
rect 24032 26580 24084 26586
rect 24032 26522 24084 26528
rect 23940 26240 23992 26246
rect 23940 26182 23992 26188
rect 23860 24670 24072 24698
rect 23848 24608 23900 24614
rect 23848 24550 23900 24556
rect 23662 24440 23718 24449
rect 23662 24375 23718 24384
rect 23676 24138 23704 24375
rect 23664 24132 23716 24138
rect 23664 24074 23716 24080
rect 23676 23633 23704 24074
rect 23860 24070 23888 24550
rect 23848 24064 23900 24070
rect 23848 24006 23900 24012
rect 23846 23896 23902 23905
rect 23846 23831 23902 23840
rect 23860 23730 23888 23831
rect 23848 23724 23900 23730
rect 23848 23666 23900 23672
rect 23662 23624 23718 23633
rect 23662 23559 23718 23568
rect 23756 23520 23808 23526
rect 23570 23488 23626 23497
rect 23756 23462 23808 23468
rect 23570 23423 23626 23432
rect 23662 23216 23718 23225
rect 23662 23151 23718 23160
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 23400 22817 23428 23054
rect 23572 22976 23624 22982
rect 23492 22936 23572 22964
rect 23386 22808 23442 22817
rect 23386 22743 23442 22752
rect 23296 22024 23348 22030
rect 23296 21966 23348 21972
rect 23492 21944 23520 22936
rect 23572 22918 23624 22924
rect 23676 22778 23704 23151
rect 23664 22772 23716 22778
rect 23664 22714 23716 22720
rect 23768 22658 23796 23462
rect 23940 23316 23992 23322
rect 23940 23258 23992 23264
rect 23676 22630 23796 22658
rect 23570 22400 23626 22409
rect 23570 22335 23626 22344
rect 23584 21962 23612 22335
rect 23400 21916 23520 21944
rect 23572 21956 23624 21962
rect 23204 21072 23256 21078
rect 23202 21040 23204 21049
rect 23256 21040 23258 21049
rect 23202 20975 23258 20984
rect 23112 20936 23164 20942
rect 23110 20904 23112 20913
rect 23164 20904 23166 20913
rect 23110 20839 23166 20848
rect 23400 20788 23428 21916
rect 23572 21898 23624 21904
rect 23478 21856 23534 21865
rect 23478 21791 23534 21800
rect 22940 20318 23060 20346
rect 23124 20760 23428 20788
rect 22940 19553 22968 20318
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 23032 19718 23060 20198
rect 23020 19712 23072 19718
rect 23020 19654 23072 19660
rect 22926 19544 22982 19553
rect 22926 19479 22982 19488
rect 22836 18828 22888 18834
rect 22836 18770 22888 18776
rect 22664 17926 22784 17954
rect 22650 17232 22706 17241
rect 22756 17202 22784 17926
rect 22836 17604 22888 17610
rect 22836 17546 22888 17552
rect 22650 17167 22652 17176
rect 22704 17167 22706 17176
rect 22744 17196 22796 17202
rect 22652 17138 22704 17144
rect 22744 17138 22796 17144
rect 22560 16992 22612 16998
rect 22560 16934 22612 16940
rect 22572 15978 22600 16934
rect 22664 16794 22692 17138
rect 22652 16788 22704 16794
rect 22652 16730 22704 16736
rect 22560 15972 22612 15978
rect 22560 15914 22612 15920
rect 22744 15700 22796 15706
rect 22744 15642 22796 15648
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 22560 14816 22612 14822
rect 22560 14758 22612 14764
rect 22572 14550 22600 14758
rect 22664 14657 22692 15438
rect 22756 15026 22784 15642
rect 22744 15020 22796 15026
rect 22744 14962 22796 14968
rect 22650 14648 22706 14657
rect 22650 14583 22706 14592
rect 22560 14544 22612 14550
rect 22560 14486 22612 14492
rect 22468 12912 22520 12918
rect 22468 12854 22520 12860
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22100 11280 22152 11286
rect 22664 11234 22692 14583
rect 22742 14512 22798 14521
rect 22742 14447 22798 14456
rect 22756 14346 22784 14447
rect 22744 14340 22796 14346
rect 22744 14282 22796 14288
rect 22848 14006 22876 17546
rect 22940 16590 22968 19479
rect 23018 17504 23074 17513
rect 23018 17439 23074 17448
rect 23032 17202 23060 17439
rect 23020 17196 23072 17202
rect 23020 17138 23072 17144
rect 22928 16584 22980 16590
rect 22928 16526 22980 16532
rect 23020 14272 23072 14278
rect 23020 14214 23072 14220
rect 22836 14000 22888 14006
rect 22836 13942 22888 13948
rect 22744 13320 22796 13326
rect 22744 13262 22796 13268
rect 22756 11801 22784 13262
rect 22848 13190 22876 13942
rect 23032 13530 23060 14214
rect 23020 13524 23072 13530
rect 23020 13466 23072 13472
rect 22836 13184 22888 13190
rect 22836 13126 22888 13132
rect 23124 12102 23152 20760
rect 23294 20632 23350 20641
rect 23294 20567 23350 20576
rect 23308 20466 23336 20567
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 23202 19680 23258 19689
rect 23202 19615 23258 19624
rect 23216 19378 23244 19615
rect 23204 19372 23256 19378
rect 23204 19314 23256 19320
rect 23204 19168 23256 19174
rect 23204 19110 23256 19116
rect 23216 18970 23244 19110
rect 23204 18964 23256 18970
rect 23204 18906 23256 18912
rect 23308 18850 23336 20402
rect 23492 20330 23520 21791
rect 23572 21616 23624 21622
rect 23572 21558 23624 21564
rect 23584 20466 23612 21558
rect 23676 21010 23704 22630
rect 23952 22506 23980 23258
rect 24044 22642 24072 24670
rect 24032 22636 24084 22642
rect 24032 22578 24084 22584
rect 23848 22500 23900 22506
rect 23848 22442 23900 22448
rect 23940 22500 23992 22506
rect 23940 22442 23992 22448
rect 23860 22094 23888 22442
rect 23768 22066 23888 22094
rect 23664 21004 23716 21010
rect 23664 20946 23716 20952
rect 23572 20460 23624 20466
rect 23572 20402 23624 20408
rect 23480 20324 23532 20330
rect 23480 20266 23532 20272
rect 23388 19712 23440 19718
rect 23388 19654 23440 19660
rect 23216 18822 23336 18850
rect 23216 17270 23244 18822
rect 23400 18766 23428 19654
rect 23584 19378 23612 20402
rect 23676 19530 23704 20946
rect 23768 19666 23796 22066
rect 23952 22030 23980 22442
rect 23940 22024 23992 22030
rect 23940 21966 23992 21972
rect 23848 21956 23900 21962
rect 23848 21898 23900 21904
rect 23860 21690 23888 21898
rect 23848 21684 23900 21690
rect 23848 21626 23900 21632
rect 23848 21548 23900 21554
rect 23848 21490 23900 21496
rect 23860 19854 23888 21490
rect 23940 21344 23992 21350
rect 23940 21286 23992 21292
rect 23952 20942 23980 21286
rect 23940 20936 23992 20942
rect 23940 20878 23992 20884
rect 24044 19854 24072 22578
rect 24136 22166 24164 31282
rect 24308 31272 24360 31278
rect 24308 31214 24360 31220
rect 24216 30932 24268 30938
rect 24216 30874 24268 30880
rect 24228 29170 24256 30874
rect 24320 30190 24348 31214
rect 24412 30938 24440 32302
rect 24504 31890 24532 35448
rect 24584 35430 24636 35436
rect 24584 35216 24636 35222
rect 24582 35184 24584 35193
rect 24636 35184 24638 35193
rect 24582 35119 24638 35128
rect 24596 35086 24624 35119
rect 24584 35080 24636 35086
rect 24584 35022 24636 35028
rect 24582 34640 24638 34649
rect 24688 34626 24716 35634
rect 24780 35630 24808 36858
rect 24872 35630 24900 37454
rect 24952 37392 25004 37398
rect 25056 37380 25084 38218
rect 25320 38208 25372 38214
rect 25320 38150 25372 38156
rect 25332 38010 25360 38150
rect 25320 38004 25372 38010
rect 25320 37946 25372 37952
rect 25504 37800 25556 37806
rect 25504 37742 25556 37748
rect 25004 37352 25084 37380
rect 24952 37334 25004 37340
rect 25228 37324 25280 37330
rect 25228 37266 25280 37272
rect 25240 36922 25268 37266
rect 25516 37194 25544 37742
rect 25608 37670 25636 38898
rect 25688 37936 25740 37942
rect 25688 37878 25740 37884
rect 25596 37664 25648 37670
rect 25596 37606 25648 37612
rect 25504 37188 25556 37194
rect 25504 37130 25556 37136
rect 25228 36916 25280 36922
rect 25228 36858 25280 36864
rect 25042 35864 25098 35873
rect 24964 35834 25042 35850
rect 24952 35828 25042 35834
rect 25004 35822 25042 35828
rect 25042 35799 25098 35808
rect 25320 35828 25372 35834
rect 24952 35770 25004 35776
rect 25320 35770 25372 35776
rect 25228 35760 25280 35766
rect 25056 35720 25228 35748
rect 24768 35624 24820 35630
rect 24768 35566 24820 35572
rect 24860 35624 24912 35630
rect 24860 35566 24912 35572
rect 24780 34746 24808 35566
rect 24768 34740 24820 34746
rect 24768 34682 24820 34688
rect 24638 34598 24716 34626
rect 24582 34575 24638 34584
rect 24584 34468 24636 34474
rect 24584 34410 24636 34416
rect 24492 31884 24544 31890
rect 24492 31826 24544 31832
rect 24596 31346 24624 34410
rect 24872 34134 24900 35566
rect 24950 35320 25006 35329
rect 24950 35255 25006 35264
rect 24860 34128 24912 34134
rect 24860 34070 24912 34076
rect 24860 33992 24912 33998
rect 24860 33934 24912 33940
rect 24964 33946 24992 35255
rect 25056 35086 25084 35720
rect 25228 35702 25280 35708
rect 25136 35488 25188 35494
rect 25136 35430 25188 35436
rect 25148 35290 25176 35430
rect 25136 35284 25188 35290
rect 25136 35226 25188 35232
rect 25332 35086 25360 35770
rect 25516 35476 25544 37130
rect 25596 36168 25648 36174
rect 25596 36110 25648 36116
rect 25608 35698 25636 36110
rect 25700 35698 25728 37878
rect 25792 37126 25820 38898
rect 26068 37262 26096 38898
rect 26160 38418 26188 39442
rect 27632 38554 27660 43982
rect 27710 43893 27766 43982
rect 30930 43893 30986 44693
rect 34794 44010 34850 44693
rect 34794 43982 35112 44010
rect 34794 43893 34850 43982
rect 30944 42226 30972 43893
rect 35084 42362 35112 43982
rect 38658 43893 38714 44693
rect 41878 43893 41934 44693
rect 35072 42356 35124 42362
rect 35072 42298 35124 42304
rect 34518 42256 34574 42265
rect 30932 42220 30984 42226
rect 38672 42226 38700 43893
rect 34518 42191 34520 42200
rect 30932 42162 30984 42168
rect 34572 42191 34574 42200
rect 38660 42220 38712 42226
rect 34520 42162 34572 42168
rect 38660 42162 38712 42168
rect 31300 42152 31352 42158
rect 31300 42094 31352 42100
rect 37188 42152 37240 42158
rect 37188 42094 37240 42100
rect 31312 41449 31340 42094
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 31298 41440 31354 41449
rect 37200 41414 37228 42094
rect 31298 41375 31354 41384
rect 36924 41386 37228 41414
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 27712 39364 27764 39370
rect 27712 39306 27764 39312
rect 27620 38548 27672 38554
rect 27620 38490 27672 38496
rect 26148 38412 26200 38418
rect 26148 38354 26200 38360
rect 26160 37806 26188 38354
rect 26424 38208 26476 38214
rect 26424 38150 26476 38156
rect 26436 37942 26464 38150
rect 27724 37942 27752 39306
rect 27804 39296 27856 39302
rect 27804 39238 27856 39244
rect 27816 38962 27844 39238
rect 27804 38956 27856 38962
rect 27856 38916 28028 38944
rect 27804 38898 27856 38904
rect 27896 38276 27948 38282
rect 27896 38218 27948 38224
rect 27804 38208 27856 38214
rect 27804 38150 27856 38156
rect 26424 37936 26476 37942
rect 26424 37878 26476 37884
rect 27712 37936 27764 37942
rect 27712 37878 27764 37884
rect 26148 37800 26200 37806
rect 26148 37742 26200 37748
rect 27252 37800 27304 37806
rect 27252 37742 27304 37748
rect 27264 37466 27292 37742
rect 27252 37460 27304 37466
rect 27252 37402 27304 37408
rect 27620 37392 27672 37398
rect 27620 37334 27672 37340
rect 27528 37324 27580 37330
rect 27528 37266 27580 37272
rect 25964 37256 26016 37262
rect 25964 37198 26016 37204
rect 26056 37256 26108 37262
rect 26056 37198 26108 37204
rect 25780 37120 25832 37126
rect 25780 37062 25832 37068
rect 25976 36310 26004 37198
rect 26240 37188 26292 37194
rect 26240 37130 26292 37136
rect 27436 37188 27488 37194
rect 27436 37130 27488 37136
rect 25964 36304 26016 36310
rect 25964 36246 26016 36252
rect 25872 36100 25924 36106
rect 25872 36042 25924 36048
rect 25964 36100 26016 36106
rect 25964 36042 26016 36048
rect 25596 35692 25648 35698
rect 25596 35634 25648 35640
rect 25688 35692 25740 35698
rect 25688 35634 25740 35640
rect 25884 35630 25912 36042
rect 25872 35624 25924 35630
rect 25872 35566 25924 35572
rect 25688 35488 25740 35494
rect 25516 35448 25688 35476
rect 25688 35430 25740 35436
rect 25044 35080 25096 35086
rect 25044 35022 25096 35028
rect 25136 35080 25188 35086
rect 25136 35022 25188 35028
rect 25320 35080 25372 35086
rect 25412 35080 25464 35086
rect 25320 35022 25372 35028
rect 25410 35048 25412 35057
rect 25504 35080 25556 35086
rect 25464 35048 25466 35057
rect 25044 34944 25096 34950
rect 25044 34886 25096 34892
rect 25056 34202 25084 34886
rect 25044 34196 25096 34202
rect 25044 34138 25096 34144
rect 24676 33856 24728 33862
rect 24676 33798 24728 33804
rect 24766 33824 24822 33833
rect 24688 32978 24716 33798
rect 24766 33759 24822 33768
rect 24780 33114 24808 33759
rect 24872 33522 24900 33934
rect 24964 33918 25084 33946
rect 24860 33516 24912 33522
rect 24860 33458 24912 33464
rect 24768 33108 24820 33114
rect 24768 33050 24820 33056
rect 24676 32972 24728 32978
rect 24676 32914 24728 32920
rect 24688 32858 24716 32914
rect 24688 32830 24808 32858
rect 24676 32768 24728 32774
rect 24676 32710 24728 32716
rect 24688 32230 24716 32710
rect 24780 32570 24808 32830
rect 24860 32836 24912 32842
rect 24860 32778 24912 32784
rect 24768 32564 24820 32570
rect 24768 32506 24820 32512
rect 24872 32502 24900 32778
rect 24860 32496 24912 32502
rect 24860 32438 24912 32444
rect 24768 32292 24820 32298
rect 24768 32234 24820 32240
rect 24676 32224 24728 32230
rect 24676 32166 24728 32172
rect 24780 31822 24808 32234
rect 24860 31884 24912 31890
rect 24860 31826 24912 31832
rect 24768 31816 24820 31822
rect 24872 31793 24900 31826
rect 24768 31758 24820 31764
rect 24858 31784 24914 31793
rect 25056 31754 25084 33918
rect 25148 33658 25176 35022
rect 25504 35022 25556 35028
rect 25410 34983 25466 34992
rect 25412 34944 25464 34950
rect 25412 34886 25464 34892
rect 25228 34060 25280 34066
rect 25228 34002 25280 34008
rect 25136 33652 25188 33658
rect 25136 33594 25188 33600
rect 25240 33318 25268 34002
rect 25424 33969 25452 34886
rect 25516 34610 25544 35022
rect 25700 35000 25728 35430
rect 25976 35154 26004 36042
rect 26252 36038 26280 37130
rect 27344 37120 27396 37126
rect 27344 37062 27396 37068
rect 27356 36786 27384 37062
rect 27448 36922 27476 37130
rect 27436 36916 27488 36922
rect 27436 36858 27488 36864
rect 27540 36786 27568 37266
rect 27632 37194 27660 37334
rect 27620 37188 27672 37194
rect 27620 37130 27672 37136
rect 27252 36780 27304 36786
rect 27252 36722 27304 36728
rect 27344 36780 27396 36786
rect 27344 36722 27396 36728
rect 27528 36780 27580 36786
rect 27528 36722 27580 36728
rect 26516 36100 26568 36106
rect 26516 36042 26568 36048
rect 26240 36032 26292 36038
rect 26240 35974 26292 35980
rect 26238 35864 26294 35873
rect 26238 35799 26240 35808
rect 26292 35799 26294 35808
rect 26240 35770 26292 35776
rect 26424 35692 26476 35698
rect 26424 35634 26476 35640
rect 26056 35624 26108 35630
rect 26330 35592 26386 35601
rect 26056 35566 26108 35572
rect 25964 35148 26016 35154
rect 25964 35090 26016 35096
rect 25780 35012 25832 35018
rect 25700 34972 25780 35000
rect 25504 34604 25556 34610
rect 25504 34546 25556 34552
rect 25596 34128 25648 34134
rect 25596 34070 25648 34076
rect 25410 33960 25466 33969
rect 25410 33895 25466 33904
rect 25424 33368 25452 33895
rect 25608 33522 25636 34070
rect 25700 33998 25728 34972
rect 25780 34954 25832 34960
rect 25688 33992 25740 33998
rect 25688 33934 25740 33940
rect 25688 33856 25740 33862
rect 25688 33798 25740 33804
rect 25596 33516 25648 33522
rect 25596 33458 25648 33464
rect 25700 33386 25728 33798
rect 25504 33380 25556 33386
rect 25424 33340 25504 33368
rect 25504 33322 25556 33328
rect 25688 33380 25740 33386
rect 25688 33322 25740 33328
rect 25228 33312 25280 33318
rect 25228 33254 25280 33260
rect 25320 33312 25372 33318
rect 25320 33254 25372 33260
rect 25780 33312 25832 33318
rect 25780 33254 25832 33260
rect 25332 32910 25360 33254
rect 25320 32904 25372 32910
rect 25320 32846 25372 32852
rect 25412 32428 25464 32434
rect 25412 32370 25464 32376
rect 25320 32224 25372 32230
rect 25320 32166 25372 32172
rect 25332 32026 25360 32166
rect 25320 32020 25372 32026
rect 25320 31962 25372 31968
rect 25320 31884 25372 31890
rect 25320 31826 25372 31832
rect 24858 31719 24914 31728
rect 24952 31748 25004 31754
rect 25056 31726 25268 31754
rect 24952 31690 25004 31696
rect 24860 31680 24912 31686
rect 24860 31622 24912 31628
rect 24676 31408 24728 31414
rect 24676 31350 24728 31356
rect 24584 31340 24636 31346
rect 24584 31282 24636 31288
rect 24400 30932 24452 30938
rect 24400 30874 24452 30880
rect 24492 30864 24544 30870
rect 24492 30806 24544 30812
rect 24308 30184 24360 30190
rect 24398 30152 24454 30161
rect 24360 30132 24398 30138
rect 24308 30126 24398 30132
rect 24320 30110 24398 30126
rect 24398 30087 24454 30096
rect 24400 29844 24452 29850
rect 24400 29786 24452 29792
rect 24308 29572 24360 29578
rect 24308 29514 24360 29520
rect 24216 29164 24268 29170
rect 24216 29106 24268 29112
rect 24320 28966 24348 29514
rect 24308 28960 24360 28966
rect 24308 28902 24360 28908
rect 24412 28762 24440 29786
rect 24504 29102 24532 30806
rect 24596 29850 24624 31282
rect 24688 30734 24716 31350
rect 24768 31272 24820 31278
rect 24766 31240 24768 31249
rect 24820 31240 24822 31249
rect 24766 31175 24822 31184
rect 24676 30728 24728 30734
rect 24676 30670 24728 30676
rect 24676 30388 24728 30394
rect 24676 30330 24728 30336
rect 24584 29844 24636 29850
rect 24584 29786 24636 29792
rect 24688 29730 24716 30330
rect 24768 30048 24820 30054
rect 24768 29990 24820 29996
rect 24596 29702 24716 29730
rect 24492 29096 24544 29102
rect 24490 29064 24492 29073
rect 24544 29064 24546 29073
rect 24490 28999 24546 29008
rect 24490 28928 24546 28937
rect 24490 28863 24546 28872
rect 24400 28756 24452 28762
rect 24400 28698 24452 28704
rect 24306 28520 24362 28529
rect 24306 28455 24362 28464
rect 24216 26784 24268 26790
rect 24216 26726 24268 26732
rect 24228 26518 24256 26726
rect 24216 26512 24268 26518
rect 24216 26454 24268 26460
rect 24228 22710 24256 26454
rect 24320 26382 24348 28455
rect 24412 27538 24440 28698
rect 24504 28694 24532 28863
rect 24492 28688 24544 28694
rect 24492 28630 24544 28636
rect 24492 28484 24544 28490
rect 24596 28472 24624 29702
rect 24676 29640 24728 29646
rect 24676 29582 24728 29588
rect 24544 28444 24624 28472
rect 24492 28426 24544 28432
rect 24400 27532 24452 27538
rect 24400 27474 24452 27480
rect 24400 26580 24452 26586
rect 24400 26522 24452 26528
rect 24308 26376 24360 26382
rect 24308 26318 24360 26324
rect 24216 22704 24268 22710
rect 24216 22646 24268 22652
rect 24216 22432 24268 22438
rect 24216 22374 24268 22380
rect 24124 22160 24176 22166
rect 24124 22102 24176 22108
rect 23848 19848 23900 19854
rect 23848 19790 23900 19796
rect 24032 19848 24084 19854
rect 24032 19790 24084 19796
rect 23940 19780 23992 19786
rect 23940 19722 23992 19728
rect 23768 19638 23888 19666
rect 23676 19502 23796 19530
rect 23572 19372 23624 19378
rect 23572 19314 23624 19320
rect 23664 19372 23716 19378
rect 23664 19314 23716 19320
rect 23478 19272 23534 19281
rect 23478 19207 23534 19216
rect 23492 18766 23520 19207
rect 23388 18760 23440 18766
rect 23388 18702 23440 18708
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23296 18624 23348 18630
rect 23296 18566 23348 18572
rect 23388 18624 23440 18630
rect 23388 18566 23440 18572
rect 23308 18358 23336 18566
rect 23296 18352 23348 18358
rect 23296 18294 23348 18300
rect 23204 17264 23256 17270
rect 23204 17206 23256 17212
rect 23400 17202 23428 18566
rect 23492 17542 23520 18702
rect 23570 17912 23626 17921
rect 23570 17847 23626 17856
rect 23584 17746 23612 17847
rect 23572 17740 23624 17746
rect 23572 17682 23624 17688
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 23572 17264 23624 17270
rect 23572 17206 23624 17212
rect 23388 17196 23440 17202
rect 23388 17138 23440 17144
rect 23584 17082 23612 17206
rect 23400 17054 23612 17082
rect 23676 17066 23704 19314
rect 23768 18970 23796 19502
rect 23860 19378 23888 19638
rect 23848 19372 23900 19378
rect 23848 19314 23900 19320
rect 23756 18964 23808 18970
rect 23756 18906 23808 18912
rect 23756 18692 23808 18698
rect 23756 18634 23808 18640
rect 23768 18290 23796 18634
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 23768 17338 23796 17614
rect 23756 17332 23808 17338
rect 23756 17274 23808 17280
rect 23768 17066 23796 17274
rect 23664 17060 23716 17066
rect 23296 14816 23348 14822
rect 23296 14758 23348 14764
rect 23308 14414 23336 14758
rect 23296 14408 23348 14414
rect 23296 14350 23348 14356
rect 23400 12889 23428 17054
rect 23664 17002 23716 17008
rect 23756 17060 23808 17066
rect 23756 17002 23808 17008
rect 23676 16794 23704 17002
rect 23768 16833 23796 17002
rect 23754 16824 23810 16833
rect 23664 16788 23716 16794
rect 23754 16759 23810 16768
rect 23664 16730 23716 16736
rect 23570 16688 23626 16697
rect 23492 16646 23570 16674
rect 23492 16590 23520 16646
rect 23626 16646 23704 16674
rect 23570 16623 23626 16632
rect 23480 16584 23532 16590
rect 23480 16526 23532 16532
rect 23572 16516 23624 16522
rect 23572 16458 23624 16464
rect 23584 14822 23612 16458
rect 23676 15450 23704 16646
rect 23756 16516 23808 16522
rect 23756 16458 23808 16464
rect 23768 16250 23796 16458
rect 23756 16244 23808 16250
rect 23756 16186 23808 16192
rect 23860 15706 23888 19314
rect 23952 18154 23980 19722
rect 24044 19446 24072 19790
rect 24032 19440 24084 19446
rect 24032 19382 24084 19388
rect 24136 18426 24164 22102
rect 24228 21350 24256 22374
rect 24216 21344 24268 21350
rect 24216 21286 24268 21292
rect 24216 21140 24268 21146
rect 24216 21082 24268 21088
rect 24124 18420 24176 18426
rect 24124 18362 24176 18368
rect 23940 18148 23992 18154
rect 23940 18090 23992 18096
rect 24136 17746 24164 18362
rect 24124 17740 24176 17746
rect 24124 17682 24176 17688
rect 24124 17536 24176 17542
rect 23938 17504 23994 17513
rect 23994 17462 24072 17490
rect 24124 17478 24176 17484
rect 23938 17439 23994 17448
rect 23940 16992 23992 16998
rect 23940 16934 23992 16940
rect 23952 15910 23980 16934
rect 23940 15904 23992 15910
rect 23940 15846 23992 15852
rect 23848 15700 23900 15706
rect 23848 15642 23900 15648
rect 24044 15502 24072 17462
rect 24136 17202 24164 17478
rect 24124 17196 24176 17202
rect 24124 17138 24176 17144
rect 24228 16810 24256 21082
rect 24320 19446 24348 26318
rect 24412 24410 24440 26522
rect 24504 25226 24532 28426
rect 24584 26784 24636 26790
rect 24582 26752 24584 26761
rect 24636 26752 24638 26761
rect 24582 26687 24638 26696
rect 24584 26580 24636 26586
rect 24584 26522 24636 26528
rect 24596 26246 24624 26522
rect 24584 26240 24636 26246
rect 24584 26182 24636 26188
rect 24492 25220 24544 25226
rect 24492 25162 24544 25168
rect 24688 24750 24716 29582
rect 24780 28994 24808 29990
rect 24872 29170 24900 31622
rect 24964 31482 24992 31690
rect 24952 31476 25004 31482
rect 24952 31418 25004 31424
rect 25240 31346 25268 31726
rect 25228 31340 25280 31346
rect 25148 31300 25228 31328
rect 24950 31104 25006 31113
rect 24950 31039 25006 31048
rect 24964 30870 24992 31039
rect 24952 30864 25004 30870
rect 24952 30806 25004 30812
rect 25044 30728 25096 30734
rect 25044 30670 25096 30676
rect 25056 30569 25084 30670
rect 25042 30560 25098 30569
rect 25042 30495 25098 30504
rect 24952 29232 25004 29238
rect 24952 29174 25004 29180
rect 24860 29164 24912 29170
rect 24860 29106 24912 29112
rect 24780 28966 24900 28994
rect 24872 28558 24900 28966
rect 24964 28762 24992 29174
rect 24952 28756 25004 28762
rect 24952 28698 25004 28704
rect 24860 28552 24912 28558
rect 24860 28494 24912 28500
rect 25044 28552 25096 28558
rect 25044 28494 25096 28500
rect 24768 28416 24820 28422
rect 24768 28358 24820 28364
rect 24780 27860 24808 28358
rect 24872 28014 24900 28494
rect 24952 28484 25004 28490
rect 24952 28426 25004 28432
rect 24964 28218 24992 28426
rect 24952 28212 25004 28218
rect 24952 28154 25004 28160
rect 24860 28008 24912 28014
rect 24860 27950 24912 27956
rect 24780 27832 24900 27860
rect 24766 27568 24822 27577
rect 24766 27503 24822 27512
rect 24780 27470 24808 27503
rect 24768 27464 24820 27470
rect 24768 27406 24820 27412
rect 24780 26926 24808 27406
rect 24768 26920 24820 26926
rect 24768 26862 24820 26868
rect 24768 26376 24820 26382
rect 24768 26318 24820 26324
rect 24780 26246 24808 26318
rect 24768 26240 24820 26246
rect 24768 26182 24820 26188
rect 24676 24744 24728 24750
rect 24676 24686 24728 24692
rect 24492 24608 24544 24614
rect 24492 24550 24544 24556
rect 24400 24404 24452 24410
rect 24400 24346 24452 24352
rect 24400 24132 24452 24138
rect 24400 24074 24452 24080
rect 24412 22094 24440 24074
rect 24504 23730 24532 24550
rect 24584 24268 24636 24274
rect 24584 24210 24636 24216
rect 24596 23730 24624 24210
rect 24676 24200 24728 24206
rect 24872 24188 24900 27832
rect 24964 26382 24992 28154
rect 25056 27946 25084 28494
rect 25148 27946 25176 31300
rect 25228 31282 25280 31288
rect 25228 29164 25280 29170
rect 25228 29106 25280 29112
rect 25240 29073 25268 29106
rect 25226 29064 25282 29073
rect 25226 28999 25282 29008
rect 25332 28937 25360 31826
rect 25424 31210 25452 32370
rect 25792 31346 25820 33254
rect 26068 33028 26096 35566
rect 26252 35550 26330 35578
rect 26252 35086 26280 35550
rect 26330 35527 26386 35536
rect 26436 35290 26464 35634
rect 26424 35284 26476 35290
rect 26424 35226 26476 35232
rect 26148 35080 26200 35086
rect 26148 35022 26200 35028
rect 26240 35080 26292 35086
rect 26240 35022 26292 35028
rect 26160 34921 26188 35022
rect 26252 34950 26280 35022
rect 26240 34944 26292 34950
rect 26146 34912 26202 34921
rect 26240 34886 26292 34892
rect 26332 34944 26384 34950
rect 26332 34886 26384 34892
rect 26146 34847 26202 34856
rect 26160 34746 26188 34847
rect 26148 34740 26200 34746
rect 26148 34682 26200 34688
rect 26344 33318 26372 34886
rect 26436 34746 26464 35226
rect 26424 34740 26476 34746
rect 26424 34682 26476 34688
rect 26528 34610 26556 36042
rect 27264 36038 27292 36722
rect 27540 36174 27568 36722
rect 27528 36168 27580 36174
rect 27528 36110 27580 36116
rect 27252 36032 27304 36038
rect 27252 35974 27304 35980
rect 27540 35766 27568 36110
rect 27528 35760 27580 35766
rect 27528 35702 27580 35708
rect 27528 35624 27580 35630
rect 27528 35566 27580 35572
rect 26896 35414 27200 35442
rect 26792 35284 26844 35290
rect 26792 35226 26844 35232
rect 26698 35184 26754 35193
rect 26698 35119 26754 35128
rect 26608 35012 26660 35018
rect 26608 34954 26660 34960
rect 26620 34785 26648 34954
rect 26606 34776 26662 34785
rect 26606 34711 26662 34720
rect 26712 34610 26740 35119
rect 26804 34746 26832 35226
rect 26792 34740 26844 34746
rect 26792 34682 26844 34688
rect 26424 34604 26476 34610
rect 26424 34546 26476 34552
rect 26516 34604 26568 34610
rect 26516 34546 26568 34552
rect 26700 34604 26752 34610
rect 26700 34546 26752 34552
rect 26332 33312 26384 33318
rect 26332 33254 26384 33260
rect 26436 33153 26464 34546
rect 26608 34400 26660 34406
rect 26608 34342 26660 34348
rect 26516 33856 26568 33862
rect 26516 33798 26568 33804
rect 26422 33144 26478 33153
rect 26528 33114 26556 33798
rect 26422 33079 26478 33088
rect 26516 33108 26568 33114
rect 26516 33050 26568 33056
rect 26068 33000 26464 33028
rect 25872 32972 25924 32978
rect 25872 32914 25924 32920
rect 25884 32026 25912 32914
rect 26056 32904 26108 32910
rect 26056 32846 26108 32852
rect 25872 32020 25924 32026
rect 25872 31962 25924 31968
rect 25884 31890 25912 31962
rect 25964 31952 26016 31958
rect 25964 31894 26016 31900
rect 25872 31884 25924 31890
rect 25872 31826 25924 31832
rect 25780 31340 25832 31346
rect 25516 31300 25780 31328
rect 25412 31204 25464 31210
rect 25412 31146 25464 31152
rect 25516 31090 25544 31300
rect 25780 31282 25832 31288
rect 25872 31340 25924 31346
rect 25976 31328 26004 31894
rect 25924 31300 26004 31328
rect 25872 31282 25924 31288
rect 25424 31062 25544 31090
rect 25688 31136 25740 31142
rect 25688 31078 25740 31084
rect 25780 31136 25832 31142
rect 25780 31078 25832 31084
rect 25424 29345 25452 31062
rect 25700 30598 25728 31078
rect 25792 30666 25820 31078
rect 25780 30660 25832 30666
rect 25780 30602 25832 30608
rect 25596 30592 25648 30598
rect 25596 30534 25648 30540
rect 25688 30592 25740 30598
rect 25688 30534 25740 30540
rect 25410 29336 25466 29345
rect 25410 29271 25466 29280
rect 25318 28928 25374 28937
rect 25318 28863 25374 28872
rect 25332 28762 25360 28863
rect 25320 28756 25372 28762
rect 25320 28698 25372 28704
rect 25320 28552 25372 28558
rect 25320 28494 25372 28500
rect 25228 28416 25280 28422
rect 25228 28358 25280 28364
rect 25044 27940 25096 27946
rect 25044 27882 25096 27888
rect 25136 27940 25188 27946
rect 25136 27882 25188 27888
rect 25240 27690 25268 28358
rect 25332 28150 25360 28494
rect 25320 28144 25372 28150
rect 25320 28086 25372 28092
rect 25318 27704 25374 27713
rect 25240 27662 25318 27690
rect 25318 27639 25374 27648
rect 25044 27532 25096 27538
rect 25044 27474 25096 27480
rect 25056 26994 25084 27474
rect 25228 27464 25280 27470
rect 25228 27406 25280 27412
rect 25044 26988 25096 26994
rect 25044 26930 25096 26936
rect 25136 26988 25188 26994
rect 25136 26930 25188 26936
rect 25148 26874 25176 26930
rect 25056 26846 25176 26874
rect 25056 26586 25084 26846
rect 25136 26784 25188 26790
rect 25136 26726 25188 26732
rect 25044 26580 25096 26586
rect 25044 26522 25096 26528
rect 25056 26489 25084 26522
rect 25042 26480 25098 26489
rect 25042 26415 25098 26424
rect 25148 26382 25176 26726
rect 25240 26382 25268 27406
rect 25332 26586 25360 27639
rect 25320 26580 25372 26586
rect 25320 26522 25372 26528
rect 24952 26376 25004 26382
rect 24952 26318 25004 26324
rect 25136 26376 25188 26382
rect 25136 26318 25188 26324
rect 25228 26376 25280 26382
rect 25228 26318 25280 26324
rect 24964 25770 24992 26318
rect 24952 25764 25004 25770
rect 24952 25706 25004 25712
rect 25136 25288 25188 25294
rect 25136 25230 25188 25236
rect 24952 25152 25004 25158
rect 24952 25094 25004 25100
rect 24964 24410 24992 25094
rect 25148 24993 25176 25230
rect 25240 25140 25268 26318
rect 25424 26024 25452 29271
rect 25504 29164 25556 29170
rect 25504 29106 25556 29112
rect 25516 28665 25544 29106
rect 25502 28656 25558 28665
rect 25502 28591 25558 28600
rect 25504 28552 25556 28558
rect 25504 28494 25556 28500
rect 25332 25996 25452 26024
rect 25332 25294 25360 25996
rect 25412 25900 25464 25906
rect 25412 25842 25464 25848
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25240 25112 25360 25140
rect 25134 24984 25190 24993
rect 25134 24919 25190 24928
rect 24952 24404 25004 24410
rect 24952 24346 25004 24352
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 24952 24200 25004 24206
rect 24728 24160 24808 24188
rect 24872 24160 24952 24188
rect 24676 24142 24728 24148
rect 24674 23760 24730 23769
rect 24492 23724 24544 23730
rect 24492 23666 24544 23672
rect 24584 23724 24636 23730
rect 24674 23695 24730 23704
rect 24584 23666 24636 23672
rect 24504 22710 24532 23666
rect 24582 23624 24638 23633
rect 24582 23559 24638 23568
rect 24492 22704 24544 22710
rect 24492 22646 24544 22652
rect 24596 22624 24624 23559
rect 24688 23254 24716 23695
rect 24676 23248 24728 23254
rect 24676 23190 24728 23196
rect 24688 22778 24716 23190
rect 24676 22772 24728 22778
rect 24676 22714 24728 22720
rect 24596 22596 24716 22624
rect 24492 22568 24544 22574
rect 24492 22510 24544 22516
rect 24504 22386 24532 22510
rect 24504 22358 24624 22386
rect 24412 22066 24532 22094
rect 24400 22024 24452 22030
rect 24398 21992 24400 22001
rect 24452 21992 24454 22001
rect 24398 21927 24454 21936
rect 24400 21888 24452 21894
rect 24400 21830 24452 21836
rect 24412 21690 24440 21830
rect 24400 21684 24452 21690
rect 24400 21626 24452 21632
rect 24400 21480 24452 21486
rect 24398 21448 24400 21457
rect 24452 21448 24454 21457
rect 24398 21383 24454 21392
rect 24400 21344 24452 21350
rect 24400 21286 24452 21292
rect 24412 21146 24440 21286
rect 24400 21140 24452 21146
rect 24400 21082 24452 21088
rect 24400 20460 24452 20466
rect 24400 20402 24452 20408
rect 24308 19440 24360 19446
rect 24308 19382 24360 19388
rect 24412 19378 24440 20402
rect 24400 19372 24452 19378
rect 24400 19314 24452 19320
rect 24400 18284 24452 18290
rect 24400 18226 24452 18232
rect 24136 16782 24256 16810
rect 24032 15496 24084 15502
rect 23952 15456 24032 15484
rect 23676 15422 23888 15450
rect 23664 15360 23716 15366
rect 23664 15302 23716 15308
rect 23676 15162 23704 15302
rect 23664 15156 23716 15162
rect 23664 15098 23716 15104
rect 23664 15020 23716 15026
rect 23664 14962 23716 14968
rect 23676 14822 23704 14962
rect 23572 14816 23624 14822
rect 23572 14758 23624 14764
rect 23664 14816 23716 14822
rect 23664 14758 23716 14764
rect 23756 14816 23808 14822
rect 23756 14758 23808 14764
rect 23584 14550 23612 14758
rect 23676 14618 23704 14758
rect 23664 14612 23716 14618
rect 23664 14554 23716 14560
rect 23572 14544 23624 14550
rect 23572 14486 23624 14492
rect 23768 14482 23796 14758
rect 23756 14476 23808 14482
rect 23756 14418 23808 14424
rect 23386 12880 23442 12889
rect 23386 12815 23442 12824
rect 23480 12776 23532 12782
rect 23860 12730 23888 15422
rect 23952 15026 23980 15456
rect 24032 15438 24084 15444
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 24136 14822 24164 16782
rect 24216 15904 24268 15910
rect 24216 15846 24268 15852
rect 24308 15904 24360 15910
rect 24308 15846 24360 15852
rect 24228 15638 24256 15846
rect 24216 15632 24268 15638
rect 24216 15574 24268 15580
rect 24320 15026 24348 15846
rect 24412 15502 24440 18226
rect 24504 17882 24532 22066
rect 24596 19514 24624 22358
rect 24688 20058 24716 22596
rect 24780 20346 24808 24160
rect 24952 24142 25004 24148
rect 24860 23724 24912 23730
rect 24860 23666 24912 23672
rect 24872 22982 24900 23666
rect 24860 22976 24912 22982
rect 24860 22918 24912 22924
rect 24858 22672 24914 22681
rect 24858 22607 24914 22616
rect 24872 22166 24900 22607
rect 24860 22160 24912 22166
rect 24860 22102 24912 22108
rect 24964 21468 24992 24142
rect 25042 24032 25098 24041
rect 25042 23967 25098 23976
rect 25056 23730 25084 23967
rect 25044 23724 25096 23730
rect 25044 23666 25096 23672
rect 25042 23216 25098 23225
rect 25042 23151 25044 23160
rect 25096 23151 25098 23160
rect 25044 23122 25096 23128
rect 25044 22704 25096 22710
rect 25044 22646 25096 22652
rect 25056 21865 25084 22646
rect 25042 21856 25098 21865
rect 25042 21791 25098 21800
rect 25148 21536 25176 24346
rect 25332 24138 25360 25112
rect 25424 24410 25452 25842
rect 25516 25498 25544 28494
rect 25608 27538 25636 30534
rect 25596 27532 25648 27538
rect 25596 27474 25648 27480
rect 25594 26344 25650 26353
rect 25594 26279 25596 26288
rect 25648 26279 25650 26288
rect 25596 26250 25648 26256
rect 25504 25492 25556 25498
rect 25504 25434 25556 25440
rect 25504 24948 25556 24954
rect 25504 24890 25556 24896
rect 25412 24404 25464 24410
rect 25412 24346 25464 24352
rect 25516 24138 25544 24890
rect 25228 24132 25280 24138
rect 25228 24074 25280 24080
rect 25320 24132 25372 24138
rect 25320 24074 25372 24080
rect 25504 24132 25556 24138
rect 25504 24074 25556 24080
rect 25240 23866 25268 24074
rect 25608 24018 25636 26250
rect 25700 24138 25728 30534
rect 25884 30433 25912 31282
rect 25964 31204 26016 31210
rect 25964 31146 26016 31152
rect 25976 30666 26004 31146
rect 25964 30660 26016 30666
rect 25964 30602 26016 30608
rect 25870 30424 25926 30433
rect 25870 30359 25926 30368
rect 25976 30258 26004 30602
rect 25964 30252 26016 30258
rect 25964 30194 26016 30200
rect 26068 29850 26096 32846
rect 26240 32768 26292 32774
rect 26240 32710 26292 32716
rect 26332 32768 26384 32774
rect 26332 32710 26384 32716
rect 26146 32328 26202 32337
rect 26146 32263 26202 32272
rect 26056 29844 26108 29850
rect 26056 29786 26108 29792
rect 26160 29730 26188 32263
rect 25884 29702 26188 29730
rect 25884 29481 25912 29702
rect 25870 29472 25926 29481
rect 25870 29407 25926 29416
rect 25780 29028 25832 29034
rect 25780 28970 25832 28976
rect 25688 24132 25740 24138
rect 25688 24074 25740 24080
rect 25332 23990 25636 24018
rect 25228 23860 25280 23866
rect 25228 23802 25280 23808
rect 25332 23746 25360 23990
rect 25240 23718 25360 23746
rect 25412 23724 25464 23730
rect 25240 21962 25268 23718
rect 25412 23666 25464 23672
rect 25320 23656 25372 23662
rect 25320 23598 25372 23604
rect 25332 22166 25360 23598
rect 25424 22545 25452 23666
rect 25792 23526 25820 28970
rect 25884 28422 25912 29407
rect 26252 29016 26280 32710
rect 26344 32298 26372 32710
rect 26332 32292 26384 32298
rect 26332 32234 26384 32240
rect 26332 31952 26384 31958
rect 26330 31920 26332 31929
rect 26384 31920 26386 31929
rect 26330 31855 26386 31864
rect 26436 31822 26464 33000
rect 26620 32858 26648 34342
rect 26804 33862 26832 34682
rect 26896 34610 26924 35414
rect 27172 35290 27200 35414
rect 27068 35284 27120 35290
rect 27068 35226 27120 35232
rect 27160 35284 27212 35290
rect 27160 35226 27212 35232
rect 26976 35080 27028 35086
rect 26976 35022 27028 35028
rect 26884 34604 26936 34610
rect 26884 34546 26936 34552
rect 26700 33856 26752 33862
rect 26700 33798 26752 33804
rect 26792 33856 26844 33862
rect 26792 33798 26844 33804
rect 26712 33658 26740 33798
rect 26700 33652 26752 33658
rect 26700 33594 26752 33600
rect 26712 33289 26740 33594
rect 26988 33454 27016 35022
rect 27080 33833 27108 35226
rect 27344 35216 27396 35222
rect 27344 35158 27396 35164
rect 27252 34944 27304 34950
rect 27252 34886 27304 34892
rect 27160 34400 27212 34406
rect 27160 34342 27212 34348
rect 27172 33998 27200 34342
rect 27160 33992 27212 33998
rect 27160 33934 27212 33940
rect 27066 33824 27122 33833
rect 27066 33759 27122 33768
rect 26976 33448 27028 33454
rect 26976 33390 27028 33396
rect 26792 33312 26844 33318
rect 26698 33280 26754 33289
rect 26792 33254 26844 33260
rect 26698 33215 26754 33224
rect 26528 32842 26648 32858
rect 26700 32904 26752 32910
rect 26700 32846 26752 32852
rect 26528 32836 26660 32842
rect 26528 32830 26608 32836
rect 26424 31816 26476 31822
rect 26424 31758 26476 31764
rect 26332 31748 26384 31754
rect 26332 31690 26384 31696
rect 26344 31210 26372 31690
rect 26424 31680 26476 31686
rect 26424 31622 26476 31628
rect 26436 31210 26464 31622
rect 26528 31346 26556 32830
rect 26608 32778 26660 32784
rect 26712 32434 26740 32846
rect 26700 32428 26752 32434
rect 26700 32370 26752 32376
rect 26608 32360 26660 32366
rect 26608 32302 26660 32308
rect 26620 32026 26648 32302
rect 26608 32020 26660 32026
rect 26608 31962 26660 31968
rect 26712 31906 26740 32370
rect 26620 31878 26740 31906
rect 26516 31340 26568 31346
rect 26516 31282 26568 31288
rect 26332 31204 26384 31210
rect 26332 31146 26384 31152
rect 26424 31204 26476 31210
rect 26424 31146 26476 31152
rect 26424 30932 26476 30938
rect 26424 30874 26476 30880
rect 26332 30660 26384 30666
rect 26332 30602 26384 30608
rect 26344 30394 26372 30602
rect 26332 30388 26384 30394
rect 26332 30330 26384 30336
rect 26332 29776 26384 29782
rect 26332 29718 26384 29724
rect 26068 28988 26280 29016
rect 25964 28960 26016 28966
rect 25964 28902 26016 28908
rect 25976 28762 26004 28902
rect 25964 28756 26016 28762
rect 25964 28698 26016 28704
rect 25962 28656 26018 28665
rect 25962 28591 26018 28600
rect 25872 28416 25924 28422
rect 25872 28358 25924 28364
rect 25872 28212 25924 28218
rect 25872 28154 25924 28160
rect 25884 27538 25912 28154
rect 25976 27878 26004 28591
rect 25964 27872 26016 27878
rect 25964 27814 26016 27820
rect 25964 27668 26016 27674
rect 25964 27610 26016 27616
rect 25872 27532 25924 27538
rect 25872 27474 25924 27480
rect 25976 26246 26004 27610
rect 26068 27470 26096 28988
rect 26240 28484 26292 28490
rect 26160 28444 26240 28472
rect 26160 28393 26188 28444
rect 26240 28426 26292 28432
rect 26146 28384 26202 28393
rect 26146 28319 26202 28328
rect 26148 27872 26200 27878
rect 26148 27814 26200 27820
rect 26056 27464 26108 27470
rect 26056 27406 26108 27412
rect 26056 26784 26108 26790
rect 26056 26726 26108 26732
rect 25964 26240 26016 26246
rect 25964 26182 26016 26188
rect 26068 25906 26096 26726
rect 26160 26450 26188 27814
rect 26344 27690 26372 29718
rect 26436 29646 26464 30874
rect 26620 30802 26648 31878
rect 26700 31816 26752 31822
rect 26700 31758 26752 31764
rect 26712 30938 26740 31758
rect 26804 31142 26832 33254
rect 27172 32910 27200 33934
rect 27264 32978 27292 34886
rect 27356 34610 27384 35158
rect 27540 35086 27568 35566
rect 27528 35080 27580 35086
rect 27528 35022 27580 35028
rect 27632 34898 27660 37130
rect 27724 36854 27752 37878
rect 27816 37670 27844 38150
rect 27804 37664 27856 37670
rect 27804 37606 27856 37612
rect 27712 36848 27764 36854
rect 27712 36790 27764 36796
rect 27816 36718 27844 37606
rect 27908 37466 27936 38218
rect 27896 37460 27948 37466
rect 27896 37402 27948 37408
rect 27804 36712 27856 36718
rect 27804 36654 27856 36660
rect 27632 34870 27752 34898
rect 27618 34776 27674 34785
rect 27618 34711 27620 34720
rect 27672 34711 27674 34720
rect 27620 34682 27672 34688
rect 27344 34604 27396 34610
rect 27344 34546 27396 34552
rect 27620 34196 27672 34202
rect 27620 34138 27672 34144
rect 27436 34128 27488 34134
rect 27436 34070 27488 34076
rect 27448 33930 27476 34070
rect 27528 33992 27580 33998
rect 27528 33934 27580 33940
rect 27436 33924 27488 33930
rect 27436 33866 27488 33872
rect 27344 33856 27396 33862
rect 27344 33798 27396 33804
rect 27356 33522 27384 33798
rect 27344 33516 27396 33522
rect 27344 33458 27396 33464
rect 27448 33318 27476 33866
rect 27540 33658 27568 33934
rect 27528 33652 27580 33658
rect 27528 33594 27580 33600
rect 27632 33318 27660 34138
rect 27724 33862 27752 34870
rect 27712 33856 27764 33862
rect 27712 33798 27764 33804
rect 27436 33312 27488 33318
rect 27436 33254 27488 33260
rect 27620 33312 27672 33318
rect 27620 33254 27672 33260
rect 27252 32972 27304 32978
rect 27252 32914 27304 32920
rect 27160 32904 27212 32910
rect 27160 32846 27212 32852
rect 27528 32904 27580 32910
rect 27528 32846 27580 32852
rect 27436 32836 27488 32842
rect 27436 32778 27488 32784
rect 26884 32768 26936 32774
rect 26884 32710 26936 32716
rect 26896 31958 26924 32710
rect 27068 32564 27120 32570
rect 27068 32506 27120 32512
rect 26974 32328 27030 32337
rect 26974 32263 27030 32272
rect 26988 31958 27016 32263
rect 27080 32230 27108 32506
rect 27068 32224 27120 32230
rect 27068 32166 27120 32172
rect 27160 32224 27212 32230
rect 27160 32166 27212 32172
rect 27344 32224 27396 32230
rect 27448 32212 27476 32778
rect 27540 32434 27568 32846
rect 27528 32428 27580 32434
rect 27528 32370 27580 32376
rect 27620 32428 27672 32434
rect 27620 32370 27672 32376
rect 27528 32224 27580 32230
rect 27448 32184 27528 32212
rect 27344 32166 27396 32172
rect 27528 32166 27580 32172
rect 26884 31952 26936 31958
rect 26884 31894 26936 31900
rect 26976 31952 27028 31958
rect 26976 31894 27028 31900
rect 27172 31754 27200 32166
rect 27356 32026 27384 32166
rect 27252 32020 27304 32026
rect 27252 31962 27304 31968
rect 27344 32020 27396 32026
rect 27344 31962 27396 31968
rect 27264 31906 27292 31962
rect 27632 31906 27660 32370
rect 27264 31878 27660 31906
rect 27252 31816 27304 31822
rect 27252 31758 27304 31764
rect 27528 31816 27580 31822
rect 27528 31758 27580 31764
rect 27160 31748 27212 31754
rect 27160 31690 27212 31696
rect 26976 31680 27028 31686
rect 26976 31622 27028 31628
rect 26792 31136 26844 31142
rect 26792 31078 26844 31084
rect 26700 30932 26752 30938
rect 26700 30874 26752 30880
rect 26804 30818 26832 31078
rect 26608 30796 26660 30802
rect 26608 30738 26660 30744
rect 26712 30790 26832 30818
rect 26516 30116 26568 30122
rect 26516 30058 26568 30064
rect 26528 29850 26556 30058
rect 26516 29844 26568 29850
rect 26516 29786 26568 29792
rect 26516 29708 26568 29714
rect 26516 29650 26568 29656
rect 26424 29640 26476 29646
rect 26424 29582 26476 29588
rect 26436 28966 26464 29582
rect 26528 29306 26556 29650
rect 26516 29300 26568 29306
rect 26516 29242 26568 29248
rect 26620 28994 26648 30738
rect 26528 28966 26648 28994
rect 26712 28994 26740 30790
rect 26792 30728 26844 30734
rect 26792 30670 26844 30676
rect 26804 29646 26832 30670
rect 26792 29640 26844 29646
rect 26792 29582 26844 29588
rect 26988 29170 27016 31622
rect 27264 31482 27292 31758
rect 27252 31476 27304 31482
rect 27252 31418 27304 31424
rect 27344 31476 27396 31482
rect 27344 31418 27396 31424
rect 27356 31249 27384 31418
rect 27342 31240 27398 31249
rect 27540 31210 27568 31758
rect 27342 31175 27398 31184
rect 27528 31204 27580 31210
rect 27528 31146 27580 31152
rect 27252 31136 27304 31142
rect 27252 31078 27304 31084
rect 27068 30728 27120 30734
rect 27068 30670 27120 30676
rect 26976 29164 27028 29170
rect 26976 29106 27028 29112
rect 26712 28966 26924 28994
rect 26424 28960 26476 28966
rect 26424 28902 26476 28908
rect 26424 28552 26476 28558
rect 26424 28494 26476 28500
rect 26436 28218 26464 28494
rect 26424 28212 26476 28218
rect 26424 28154 26476 28160
rect 26424 28076 26476 28082
rect 26424 28018 26476 28024
rect 26252 27662 26372 27690
rect 26436 27674 26464 28018
rect 26424 27668 26476 27674
rect 26148 26444 26200 26450
rect 26148 26386 26200 26392
rect 26252 25906 26280 27662
rect 26424 27610 26476 27616
rect 26332 27600 26384 27606
rect 26528 27554 26556 28966
rect 26608 28960 26660 28966
rect 26608 28902 26660 28908
rect 26792 28756 26844 28762
rect 26792 28698 26844 28704
rect 26608 28552 26660 28558
rect 26608 28494 26660 28500
rect 26700 28552 26752 28558
rect 26804 28506 26832 28698
rect 26896 28626 26924 28966
rect 26884 28620 26936 28626
rect 26936 28580 27016 28608
rect 26884 28562 26936 28568
rect 26752 28500 26832 28506
rect 26700 28494 26832 28500
rect 26620 28370 26648 28494
rect 26712 28478 26832 28494
rect 26698 28384 26754 28393
rect 26620 28342 26698 28370
rect 26698 28319 26754 28328
rect 26700 28008 26752 28014
rect 26606 27976 26662 27985
rect 26700 27950 26752 27956
rect 26606 27911 26662 27920
rect 26620 27606 26648 27911
rect 26332 27542 26384 27548
rect 26344 27402 26372 27542
rect 26436 27526 26556 27554
rect 26608 27600 26660 27606
rect 26608 27542 26660 27548
rect 26332 27396 26384 27402
rect 26332 27338 26384 27344
rect 26436 26994 26464 27526
rect 26516 27464 26568 27470
rect 26516 27406 26568 27412
rect 26424 26988 26476 26994
rect 26424 26930 26476 26936
rect 26424 26580 26476 26586
rect 26424 26522 26476 26528
rect 26332 26376 26384 26382
rect 26332 26318 26384 26324
rect 25964 25900 26016 25906
rect 25964 25842 26016 25848
rect 26056 25900 26108 25906
rect 26056 25842 26108 25848
rect 26240 25900 26292 25906
rect 26240 25842 26292 25848
rect 25872 25832 25924 25838
rect 25872 25774 25924 25780
rect 25780 23520 25832 23526
rect 25780 23462 25832 23468
rect 25884 23338 25912 25774
rect 25976 25752 26004 25842
rect 26056 25764 26108 25770
rect 25976 25724 26056 25752
rect 25976 24614 26004 25724
rect 26056 25706 26108 25712
rect 25964 24608 26016 24614
rect 25964 24550 26016 24556
rect 26238 24304 26294 24313
rect 25964 24268 26016 24274
rect 26238 24239 26294 24248
rect 25964 24210 26016 24216
rect 25976 24041 26004 24210
rect 26056 24132 26108 24138
rect 26056 24074 26108 24080
rect 25962 24032 26018 24041
rect 25962 23967 26018 23976
rect 25964 23656 26016 23662
rect 26068 23633 26096 24074
rect 26148 24064 26200 24070
rect 26148 24006 26200 24012
rect 25964 23598 26016 23604
rect 26054 23624 26110 23633
rect 25700 23310 25912 23338
rect 25504 23044 25556 23050
rect 25504 22986 25556 22992
rect 25410 22536 25466 22545
rect 25410 22471 25466 22480
rect 25516 22166 25544 22986
rect 25596 22568 25648 22574
rect 25596 22510 25648 22516
rect 25320 22160 25372 22166
rect 25320 22102 25372 22108
rect 25504 22160 25556 22166
rect 25504 22102 25556 22108
rect 25608 22012 25636 22510
rect 25516 21984 25636 22012
rect 25228 21956 25280 21962
rect 25228 21898 25280 21904
rect 25412 21548 25464 21554
rect 25148 21508 25412 21536
rect 25412 21490 25464 21496
rect 24964 21440 25360 21468
rect 24860 21412 24912 21418
rect 24860 21354 24912 21360
rect 24872 21010 24900 21354
rect 25044 21344 25096 21350
rect 25044 21286 25096 21292
rect 24950 21040 25006 21049
rect 24860 21004 24912 21010
rect 24950 20975 25006 20984
rect 24860 20946 24912 20952
rect 24964 20806 24992 20975
rect 24952 20800 25004 20806
rect 24952 20742 25004 20748
rect 24780 20318 24900 20346
rect 24766 20224 24822 20233
rect 24766 20159 24822 20168
rect 24676 20052 24728 20058
rect 24676 19994 24728 20000
rect 24780 19922 24808 20159
rect 24768 19916 24820 19922
rect 24768 19858 24820 19864
rect 24584 19508 24636 19514
rect 24584 19450 24636 19456
rect 24596 19417 24624 19450
rect 24676 19440 24728 19446
rect 24582 19408 24638 19417
rect 24676 19382 24728 19388
rect 24582 19343 24638 19352
rect 24584 19236 24636 19242
rect 24584 19178 24636 19184
rect 24596 18970 24624 19178
rect 24584 18964 24636 18970
rect 24584 18906 24636 18912
rect 24596 17882 24624 18906
rect 24492 17876 24544 17882
rect 24492 17818 24544 17824
rect 24584 17876 24636 17882
rect 24584 17818 24636 17824
rect 24584 17332 24636 17338
rect 24584 17274 24636 17280
rect 24596 17202 24624 17274
rect 24492 17196 24544 17202
rect 24492 17138 24544 17144
rect 24584 17196 24636 17202
rect 24584 17138 24636 17144
rect 24504 16794 24532 17138
rect 24492 16788 24544 16794
rect 24492 16730 24544 16736
rect 24688 16182 24716 19382
rect 24872 19310 24900 20318
rect 24860 19304 24912 19310
rect 24780 19252 24860 19258
rect 24780 19246 24912 19252
rect 24780 19230 24900 19246
rect 24780 18766 24808 19230
rect 24952 19168 25004 19174
rect 24952 19110 25004 19116
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 24766 18456 24822 18465
rect 24964 18442 24992 19110
rect 24822 18414 24992 18442
rect 24766 18391 24822 18400
rect 24860 18148 24912 18154
rect 24860 18090 24912 18096
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 24676 16176 24728 16182
rect 24676 16118 24728 16124
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24582 15192 24638 15201
rect 24582 15127 24638 15136
rect 24308 15020 24360 15026
rect 24308 14962 24360 14968
rect 24400 15020 24452 15026
rect 24400 14962 24452 14968
rect 24124 14816 24176 14822
rect 24124 14758 24176 14764
rect 24308 14816 24360 14822
rect 24308 14758 24360 14764
rect 24320 14550 24348 14758
rect 24412 14550 24440 14962
rect 24308 14544 24360 14550
rect 24308 14486 24360 14492
rect 24400 14544 24452 14550
rect 24400 14486 24452 14492
rect 24124 14476 24176 14482
rect 24124 14418 24176 14424
rect 23940 12912 23992 12918
rect 23940 12854 23992 12860
rect 24032 12912 24084 12918
rect 24032 12854 24084 12860
rect 23480 12718 23532 12724
rect 23296 12640 23348 12646
rect 23296 12582 23348 12588
rect 23308 12238 23336 12582
rect 23492 12442 23520 12718
rect 23768 12702 23888 12730
rect 23480 12436 23532 12442
rect 23480 12378 23532 12384
rect 23478 12336 23534 12345
rect 23478 12271 23480 12280
rect 23532 12271 23534 12280
rect 23480 12242 23532 12248
rect 23296 12232 23348 12238
rect 23296 12174 23348 12180
rect 23112 12096 23164 12102
rect 23112 12038 23164 12044
rect 22742 11792 22798 11801
rect 22742 11727 22798 11736
rect 23492 11694 23520 12242
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 23676 11898 23704 12174
rect 23664 11892 23716 11898
rect 23664 11834 23716 11840
rect 23768 11762 23796 12702
rect 23848 12640 23900 12646
rect 23848 12582 23900 12588
rect 23860 12306 23888 12582
rect 23952 12442 23980 12854
rect 23940 12436 23992 12442
rect 23940 12378 23992 12384
rect 24044 12306 24072 12854
rect 24136 12646 24164 14418
rect 24492 14340 24544 14346
rect 24492 14282 24544 14288
rect 24306 13696 24362 13705
rect 24306 13631 24362 13640
rect 24320 12986 24348 13631
rect 24308 12980 24360 12986
rect 24308 12922 24360 12928
rect 24124 12640 24176 12646
rect 24124 12582 24176 12588
rect 24398 12472 24454 12481
rect 24398 12407 24454 12416
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 24032 12300 24084 12306
rect 24032 12242 24084 12248
rect 23756 11756 23808 11762
rect 23756 11698 23808 11704
rect 23480 11688 23532 11694
rect 23480 11630 23532 11636
rect 24044 11626 24072 12242
rect 24412 12238 24440 12407
rect 24400 12232 24452 12238
rect 24400 12174 24452 12180
rect 24504 12084 24532 14282
rect 24596 12918 24624 15127
rect 24676 14884 24728 14890
rect 24676 14826 24728 14832
rect 24688 14414 24716 14826
rect 24676 14408 24728 14414
rect 24676 14350 24728 14356
rect 24780 14346 24808 17818
rect 24872 16454 24900 18090
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 24964 14498 24992 17614
rect 25056 16590 25084 21286
rect 25228 20596 25280 20602
rect 25228 20538 25280 20544
rect 25136 19848 25188 19854
rect 25136 19790 25188 19796
rect 25148 19514 25176 19790
rect 25136 19508 25188 19514
rect 25136 19450 25188 19456
rect 25240 19446 25268 20538
rect 25228 19440 25280 19446
rect 25228 19382 25280 19388
rect 25136 19372 25188 19378
rect 25136 19314 25188 19320
rect 25148 19174 25176 19314
rect 25136 19168 25188 19174
rect 25136 19110 25188 19116
rect 25134 19000 25190 19009
rect 25134 18935 25190 18944
rect 25148 18766 25176 18935
rect 25136 18760 25188 18766
rect 25136 18702 25188 18708
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 25056 15978 25084 16050
rect 25044 15972 25096 15978
rect 25044 15914 25096 15920
rect 24872 14470 24992 14498
rect 24768 14340 24820 14346
rect 24768 14282 24820 14288
rect 24584 12912 24636 12918
rect 24584 12854 24636 12860
rect 24872 12850 24900 14470
rect 24952 14408 25004 14414
rect 24952 14350 25004 14356
rect 24964 14074 24992 14350
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 25056 14006 25084 15914
rect 25148 14958 25176 18702
rect 25240 17746 25268 19382
rect 25332 18698 25360 21440
rect 25424 20924 25452 21490
rect 25516 21486 25544 21984
rect 25596 21888 25648 21894
rect 25596 21830 25648 21836
rect 25504 21480 25556 21486
rect 25504 21422 25556 21428
rect 25424 20896 25544 20924
rect 25412 19712 25464 19718
rect 25412 19654 25464 19660
rect 25424 19310 25452 19654
rect 25412 19304 25464 19310
rect 25412 19246 25464 19252
rect 25320 18692 25372 18698
rect 25320 18634 25372 18640
rect 25228 17740 25280 17746
rect 25280 17700 25360 17728
rect 25228 17682 25280 17688
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 25240 16250 25268 16526
rect 25228 16244 25280 16250
rect 25228 16186 25280 16192
rect 25332 16046 25360 17700
rect 25424 16046 25452 19246
rect 25516 18850 25544 20896
rect 25608 19854 25636 21830
rect 25596 19848 25648 19854
rect 25596 19790 25648 19796
rect 25594 19544 25650 19553
rect 25594 19479 25596 19488
rect 25648 19479 25650 19488
rect 25596 19450 25648 19456
rect 25700 19446 25728 23310
rect 25976 22094 26004 23598
rect 26054 23559 26110 23568
rect 26056 23112 26108 23118
rect 26056 23054 26108 23060
rect 26068 22681 26096 23054
rect 26054 22672 26110 22681
rect 26054 22607 26110 22616
rect 26160 22250 26188 24006
rect 26252 23798 26280 24239
rect 26240 23792 26292 23798
rect 26240 23734 26292 23740
rect 26344 23594 26372 26318
rect 26332 23588 26384 23594
rect 26332 23530 26384 23536
rect 26436 23322 26464 26522
rect 26528 24818 26556 27406
rect 26608 27056 26660 27062
rect 26608 26998 26660 27004
rect 26620 26058 26648 26998
rect 26712 26382 26740 27950
rect 26700 26376 26752 26382
rect 26700 26318 26752 26324
rect 26620 26030 26740 26058
rect 26608 25968 26660 25974
rect 26608 25910 26660 25916
rect 26516 24812 26568 24818
rect 26516 24754 26568 24760
rect 26424 23316 26476 23322
rect 26424 23258 26476 23264
rect 26528 23186 26556 24754
rect 26620 23866 26648 25910
rect 26712 24070 26740 26030
rect 26700 24064 26752 24070
rect 26700 24006 26752 24012
rect 26608 23860 26660 23866
rect 26608 23802 26660 23808
rect 26700 23792 26752 23798
rect 26700 23734 26752 23740
rect 26608 23724 26660 23730
rect 26608 23666 26660 23672
rect 26516 23180 26568 23186
rect 26516 23122 26568 23128
rect 26620 22930 26648 23666
rect 26712 23497 26740 23734
rect 26698 23488 26754 23497
rect 26698 23423 26754 23432
rect 26436 22902 26648 22930
rect 26240 22568 26292 22574
rect 26240 22510 26292 22516
rect 26068 22222 26188 22250
rect 26068 22166 26096 22222
rect 26056 22160 26108 22166
rect 26252 22148 26280 22510
rect 26056 22102 26108 22108
rect 26160 22120 26280 22148
rect 25884 22066 26004 22094
rect 25780 22024 25832 22030
rect 25780 21966 25832 21972
rect 25792 21350 25820 21966
rect 25780 21344 25832 21350
rect 25780 21286 25832 21292
rect 25780 21004 25832 21010
rect 25780 20946 25832 20952
rect 25792 20777 25820 20946
rect 25778 20768 25834 20777
rect 25778 20703 25834 20712
rect 25884 19938 25912 22066
rect 25964 22024 26016 22030
rect 25962 21992 25964 22001
rect 26016 21992 26018 22001
rect 25962 21927 26018 21936
rect 26056 21956 26108 21962
rect 26056 21898 26108 21904
rect 25962 21856 26018 21865
rect 25962 21791 26018 21800
rect 25976 21622 26004 21791
rect 25964 21616 26016 21622
rect 25964 21558 26016 21564
rect 25976 20602 26004 21558
rect 25964 20596 26016 20602
rect 25964 20538 26016 20544
rect 26068 20262 26096 21898
rect 26160 20534 26188 22120
rect 26436 22030 26464 22902
rect 26804 22658 26832 28478
rect 26884 28518 26936 28524
rect 26884 28460 26936 28466
rect 26896 28422 26924 28460
rect 26884 28416 26936 28422
rect 26884 28358 26936 28364
rect 26896 28257 26924 28358
rect 26882 28248 26938 28257
rect 26882 28183 26938 28192
rect 26884 27872 26936 27878
rect 26884 27814 26936 27820
rect 26896 27713 26924 27814
rect 26882 27704 26938 27713
rect 26882 27639 26938 27648
rect 26988 26382 27016 28580
rect 27080 28370 27108 30670
rect 27264 30394 27292 31078
rect 27528 30728 27580 30734
rect 27528 30670 27580 30676
rect 27436 30592 27488 30598
rect 27436 30534 27488 30540
rect 27252 30388 27304 30394
rect 27252 30330 27304 30336
rect 27344 29028 27396 29034
rect 27344 28970 27396 28976
rect 27252 28960 27304 28966
rect 27252 28902 27304 28908
rect 27264 28558 27292 28902
rect 27160 28552 27212 28558
rect 27158 28520 27160 28529
rect 27252 28552 27304 28558
rect 27212 28520 27214 28529
rect 27252 28494 27304 28500
rect 27158 28455 27214 28464
rect 27252 28416 27304 28422
rect 27080 28342 27200 28370
rect 27252 28358 27304 28364
rect 27172 27010 27200 28342
rect 27264 28218 27292 28358
rect 27252 28212 27304 28218
rect 27252 28154 27304 28160
rect 27252 28076 27304 28082
rect 27252 28018 27304 28024
rect 27264 27674 27292 28018
rect 27356 27674 27384 28970
rect 27448 28801 27476 30534
rect 27540 30258 27568 30670
rect 27528 30252 27580 30258
rect 27528 30194 27580 30200
rect 27540 29730 27568 30194
rect 27632 29850 27660 31878
rect 27620 29844 27672 29850
rect 27620 29786 27672 29792
rect 27540 29702 27660 29730
rect 27528 29504 27580 29510
rect 27528 29446 27580 29452
rect 27434 28792 27490 28801
rect 27434 28727 27490 28736
rect 27540 28558 27568 29446
rect 27436 28552 27488 28558
rect 27436 28494 27488 28500
rect 27528 28552 27580 28558
rect 27528 28494 27580 28500
rect 27252 27668 27304 27674
rect 27252 27610 27304 27616
rect 27344 27668 27396 27674
rect 27344 27610 27396 27616
rect 27252 27532 27304 27538
rect 27252 27474 27304 27480
rect 27080 26982 27200 27010
rect 26976 26376 27028 26382
rect 26976 26318 27028 26324
rect 27080 26246 27108 26982
rect 27160 26920 27212 26926
rect 27160 26862 27212 26868
rect 27068 26240 27120 26246
rect 27068 26182 27120 26188
rect 26974 25936 27030 25945
rect 26884 25900 26936 25906
rect 27080 25906 27108 26182
rect 26974 25871 27030 25880
rect 27068 25900 27120 25906
rect 26884 25842 26936 25848
rect 26896 23882 26924 25842
rect 26988 25786 27016 25871
rect 27068 25842 27120 25848
rect 26988 25758 27108 25786
rect 26976 25152 27028 25158
rect 26976 25094 27028 25100
rect 26988 24954 27016 25094
rect 26976 24948 27028 24954
rect 26976 24890 27028 24896
rect 26976 24200 27028 24206
rect 26974 24168 26976 24177
rect 27028 24168 27030 24177
rect 26974 24103 27030 24112
rect 26896 23854 27016 23882
rect 26884 23520 26936 23526
rect 26884 23462 26936 23468
rect 26896 23322 26924 23462
rect 26884 23316 26936 23322
rect 26884 23258 26936 23264
rect 26896 23118 26924 23258
rect 26884 23112 26936 23118
rect 26884 23054 26936 23060
rect 26884 22976 26936 22982
rect 26884 22918 26936 22924
rect 26528 22630 26832 22658
rect 26332 22024 26384 22030
rect 26332 21966 26384 21972
rect 26424 22024 26476 22030
rect 26424 21966 26476 21972
rect 26344 21486 26372 21966
rect 26332 21480 26384 21486
rect 26332 21422 26384 21428
rect 26148 20528 26200 20534
rect 26148 20470 26200 20476
rect 26240 20528 26292 20534
rect 26240 20470 26292 20476
rect 26252 20330 26280 20470
rect 26240 20324 26292 20330
rect 26240 20266 26292 20272
rect 26056 20256 26108 20262
rect 26056 20198 26108 20204
rect 25792 19922 25912 19938
rect 25780 19916 25912 19922
rect 25832 19910 25912 19916
rect 25780 19858 25832 19864
rect 25688 19440 25740 19446
rect 25688 19382 25740 19388
rect 25596 19372 25648 19378
rect 25596 19314 25648 19320
rect 25608 18970 25636 19314
rect 25792 19174 25820 19858
rect 25872 19848 25924 19854
rect 25872 19790 25924 19796
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 25596 18964 25648 18970
rect 25596 18906 25648 18912
rect 25688 18964 25740 18970
rect 25688 18906 25740 18912
rect 25700 18850 25728 18906
rect 25516 18822 25728 18850
rect 25504 18692 25556 18698
rect 25504 18634 25556 18640
rect 25516 17678 25544 18634
rect 25504 17672 25556 17678
rect 25504 17614 25556 17620
rect 25516 16590 25544 17614
rect 25504 16584 25556 16590
rect 25504 16526 25556 16532
rect 25516 16114 25544 16526
rect 25504 16108 25556 16114
rect 25504 16050 25556 16056
rect 25320 16040 25372 16046
rect 25320 15982 25372 15988
rect 25412 16040 25464 16046
rect 25412 15982 25464 15988
rect 25136 14952 25188 14958
rect 25136 14894 25188 14900
rect 25044 14000 25096 14006
rect 25044 13942 25096 13948
rect 25148 12850 25176 14894
rect 25228 14340 25280 14346
rect 25228 14282 25280 14288
rect 25240 14113 25268 14282
rect 25424 14278 25452 15982
rect 25504 14408 25556 14414
rect 25502 14376 25504 14385
rect 25556 14376 25558 14385
rect 25502 14311 25558 14320
rect 25412 14272 25464 14278
rect 25412 14214 25464 14220
rect 25226 14104 25282 14113
rect 25226 14039 25282 14048
rect 25240 13802 25268 14039
rect 25228 13796 25280 13802
rect 25228 13738 25280 13744
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 25136 12844 25188 12850
rect 25136 12786 25188 12792
rect 24872 12442 24900 12786
rect 24952 12640 25004 12646
rect 24952 12582 25004 12588
rect 24860 12436 24912 12442
rect 24860 12378 24912 12384
rect 24676 12096 24728 12102
rect 24504 12056 24676 12084
rect 24676 12038 24728 12044
rect 24964 11762 24992 12582
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24032 11620 24084 11626
rect 24032 11562 24084 11568
rect 22100 11222 22152 11228
rect 22572 11206 22692 11234
rect 22376 11144 22428 11150
rect 22376 11086 22428 11092
rect 22388 10266 22416 11086
rect 22468 11076 22520 11082
rect 22468 11018 22520 11024
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 22376 10260 22428 10266
rect 22376 10202 22428 10208
rect 22100 10192 22152 10198
rect 22100 10134 22152 10140
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 22020 9586 22048 9998
rect 22008 9580 22060 9586
rect 22008 9522 22060 9528
rect 22112 9042 22140 10134
rect 22204 9586 22232 10202
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 22480 9500 22508 11018
rect 22572 10266 22600 11206
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 23112 11144 23164 11150
rect 23112 11086 23164 11092
rect 22560 10260 22612 10266
rect 22560 10202 22612 10208
rect 22560 10056 22612 10062
rect 22558 10024 22560 10033
rect 22664 10044 22692 11086
rect 23124 10062 23152 11086
rect 25148 11014 25176 12786
rect 25424 12646 25452 14214
rect 25608 13938 25636 18822
rect 25792 17218 25820 19110
rect 25884 18698 25912 19790
rect 25964 19440 26016 19446
rect 25964 19382 26016 19388
rect 25976 18748 26004 19382
rect 26068 19378 26096 20198
rect 26238 19408 26294 19417
rect 26056 19372 26108 19378
rect 26238 19343 26294 19352
rect 26056 19314 26108 19320
rect 26148 19304 26200 19310
rect 26252 19258 26280 19343
rect 26200 19252 26280 19258
rect 26148 19246 26280 19252
rect 26160 19230 26280 19246
rect 26056 18760 26108 18766
rect 25976 18720 26056 18748
rect 25872 18692 25924 18698
rect 25872 18634 25924 18640
rect 25884 18057 25912 18634
rect 25870 18048 25926 18057
rect 25870 17983 25926 17992
rect 25700 17190 25820 17218
rect 25700 16590 25728 17190
rect 25780 17128 25832 17134
rect 25780 17070 25832 17076
rect 25792 16794 25820 17070
rect 25780 16788 25832 16794
rect 25780 16730 25832 16736
rect 25870 16688 25926 16697
rect 25870 16623 25926 16632
rect 25884 16590 25912 16623
rect 25688 16584 25740 16590
rect 25872 16584 25924 16590
rect 25688 16526 25740 16532
rect 25792 16544 25872 16572
rect 25792 16454 25820 16544
rect 25872 16526 25924 16532
rect 25780 16448 25832 16454
rect 25780 16390 25832 16396
rect 25872 16448 25924 16454
rect 25872 16390 25924 16396
rect 25688 16040 25740 16046
rect 25688 15982 25740 15988
rect 25700 15706 25728 15982
rect 25884 15978 25912 16390
rect 25872 15972 25924 15978
rect 25872 15914 25924 15920
rect 25688 15700 25740 15706
rect 25688 15642 25740 15648
rect 25976 15586 26004 18720
rect 26056 18702 26108 18708
rect 26148 18692 26200 18698
rect 26148 18634 26200 18640
rect 26160 18154 26188 18634
rect 26148 18148 26200 18154
rect 26148 18090 26200 18096
rect 26056 17808 26108 17814
rect 26056 17750 26108 17756
rect 26068 16969 26096 17750
rect 26148 17536 26200 17542
rect 26148 17478 26200 17484
rect 26160 17338 26188 17478
rect 26148 17332 26200 17338
rect 26148 17274 26200 17280
rect 26252 16998 26280 19230
rect 26330 19000 26386 19009
rect 26330 18935 26386 18944
rect 26344 18698 26372 18935
rect 26332 18692 26384 18698
rect 26332 18634 26384 18640
rect 26344 17746 26372 18634
rect 26332 17740 26384 17746
rect 26332 17682 26384 17688
rect 26332 17128 26384 17134
rect 26330 17096 26332 17105
rect 26384 17096 26386 17105
rect 26330 17031 26386 17040
rect 26240 16992 26292 16998
rect 26054 16960 26110 16969
rect 26240 16934 26292 16940
rect 26054 16895 26110 16904
rect 26330 16688 26386 16697
rect 26330 16623 26386 16632
rect 26146 16552 26202 16561
rect 26056 16516 26108 16522
rect 26344 16522 26372 16623
rect 26146 16487 26202 16496
rect 26332 16516 26384 16522
rect 26056 16458 26108 16464
rect 25700 15558 26004 15586
rect 25596 13932 25648 13938
rect 25596 13874 25648 13880
rect 25412 12640 25464 12646
rect 25412 12582 25464 12588
rect 25608 12442 25636 13874
rect 25596 12436 25648 12442
rect 25596 12378 25648 12384
rect 25608 12345 25636 12378
rect 25594 12336 25650 12345
rect 25594 12271 25650 12280
rect 25596 12232 25648 12238
rect 25596 12174 25648 12180
rect 25608 11830 25636 12174
rect 25700 12170 25728 15558
rect 25780 15496 25832 15502
rect 25964 15496 26016 15502
rect 25832 15456 25912 15484
rect 25780 15438 25832 15444
rect 25778 15192 25834 15201
rect 25778 15127 25834 15136
rect 25792 14618 25820 15127
rect 25780 14612 25832 14618
rect 25780 14554 25832 14560
rect 25780 14408 25832 14414
rect 25780 14350 25832 14356
rect 25792 14074 25820 14350
rect 25884 14278 25912 15456
rect 25964 15438 26016 15444
rect 25976 15094 26004 15438
rect 25964 15088 26016 15094
rect 25964 15030 26016 15036
rect 25964 14952 26016 14958
rect 25964 14894 26016 14900
rect 25976 14414 26004 14894
rect 25964 14408 26016 14414
rect 25964 14350 26016 14356
rect 25872 14272 25924 14278
rect 25872 14214 25924 14220
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 25780 13932 25832 13938
rect 25780 13874 25832 13880
rect 25688 12164 25740 12170
rect 25688 12106 25740 12112
rect 25792 11898 25820 13874
rect 25872 12776 25924 12782
rect 25872 12718 25924 12724
rect 25884 12442 25912 12718
rect 26068 12442 26096 16458
rect 26160 15570 26188 16487
rect 26332 16458 26384 16464
rect 26332 16040 26384 16046
rect 26332 15982 26384 15988
rect 26240 15972 26292 15978
rect 26240 15914 26292 15920
rect 26252 15570 26280 15914
rect 26148 15564 26200 15570
rect 26148 15506 26200 15512
rect 26240 15564 26292 15570
rect 26240 15506 26292 15512
rect 26148 15428 26200 15434
rect 26148 15370 26200 15376
rect 26160 14890 26188 15370
rect 26344 15366 26372 15982
rect 26332 15360 26384 15366
rect 26238 15328 26294 15337
rect 26332 15302 26384 15308
rect 26238 15263 26294 15272
rect 26252 15162 26280 15263
rect 26240 15156 26292 15162
rect 26240 15098 26292 15104
rect 26240 15020 26292 15026
rect 26240 14962 26292 14968
rect 26148 14884 26200 14890
rect 26148 14826 26200 14832
rect 26252 13326 26280 14962
rect 26436 13802 26464 21966
rect 26528 20942 26556 22630
rect 26700 21480 26752 21486
rect 26606 21448 26662 21457
rect 26896 21434 26924 22918
rect 26700 21422 26752 21428
rect 26606 21383 26662 21392
rect 26516 20936 26568 20942
rect 26516 20878 26568 20884
rect 26528 19378 26556 20878
rect 26620 20602 26648 21383
rect 26608 20596 26660 20602
rect 26608 20538 26660 20544
rect 26620 19378 26648 20538
rect 26516 19372 26568 19378
rect 26516 19314 26568 19320
rect 26608 19372 26660 19378
rect 26608 19314 26660 19320
rect 26606 19272 26662 19281
rect 26606 19207 26608 19216
rect 26660 19207 26662 19216
rect 26608 19178 26660 19184
rect 26608 18964 26660 18970
rect 26608 18906 26660 18912
rect 26620 18737 26648 18906
rect 26606 18728 26662 18737
rect 26606 18663 26662 18672
rect 26516 18624 26568 18630
rect 26516 18566 26568 18572
rect 26528 18426 26556 18566
rect 26516 18420 26568 18426
rect 26516 18362 26568 18368
rect 26514 17912 26570 17921
rect 26514 17847 26570 17856
rect 26528 17202 26556 17847
rect 26712 17490 26740 21422
rect 26620 17462 26740 17490
rect 26804 21406 26924 21434
rect 26516 17196 26568 17202
rect 26516 17138 26568 17144
rect 26516 16992 26568 16998
rect 26516 16934 26568 16940
rect 26528 14958 26556 16934
rect 26620 16114 26648 17462
rect 26698 17368 26754 17377
rect 26698 17303 26700 17312
rect 26752 17303 26754 17312
rect 26700 17274 26752 17280
rect 26700 16176 26752 16182
rect 26700 16118 26752 16124
rect 26608 16108 26660 16114
rect 26608 16050 26660 16056
rect 26608 15496 26660 15502
rect 26608 15438 26660 15444
rect 26516 14952 26568 14958
rect 26516 14894 26568 14900
rect 26516 13932 26568 13938
rect 26516 13874 26568 13880
rect 26424 13796 26476 13802
rect 26424 13738 26476 13744
rect 26240 13320 26292 13326
rect 26240 13262 26292 13268
rect 26240 12844 26292 12850
rect 26240 12786 26292 12792
rect 25872 12436 25924 12442
rect 25872 12378 25924 12384
rect 26056 12436 26108 12442
rect 26056 12378 26108 12384
rect 26252 12434 26280 12786
rect 26252 12406 26372 12434
rect 26056 12300 26108 12306
rect 26252 12288 26280 12406
rect 26108 12260 26280 12288
rect 26056 12242 26108 12248
rect 26344 12238 26372 12406
rect 26528 12345 26556 13874
rect 26620 13802 26648 15438
rect 26712 14346 26740 16118
rect 26804 15978 26832 21406
rect 26884 20392 26936 20398
rect 26884 20334 26936 20340
rect 26896 19310 26924 20334
rect 26988 19334 27016 23854
rect 27080 22166 27108 25758
rect 27068 22160 27120 22166
rect 27068 22102 27120 22108
rect 27068 22024 27120 22030
rect 27068 21966 27120 21972
rect 27080 21622 27108 21966
rect 27172 21690 27200 26862
rect 27264 25974 27292 27474
rect 27356 26858 27384 27610
rect 27448 27470 27476 28494
rect 27528 28416 27580 28422
rect 27528 28358 27580 28364
rect 27540 28150 27568 28358
rect 27528 28144 27580 28150
rect 27528 28086 27580 28092
rect 27632 28014 27660 29702
rect 27724 28762 27752 33798
rect 27816 31414 27844 36654
rect 28000 36242 28028 38916
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 31208 38276 31260 38282
rect 31208 38218 31260 38224
rect 30012 38208 30064 38214
rect 30012 38150 30064 38156
rect 29368 37664 29420 37670
rect 29368 37606 29420 37612
rect 28448 37256 28500 37262
rect 28448 37198 28500 37204
rect 28172 36916 28224 36922
rect 28172 36858 28224 36864
rect 28184 36718 28212 36858
rect 28172 36712 28224 36718
rect 28172 36654 28224 36660
rect 28460 36378 28488 37198
rect 29380 36582 29408 37606
rect 30024 36786 30052 38150
rect 31220 37330 31248 38218
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 31208 37324 31260 37330
rect 31208 37266 31260 37272
rect 31852 37188 31904 37194
rect 31852 37130 31904 37136
rect 35624 37188 35676 37194
rect 35624 37130 35676 37136
rect 31484 37120 31536 37126
rect 31484 37062 31536 37068
rect 30012 36780 30064 36786
rect 30012 36722 30064 36728
rect 29828 36712 29880 36718
rect 29828 36654 29880 36660
rect 28724 36576 28776 36582
rect 28724 36518 28776 36524
rect 29368 36576 29420 36582
rect 29368 36518 29420 36524
rect 28736 36378 28764 36518
rect 28356 36372 28408 36378
rect 28356 36314 28408 36320
rect 28448 36372 28500 36378
rect 28448 36314 28500 36320
rect 28724 36372 28776 36378
rect 28724 36314 28776 36320
rect 27988 36236 28040 36242
rect 27988 36178 28040 36184
rect 28264 36168 28316 36174
rect 28262 36136 28264 36145
rect 28316 36136 28318 36145
rect 28262 36071 28318 36080
rect 28080 36032 28132 36038
rect 28080 35974 28132 35980
rect 27988 33652 28040 33658
rect 27988 33594 28040 33600
rect 28000 32609 28028 33594
rect 28092 32910 28120 35974
rect 28172 35760 28224 35766
rect 28172 35702 28224 35708
rect 28080 32904 28132 32910
rect 28080 32846 28132 32852
rect 27986 32600 28042 32609
rect 27986 32535 28042 32544
rect 27988 32360 28040 32366
rect 27988 32302 28040 32308
rect 27896 32292 27948 32298
rect 27896 32234 27948 32240
rect 27908 32026 27936 32234
rect 28000 32026 28028 32302
rect 27896 32020 27948 32026
rect 27896 31962 27948 31968
rect 27988 32020 28040 32026
rect 27988 31962 28040 31968
rect 28092 31906 28120 32846
rect 28184 32348 28212 35702
rect 28264 34672 28316 34678
rect 28264 34614 28316 34620
rect 28276 32842 28304 34614
rect 28264 32836 28316 32842
rect 28264 32778 28316 32784
rect 28276 32502 28304 32778
rect 28264 32496 28316 32502
rect 28264 32438 28316 32444
rect 28184 32320 28304 32348
rect 28000 31878 28120 31906
rect 27896 31680 27948 31686
rect 27894 31648 27896 31657
rect 27948 31648 27950 31657
rect 27894 31583 27950 31592
rect 27804 31408 27856 31414
rect 27804 31350 27856 31356
rect 27896 31340 27948 31346
rect 27896 31282 27948 31288
rect 27908 30394 27936 31282
rect 27896 30388 27948 30394
rect 27896 30330 27948 30336
rect 27804 29504 27856 29510
rect 27804 29446 27856 29452
rect 27712 28756 27764 28762
rect 27712 28698 27764 28704
rect 27724 28422 27752 28698
rect 27712 28416 27764 28422
rect 27712 28358 27764 28364
rect 27710 28248 27766 28257
rect 27710 28183 27766 28192
rect 27620 28008 27672 28014
rect 27620 27950 27672 27956
rect 27528 27940 27580 27946
rect 27528 27882 27580 27888
rect 27436 27464 27488 27470
rect 27436 27406 27488 27412
rect 27344 26852 27396 26858
rect 27344 26794 27396 26800
rect 27356 26364 27384 26794
rect 27540 26382 27568 27882
rect 27724 27878 27752 28183
rect 27712 27872 27764 27878
rect 27712 27814 27764 27820
rect 27816 27606 27844 29446
rect 27894 29336 27950 29345
rect 27894 29271 27950 29280
rect 27804 27600 27856 27606
rect 27804 27542 27856 27548
rect 27804 26580 27856 26586
rect 27804 26522 27856 26528
rect 27816 26382 27844 26522
rect 27908 26432 27936 29271
rect 28000 28257 28028 31878
rect 28080 31816 28132 31822
rect 28080 31758 28132 31764
rect 27986 28248 28042 28257
rect 27986 28183 28042 28192
rect 27988 28076 28040 28082
rect 27988 28018 28040 28024
rect 28000 27577 28028 28018
rect 28092 28014 28120 31758
rect 28172 31748 28224 31754
rect 28172 31690 28224 31696
rect 28184 31521 28212 31690
rect 28170 31512 28226 31521
rect 28170 31447 28226 31456
rect 28276 31142 28304 32320
rect 28264 31136 28316 31142
rect 28264 31078 28316 31084
rect 28262 30288 28318 30297
rect 28262 30223 28318 30232
rect 28276 30190 28304 30223
rect 28264 30184 28316 30190
rect 28264 30126 28316 30132
rect 28170 29472 28226 29481
rect 28170 29407 28226 29416
rect 28184 28762 28212 29407
rect 28276 29073 28304 30126
rect 28262 29064 28318 29073
rect 28262 28999 28318 29008
rect 28264 28960 28316 28966
rect 28264 28902 28316 28908
rect 28172 28756 28224 28762
rect 28172 28698 28224 28704
rect 28276 28506 28304 28902
rect 28368 28801 28396 36314
rect 29380 36242 29408 36518
rect 29736 36372 29788 36378
rect 29736 36314 29788 36320
rect 29368 36236 29420 36242
rect 29368 36178 29420 36184
rect 29000 36168 29052 36174
rect 29000 36110 29052 36116
rect 28632 36100 28684 36106
rect 28632 36042 28684 36048
rect 28644 36009 28672 36042
rect 28908 36032 28960 36038
rect 28630 36000 28686 36009
rect 28908 35974 28960 35980
rect 28630 35935 28686 35944
rect 28920 35086 28948 35974
rect 29012 35086 29040 36110
rect 29276 35624 29328 35630
rect 29276 35566 29328 35572
rect 29184 35284 29236 35290
rect 29184 35226 29236 35232
rect 28908 35080 28960 35086
rect 28908 35022 28960 35028
rect 29000 35080 29052 35086
rect 29000 35022 29052 35028
rect 28816 35012 28868 35018
rect 28816 34954 28868 34960
rect 28828 34610 28856 34954
rect 28908 34672 28960 34678
rect 28908 34614 28960 34620
rect 28816 34604 28868 34610
rect 28816 34546 28868 34552
rect 28540 34468 28592 34474
rect 28540 34410 28592 34416
rect 28552 34202 28580 34410
rect 28724 34400 28776 34406
rect 28724 34342 28776 34348
rect 28540 34196 28592 34202
rect 28540 34138 28592 34144
rect 28736 34134 28764 34342
rect 28724 34128 28776 34134
rect 28724 34070 28776 34076
rect 28828 33998 28856 34546
rect 28920 34542 28948 34614
rect 28908 34536 28960 34542
rect 28908 34478 28960 34484
rect 29012 34388 29040 35022
rect 29092 34740 29144 34746
rect 29092 34682 29144 34688
rect 28920 34360 29040 34388
rect 28540 33992 28592 33998
rect 28540 33934 28592 33940
rect 28816 33992 28868 33998
rect 28816 33934 28868 33940
rect 28446 31376 28502 31385
rect 28446 31311 28502 31320
rect 28460 30802 28488 31311
rect 28552 31278 28580 33934
rect 28828 33386 28856 33934
rect 28920 33930 28948 34360
rect 29000 33992 29052 33998
rect 29000 33934 29052 33940
rect 28908 33924 28960 33930
rect 28908 33866 28960 33872
rect 28920 33454 28948 33866
rect 29012 33590 29040 33934
rect 29000 33584 29052 33590
rect 29000 33526 29052 33532
rect 28908 33448 28960 33454
rect 28908 33390 28960 33396
rect 28816 33380 28868 33386
rect 28816 33322 28868 33328
rect 28814 33144 28870 33153
rect 28814 33079 28870 33088
rect 28828 32745 28856 33079
rect 28814 32736 28870 32745
rect 28814 32671 28870 32680
rect 28632 32496 28684 32502
rect 28632 32438 28684 32444
rect 28540 31272 28592 31278
rect 28540 31214 28592 31220
rect 28540 31136 28592 31142
rect 28540 31078 28592 31084
rect 28448 30796 28500 30802
rect 28448 30738 28500 30744
rect 28448 30116 28500 30122
rect 28448 30058 28500 30064
rect 28354 28792 28410 28801
rect 28354 28727 28410 28736
rect 28460 28665 28488 30058
rect 28552 28994 28580 31078
rect 28644 29714 28672 32438
rect 28828 32434 28856 32671
rect 28816 32428 28868 32434
rect 28816 32370 28868 32376
rect 28920 31958 28948 33390
rect 29000 32428 29052 32434
rect 29000 32370 29052 32376
rect 29012 32230 29040 32370
rect 29000 32224 29052 32230
rect 29000 32166 29052 32172
rect 28908 31952 28960 31958
rect 28908 31894 28960 31900
rect 29012 31822 29040 32166
rect 29104 31958 29132 34682
rect 29196 33946 29224 35226
rect 29288 34678 29316 35566
rect 29276 34672 29328 34678
rect 29276 34614 29328 34620
rect 29288 34134 29316 34614
rect 29380 34474 29408 36178
rect 29748 35766 29776 36314
rect 29840 36174 29868 36654
rect 30024 36242 30052 36722
rect 30196 36644 30248 36650
rect 30196 36586 30248 36592
rect 30012 36236 30064 36242
rect 30012 36178 30064 36184
rect 29828 36168 29880 36174
rect 29828 36110 29880 36116
rect 29736 35760 29788 35766
rect 29736 35702 29788 35708
rect 29840 35630 29868 36110
rect 29920 35692 29972 35698
rect 29920 35634 29972 35640
rect 30104 35692 30156 35698
rect 30104 35634 30156 35640
rect 29828 35624 29880 35630
rect 29828 35566 29880 35572
rect 29552 35148 29604 35154
rect 29552 35090 29604 35096
rect 29460 34944 29512 34950
rect 29460 34886 29512 34892
rect 29472 34610 29500 34886
rect 29564 34746 29592 35090
rect 29736 35012 29788 35018
rect 29736 34954 29788 34960
rect 29552 34740 29604 34746
rect 29552 34682 29604 34688
rect 29748 34678 29776 34954
rect 29736 34672 29788 34678
rect 29932 34649 29960 35634
rect 30012 34944 30064 34950
rect 30012 34886 30064 34892
rect 30024 34785 30052 34886
rect 30010 34776 30066 34785
rect 30116 34746 30144 35634
rect 30010 34711 30066 34720
rect 30104 34740 30156 34746
rect 30104 34682 30156 34688
rect 30208 34678 30236 36586
rect 31116 36100 31168 36106
rect 31116 36042 31168 36048
rect 31128 35698 31156 36042
rect 30288 35692 30340 35698
rect 30288 35634 30340 35640
rect 31116 35692 31168 35698
rect 31116 35634 31168 35640
rect 30012 34672 30064 34678
rect 29736 34614 29788 34620
rect 29918 34640 29974 34649
rect 29460 34604 29512 34610
rect 29460 34546 29512 34552
rect 29552 34604 29604 34610
rect 30012 34614 30064 34620
rect 30196 34672 30248 34678
rect 30196 34614 30248 34620
rect 29918 34575 29974 34584
rect 29552 34546 29604 34552
rect 29368 34468 29420 34474
rect 29368 34410 29420 34416
rect 29564 34241 29592 34546
rect 30024 34524 30052 34614
rect 29734 34504 29790 34513
rect 29734 34439 29736 34448
rect 29788 34439 29790 34448
rect 29840 34496 30052 34524
rect 29736 34410 29788 34416
rect 29550 34232 29606 34241
rect 29550 34167 29606 34176
rect 29276 34128 29328 34134
rect 29276 34070 29328 34076
rect 29644 33992 29696 33998
rect 29196 33918 29316 33946
rect 29644 33934 29696 33940
rect 29184 33856 29236 33862
rect 29184 33798 29236 33804
rect 29092 31952 29144 31958
rect 29092 31894 29144 31900
rect 29000 31816 29052 31822
rect 29000 31758 29052 31764
rect 29092 31748 29144 31754
rect 29092 31690 29144 31696
rect 29000 31476 29052 31482
rect 29000 31418 29052 31424
rect 28816 30796 28868 30802
rect 28816 30738 28868 30744
rect 28632 29708 28684 29714
rect 28632 29650 28684 29656
rect 28828 29345 28856 30738
rect 28908 30728 28960 30734
rect 28908 30670 28960 30676
rect 28920 30569 28948 30670
rect 28906 30560 28962 30569
rect 28906 30495 28962 30504
rect 28814 29336 28870 29345
rect 28814 29271 28870 29280
rect 28828 29073 28856 29271
rect 28814 29064 28870 29073
rect 28814 28999 28870 29008
rect 28552 28966 28672 28994
rect 28644 28937 28672 28966
rect 28630 28928 28686 28937
rect 28630 28863 28686 28872
rect 28724 28756 28776 28762
rect 28552 28716 28724 28744
rect 28446 28656 28502 28665
rect 28446 28591 28502 28600
rect 28184 28490 28304 28506
rect 28356 28552 28408 28558
rect 28552 28540 28580 28716
rect 28724 28698 28776 28704
rect 28630 28656 28686 28665
rect 29012 28642 29040 31418
rect 29104 31346 29132 31690
rect 29092 31340 29144 31346
rect 29092 31282 29144 31288
rect 29196 28762 29224 33798
rect 29288 32774 29316 33918
rect 29460 33924 29512 33930
rect 29460 33866 29512 33872
rect 29368 33856 29420 33862
rect 29368 33798 29420 33804
rect 29276 32768 29328 32774
rect 29276 32710 29328 32716
rect 29288 32434 29316 32710
rect 29276 32428 29328 32434
rect 29276 32370 29328 32376
rect 29288 31226 29316 32370
rect 29380 31482 29408 33798
rect 29472 33454 29500 33866
rect 29460 33448 29512 33454
rect 29460 33390 29512 33396
rect 29656 32434 29684 33934
rect 29460 32428 29512 32434
rect 29644 32428 29696 32434
rect 29460 32370 29512 32376
rect 29564 32388 29644 32416
rect 29472 31686 29500 32370
rect 29564 31754 29592 32388
rect 29644 32370 29696 32376
rect 29644 32224 29696 32230
rect 29644 32166 29696 32172
rect 29656 31890 29684 32166
rect 29644 31884 29696 31890
rect 29644 31826 29696 31832
rect 29552 31748 29604 31754
rect 29552 31690 29604 31696
rect 29460 31680 29512 31686
rect 29460 31622 29512 31628
rect 29368 31476 29420 31482
rect 29368 31418 29420 31424
rect 29472 31260 29500 31622
rect 29552 31272 29604 31278
rect 29472 31232 29552 31260
rect 29288 31198 29408 31226
rect 29552 31214 29604 31220
rect 29276 31136 29328 31142
rect 29276 31078 29328 31084
rect 29184 28756 29236 28762
rect 29184 28698 29236 28704
rect 28630 28591 28686 28600
rect 28736 28614 29040 28642
rect 29092 28688 29144 28694
rect 29092 28630 29144 28636
rect 28408 28512 28580 28540
rect 28356 28494 28408 28500
rect 28172 28484 28304 28490
rect 28224 28478 28304 28484
rect 28172 28426 28224 28432
rect 28264 28416 28316 28422
rect 28264 28358 28316 28364
rect 28356 28416 28408 28422
rect 28356 28358 28408 28364
rect 28276 28257 28304 28358
rect 28262 28248 28318 28257
rect 28368 28218 28396 28358
rect 28552 28218 28580 28512
rect 28262 28183 28318 28192
rect 28356 28212 28408 28218
rect 28356 28154 28408 28160
rect 28540 28212 28592 28218
rect 28540 28154 28592 28160
rect 28538 28112 28594 28121
rect 28172 28076 28224 28082
rect 28224 28036 28396 28064
rect 28538 28047 28594 28056
rect 28172 28018 28224 28024
rect 28080 28008 28132 28014
rect 28080 27950 28132 27956
rect 27986 27568 28042 27577
rect 27986 27503 28042 27512
rect 28092 26926 28120 27950
rect 28184 27713 28212 28018
rect 28368 27946 28396 28036
rect 28552 28014 28580 28047
rect 28540 28008 28592 28014
rect 28540 27950 28592 27956
rect 28356 27940 28408 27946
rect 28356 27882 28408 27888
rect 28264 27872 28316 27878
rect 28264 27814 28316 27820
rect 28170 27704 28226 27713
rect 28170 27639 28226 27648
rect 28184 27538 28212 27639
rect 28172 27532 28224 27538
rect 28172 27474 28224 27480
rect 28172 26988 28224 26994
rect 28172 26930 28224 26936
rect 28080 26920 28132 26926
rect 28080 26862 28132 26868
rect 27908 26404 28028 26432
rect 27528 26376 27580 26382
rect 27356 26336 27476 26364
rect 27344 26240 27396 26246
rect 27344 26182 27396 26188
rect 27252 25968 27304 25974
rect 27252 25910 27304 25916
rect 27356 25906 27384 26182
rect 27448 26042 27476 26336
rect 27804 26376 27856 26382
rect 27580 26324 27752 26330
rect 27528 26318 27752 26324
rect 27804 26318 27856 26324
rect 27540 26302 27752 26318
rect 27620 26240 27672 26246
rect 27620 26182 27672 26188
rect 27436 26036 27488 26042
rect 27436 25978 27488 25984
rect 27344 25900 27396 25906
rect 27344 25842 27396 25848
rect 27632 25838 27660 26182
rect 27620 25832 27672 25838
rect 27620 25774 27672 25780
rect 27436 25696 27488 25702
rect 27436 25638 27488 25644
rect 27448 24886 27476 25638
rect 27528 25356 27580 25362
rect 27528 25298 27580 25304
rect 27344 24880 27396 24886
rect 27344 24822 27396 24828
rect 27436 24880 27488 24886
rect 27436 24822 27488 24828
rect 27252 24608 27304 24614
rect 27252 24550 27304 24556
rect 27264 24070 27292 24550
rect 27356 24392 27384 24822
rect 27436 24404 27488 24410
rect 27356 24364 27436 24392
rect 27436 24346 27488 24352
rect 27540 24206 27568 25298
rect 27632 25294 27660 25774
rect 27620 25288 27672 25294
rect 27620 25230 27672 25236
rect 27620 24948 27672 24954
rect 27620 24890 27672 24896
rect 27632 24342 27660 24890
rect 27620 24336 27672 24342
rect 27620 24278 27672 24284
rect 27528 24200 27580 24206
rect 27528 24142 27580 24148
rect 27620 24200 27672 24206
rect 27620 24142 27672 24148
rect 27252 24064 27304 24070
rect 27252 24006 27304 24012
rect 27344 24064 27396 24070
rect 27344 24006 27396 24012
rect 27264 23118 27292 24006
rect 27356 23322 27384 24006
rect 27436 23520 27488 23526
rect 27436 23462 27488 23468
rect 27344 23316 27396 23322
rect 27344 23258 27396 23264
rect 27252 23112 27304 23118
rect 27252 23054 27304 23060
rect 27448 22094 27476 23462
rect 27540 22778 27568 24142
rect 27632 23322 27660 24142
rect 27724 23730 27752 26302
rect 28000 26246 28028 26404
rect 27896 26240 27948 26246
rect 27988 26240 28040 26246
rect 27896 26182 27948 26188
rect 27986 26208 27988 26217
rect 28040 26208 28042 26217
rect 27804 25696 27856 25702
rect 27804 25638 27856 25644
rect 27816 25498 27844 25638
rect 27804 25492 27856 25498
rect 27804 25434 27856 25440
rect 27908 25344 27936 26182
rect 27986 26143 28042 26152
rect 27816 25316 27936 25344
rect 27816 25158 27844 25316
rect 27896 25220 27948 25226
rect 27948 25180 28028 25208
rect 27896 25162 27948 25168
rect 27804 25152 27856 25158
rect 27804 25094 27856 25100
rect 27712 23724 27764 23730
rect 27712 23666 27764 23672
rect 27712 23588 27764 23594
rect 27712 23530 27764 23536
rect 27620 23316 27672 23322
rect 27620 23258 27672 23264
rect 27620 23112 27672 23118
rect 27620 23054 27672 23060
rect 27528 22772 27580 22778
rect 27528 22714 27580 22720
rect 27632 22658 27660 23054
rect 27264 22066 27476 22094
rect 27540 22630 27660 22658
rect 27160 21684 27212 21690
rect 27160 21626 27212 21632
rect 27068 21616 27120 21622
rect 27068 21558 27120 21564
rect 27068 21344 27120 21350
rect 27068 21286 27120 21292
rect 27080 20942 27108 21286
rect 27068 20936 27120 20942
rect 27068 20878 27120 20884
rect 26884 19304 26936 19310
rect 26988 19306 27108 19334
rect 26884 19246 26936 19252
rect 26882 19136 26938 19145
rect 26882 19071 26938 19080
rect 26792 15972 26844 15978
rect 26792 15914 26844 15920
rect 26896 15706 26924 19071
rect 26884 15700 26936 15706
rect 26884 15642 26936 15648
rect 26976 15564 27028 15570
rect 26976 15506 27028 15512
rect 26792 15496 26844 15502
rect 26792 15438 26844 15444
rect 26804 15162 26832 15438
rect 26884 15360 26936 15366
rect 26882 15328 26884 15337
rect 26936 15328 26938 15337
rect 26882 15263 26938 15272
rect 26882 15192 26938 15201
rect 26792 15156 26844 15162
rect 26882 15127 26938 15136
rect 26792 15098 26844 15104
rect 26896 14618 26924 15127
rect 26884 14612 26936 14618
rect 26884 14554 26936 14560
rect 26700 14340 26752 14346
rect 26700 14282 26752 14288
rect 26882 14240 26938 14249
rect 26712 14198 26882 14226
rect 26608 13796 26660 13802
rect 26608 13738 26660 13744
rect 26620 12986 26648 13738
rect 26608 12980 26660 12986
rect 26608 12922 26660 12928
rect 26712 12866 26740 14198
rect 26882 14175 26938 14184
rect 26988 14056 27016 15506
rect 27080 15162 27108 19306
rect 27172 17202 27200 21626
rect 27264 17354 27292 22066
rect 27344 22024 27396 22030
rect 27344 21966 27396 21972
rect 27356 21146 27384 21966
rect 27436 21956 27488 21962
rect 27436 21898 27488 21904
rect 27448 21690 27476 21898
rect 27436 21684 27488 21690
rect 27436 21626 27488 21632
rect 27540 21570 27568 22630
rect 27620 21956 27672 21962
rect 27724 21944 27752 23530
rect 27672 21916 27752 21944
rect 27620 21898 27672 21904
rect 27448 21542 27568 21570
rect 27344 21140 27396 21146
rect 27344 21082 27396 21088
rect 27448 20466 27476 21542
rect 27632 21185 27660 21898
rect 27816 21622 27844 25094
rect 27896 24200 27948 24206
rect 27896 24142 27948 24148
rect 27908 23118 27936 24142
rect 28000 23526 28028 25180
rect 28080 24812 28132 24818
rect 28080 24754 28132 24760
rect 28092 23905 28120 24754
rect 28184 24206 28212 26930
rect 28276 24732 28304 27814
rect 28540 27464 28592 27470
rect 28540 27406 28592 27412
rect 28552 26994 28580 27406
rect 28644 27130 28672 28591
rect 28736 27878 28764 28614
rect 28908 28552 28960 28558
rect 28908 28494 28960 28500
rect 28814 28248 28870 28257
rect 28814 28183 28870 28192
rect 28724 27872 28776 27878
rect 28724 27814 28776 27820
rect 28632 27124 28684 27130
rect 28632 27066 28684 27072
rect 28540 26988 28592 26994
rect 28540 26930 28592 26936
rect 28828 26586 28856 28183
rect 28920 28082 28948 28494
rect 29000 28484 29052 28490
rect 29000 28426 29052 28432
rect 28908 28076 28960 28082
rect 28908 28018 28960 28024
rect 29012 27713 29040 28426
rect 29104 28218 29132 28630
rect 29184 28552 29236 28558
rect 29182 28520 29184 28529
rect 29236 28520 29238 28529
rect 29182 28455 29238 28464
rect 29184 28416 29236 28422
rect 29184 28358 29236 28364
rect 29092 28212 29144 28218
rect 29092 28154 29144 28160
rect 29090 28112 29146 28121
rect 29196 28098 29224 28358
rect 29146 28070 29224 28098
rect 29288 28082 29316 31078
rect 29380 30258 29408 31198
rect 29460 31136 29512 31142
rect 29458 31104 29460 31113
rect 29512 31104 29514 31113
rect 29458 31039 29514 31048
rect 29458 30424 29514 30433
rect 29458 30359 29514 30368
rect 29472 30258 29500 30359
rect 29368 30252 29420 30258
rect 29368 30194 29420 30200
rect 29460 30252 29512 30258
rect 29460 30194 29512 30200
rect 29368 29640 29420 29646
rect 29368 29582 29420 29588
rect 29460 29640 29512 29646
rect 29460 29582 29512 29588
rect 29380 29345 29408 29582
rect 29366 29336 29422 29345
rect 29366 29271 29422 29280
rect 29472 28966 29500 29582
rect 29368 28960 29420 28966
rect 29368 28902 29420 28908
rect 29460 28960 29512 28966
rect 29460 28902 29512 28908
rect 29380 28626 29408 28902
rect 29472 28762 29500 28902
rect 29460 28756 29512 28762
rect 29460 28698 29512 28704
rect 29368 28620 29420 28626
rect 29368 28562 29420 28568
rect 29458 28248 29514 28257
rect 29458 28183 29514 28192
rect 29276 28076 29328 28082
rect 29090 28047 29146 28056
rect 29328 28036 29408 28064
rect 29276 28018 29328 28024
rect 29092 27940 29144 27946
rect 29092 27882 29144 27888
rect 28998 27704 29054 27713
rect 28998 27639 29054 27648
rect 29104 27062 29132 27882
rect 29184 27668 29236 27674
rect 29184 27610 29236 27616
rect 29092 27056 29144 27062
rect 29092 26998 29144 27004
rect 28816 26580 28868 26586
rect 28816 26522 28868 26528
rect 28908 26444 28960 26450
rect 28960 26404 29040 26432
rect 28908 26386 28960 26392
rect 28632 26308 28684 26314
rect 28632 26250 28684 26256
rect 28448 26240 28500 26246
rect 28448 26182 28500 26188
rect 28460 25906 28488 26182
rect 28644 26042 28672 26250
rect 28632 26036 28684 26042
rect 28632 25978 28684 25984
rect 28724 26036 28776 26042
rect 28724 25978 28776 25984
rect 28448 25900 28500 25906
rect 28448 25842 28500 25848
rect 28644 24818 28672 25978
rect 28736 25362 28764 25978
rect 28814 25664 28870 25673
rect 28814 25599 28870 25608
rect 28724 25356 28776 25362
rect 28724 25298 28776 25304
rect 28540 24812 28592 24818
rect 28540 24754 28592 24760
rect 28632 24812 28684 24818
rect 28632 24754 28684 24760
rect 28724 24812 28776 24818
rect 28724 24754 28776 24760
rect 28276 24704 28396 24732
rect 28264 24608 28316 24614
rect 28264 24550 28316 24556
rect 28276 24342 28304 24550
rect 28264 24336 28316 24342
rect 28264 24278 28316 24284
rect 28172 24200 28224 24206
rect 28172 24142 28224 24148
rect 28264 24200 28316 24206
rect 28264 24142 28316 24148
rect 28078 23896 28134 23905
rect 28184 23866 28212 24142
rect 28276 23866 28304 24142
rect 28368 24070 28396 24704
rect 28448 24676 28500 24682
rect 28448 24618 28500 24624
rect 28460 24313 28488 24618
rect 28552 24410 28580 24754
rect 28540 24404 28592 24410
rect 28540 24346 28592 24352
rect 28446 24304 28502 24313
rect 28736 24274 28764 24754
rect 28828 24410 28856 25599
rect 28908 25288 28960 25294
rect 28908 25230 28960 25236
rect 28920 24954 28948 25230
rect 28908 24948 28960 24954
rect 28908 24890 28960 24896
rect 28816 24404 28868 24410
rect 28816 24346 28868 24352
rect 28446 24239 28502 24248
rect 28724 24268 28776 24274
rect 28724 24210 28776 24216
rect 28448 24200 28500 24206
rect 28448 24142 28500 24148
rect 28356 24064 28408 24070
rect 28356 24006 28408 24012
rect 28078 23831 28134 23840
rect 28172 23860 28224 23866
rect 28092 23798 28120 23831
rect 28172 23802 28224 23808
rect 28264 23860 28316 23866
rect 28264 23802 28316 23808
rect 28460 23798 28488 24142
rect 28080 23792 28132 23798
rect 28080 23734 28132 23740
rect 28448 23792 28500 23798
rect 28448 23734 28500 23740
rect 27988 23520 28040 23526
rect 27988 23462 28040 23468
rect 27896 23112 27948 23118
rect 27896 23054 27948 23060
rect 28000 22094 28028 23462
rect 28092 22982 28120 23734
rect 28172 23724 28224 23730
rect 28172 23666 28224 23672
rect 28080 22976 28132 22982
rect 28080 22918 28132 22924
rect 27908 22066 28028 22094
rect 27804 21616 27856 21622
rect 27804 21558 27856 21564
rect 27712 21548 27764 21554
rect 27712 21490 27764 21496
rect 27618 21176 27674 21185
rect 27528 21140 27580 21146
rect 27618 21111 27674 21120
rect 27528 21082 27580 21088
rect 27436 20460 27488 20466
rect 27436 20402 27488 20408
rect 27342 19952 27398 19961
rect 27342 19887 27398 19896
rect 27356 19310 27384 19887
rect 27540 19786 27568 21082
rect 27620 20324 27672 20330
rect 27620 20266 27672 20272
rect 27632 19990 27660 20266
rect 27620 19984 27672 19990
rect 27620 19926 27672 19932
rect 27724 19836 27752 21490
rect 27804 21344 27856 21350
rect 27804 21286 27856 21292
rect 27816 20262 27844 21286
rect 27908 20369 27936 22066
rect 27988 22024 28040 22030
rect 27988 21966 28040 21972
rect 28000 21622 28028 21966
rect 28080 21888 28132 21894
rect 28080 21830 28132 21836
rect 27988 21616 28040 21622
rect 27988 21558 28040 21564
rect 28092 21554 28120 21830
rect 28080 21548 28132 21554
rect 28080 21490 28132 21496
rect 28184 21146 28212 23666
rect 28264 23656 28316 23662
rect 28264 23598 28316 23604
rect 28276 22642 28304 23598
rect 28356 23520 28408 23526
rect 28356 23462 28408 23468
rect 28538 23488 28594 23497
rect 28368 23118 28396 23462
rect 28538 23423 28594 23432
rect 28446 23352 28502 23361
rect 28446 23287 28502 23296
rect 28356 23112 28408 23118
rect 28356 23054 28408 23060
rect 28460 22710 28488 23287
rect 28552 23118 28580 23423
rect 28540 23112 28592 23118
rect 28540 23054 28592 23060
rect 28538 22944 28594 22953
rect 28538 22879 28594 22888
rect 28448 22704 28500 22710
rect 28448 22646 28500 22652
rect 28264 22636 28316 22642
rect 28264 22578 28316 22584
rect 28264 22024 28316 22030
rect 28264 21966 28316 21972
rect 28276 21486 28304 21966
rect 28264 21480 28316 21486
rect 28264 21422 28316 21428
rect 28460 21418 28488 22646
rect 28552 22030 28580 22879
rect 28736 22658 28764 24210
rect 28828 23798 28856 24346
rect 28816 23792 28868 23798
rect 28816 23734 28868 23740
rect 28920 23730 28948 24890
rect 29012 23730 29040 26404
rect 29092 24132 29144 24138
rect 29092 24074 29144 24080
rect 28908 23724 28960 23730
rect 28908 23666 28960 23672
rect 29000 23724 29052 23730
rect 29000 23666 29052 23672
rect 28632 22636 28684 22642
rect 28736 22630 28856 22658
rect 28632 22578 28684 22584
rect 28644 22409 28672 22578
rect 28724 22568 28776 22574
rect 28724 22510 28776 22516
rect 28630 22400 28686 22409
rect 28630 22335 28686 22344
rect 28540 22024 28592 22030
rect 28540 21966 28592 21972
rect 28632 22024 28684 22030
rect 28632 21966 28684 21972
rect 28644 21690 28672 21966
rect 28736 21962 28764 22510
rect 28724 21956 28776 21962
rect 28724 21898 28776 21904
rect 28632 21684 28684 21690
rect 28632 21626 28684 21632
rect 28540 21548 28592 21554
rect 28540 21490 28592 21496
rect 28448 21412 28500 21418
rect 28448 21354 28500 21360
rect 28172 21140 28224 21146
rect 28172 21082 28224 21088
rect 28354 21040 28410 21049
rect 27988 21004 28040 21010
rect 28354 20975 28410 20984
rect 27988 20946 28040 20952
rect 27894 20360 27950 20369
rect 27894 20295 27896 20304
rect 27948 20295 27950 20304
rect 27896 20266 27948 20272
rect 27804 20256 27856 20262
rect 27804 20198 27856 20204
rect 27632 19808 27752 19836
rect 27528 19780 27580 19786
rect 27528 19722 27580 19728
rect 27436 19712 27488 19718
rect 27436 19654 27488 19660
rect 27344 19304 27396 19310
rect 27344 19246 27396 19252
rect 27344 18624 27396 18630
rect 27344 18566 27396 18572
rect 27356 18426 27384 18566
rect 27344 18420 27396 18426
rect 27344 18362 27396 18368
rect 27264 17326 27384 17354
rect 27356 17202 27384 17326
rect 27160 17196 27212 17202
rect 27160 17138 27212 17144
rect 27344 17196 27396 17202
rect 27344 17138 27396 17144
rect 27252 17128 27304 17134
rect 27252 17070 27304 17076
rect 27264 15502 27292 17070
rect 27356 16454 27384 17138
rect 27448 16980 27476 19654
rect 27540 19281 27568 19722
rect 27526 19272 27582 19281
rect 27526 19207 27582 19216
rect 27528 17604 27580 17610
rect 27528 17546 27580 17552
rect 27540 17338 27568 17546
rect 27528 17332 27580 17338
rect 27528 17274 27580 17280
rect 27632 17082 27660 19808
rect 27712 19712 27764 19718
rect 27710 19680 27712 19689
rect 27764 19680 27766 19689
rect 27710 19615 27766 19624
rect 27710 19544 27766 19553
rect 27710 19479 27712 19488
rect 27764 19479 27766 19488
rect 27712 19450 27764 19456
rect 27710 19408 27766 19417
rect 27710 19343 27712 19352
rect 27764 19343 27766 19352
rect 27712 19314 27764 19320
rect 27712 19168 27764 19174
rect 27712 19110 27764 19116
rect 27724 17746 27752 19110
rect 27712 17740 27764 17746
rect 27712 17682 27764 17688
rect 27816 17678 27844 20198
rect 27894 20088 27950 20097
rect 27894 20023 27950 20032
rect 27908 19514 27936 20023
rect 27896 19508 27948 19514
rect 27896 19450 27948 19456
rect 27896 19372 27948 19378
rect 27896 19314 27948 19320
rect 27908 18290 27936 19314
rect 27896 18284 27948 18290
rect 27896 18226 27948 18232
rect 27804 17672 27856 17678
rect 27804 17614 27856 17620
rect 27908 17270 27936 18226
rect 27896 17264 27948 17270
rect 27896 17206 27948 17212
rect 27632 17054 27752 17082
rect 27528 16992 27580 16998
rect 27448 16952 27528 16980
rect 27528 16934 27580 16940
rect 27620 16992 27672 16998
rect 27620 16934 27672 16940
rect 27344 16448 27396 16454
rect 27344 16390 27396 16396
rect 27252 15496 27304 15502
rect 27252 15438 27304 15444
rect 27068 15156 27120 15162
rect 27068 15098 27120 15104
rect 27080 14618 27108 15098
rect 27160 14884 27212 14890
rect 27160 14826 27212 14832
rect 27068 14612 27120 14618
rect 27068 14554 27120 14560
rect 26896 14028 27016 14056
rect 26792 13796 26844 13802
rect 26792 13738 26844 13744
rect 26804 13462 26832 13738
rect 26792 13456 26844 13462
rect 26792 13398 26844 13404
rect 26620 12838 26740 12866
rect 26620 12442 26648 12838
rect 26700 12776 26752 12782
rect 26700 12718 26752 12724
rect 26608 12436 26660 12442
rect 26608 12378 26660 12384
rect 26514 12336 26570 12345
rect 26514 12271 26570 12280
rect 25872 12232 25924 12238
rect 25872 12174 25924 12180
rect 26332 12232 26384 12238
rect 26332 12174 26384 12180
rect 26608 12232 26660 12238
rect 26608 12174 26660 12180
rect 25780 11892 25832 11898
rect 25780 11834 25832 11840
rect 25596 11824 25648 11830
rect 25884 11778 25912 12174
rect 26056 12164 26108 12170
rect 26056 12106 26108 12112
rect 25596 11766 25648 11772
rect 25792 11750 25912 11778
rect 25136 11008 25188 11014
rect 25136 10950 25188 10956
rect 23572 10600 23624 10606
rect 23572 10542 23624 10548
rect 23388 10192 23440 10198
rect 23388 10134 23440 10140
rect 22612 10024 22692 10044
rect 22614 10016 22692 10024
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 22558 9959 22614 9968
rect 23124 9722 23152 9998
rect 23112 9716 23164 9722
rect 23112 9658 23164 9664
rect 22560 9512 22612 9518
rect 22480 9472 22560 9500
rect 22560 9454 22612 9460
rect 22100 9036 22152 9042
rect 22100 8978 22152 8984
rect 22572 8906 22600 9454
rect 21916 8900 21968 8906
rect 21916 8842 21968 8848
rect 22100 8900 22152 8906
rect 22100 8842 22152 8848
rect 22560 8900 22612 8906
rect 22560 8842 22612 8848
rect 21088 8832 21140 8838
rect 21088 8774 21140 8780
rect 20812 8084 20864 8090
rect 20812 8026 20864 8032
rect 20720 7812 20772 7818
rect 20720 7754 20772 7760
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20260 6112 20312 6118
rect 20260 6054 20312 6060
rect 20272 5914 20300 6054
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20732 5710 20760 7754
rect 20824 7410 20852 8026
rect 21824 7948 21876 7954
rect 21824 7890 21876 7896
rect 20904 7744 20956 7750
rect 20904 7686 20956 7692
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20810 7304 20866 7313
rect 20810 7239 20866 7248
rect 20824 6254 20852 7239
rect 20916 6866 20944 7686
rect 21836 6866 21864 7890
rect 21916 7812 21968 7818
rect 21916 7754 21968 7760
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 21824 6860 21876 6866
rect 21824 6802 21876 6808
rect 21088 6792 21140 6798
rect 21088 6734 21140 6740
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 20824 5914 20852 6190
rect 21100 6118 21128 6734
rect 20996 6112 21048 6118
rect 20996 6054 21048 6060
rect 21088 6112 21140 6118
rect 21088 6054 21140 6060
rect 21008 5914 21036 6054
rect 21100 5914 21128 6054
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 20996 5908 21048 5914
rect 20996 5850 21048 5856
rect 21088 5908 21140 5914
rect 21088 5850 21140 5856
rect 21836 5778 21864 6802
rect 21928 5778 21956 7754
rect 22112 7410 22140 8842
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22572 6730 22600 8842
rect 23400 7886 23428 10134
rect 23584 10062 23612 10542
rect 23756 10464 23808 10470
rect 23756 10406 23808 10412
rect 23848 10464 23900 10470
rect 25136 10464 25188 10470
rect 23848 10406 23900 10412
rect 24490 10432 24546 10441
rect 23572 10056 23624 10062
rect 23572 9998 23624 10004
rect 23768 9042 23796 10406
rect 23860 10266 23888 10406
rect 25136 10406 25188 10412
rect 24490 10367 24546 10376
rect 24504 10266 24532 10367
rect 23848 10260 23900 10266
rect 23848 10202 23900 10208
rect 24492 10260 24544 10266
rect 24492 10202 24544 10208
rect 25148 9994 25176 10406
rect 25228 10124 25280 10130
rect 25228 10066 25280 10072
rect 24952 9988 25004 9994
rect 24952 9930 25004 9936
rect 25136 9988 25188 9994
rect 25136 9930 25188 9936
rect 24124 9920 24176 9926
rect 24124 9862 24176 9868
rect 24136 9518 24164 9862
rect 24860 9716 24912 9722
rect 24860 9658 24912 9664
rect 24124 9512 24176 9518
rect 24124 9454 24176 9460
rect 24216 9512 24268 9518
rect 24216 9454 24268 9460
rect 24492 9512 24544 9518
rect 24492 9454 24544 9460
rect 23756 9036 23808 9042
rect 23756 8978 23808 8984
rect 23572 8016 23624 8022
rect 23572 7958 23624 7964
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 23584 7750 23612 7958
rect 24228 7954 24256 9454
rect 24504 9178 24532 9454
rect 24492 9172 24544 9178
rect 24492 9114 24544 9120
rect 24216 7948 24268 7954
rect 24136 7908 24216 7936
rect 23572 7744 23624 7750
rect 23572 7686 23624 7692
rect 23584 7546 23612 7686
rect 24136 7546 24164 7908
rect 24216 7890 24268 7896
rect 24872 7800 24900 9658
rect 24964 9518 24992 9930
rect 25148 9722 25176 9930
rect 25136 9716 25188 9722
rect 25136 9658 25188 9664
rect 24952 9512 25004 9518
rect 24952 9454 25004 9460
rect 25240 9042 25268 10066
rect 25228 9036 25280 9042
rect 25228 8978 25280 8984
rect 24952 7812 25004 7818
rect 24872 7772 24952 7800
rect 23572 7540 23624 7546
rect 23572 7482 23624 7488
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 24872 7410 24900 7772
rect 24952 7754 25004 7760
rect 25792 7546 25820 11750
rect 25964 11688 26016 11694
rect 25964 11630 26016 11636
rect 25872 11552 25924 11558
rect 25872 11494 25924 11500
rect 25884 11218 25912 11494
rect 25872 11212 25924 11218
rect 25872 11154 25924 11160
rect 25976 11082 26004 11630
rect 26068 11354 26096 12106
rect 26056 11348 26108 11354
rect 26056 11290 26108 11296
rect 25964 11076 26016 11082
rect 25964 11018 26016 11024
rect 25976 9722 26004 11018
rect 26240 10668 26292 10674
rect 26240 10610 26292 10616
rect 26252 10266 26280 10610
rect 26240 10260 26292 10266
rect 26240 10202 26292 10208
rect 26344 10146 26372 12174
rect 26516 12096 26568 12102
rect 26516 12038 26568 12044
rect 26424 11756 26476 11762
rect 26424 11698 26476 11704
rect 26436 10470 26464 11698
rect 26528 11694 26556 12038
rect 26620 11830 26648 12174
rect 26608 11824 26660 11830
rect 26608 11766 26660 11772
rect 26712 11762 26740 12718
rect 26804 11898 26832 13398
rect 26896 12442 26924 14028
rect 27066 13968 27122 13977
rect 26976 13932 27028 13938
rect 27066 13903 27068 13912
rect 26976 13874 27028 13880
rect 27120 13903 27122 13912
rect 27068 13874 27120 13880
rect 26988 13530 27016 13874
rect 26976 13524 27028 13530
rect 26976 13466 27028 13472
rect 27080 13258 27108 13874
rect 27068 13252 27120 13258
rect 27068 13194 27120 13200
rect 26884 12436 26936 12442
rect 26884 12378 26936 12384
rect 26976 12232 27028 12238
rect 26976 12174 27028 12180
rect 27068 12232 27120 12238
rect 27068 12174 27120 12180
rect 26792 11892 26844 11898
rect 26792 11834 26844 11840
rect 26884 11892 26936 11898
rect 26988 11880 27016 12174
rect 27080 12102 27108 12174
rect 27068 12096 27120 12102
rect 27068 12038 27120 12044
rect 26936 11852 27016 11880
rect 26884 11834 26936 11840
rect 26700 11756 26752 11762
rect 26700 11698 26752 11704
rect 26516 11688 26568 11694
rect 26516 11630 26568 11636
rect 26792 11688 26844 11694
rect 26792 11630 26844 11636
rect 26424 10464 26476 10470
rect 26424 10406 26476 10412
rect 26252 10118 26372 10146
rect 25964 9716 26016 9722
rect 25964 9658 26016 9664
rect 26056 9580 26108 9586
rect 26056 9522 26108 9528
rect 26068 7818 26096 9522
rect 26056 7812 26108 7818
rect 26056 7754 26108 7760
rect 25780 7540 25832 7546
rect 25780 7482 25832 7488
rect 26068 7460 26096 7754
rect 26148 7472 26200 7478
rect 26068 7432 26148 7460
rect 26148 7414 26200 7420
rect 24860 7404 24912 7410
rect 24860 7346 24912 7352
rect 25228 7404 25280 7410
rect 25228 7346 25280 7352
rect 24492 6792 24544 6798
rect 24492 6734 24544 6740
rect 22560 6724 22612 6730
rect 22560 6666 22612 6672
rect 23848 6724 23900 6730
rect 23848 6666 23900 6672
rect 22376 6656 22428 6662
rect 22376 6598 22428 6604
rect 22388 6390 22416 6598
rect 22376 6384 22428 6390
rect 22376 6326 22428 6332
rect 22284 6316 22336 6322
rect 22284 6258 22336 6264
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 22020 5914 22048 6054
rect 22008 5908 22060 5914
rect 22008 5850 22060 5856
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 21824 5772 21876 5778
rect 21824 5714 21876 5720
rect 21916 5772 21968 5778
rect 21916 5714 21968 5720
rect 20720 5704 20772 5710
rect 20720 5646 20772 5652
rect 20732 5556 20760 5646
rect 20640 5528 20760 5556
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 20640 5302 20668 5528
rect 20628 5296 20680 5302
rect 20628 5238 20680 5244
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 20640 2514 20668 4966
rect 20628 2508 20680 2514
rect 20628 2450 20680 2456
rect 22112 2446 22140 5850
rect 22296 5234 22324 6258
rect 22572 5710 22600 6666
rect 23860 6390 23888 6666
rect 23848 6384 23900 6390
rect 23848 6326 23900 6332
rect 24504 6322 24532 6734
rect 25240 6390 25268 7346
rect 26056 6860 26108 6866
rect 26056 6802 26108 6808
rect 25780 6724 25832 6730
rect 25780 6666 25832 6672
rect 25228 6384 25280 6390
rect 25228 6326 25280 6332
rect 24492 6316 24544 6322
rect 24492 6258 24544 6264
rect 22560 5704 22612 5710
rect 22560 5646 22612 5652
rect 23204 5636 23256 5642
rect 23204 5578 23256 5584
rect 22468 5568 22520 5574
rect 22468 5510 22520 5516
rect 22480 5370 22508 5510
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 23216 5166 23244 5578
rect 23204 5160 23256 5166
rect 23204 5102 23256 5108
rect 23216 3466 23244 5102
rect 23204 3460 23256 3466
rect 23204 3402 23256 3408
rect 22100 2440 22152 2446
rect 21928 2366 22048 2394
rect 22100 2382 22152 2388
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 21928 800 21956 2366
rect 22020 2310 22048 2366
rect 22008 2304 22060 2310
rect 22008 2246 22060 2252
rect 25792 800 25820 6666
rect 26068 5574 26096 6802
rect 26252 6730 26280 10118
rect 26436 10044 26464 10406
rect 26528 10266 26556 11630
rect 26804 11354 26832 11630
rect 27172 11558 27200 14826
rect 27264 13841 27292 15438
rect 27344 14884 27396 14890
rect 27344 14826 27396 14832
rect 27356 14074 27384 14826
rect 27434 14648 27490 14657
rect 27434 14583 27436 14592
rect 27488 14583 27490 14592
rect 27436 14554 27488 14560
rect 27436 14272 27488 14278
rect 27436 14214 27488 14220
rect 27344 14068 27396 14074
rect 27344 14010 27396 14016
rect 27250 13832 27306 13841
rect 27250 13767 27306 13776
rect 27250 13696 27306 13705
rect 27250 13631 27306 13640
rect 27264 13258 27292 13631
rect 27448 13569 27476 14214
rect 27540 13716 27568 16934
rect 27632 16726 27660 16934
rect 27620 16720 27672 16726
rect 27620 16662 27672 16668
rect 27620 14884 27672 14890
rect 27724 14872 27752 17054
rect 27804 16448 27856 16454
rect 27804 16390 27856 16396
rect 27672 14844 27752 14872
rect 27620 14826 27672 14832
rect 27632 13954 27660 14826
rect 27816 14498 27844 16390
rect 27894 15192 27950 15201
rect 27894 15127 27950 15136
rect 27908 15026 27936 15127
rect 27896 15020 27948 15026
rect 27896 14962 27948 14968
rect 27908 14618 27936 14962
rect 27896 14612 27948 14618
rect 27896 14554 27948 14560
rect 27816 14482 27936 14498
rect 27816 14476 27948 14482
rect 27816 14470 27896 14476
rect 27896 14418 27948 14424
rect 27712 14408 27764 14414
rect 27712 14350 27764 14356
rect 27802 14376 27858 14385
rect 27724 14074 27752 14350
rect 27802 14311 27804 14320
rect 27856 14311 27858 14320
rect 27804 14282 27856 14288
rect 27802 14240 27858 14249
rect 27802 14175 27858 14184
rect 27816 14074 27844 14175
rect 27712 14068 27764 14074
rect 27712 14010 27764 14016
rect 27804 14068 27856 14074
rect 27804 14010 27856 14016
rect 27632 13926 27844 13954
rect 27620 13864 27672 13870
rect 27618 13832 27620 13841
rect 27712 13864 27764 13870
rect 27672 13832 27674 13841
rect 27712 13806 27764 13812
rect 27618 13767 27674 13776
rect 27540 13688 27660 13716
rect 27434 13560 27490 13569
rect 27434 13495 27490 13504
rect 27436 13320 27488 13326
rect 27436 13262 27488 13268
rect 27252 13252 27304 13258
rect 27252 13194 27304 13200
rect 27448 12434 27476 13262
rect 27528 13252 27580 13258
rect 27528 13194 27580 13200
rect 27264 12406 27476 12434
rect 27540 12434 27568 13194
rect 27632 12782 27660 13688
rect 27724 13530 27752 13806
rect 27712 13524 27764 13530
rect 27712 13466 27764 13472
rect 27712 12844 27764 12850
rect 27712 12786 27764 12792
rect 27620 12776 27672 12782
rect 27620 12718 27672 12724
rect 27540 12406 27660 12434
rect 27264 11762 27292 12406
rect 27526 12336 27582 12345
rect 27526 12271 27582 12280
rect 27540 12238 27568 12271
rect 27632 12238 27660 12406
rect 27724 12238 27752 12786
rect 27528 12232 27580 12238
rect 27528 12174 27580 12180
rect 27620 12232 27672 12238
rect 27620 12174 27672 12180
rect 27712 12232 27764 12238
rect 27712 12174 27764 12180
rect 27252 11756 27304 11762
rect 27252 11698 27304 11704
rect 27344 11756 27396 11762
rect 27344 11698 27396 11704
rect 27160 11552 27212 11558
rect 27160 11494 27212 11500
rect 26792 11348 26844 11354
rect 26792 11290 26844 11296
rect 26700 11076 26752 11082
rect 26700 11018 26752 11024
rect 26712 10674 26740 11018
rect 26700 10668 26752 10674
rect 26700 10610 26752 10616
rect 26516 10260 26568 10266
rect 26516 10202 26568 10208
rect 26804 10062 26832 11290
rect 27172 11082 27200 11494
rect 27160 11076 27212 11082
rect 27160 11018 27212 11024
rect 26976 10260 27028 10266
rect 26976 10202 27028 10208
rect 26344 10016 26464 10044
rect 26792 10056 26844 10062
rect 26344 9654 26372 10016
rect 26792 9998 26844 10004
rect 26424 9920 26476 9926
rect 26424 9862 26476 9868
rect 26332 9648 26384 9654
rect 26332 9590 26384 9596
rect 26436 9178 26464 9862
rect 26424 9172 26476 9178
rect 26424 9114 26476 9120
rect 26988 8430 27016 10202
rect 27068 10124 27120 10130
rect 27068 10066 27120 10072
rect 27080 9926 27108 10066
rect 27068 9920 27120 9926
rect 27068 9862 27120 9868
rect 27160 9580 27212 9586
rect 27160 9522 27212 9528
rect 27252 9580 27304 9586
rect 27252 9522 27304 9528
rect 27172 8634 27200 9522
rect 27264 8838 27292 9522
rect 27356 9450 27384 11698
rect 27540 11354 27568 12174
rect 27632 11558 27660 12174
rect 27620 11552 27672 11558
rect 27620 11494 27672 11500
rect 27528 11348 27580 11354
rect 27528 11290 27580 11296
rect 27434 10976 27490 10985
rect 27434 10911 27490 10920
rect 27448 10674 27476 10911
rect 27436 10668 27488 10674
rect 27436 10610 27488 10616
rect 27436 10260 27488 10266
rect 27436 10202 27488 10208
rect 27344 9444 27396 9450
rect 27344 9386 27396 9392
rect 27344 8900 27396 8906
rect 27448 8888 27476 10202
rect 27618 10160 27674 10169
rect 27618 10095 27674 10104
rect 27632 10062 27660 10095
rect 27620 10056 27672 10062
rect 27620 9998 27672 10004
rect 27528 9512 27580 9518
rect 27528 9454 27580 9460
rect 27396 8860 27476 8888
rect 27344 8842 27396 8848
rect 27252 8832 27304 8838
rect 27252 8774 27304 8780
rect 27160 8628 27212 8634
rect 27160 8570 27212 8576
rect 27264 8566 27292 8774
rect 27252 8560 27304 8566
rect 27252 8502 27304 8508
rect 26976 8424 27028 8430
rect 26976 8366 27028 8372
rect 26988 8090 27016 8366
rect 26976 8084 27028 8090
rect 26976 8026 27028 8032
rect 27160 7812 27212 7818
rect 27160 7754 27212 7760
rect 27172 7478 27200 7754
rect 27160 7472 27212 7478
rect 27160 7414 27212 7420
rect 26792 7336 26844 7342
rect 26792 7278 26844 7284
rect 26804 6866 26832 7278
rect 27252 7200 27304 7206
rect 27252 7142 27304 7148
rect 26792 6860 26844 6866
rect 26792 6802 26844 6808
rect 26240 6724 26292 6730
rect 26240 6666 26292 6672
rect 26252 6458 26280 6666
rect 26700 6656 26752 6662
rect 26700 6598 26752 6604
rect 26712 6458 26740 6598
rect 26240 6452 26292 6458
rect 26240 6394 26292 6400
rect 26700 6452 26752 6458
rect 26700 6394 26752 6400
rect 26056 5568 26108 5574
rect 26056 5510 26108 5516
rect 26068 4690 26096 5510
rect 27264 5234 27292 7142
rect 27356 6746 27384 8842
rect 27436 8288 27488 8294
rect 27434 8256 27436 8265
rect 27488 8256 27490 8265
rect 27434 8191 27490 8200
rect 27436 7404 27488 7410
rect 27540 7392 27568 9454
rect 27620 9376 27672 9382
rect 27620 9318 27672 9324
rect 27632 9178 27660 9318
rect 27620 9172 27672 9178
rect 27620 9114 27672 9120
rect 27724 9058 27752 12174
rect 27632 9030 27752 9058
rect 27632 7410 27660 9030
rect 27712 8288 27764 8294
rect 27712 8230 27764 8236
rect 27724 8022 27752 8230
rect 27712 8016 27764 8022
rect 27712 7958 27764 7964
rect 27488 7364 27568 7392
rect 27620 7404 27672 7410
rect 27436 7346 27488 7352
rect 27620 7346 27672 7352
rect 27448 6882 27476 7346
rect 27528 7200 27580 7206
rect 27528 7142 27580 7148
rect 27540 7002 27568 7142
rect 27632 7002 27660 7346
rect 27528 6996 27580 7002
rect 27528 6938 27580 6944
rect 27620 6996 27672 7002
rect 27620 6938 27672 6944
rect 27712 6928 27764 6934
rect 27448 6854 27568 6882
rect 27712 6870 27764 6876
rect 27436 6792 27488 6798
rect 27356 6740 27436 6746
rect 27356 6734 27488 6740
rect 27356 6718 27476 6734
rect 27252 5228 27304 5234
rect 27252 5170 27304 5176
rect 26976 5024 27028 5030
rect 26976 4966 27028 4972
rect 26988 4690 27016 4966
rect 26056 4684 26108 4690
rect 26056 4626 26108 4632
rect 26976 4684 27028 4690
rect 26976 4626 27028 4632
rect 27448 4622 27476 6718
rect 27540 6322 27568 6854
rect 27528 6316 27580 6322
rect 27528 6258 27580 6264
rect 27540 5846 27568 6258
rect 27528 5840 27580 5846
rect 27528 5782 27580 5788
rect 27724 5658 27752 6870
rect 27816 5914 27844 13926
rect 27908 13326 27936 14418
rect 28000 14056 28028 20946
rect 28368 20534 28396 20975
rect 28172 20528 28224 20534
rect 28092 20488 28172 20516
rect 28092 19310 28120 20488
rect 28172 20470 28224 20476
rect 28356 20528 28408 20534
rect 28356 20470 28408 20476
rect 28448 20324 28500 20330
rect 28448 20266 28500 20272
rect 28172 20052 28224 20058
rect 28172 19994 28224 20000
rect 28184 19446 28212 19994
rect 28460 19854 28488 20266
rect 28448 19848 28500 19854
rect 28448 19790 28500 19796
rect 28356 19712 28408 19718
rect 28356 19654 28408 19660
rect 28172 19440 28224 19446
rect 28172 19382 28224 19388
rect 28080 19304 28132 19310
rect 28080 19246 28132 19252
rect 28092 17202 28120 19246
rect 28262 17776 28318 17785
rect 28262 17711 28318 17720
rect 28276 17678 28304 17711
rect 28264 17672 28316 17678
rect 28264 17614 28316 17620
rect 28080 17196 28132 17202
rect 28080 17138 28132 17144
rect 28092 17105 28120 17138
rect 28172 17128 28224 17134
rect 28078 17096 28134 17105
rect 28172 17070 28224 17076
rect 28078 17031 28134 17040
rect 28184 14278 28212 17070
rect 28368 16182 28396 19654
rect 28356 16176 28408 16182
rect 28356 16118 28408 16124
rect 28460 16130 28488 19790
rect 28552 19417 28580 21490
rect 28828 19854 28856 22630
rect 28998 22536 29054 22545
rect 29104 22522 29132 24074
rect 29196 22642 29224 27610
rect 29276 26784 29328 26790
rect 29276 26726 29328 26732
rect 29288 26450 29316 26726
rect 29380 26586 29408 28036
rect 29472 27441 29500 28183
rect 29458 27432 29514 27441
rect 29458 27367 29514 27376
rect 29460 26784 29512 26790
rect 29460 26726 29512 26732
rect 29368 26580 29420 26586
rect 29368 26522 29420 26528
rect 29276 26444 29328 26450
rect 29276 26386 29328 26392
rect 29472 26353 29500 26726
rect 29458 26344 29514 26353
rect 29368 26308 29420 26314
rect 29458 26279 29514 26288
rect 29368 26250 29420 26256
rect 29276 26240 29328 26246
rect 29276 26182 29328 26188
rect 29288 24177 29316 26182
rect 29380 25906 29408 26250
rect 29368 25900 29420 25906
rect 29368 25842 29420 25848
rect 29460 24200 29512 24206
rect 29274 24168 29330 24177
rect 29274 24103 29330 24112
rect 29458 24168 29460 24177
rect 29512 24168 29514 24177
rect 29458 24103 29514 24112
rect 29184 22636 29236 22642
rect 29184 22578 29236 22584
rect 29054 22494 29132 22522
rect 28998 22471 29054 22480
rect 29092 22228 29144 22234
rect 29092 22170 29144 22176
rect 29104 21962 29132 22170
rect 29092 21956 29144 21962
rect 29092 21898 29144 21904
rect 29196 21690 29224 22578
rect 29288 22234 29316 24103
rect 29368 23724 29420 23730
rect 29368 23666 29420 23672
rect 29460 23724 29512 23730
rect 29460 23666 29512 23672
rect 29276 22228 29328 22234
rect 29276 22170 29328 22176
rect 29276 22092 29328 22098
rect 29276 22034 29328 22040
rect 29184 21684 29236 21690
rect 29184 21626 29236 21632
rect 29288 21570 29316 22034
rect 29196 21542 29316 21570
rect 28908 21344 28960 21350
rect 28908 21286 28960 21292
rect 28920 20058 28948 21286
rect 29000 20256 29052 20262
rect 29000 20198 29052 20204
rect 28908 20052 28960 20058
rect 28908 19994 28960 20000
rect 29012 19990 29040 20198
rect 29000 19984 29052 19990
rect 28998 19952 29000 19961
rect 29052 19952 29054 19961
rect 28998 19887 29054 19896
rect 28816 19848 28868 19854
rect 29196 19802 29224 21542
rect 29276 20256 29328 20262
rect 29276 20198 29328 20204
rect 28816 19790 28868 19796
rect 28538 19408 28594 19417
rect 28538 19343 28594 19352
rect 28828 19334 28856 19790
rect 28736 19306 28856 19334
rect 29012 19774 29224 19802
rect 29288 19786 29316 20198
rect 29380 19854 29408 23666
rect 29472 23254 29500 23666
rect 29460 23248 29512 23254
rect 29460 23190 29512 23196
rect 29460 22568 29512 22574
rect 29460 22510 29512 22516
rect 29472 22234 29500 22510
rect 29460 22228 29512 22234
rect 29460 22170 29512 22176
rect 29564 22166 29592 31214
rect 29656 30258 29684 31826
rect 29736 31476 29788 31482
rect 29736 31418 29788 31424
rect 29748 30938 29776 31418
rect 29736 30932 29788 30938
rect 29736 30874 29788 30880
rect 29840 30734 29868 34496
rect 30300 34406 30328 35634
rect 31116 35556 31168 35562
rect 31116 35498 31168 35504
rect 30472 35488 30524 35494
rect 30472 35430 30524 35436
rect 31024 35488 31076 35494
rect 31024 35430 31076 35436
rect 30484 34746 30512 35430
rect 31036 35290 31064 35430
rect 31128 35290 31156 35498
rect 31392 35488 31444 35494
rect 31392 35430 31444 35436
rect 31024 35284 31076 35290
rect 31024 35226 31076 35232
rect 31116 35284 31168 35290
rect 31116 35226 31168 35232
rect 31404 35193 31432 35430
rect 31390 35184 31446 35193
rect 31024 35148 31076 35154
rect 31390 35119 31446 35128
rect 31024 35090 31076 35096
rect 30472 34740 30524 34746
rect 30472 34682 30524 34688
rect 30564 34468 30616 34474
rect 30564 34410 30616 34416
rect 30288 34400 30340 34406
rect 30288 34342 30340 34348
rect 30288 34060 30340 34066
rect 30288 34002 30340 34008
rect 30012 33992 30064 33998
rect 30012 33934 30064 33940
rect 30024 33658 30052 33934
rect 30012 33652 30064 33658
rect 30012 33594 30064 33600
rect 30300 33454 30328 34002
rect 30576 33998 30604 34410
rect 30654 34096 30710 34105
rect 30654 34031 30710 34040
rect 30668 33998 30696 34031
rect 30564 33992 30616 33998
rect 30564 33934 30616 33940
rect 30656 33992 30708 33998
rect 30656 33934 30708 33940
rect 30472 33856 30524 33862
rect 30472 33798 30524 33804
rect 30484 33522 30512 33798
rect 30472 33516 30524 33522
rect 30472 33458 30524 33464
rect 30288 33448 30340 33454
rect 30288 33390 30340 33396
rect 30288 33040 30340 33046
rect 30288 32982 30340 32988
rect 30300 32434 30328 32982
rect 30380 32904 30432 32910
rect 30380 32846 30432 32852
rect 30392 32434 30420 32846
rect 30288 32428 30340 32434
rect 30288 32370 30340 32376
rect 30380 32428 30432 32434
rect 30380 32370 30432 32376
rect 29920 32360 29972 32366
rect 29920 32302 29972 32308
rect 29828 30728 29880 30734
rect 29828 30670 29880 30676
rect 29644 30252 29696 30258
rect 29644 30194 29696 30200
rect 29736 29776 29788 29782
rect 29736 29718 29788 29724
rect 29748 29170 29776 29718
rect 29840 29510 29868 30670
rect 29828 29504 29880 29510
rect 29828 29446 29880 29452
rect 29826 29336 29882 29345
rect 29826 29271 29882 29280
rect 29840 29170 29868 29271
rect 29736 29164 29788 29170
rect 29736 29106 29788 29112
rect 29828 29164 29880 29170
rect 29828 29106 29880 29112
rect 29840 29073 29868 29106
rect 29826 29064 29882 29073
rect 29736 29028 29788 29034
rect 29826 28999 29882 29008
rect 29736 28970 29788 28976
rect 29644 28484 29696 28490
rect 29644 28426 29696 28432
rect 29656 27538 29684 28426
rect 29644 27532 29696 27538
rect 29644 27474 29696 27480
rect 29644 26444 29696 26450
rect 29644 26386 29696 26392
rect 29656 25498 29684 26386
rect 29644 25492 29696 25498
rect 29644 25434 29696 25440
rect 29644 25288 29696 25294
rect 29644 25230 29696 25236
rect 29656 24886 29684 25230
rect 29644 24880 29696 24886
rect 29644 24822 29696 24828
rect 29644 24608 29696 24614
rect 29644 24550 29696 24556
rect 29656 24410 29684 24550
rect 29644 24404 29696 24410
rect 29644 24346 29696 24352
rect 29748 24206 29776 28970
rect 29828 28960 29880 28966
rect 29828 28902 29880 28908
rect 29840 28558 29868 28902
rect 29828 28552 29880 28558
rect 29828 28494 29880 28500
rect 29828 26920 29880 26926
rect 29828 26862 29880 26868
rect 29736 24200 29788 24206
rect 29736 24142 29788 24148
rect 29644 23724 29696 23730
rect 29644 23666 29696 23672
rect 29656 22642 29684 23666
rect 29748 23526 29776 24142
rect 29736 23520 29788 23526
rect 29736 23462 29788 23468
rect 29644 22636 29696 22642
rect 29748 22624 29776 23462
rect 29840 23254 29868 26862
rect 29932 26024 29960 32302
rect 30196 32224 30248 32230
rect 30196 32166 30248 32172
rect 30012 31952 30064 31958
rect 30012 31894 30064 31900
rect 30024 30054 30052 31894
rect 30104 31136 30156 31142
rect 30104 31078 30156 31084
rect 30116 30394 30144 31078
rect 30104 30388 30156 30394
rect 30104 30330 30156 30336
rect 30012 30048 30064 30054
rect 30012 29990 30064 29996
rect 30024 29714 30052 29990
rect 30012 29708 30064 29714
rect 30012 29650 30064 29656
rect 30024 28994 30052 29650
rect 30024 28966 30144 28994
rect 30012 28756 30064 28762
rect 30012 28698 30064 28704
rect 30024 26738 30052 28698
rect 30116 27674 30144 28966
rect 30104 27668 30156 27674
rect 30104 27610 30156 27616
rect 30024 26710 30144 26738
rect 30010 26616 30066 26625
rect 30010 26551 30012 26560
rect 30064 26551 30066 26560
rect 30012 26522 30064 26528
rect 29932 25996 30052 26024
rect 29920 25900 29972 25906
rect 29920 25842 29972 25848
rect 29932 25498 29960 25842
rect 29920 25492 29972 25498
rect 29920 25434 29972 25440
rect 30024 25378 30052 25996
rect 29932 25350 30052 25378
rect 29932 25294 29960 25350
rect 29920 25288 29972 25294
rect 29920 25230 29972 25236
rect 30012 25288 30064 25294
rect 30012 25230 30064 25236
rect 29932 24070 29960 25230
rect 30024 25129 30052 25230
rect 30010 25120 30066 25129
rect 30010 25055 30066 25064
rect 30012 24880 30064 24886
rect 30012 24822 30064 24828
rect 30024 24410 30052 24822
rect 30012 24404 30064 24410
rect 30012 24346 30064 24352
rect 30024 24313 30052 24346
rect 30010 24304 30066 24313
rect 30010 24239 30066 24248
rect 30116 24206 30144 26710
rect 30208 25906 30236 32166
rect 30288 31884 30340 31890
rect 30288 31826 30340 31832
rect 30300 30977 30328 31826
rect 30380 31816 30432 31822
rect 30484 31793 30512 33458
rect 30576 33318 30604 33934
rect 30564 33312 30616 33318
rect 30564 33254 30616 33260
rect 30656 32904 30708 32910
rect 30656 32846 30708 32852
rect 30668 32502 30696 32846
rect 30840 32768 30892 32774
rect 30840 32710 30892 32716
rect 30656 32496 30708 32502
rect 30656 32438 30708 32444
rect 30668 32201 30696 32438
rect 30748 32224 30800 32230
rect 30654 32192 30710 32201
rect 30748 32166 30800 32172
rect 30654 32127 30710 32136
rect 30380 31758 30432 31764
rect 30470 31784 30526 31793
rect 30286 30968 30342 30977
rect 30286 30903 30342 30912
rect 30288 30184 30340 30190
rect 30288 30126 30340 30132
rect 30300 29782 30328 30126
rect 30288 29776 30340 29782
rect 30288 29718 30340 29724
rect 30392 29646 30420 31758
rect 30470 31719 30526 31728
rect 30564 31748 30616 31754
rect 30564 31690 30616 31696
rect 30472 30796 30524 30802
rect 30472 30738 30524 30744
rect 30288 29640 30340 29646
rect 30288 29582 30340 29588
rect 30380 29640 30432 29646
rect 30380 29582 30432 29588
rect 30300 29345 30328 29582
rect 30484 29510 30512 30738
rect 30576 29850 30604 31690
rect 30564 29844 30616 29850
rect 30564 29786 30616 29792
rect 30380 29504 30432 29510
rect 30380 29446 30432 29452
rect 30472 29504 30524 29510
rect 30472 29446 30524 29452
rect 30286 29336 30342 29345
rect 30286 29271 30342 29280
rect 30392 29220 30420 29446
rect 30472 29300 30524 29306
rect 30472 29242 30524 29248
rect 30300 29192 30420 29220
rect 30300 27674 30328 29192
rect 30484 29034 30512 29242
rect 30472 29028 30524 29034
rect 30472 28970 30524 28976
rect 30564 29028 30616 29034
rect 30564 28970 30616 28976
rect 30288 27668 30340 27674
rect 30288 27610 30340 27616
rect 30288 27532 30340 27538
rect 30288 27474 30340 27480
rect 30300 26926 30328 27474
rect 30288 26920 30340 26926
rect 30288 26862 30340 26868
rect 30472 26376 30524 26382
rect 30472 26318 30524 26324
rect 30196 25900 30248 25906
rect 30196 25842 30248 25848
rect 30380 25832 30432 25838
rect 30378 25800 30380 25809
rect 30432 25800 30434 25809
rect 30378 25735 30434 25744
rect 30380 25288 30432 25294
rect 30380 25230 30432 25236
rect 30288 25220 30340 25226
rect 30288 25162 30340 25168
rect 30300 24206 30328 25162
rect 30392 24449 30420 25230
rect 30378 24440 30434 24449
rect 30378 24375 30434 24384
rect 30392 24206 30420 24375
rect 30104 24200 30156 24206
rect 30024 24160 30104 24188
rect 29920 24064 29972 24070
rect 29920 24006 29972 24012
rect 30024 23882 30052 24160
rect 30104 24142 30156 24148
rect 30288 24200 30340 24206
rect 30288 24142 30340 24148
rect 30380 24200 30432 24206
rect 30380 24142 30432 24148
rect 30104 24064 30156 24070
rect 30104 24006 30156 24012
rect 30380 24064 30432 24070
rect 30380 24006 30432 24012
rect 29932 23854 30052 23882
rect 30116 23882 30144 24006
rect 30116 23854 30236 23882
rect 29828 23248 29880 23254
rect 29828 23190 29880 23196
rect 29748 22596 29868 22624
rect 29644 22578 29696 22584
rect 29656 22488 29684 22578
rect 29656 22460 29776 22488
rect 29552 22160 29604 22166
rect 29552 22102 29604 22108
rect 29552 21888 29604 21894
rect 29552 21830 29604 21836
rect 29460 21412 29512 21418
rect 29460 21354 29512 21360
rect 29368 19848 29420 19854
rect 29368 19790 29420 19796
rect 29276 19780 29328 19786
rect 28540 17672 28592 17678
rect 28540 17614 28592 17620
rect 28552 16250 28580 17614
rect 28630 17232 28686 17241
rect 28630 17167 28632 17176
rect 28684 17167 28686 17176
rect 28632 17138 28684 17144
rect 28632 16992 28684 16998
rect 28632 16934 28684 16940
rect 28644 16658 28672 16934
rect 28736 16794 28764 19306
rect 29012 17746 29040 19774
rect 29276 19722 29328 19728
rect 29182 19544 29238 19553
rect 29182 19479 29238 19488
rect 29092 19372 29144 19378
rect 29092 19314 29144 19320
rect 29000 17740 29052 17746
rect 29000 17682 29052 17688
rect 28816 17332 28868 17338
rect 28868 17292 29040 17320
rect 28816 17274 28868 17280
rect 29012 17202 29040 17292
rect 29000 17196 29052 17202
rect 29000 17138 29052 17144
rect 28906 17096 28962 17105
rect 28906 17031 28908 17040
rect 28960 17031 28962 17040
rect 28908 17002 28960 17008
rect 29104 16998 29132 19314
rect 29196 17270 29224 19479
rect 29276 17740 29328 17746
rect 29276 17682 29328 17688
rect 29184 17264 29236 17270
rect 29184 17206 29236 17212
rect 29288 17066 29316 17682
rect 29276 17060 29328 17066
rect 29276 17002 29328 17008
rect 29092 16992 29144 16998
rect 29092 16934 29144 16940
rect 28724 16788 28776 16794
rect 28724 16730 28776 16736
rect 28632 16652 28684 16658
rect 28632 16594 28684 16600
rect 28540 16244 28592 16250
rect 28540 16186 28592 16192
rect 28460 16102 28580 16130
rect 28446 15192 28502 15201
rect 28446 15127 28448 15136
rect 28500 15127 28502 15136
rect 28448 15098 28500 15104
rect 28264 15088 28316 15094
rect 28264 15030 28316 15036
rect 28276 14550 28304 15030
rect 28356 14816 28408 14822
rect 28356 14758 28408 14764
rect 28264 14544 28316 14550
rect 28368 14521 28396 14758
rect 28264 14486 28316 14492
rect 28354 14512 28410 14521
rect 28172 14272 28224 14278
rect 28172 14214 28224 14220
rect 28080 14068 28132 14074
rect 28000 14028 28080 14056
rect 28080 14010 28132 14016
rect 28170 13968 28226 13977
rect 28170 13903 28172 13912
rect 28224 13903 28226 13912
rect 28172 13874 28224 13880
rect 28172 13728 28224 13734
rect 28172 13670 28224 13676
rect 28184 13530 28212 13670
rect 28172 13524 28224 13530
rect 28172 13466 28224 13472
rect 27896 13320 27948 13326
rect 27896 13262 27948 13268
rect 27908 12918 27936 13262
rect 28080 13184 28132 13190
rect 28080 13126 28132 13132
rect 27896 12912 27948 12918
rect 27896 12854 27948 12860
rect 28092 12238 28120 13126
rect 28080 12232 28132 12238
rect 28080 12174 28132 12180
rect 27896 12096 27948 12102
rect 27896 12038 27948 12044
rect 27908 9674 27936 12038
rect 28000 9982 28212 10010
rect 28000 9926 28028 9982
rect 27988 9920 28040 9926
rect 27988 9862 28040 9868
rect 28080 9920 28132 9926
rect 28080 9862 28132 9868
rect 27908 9646 28028 9674
rect 27896 9376 27948 9382
rect 27896 9318 27948 9324
rect 27908 9178 27936 9318
rect 27896 9172 27948 9178
rect 27896 9114 27948 9120
rect 27804 5908 27856 5914
rect 27804 5850 27856 5856
rect 28000 5710 28028 9646
rect 28092 9110 28120 9862
rect 28080 9104 28132 9110
rect 28080 9046 28132 9052
rect 28080 8492 28132 8498
rect 28080 8434 28132 8440
rect 28092 8294 28120 8434
rect 28080 8288 28132 8294
rect 28080 8230 28132 8236
rect 28184 7857 28212 9982
rect 28276 9042 28304 14486
rect 28354 14447 28410 14456
rect 28552 14278 28580 16102
rect 28632 16108 28684 16114
rect 28632 16050 28684 16056
rect 28540 14272 28592 14278
rect 28540 14214 28592 14220
rect 28354 14104 28410 14113
rect 28410 14074 28488 14090
rect 28410 14068 28500 14074
rect 28410 14062 28448 14068
rect 28354 14039 28410 14048
rect 28448 14010 28500 14016
rect 28644 12481 28672 16050
rect 28736 16046 28764 16730
rect 28724 16040 28776 16046
rect 28724 15982 28776 15988
rect 29288 15162 29316 17002
rect 29276 15156 29328 15162
rect 29276 15098 29328 15104
rect 28908 15020 28960 15026
rect 29380 15008 29408 19790
rect 29472 17762 29500 21354
rect 29564 20262 29592 21830
rect 29748 21690 29776 22460
rect 29736 21684 29788 21690
rect 29736 21626 29788 21632
rect 29840 20942 29868 22596
rect 29828 20936 29880 20942
rect 29828 20878 29880 20884
rect 29644 20800 29696 20806
rect 29932 20788 29960 23854
rect 30208 23730 30236 23854
rect 30104 23724 30156 23730
rect 30104 23666 30156 23672
rect 30196 23724 30248 23730
rect 30196 23666 30248 23672
rect 30012 23316 30064 23322
rect 30012 23258 30064 23264
rect 30024 22506 30052 23258
rect 30116 22681 30144 23666
rect 30196 23248 30248 23254
rect 30196 23190 30248 23196
rect 30102 22672 30158 22681
rect 30208 22642 30236 23190
rect 30392 23118 30420 24006
rect 30380 23112 30432 23118
rect 30380 23054 30432 23060
rect 30102 22607 30158 22616
rect 30196 22636 30248 22642
rect 30012 22500 30064 22506
rect 30012 22442 30064 22448
rect 29644 20742 29696 20748
rect 29748 20760 29960 20788
rect 29552 20256 29604 20262
rect 29552 20198 29604 20204
rect 29552 19984 29604 19990
rect 29552 19926 29604 19932
rect 29564 19514 29592 19926
rect 29552 19508 29604 19514
rect 29552 19450 29604 19456
rect 29656 17882 29684 20742
rect 29748 19334 29776 20760
rect 30024 20534 30052 22442
rect 30116 22030 30144 22607
rect 30196 22578 30248 22584
rect 30380 22636 30432 22642
rect 30380 22578 30432 22584
rect 30196 22432 30248 22438
rect 30196 22374 30248 22380
rect 30104 22024 30156 22030
rect 30104 21966 30156 21972
rect 30104 21548 30156 21554
rect 30104 21490 30156 21496
rect 30012 20528 30064 20534
rect 30012 20470 30064 20476
rect 29828 20256 29880 20262
rect 29828 20198 29880 20204
rect 29840 19854 29868 20198
rect 30024 20097 30052 20470
rect 30010 20088 30066 20097
rect 30010 20023 30066 20032
rect 30012 19984 30064 19990
rect 30012 19926 30064 19932
rect 29828 19848 29880 19854
rect 29828 19790 29880 19796
rect 29920 19848 29972 19854
rect 30024 19836 30052 19926
rect 29972 19808 30052 19836
rect 29920 19790 29972 19796
rect 29840 19718 29868 19790
rect 29828 19712 29880 19718
rect 29828 19654 29880 19660
rect 29932 19514 29960 19790
rect 30012 19712 30064 19718
rect 30012 19654 30064 19660
rect 29920 19508 29972 19514
rect 29920 19450 29972 19456
rect 29748 19306 29868 19334
rect 29736 18080 29788 18086
rect 29736 18022 29788 18028
rect 29644 17876 29696 17882
rect 29644 17818 29696 17824
rect 29472 17734 29684 17762
rect 29656 17649 29684 17734
rect 29642 17640 29698 17649
rect 29552 17604 29604 17610
rect 29642 17575 29644 17584
rect 29552 17546 29604 17552
rect 29696 17575 29698 17584
rect 29644 17546 29696 17552
rect 29460 16992 29512 16998
rect 29460 16934 29512 16940
rect 29472 16522 29500 16934
rect 29460 16516 29512 16522
rect 29460 16458 29512 16464
rect 29458 15192 29514 15201
rect 29458 15127 29514 15136
rect 28960 14980 29408 15008
rect 28908 14962 28960 14968
rect 29092 14884 29144 14890
rect 29092 14826 29144 14832
rect 29184 14884 29236 14890
rect 29184 14826 29236 14832
rect 28908 14272 28960 14278
rect 28908 14214 28960 14220
rect 28920 13938 28948 14214
rect 28908 13932 28960 13938
rect 28908 13874 28960 13880
rect 29104 12850 29132 14826
rect 29196 14618 29224 14826
rect 29184 14612 29236 14618
rect 29184 14554 29236 14560
rect 29380 14074 29408 14980
rect 29472 14958 29500 15127
rect 29460 14952 29512 14958
rect 29460 14894 29512 14900
rect 29368 14068 29420 14074
rect 29368 14010 29420 14016
rect 29380 13530 29408 14010
rect 29368 13524 29420 13530
rect 29368 13466 29420 13472
rect 29092 12844 29144 12850
rect 29092 12786 29144 12792
rect 28630 12472 28686 12481
rect 29564 12434 29592 17546
rect 29644 17332 29696 17338
rect 29644 17274 29696 17280
rect 29656 15026 29684 17274
rect 29748 15366 29776 18022
rect 29840 17954 29868 19306
rect 30024 18222 30052 19654
rect 30116 18222 30144 21490
rect 30208 21010 30236 22374
rect 30392 22030 30420 22578
rect 30484 22506 30512 26318
rect 30576 25906 30604 28970
rect 30760 26518 30788 32166
rect 30852 29345 30880 32710
rect 31036 31482 31064 35090
rect 31404 35086 31432 35119
rect 31392 35080 31444 35086
rect 31392 35022 31444 35028
rect 31116 34944 31168 34950
rect 31116 34886 31168 34892
rect 30932 31476 30984 31482
rect 30932 31418 30984 31424
rect 31024 31476 31076 31482
rect 31024 31418 31076 31424
rect 30944 31278 30972 31418
rect 30932 31272 30984 31278
rect 30932 31214 30984 31220
rect 31036 30870 31064 31418
rect 31024 30864 31076 30870
rect 31024 30806 31076 30812
rect 31128 30716 31156 34886
rect 31300 34604 31352 34610
rect 31300 34546 31352 34552
rect 31208 32564 31260 32570
rect 31208 32506 31260 32512
rect 31220 31822 31248 32506
rect 31208 31816 31260 31822
rect 31208 31758 31260 31764
rect 31220 30870 31248 31758
rect 31208 30864 31260 30870
rect 31208 30806 31260 30812
rect 31208 30728 31260 30734
rect 31128 30688 31208 30716
rect 31208 30670 31260 30676
rect 30932 29640 30984 29646
rect 30932 29582 30984 29588
rect 31024 29640 31076 29646
rect 31024 29582 31076 29588
rect 30838 29336 30894 29345
rect 30944 29306 30972 29582
rect 30838 29271 30894 29280
rect 30932 29300 30984 29306
rect 30932 29242 30984 29248
rect 31036 28762 31064 29582
rect 31116 29504 31168 29510
rect 31116 29446 31168 29452
rect 31128 29170 31156 29446
rect 31116 29164 31168 29170
rect 31116 29106 31168 29112
rect 31208 29164 31260 29170
rect 31312 29152 31340 34546
rect 31496 31822 31524 37062
rect 31864 36922 31892 37130
rect 31852 36916 31904 36922
rect 31852 36858 31904 36864
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 31852 36168 31904 36174
rect 31852 36110 31904 36116
rect 31944 36168 31996 36174
rect 31944 36110 31996 36116
rect 34152 36168 34204 36174
rect 34152 36110 34204 36116
rect 31864 35766 31892 36110
rect 31852 35760 31904 35766
rect 31852 35702 31904 35708
rect 31760 35692 31812 35698
rect 31760 35634 31812 35640
rect 31772 35018 31800 35634
rect 31956 35562 31984 36110
rect 32128 36032 32180 36038
rect 32128 35974 32180 35980
rect 33140 36032 33192 36038
rect 33140 35974 33192 35980
rect 33876 36032 33928 36038
rect 33876 35974 33928 35980
rect 33968 36032 34020 36038
rect 33968 35974 34020 35980
rect 32140 35766 32168 35974
rect 33152 35766 33180 35974
rect 32128 35760 32180 35766
rect 32128 35702 32180 35708
rect 33140 35760 33192 35766
rect 33140 35702 33192 35708
rect 32128 35624 32180 35630
rect 32128 35566 32180 35572
rect 33506 35592 33562 35601
rect 31944 35556 31996 35562
rect 31944 35498 31996 35504
rect 31576 35012 31628 35018
rect 31576 34954 31628 34960
rect 31668 35012 31720 35018
rect 31668 34954 31720 34960
rect 31760 35012 31812 35018
rect 31760 34954 31812 34960
rect 31588 34678 31616 34954
rect 31680 34921 31708 34954
rect 31666 34912 31722 34921
rect 31666 34847 31722 34856
rect 31576 34672 31628 34678
rect 31576 34614 31628 34620
rect 31680 33289 31708 34847
rect 32140 33930 32168 35566
rect 33506 35527 33562 35536
rect 33784 35556 33836 35562
rect 32310 35320 32366 35329
rect 33520 35290 33548 35527
rect 33784 35498 33836 35504
rect 32310 35255 32366 35264
rect 33508 35284 33560 35290
rect 32324 34678 32352 35255
rect 33508 35226 33560 35232
rect 33796 35154 33824 35498
rect 32588 35148 32640 35154
rect 32588 35090 32640 35096
rect 33784 35148 33836 35154
rect 33784 35090 33836 35096
rect 32600 35018 32628 35090
rect 32864 35080 32916 35086
rect 32864 35022 32916 35028
rect 33414 35048 33470 35057
rect 32588 35012 32640 35018
rect 32588 34954 32640 34960
rect 32312 34672 32364 34678
rect 32312 34614 32364 34620
rect 32220 34536 32272 34542
rect 32220 34478 32272 34484
rect 32232 34134 32260 34478
rect 32220 34128 32272 34134
rect 32220 34070 32272 34076
rect 32600 34066 32628 34954
rect 32772 34740 32824 34746
rect 32772 34682 32824 34688
rect 32680 34604 32732 34610
rect 32680 34546 32732 34552
rect 32588 34060 32640 34066
rect 32588 34002 32640 34008
rect 32128 33924 32180 33930
rect 32128 33866 32180 33872
rect 32692 33862 32720 34546
rect 32784 33998 32812 34682
rect 32772 33992 32824 33998
rect 32772 33934 32824 33940
rect 32312 33856 32364 33862
rect 32312 33798 32364 33804
rect 32680 33856 32732 33862
rect 32680 33798 32732 33804
rect 32220 33516 32272 33522
rect 32324 33504 32352 33798
rect 32272 33476 32352 33504
rect 32220 33458 32272 33464
rect 32128 33312 32180 33318
rect 31666 33280 31722 33289
rect 32128 33254 32180 33260
rect 31666 33215 31722 33224
rect 32140 32586 32168 33254
rect 31956 32558 32168 32586
rect 31760 31884 31812 31890
rect 31760 31826 31812 31832
rect 31484 31816 31536 31822
rect 31484 31758 31536 31764
rect 31484 31680 31536 31686
rect 31484 31622 31536 31628
rect 31496 31346 31524 31622
rect 31772 31346 31800 31826
rect 31392 31340 31444 31346
rect 31392 31282 31444 31288
rect 31484 31340 31536 31346
rect 31484 31282 31536 31288
rect 31760 31340 31812 31346
rect 31760 31282 31812 31288
rect 31404 31226 31432 31282
rect 31404 31198 31800 31226
rect 31484 31136 31536 31142
rect 31484 31078 31536 31084
rect 31496 30734 31524 31078
rect 31668 30864 31720 30870
rect 31668 30806 31720 30812
rect 31772 30818 31800 31198
rect 31484 30728 31536 30734
rect 31484 30670 31536 30676
rect 31576 30184 31628 30190
rect 31576 30126 31628 30132
rect 31588 29850 31616 30126
rect 31576 29844 31628 29850
rect 31576 29786 31628 29792
rect 31680 29646 31708 30806
rect 31772 30790 31892 30818
rect 31864 30394 31892 30790
rect 31852 30388 31904 30394
rect 31852 30330 31904 30336
rect 31760 30252 31812 30258
rect 31760 30194 31812 30200
rect 31668 29640 31720 29646
rect 31668 29582 31720 29588
rect 31392 29232 31444 29238
rect 31392 29174 31444 29180
rect 31260 29124 31340 29152
rect 31208 29106 31260 29112
rect 31116 29028 31168 29034
rect 31220 29016 31248 29106
rect 31168 28988 31248 29016
rect 31116 28970 31168 28976
rect 31024 28756 31076 28762
rect 31024 28698 31076 28704
rect 31036 28422 31064 28698
rect 31404 28558 31432 29174
rect 31680 29170 31708 29582
rect 31668 29164 31720 29170
rect 31668 29106 31720 29112
rect 31208 28552 31260 28558
rect 31208 28494 31260 28500
rect 31392 28552 31444 28558
rect 31392 28494 31444 28500
rect 31024 28416 31076 28422
rect 31024 28358 31076 28364
rect 31024 27872 31076 27878
rect 31024 27814 31076 27820
rect 30930 27704 30986 27713
rect 31036 27674 31064 27814
rect 30930 27639 30986 27648
rect 31024 27668 31076 27674
rect 30944 27606 30972 27639
rect 31024 27610 31076 27616
rect 30932 27600 30984 27606
rect 30932 27542 30984 27548
rect 30840 27464 30892 27470
rect 30838 27432 30840 27441
rect 30892 27432 30894 27441
rect 30838 27367 30894 27376
rect 30840 27124 30892 27130
rect 30840 27066 30892 27072
rect 30748 26512 30800 26518
rect 30748 26454 30800 26460
rect 30564 25900 30616 25906
rect 30564 25842 30616 25848
rect 30656 25288 30708 25294
rect 30656 25230 30708 25236
rect 30668 24750 30696 25230
rect 30656 24744 30708 24750
rect 30656 24686 30708 24692
rect 30562 24440 30618 24449
rect 30618 24398 30696 24426
rect 30562 24375 30618 24384
rect 30564 22976 30616 22982
rect 30564 22918 30616 22924
rect 30472 22500 30524 22506
rect 30472 22442 30524 22448
rect 30470 22264 30526 22273
rect 30470 22199 30472 22208
rect 30524 22199 30526 22208
rect 30472 22170 30524 22176
rect 30380 22024 30432 22030
rect 30380 21966 30432 21972
rect 30196 21004 30248 21010
rect 30196 20946 30248 20952
rect 30288 20936 30340 20942
rect 30208 20884 30288 20890
rect 30208 20878 30340 20884
rect 30380 20936 30432 20942
rect 30380 20878 30432 20884
rect 30208 20862 30328 20878
rect 30012 18216 30064 18222
rect 30012 18158 30064 18164
rect 30104 18216 30156 18222
rect 30104 18158 30156 18164
rect 30024 18086 30052 18158
rect 30012 18080 30064 18086
rect 30012 18022 30064 18028
rect 29840 17926 29960 17954
rect 29828 17128 29880 17134
rect 29932 17116 29960 17926
rect 30010 17368 30066 17377
rect 30010 17303 30012 17312
rect 30064 17303 30066 17312
rect 30012 17274 30064 17280
rect 29880 17088 29960 17116
rect 29828 17070 29880 17076
rect 29736 15360 29788 15366
rect 29736 15302 29788 15308
rect 29828 15088 29880 15094
rect 29828 15030 29880 15036
rect 29644 15020 29696 15026
rect 29644 14962 29696 14968
rect 29734 14376 29790 14385
rect 29734 14311 29790 14320
rect 29748 13938 29776 14311
rect 29736 13932 29788 13938
rect 29736 13874 29788 13880
rect 29736 13320 29788 13326
rect 29736 13262 29788 13268
rect 29748 12986 29776 13262
rect 29736 12980 29788 12986
rect 29736 12922 29788 12928
rect 29840 12850 29868 15030
rect 29932 14958 29960 17088
rect 30116 15706 30144 18158
rect 30208 17202 30236 20862
rect 30392 20210 30420 20878
rect 30300 20182 30420 20210
rect 30300 19394 30328 20182
rect 30378 20088 30434 20097
rect 30378 20023 30434 20032
rect 30392 19922 30420 20023
rect 30380 19916 30432 19922
rect 30380 19858 30432 19864
rect 30392 19514 30420 19858
rect 30380 19508 30432 19514
rect 30380 19450 30432 19456
rect 30484 19446 30512 22170
rect 30472 19440 30524 19446
rect 30300 19366 30420 19394
rect 30472 19382 30524 19388
rect 30392 18306 30420 19366
rect 30484 18426 30512 19382
rect 30472 18420 30524 18426
rect 30472 18362 30524 18368
rect 30300 18278 30420 18306
rect 30300 17490 30328 18278
rect 30576 18154 30604 22918
rect 30668 22642 30696 24398
rect 30760 22642 30788 26454
rect 30852 26382 30880 27066
rect 30840 26376 30892 26382
rect 30840 26318 30892 26324
rect 30852 25294 30880 26318
rect 30840 25288 30892 25294
rect 30840 25230 30892 25236
rect 30852 24698 30880 25230
rect 30944 24818 30972 27542
rect 31220 27470 31248 28494
rect 31392 28416 31444 28422
rect 31392 28358 31444 28364
rect 31300 27872 31352 27878
rect 31404 27849 31432 28358
rect 31772 28234 31800 30194
rect 31852 29776 31904 29782
rect 31852 29718 31904 29724
rect 31864 29170 31892 29718
rect 31852 29164 31904 29170
rect 31852 29106 31904 29112
rect 31772 28206 31892 28234
rect 31760 28144 31812 28150
rect 31760 28086 31812 28092
rect 31576 28076 31628 28082
rect 31576 28018 31628 28024
rect 31300 27814 31352 27820
rect 31390 27840 31446 27849
rect 31024 27464 31076 27470
rect 31024 27406 31076 27412
rect 31208 27464 31260 27470
rect 31208 27406 31260 27412
rect 31036 27169 31064 27406
rect 31116 27396 31168 27402
rect 31116 27338 31168 27344
rect 31022 27160 31078 27169
rect 31128 27130 31156 27338
rect 31022 27095 31078 27104
rect 31116 27124 31168 27130
rect 31036 26382 31064 27095
rect 31116 27066 31168 27072
rect 31220 26994 31248 27406
rect 31208 26988 31260 26994
rect 31208 26930 31260 26936
rect 31024 26376 31076 26382
rect 31024 26318 31076 26324
rect 31206 26208 31262 26217
rect 31206 26143 31262 26152
rect 31116 25900 31168 25906
rect 31116 25842 31168 25848
rect 30932 24812 30984 24818
rect 30932 24754 30984 24760
rect 30852 24670 30972 24698
rect 30840 24608 30892 24614
rect 30840 24550 30892 24556
rect 30852 24342 30880 24550
rect 30840 24336 30892 24342
rect 30840 24278 30892 24284
rect 30840 24200 30892 24206
rect 30840 24142 30892 24148
rect 30852 22778 30880 24142
rect 30944 24018 30972 24670
rect 30944 23990 31064 24018
rect 30840 22772 30892 22778
rect 30840 22714 30892 22720
rect 30656 22636 30708 22642
rect 30656 22578 30708 22584
rect 30748 22636 30800 22642
rect 30748 22578 30800 22584
rect 30746 22536 30802 22545
rect 30746 22471 30802 22480
rect 30656 22432 30708 22438
rect 30656 22374 30708 22380
rect 30668 22234 30696 22374
rect 30656 22228 30708 22234
rect 30656 22170 30708 22176
rect 30656 21956 30708 21962
rect 30656 21898 30708 21904
rect 30668 20942 30696 21898
rect 30656 20936 30708 20942
rect 30656 20878 30708 20884
rect 30656 20256 30708 20262
rect 30656 20198 30708 20204
rect 30668 20058 30696 20198
rect 30656 20052 30708 20058
rect 30656 19994 30708 20000
rect 30668 19718 30696 19994
rect 30656 19712 30708 19718
rect 30656 19654 30708 19660
rect 30654 19544 30710 19553
rect 30654 19479 30710 19488
rect 30668 18290 30696 19479
rect 30760 19242 30788 22471
rect 30852 22234 30880 22714
rect 30932 22636 30984 22642
rect 30932 22578 30984 22584
rect 30840 22228 30892 22234
rect 30840 22170 30892 22176
rect 30838 22128 30894 22137
rect 30944 22098 30972 22578
rect 31036 22574 31064 23990
rect 31024 22568 31076 22574
rect 31024 22510 31076 22516
rect 31024 22432 31076 22438
rect 31024 22374 31076 22380
rect 30838 22063 30894 22072
rect 30932 22092 30984 22098
rect 30852 21978 30880 22063
rect 30932 22034 30984 22040
rect 30852 21950 30972 21978
rect 30840 21684 30892 21690
rect 30840 21626 30892 21632
rect 30852 19854 30880 21626
rect 30944 21146 30972 21950
rect 30932 21140 30984 21146
rect 30932 21082 30984 21088
rect 30932 20936 30984 20942
rect 30932 20878 30984 20884
rect 30840 19848 30892 19854
rect 30840 19790 30892 19796
rect 30944 19378 30972 20878
rect 31036 20058 31064 22374
rect 31128 21418 31156 25842
rect 31220 24750 31248 26143
rect 31208 24744 31260 24750
rect 31208 24686 31260 24692
rect 31220 23730 31248 24686
rect 31312 24614 31340 27814
rect 31390 27775 31446 27784
rect 31300 24608 31352 24614
rect 31300 24550 31352 24556
rect 31300 24132 31352 24138
rect 31300 24074 31352 24080
rect 31312 23866 31340 24074
rect 31300 23860 31352 23866
rect 31300 23802 31352 23808
rect 31208 23724 31260 23730
rect 31208 23666 31260 23672
rect 31300 23724 31352 23730
rect 31300 23666 31352 23672
rect 31206 23624 31262 23633
rect 31206 23559 31208 23568
rect 31260 23559 31262 23568
rect 31208 23530 31260 23536
rect 31208 22704 31260 22710
rect 31312 22692 31340 23666
rect 31260 22664 31340 22692
rect 31208 22646 31260 22652
rect 31208 22228 31260 22234
rect 31208 22170 31260 22176
rect 31116 21412 31168 21418
rect 31116 21354 31168 21360
rect 31220 21298 31248 22170
rect 31312 22001 31340 22664
rect 31404 22642 31432 27775
rect 31484 27532 31536 27538
rect 31484 27474 31536 27480
rect 31496 25498 31524 27474
rect 31588 27470 31616 28018
rect 31666 27840 31722 27849
rect 31666 27775 31722 27784
rect 31680 27606 31708 27775
rect 31668 27600 31720 27606
rect 31668 27542 31720 27548
rect 31576 27464 31628 27470
rect 31576 27406 31628 27412
rect 31772 27282 31800 28086
rect 31864 27878 31892 28206
rect 31852 27872 31904 27878
rect 31852 27814 31904 27820
rect 31852 27464 31904 27470
rect 31852 27406 31904 27412
rect 31588 27254 31800 27282
rect 31484 25492 31536 25498
rect 31484 25434 31536 25440
rect 31496 24410 31524 25434
rect 31484 24404 31536 24410
rect 31484 24346 31536 24352
rect 31484 24200 31536 24206
rect 31484 24142 31536 24148
rect 31392 22636 31444 22642
rect 31392 22578 31444 22584
rect 31390 22536 31446 22545
rect 31390 22471 31446 22480
rect 31298 21992 31354 22001
rect 31298 21927 31354 21936
rect 31300 21888 31352 21894
rect 31300 21830 31352 21836
rect 31312 21418 31340 21830
rect 31404 21554 31432 22471
rect 31392 21548 31444 21554
rect 31392 21490 31444 21496
rect 31300 21412 31352 21418
rect 31300 21354 31352 21360
rect 31392 21412 31444 21418
rect 31392 21354 31444 21360
rect 31404 21298 31432 21354
rect 31128 21270 31248 21298
rect 31312 21270 31432 21298
rect 31128 20806 31156 21270
rect 31208 20936 31260 20942
rect 31312 20924 31340 21270
rect 31496 21128 31524 24142
rect 31588 22642 31616 27254
rect 31760 27124 31812 27130
rect 31760 27066 31812 27072
rect 31668 26920 31720 26926
rect 31668 26862 31720 26868
rect 31680 26586 31708 26862
rect 31668 26580 31720 26586
rect 31668 26522 31720 26528
rect 31772 26246 31800 27066
rect 31760 26240 31812 26246
rect 31760 26182 31812 26188
rect 31760 25220 31812 25226
rect 31760 25162 31812 25168
rect 31668 23860 31720 23866
rect 31668 23802 31720 23808
rect 31680 23118 31708 23802
rect 31772 23118 31800 25162
rect 31864 24410 31892 27406
rect 31956 26874 31984 32558
rect 32232 32366 32260 33458
rect 32692 33454 32720 33798
rect 32680 33448 32732 33454
rect 32680 33390 32732 33396
rect 32784 33318 32812 33934
rect 32772 33312 32824 33318
rect 32772 33254 32824 33260
rect 32876 32570 32904 35022
rect 33414 34983 33470 34992
rect 33428 34542 33456 34983
rect 33692 34604 33744 34610
rect 33692 34546 33744 34552
rect 33416 34536 33468 34542
rect 33416 34478 33468 34484
rect 32956 34128 33008 34134
rect 32956 34070 33008 34076
rect 32968 33522 32996 34070
rect 33048 34060 33100 34066
rect 33048 34002 33100 34008
rect 32956 33516 33008 33522
rect 32956 33458 33008 33464
rect 32588 32564 32640 32570
rect 32588 32506 32640 32512
rect 32864 32564 32916 32570
rect 32864 32506 32916 32512
rect 32220 32360 32272 32366
rect 32220 32302 32272 32308
rect 32036 32224 32088 32230
rect 32036 32166 32088 32172
rect 32048 28966 32076 32166
rect 32128 31816 32180 31822
rect 32128 31758 32180 31764
rect 32404 31816 32456 31822
rect 32404 31758 32456 31764
rect 32140 31142 32168 31758
rect 32416 31346 32444 31758
rect 32496 31680 32548 31686
rect 32496 31622 32548 31628
rect 32508 31346 32536 31622
rect 32404 31340 32456 31346
rect 32404 31282 32456 31288
rect 32496 31340 32548 31346
rect 32496 31282 32548 31288
rect 32128 31136 32180 31142
rect 32180 31096 32352 31124
rect 32128 31078 32180 31084
rect 32128 30728 32180 30734
rect 32128 30670 32180 30676
rect 32140 30410 32168 30670
rect 32324 30569 32352 31096
rect 32416 30682 32444 31282
rect 32600 30938 32628 32506
rect 32680 32428 32732 32434
rect 32680 32370 32732 32376
rect 32692 31754 32720 32370
rect 32680 31748 32732 31754
rect 32680 31690 32732 31696
rect 32876 31521 32904 32506
rect 33060 32434 33088 34002
rect 33600 33992 33652 33998
rect 33600 33934 33652 33940
rect 33232 33652 33284 33658
rect 33232 33594 33284 33600
rect 33048 32428 33100 32434
rect 33048 32370 33100 32376
rect 32862 31512 32918 31521
rect 32918 31470 32996 31498
rect 32862 31447 32918 31456
rect 32680 31136 32732 31142
rect 32680 31078 32732 31084
rect 32692 30938 32720 31078
rect 32588 30932 32640 30938
rect 32588 30874 32640 30880
rect 32680 30932 32732 30938
rect 32680 30874 32732 30880
rect 32680 30796 32732 30802
rect 32680 30738 32732 30744
rect 32416 30654 32536 30682
rect 32404 30592 32456 30598
rect 32310 30560 32366 30569
rect 32404 30534 32456 30540
rect 32310 30495 32366 30504
rect 32140 30382 32260 30410
rect 32232 30054 32260 30382
rect 32220 30048 32272 30054
rect 32220 29990 32272 29996
rect 32036 28960 32088 28966
rect 32036 28902 32088 28908
rect 32036 28552 32088 28558
rect 32036 28494 32088 28500
rect 32126 28520 32182 28529
rect 32048 26994 32076 28494
rect 32126 28455 32128 28464
rect 32180 28455 32182 28464
rect 32128 28426 32180 28432
rect 32126 27568 32182 27577
rect 32126 27503 32182 27512
rect 32140 27334 32168 27503
rect 32128 27328 32180 27334
rect 32128 27270 32180 27276
rect 32036 26988 32088 26994
rect 32036 26930 32088 26936
rect 31956 26846 32168 26874
rect 32034 26752 32090 26761
rect 32034 26687 32090 26696
rect 32048 26586 32076 26687
rect 32036 26580 32088 26586
rect 32036 26522 32088 26528
rect 32140 26450 32168 26846
rect 32128 26444 32180 26450
rect 32128 26386 32180 26392
rect 32036 26376 32088 26382
rect 32036 26318 32088 26324
rect 32048 26042 32076 26318
rect 32128 26240 32180 26246
rect 32128 26182 32180 26188
rect 32036 26036 32088 26042
rect 32036 25978 32088 25984
rect 32036 25900 32088 25906
rect 32036 25842 32088 25848
rect 32048 25294 32076 25842
rect 32140 25498 32168 26182
rect 32128 25492 32180 25498
rect 32128 25434 32180 25440
rect 32036 25288 32088 25294
rect 32036 25230 32088 25236
rect 32036 24744 32088 24750
rect 31956 24704 32036 24732
rect 31852 24404 31904 24410
rect 31852 24346 31904 24352
rect 31668 23112 31720 23118
rect 31668 23054 31720 23060
rect 31760 23112 31812 23118
rect 31760 23054 31812 23060
rect 31852 22976 31904 22982
rect 31852 22918 31904 22924
rect 31760 22772 31812 22778
rect 31760 22714 31812 22720
rect 31668 22704 31720 22710
rect 31668 22646 31720 22652
rect 31576 22636 31628 22642
rect 31576 22578 31628 22584
rect 31588 22234 31616 22578
rect 31576 22228 31628 22234
rect 31576 22170 31628 22176
rect 31680 22094 31708 22646
rect 31588 22066 31708 22094
rect 31588 22030 31616 22066
rect 31576 22024 31628 22030
rect 31576 21966 31628 21972
rect 31666 21992 31722 22001
rect 31666 21927 31722 21936
rect 31260 20896 31340 20924
rect 31404 21100 31524 21128
rect 31208 20878 31260 20884
rect 31116 20800 31168 20806
rect 31116 20742 31168 20748
rect 31024 20052 31076 20058
rect 31024 19994 31076 20000
rect 31128 19938 31156 20742
rect 31036 19910 31156 19938
rect 30932 19372 30984 19378
rect 30932 19314 30984 19320
rect 30748 19236 30800 19242
rect 30748 19178 30800 19184
rect 30760 18290 30788 19178
rect 30932 19168 30984 19174
rect 30932 19110 30984 19116
rect 30944 18970 30972 19110
rect 30932 18964 30984 18970
rect 30932 18906 30984 18912
rect 30656 18284 30708 18290
rect 30656 18226 30708 18232
rect 30748 18284 30800 18290
rect 30748 18226 30800 18232
rect 30380 18148 30432 18154
rect 30380 18090 30432 18096
rect 30564 18148 30616 18154
rect 30564 18090 30616 18096
rect 30392 17678 30420 18090
rect 30472 18080 30524 18086
rect 30472 18022 30524 18028
rect 30656 18080 30708 18086
rect 30656 18022 30708 18028
rect 30484 17678 30512 18022
rect 30380 17672 30432 17678
rect 30380 17614 30432 17620
rect 30472 17672 30524 17678
rect 30472 17614 30524 17620
rect 30300 17462 30512 17490
rect 30196 17196 30248 17202
rect 30196 17138 30248 17144
rect 30380 16448 30432 16454
rect 30300 16408 30380 16436
rect 30300 15910 30328 16408
rect 30380 16390 30432 16396
rect 30380 16108 30432 16114
rect 30380 16050 30432 16056
rect 30288 15904 30340 15910
rect 30288 15846 30340 15852
rect 30300 15706 30328 15846
rect 30104 15700 30156 15706
rect 30104 15642 30156 15648
rect 30288 15700 30340 15706
rect 30288 15642 30340 15648
rect 30196 15632 30248 15638
rect 30196 15574 30248 15580
rect 30104 15496 30156 15502
rect 30104 15438 30156 15444
rect 29920 14952 29972 14958
rect 29920 14894 29972 14900
rect 29920 14816 29972 14822
rect 29920 14758 29972 14764
rect 29932 14074 29960 14758
rect 29920 14068 29972 14074
rect 29920 14010 29972 14016
rect 29932 13938 29960 14010
rect 29920 13932 29972 13938
rect 29920 13874 29972 13880
rect 30012 13864 30064 13870
rect 30012 13806 30064 13812
rect 29828 12844 29880 12850
rect 29828 12786 29880 12792
rect 28630 12407 28686 12416
rect 28644 12306 28672 12407
rect 29380 12406 29592 12434
rect 28632 12300 28684 12306
rect 28632 12242 28684 12248
rect 29380 12238 29408 12406
rect 29368 12232 29420 12238
rect 29368 12174 29420 12180
rect 29920 12232 29972 12238
rect 29920 12174 29972 12180
rect 29274 11928 29330 11937
rect 29274 11863 29330 11872
rect 29000 11756 29052 11762
rect 29000 11698 29052 11704
rect 29012 11286 29040 11698
rect 29288 11694 29316 11863
rect 29380 11762 29408 12174
rect 29736 12164 29788 12170
rect 29736 12106 29788 12112
rect 29748 11830 29776 12106
rect 29736 11824 29788 11830
rect 29736 11766 29788 11772
rect 29368 11756 29420 11762
rect 29368 11698 29420 11704
rect 29932 11694 29960 12174
rect 29276 11688 29328 11694
rect 29276 11630 29328 11636
rect 29920 11688 29972 11694
rect 29920 11630 29972 11636
rect 29000 11280 29052 11286
rect 29000 11222 29052 11228
rect 29184 11008 29236 11014
rect 29184 10950 29236 10956
rect 29196 10674 29224 10950
rect 28724 10668 28776 10674
rect 28724 10610 28776 10616
rect 29184 10668 29236 10674
rect 29184 10610 29236 10616
rect 28448 10464 28500 10470
rect 28448 10406 28500 10412
rect 28460 9926 28488 10406
rect 28736 10266 28764 10610
rect 28998 10296 29054 10305
rect 28724 10260 28776 10266
rect 29054 10254 29132 10282
rect 28998 10231 29054 10240
rect 28724 10202 28776 10208
rect 28538 10160 28594 10169
rect 28538 10095 28540 10104
rect 28592 10095 28594 10104
rect 28540 10066 28592 10072
rect 28448 9920 28500 9926
rect 28448 9862 28500 9868
rect 29000 9920 29052 9926
rect 29000 9862 29052 9868
rect 28356 9512 28408 9518
rect 28356 9454 28408 9460
rect 28264 9036 28316 9042
rect 28264 8978 28316 8984
rect 28368 8566 28396 9454
rect 28552 8906 28764 8922
rect 28540 8900 28764 8906
rect 28592 8894 28764 8900
rect 28540 8842 28592 8848
rect 28632 8832 28684 8838
rect 28632 8774 28684 8780
rect 28644 8634 28672 8774
rect 28736 8634 28764 8894
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 28724 8628 28776 8634
rect 28724 8570 28776 8576
rect 28356 8560 28408 8566
rect 28356 8502 28408 8508
rect 28632 8492 28684 8498
rect 28632 8434 28684 8440
rect 28356 8424 28408 8430
rect 28356 8366 28408 8372
rect 28368 8265 28396 8366
rect 28644 8294 28672 8434
rect 28632 8288 28684 8294
rect 28354 8256 28410 8265
rect 28632 8230 28684 8236
rect 28354 8191 28410 8200
rect 28170 7848 28226 7857
rect 28170 7783 28226 7792
rect 28184 7002 28212 7783
rect 28356 7744 28408 7750
rect 28356 7686 28408 7692
rect 28368 7478 28396 7686
rect 28356 7472 28408 7478
rect 28356 7414 28408 7420
rect 28630 7440 28686 7449
rect 28630 7375 28686 7384
rect 28644 7342 28672 7375
rect 28632 7336 28684 7342
rect 28632 7278 28684 7284
rect 28632 7200 28684 7206
rect 28632 7142 28684 7148
rect 28172 6996 28224 7002
rect 28172 6938 28224 6944
rect 28644 6934 28672 7142
rect 28632 6928 28684 6934
rect 28632 6870 28684 6876
rect 28736 6798 28764 8570
rect 28908 7200 28960 7206
rect 29012 7188 29040 9862
rect 29104 9674 29132 10254
rect 29288 10130 29316 11630
rect 29736 11620 29788 11626
rect 29736 11562 29788 11568
rect 29368 11552 29420 11558
rect 29368 11494 29420 11500
rect 29276 10124 29328 10130
rect 29276 10066 29328 10072
rect 29104 9646 29316 9674
rect 29288 7886 29316 9646
rect 29276 7880 29328 7886
rect 29276 7822 29328 7828
rect 29092 7744 29144 7750
rect 29092 7686 29144 7692
rect 29104 7342 29132 7686
rect 29288 7410 29316 7822
rect 29184 7404 29236 7410
rect 29184 7346 29236 7352
rect 29276 7404 29328 7410
rect 29276 7346 29328 7352
rect 29092 7336 29144 7342
rect 29092 7278 29144 7284
rect 29012 7160 29132 7188
rect 28908 7142 28960 7148
rect 28920 6798 28948 7142
rect 28724 6792 28776 6798
rect 28724 6734 28776 6740
rect 28908 6792 28960 6798
rect 28908 6734 28960 6740
rect 29000 6656 29052 6662
rect 29000 6598 29052 6604
rect 29012 6390 29040 6598
rect 29000 6384 29052 6390
rect 29000 6326 29052 6332
rect 28724 6112 28776 6118
rect 28724 6054 28776 6060
rect 28736 5710 28764 6054
rect 27632 5630 27752 5658
rect 27988 5704 28040 5710
rect 27988 5646 28040 5652
rect 28172 5704 28224 5710
rect 28172 5646 28224 5652
rect 28724 5704 28776 5710
rect 28724 5646 28776 5652
rect 27528 5228 27580 5234
rect 27528 5170 27580 5176
rect 27540 4826 27568 5170
rect 27632 5098 27660 5630
rect 27710 5536 27766 5545
rect 27710 5471 27766 5480
rect 27620 5092 27672 5098
rect 27620 5034 27672 5040
rect 27724 5030 27752 5471
rect 28184 5234 28212 5646
rect 28264 5568 28316 5574
rect 28264 5510 28316 5516
rect 28276 5234 28304 5510
rect 29104 5386 29132 7160
rect 29196 7002 29224 7346
rect 29184 6996 29236 7002
rect 29184 6938 29236 6944
rect 29196 6322 29224 6938
rect 29288 6798 29316 7346
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 29184 6316 29236 6322
rect 29184 6258 29236 6264
rect 29380 5710 29408 11494
rect 29552 11008 29604 11014
rect 29552 10950 29604 10956
rect 29564 10674 29592 10950
rect 29642 10840 29698 10849
rect 29642 10775 29698 10784
rect 29656 10674 29684 10775
rect 29552 10668 29604 10674
rect 29552 10610 29604 10616
rect 29644 10668 29696 10674
rect 29644 10610 29696 10616
rect 29564 10470 29592 10610
rect 29552 10464 29604 10470
rect 29552 10406 29604 10412
rect 29748 10062 29776 11562
rect 29932 10554 29960 11630
rect 29840 10526 29960 10554
rect 29736 10056 29788 10062
rect 29736 9998 29788 10004
rect 29644 9512 29696 9518
rect 29644 9454 29696 9460
rect 29552 9104 29604 9110
rect 29552 9046 29604 9052
rect 29460 8492 29512 8498
rect 29460 8434 29512 8440
rect 29472 7818 29500 8434
rect 29564 8090 29592 9046
rect 29656 8498 29684 9454
rect 29736 8968 29788 8974
rect 29736 8910 29788 8916
rect 29644 8492 29696 8498
rect 29644 8434 29696 8440
rect 29552 8084 29604 8090
rect 29552 8026 29604 8032
rect 29564 7818 29592 8026
rect 29748 7954 29776 8910
rect 29840 8090 29868 10526
rect 29920 10464 29972 10470
rect 29920 10406 29972 10412
rect 29932 8974 29960 10406
rect 30024 9024 30052 13806
rect 30116 13802 30144 15438
rect 30208 15366 30236 15574
rect 30392 15502 30420 16050
rect 30380 15496 30432 15502
rect 30380 15438 30432 15444
rect 30196 15360 30248 15366
rect 30196 15302 30248 15308
rect 30208 14793 30236 15302
rect 30194 14784 30250 14793
rect 30194 14719 30250 14728
rect 30380 14408 30432 14414
rect 30380 14350 30432 14356
rect 30196 14272 30248 14278
rect 30196 14214 30248 14220
rect 30104 13796 30156 13802
rect 30104 13738 30156 13744
rect 30116 12918 30144 13738
rect 30104 12912 30156 12918
rect 30104 12854 30156 12860
rect 30104 12776 30156 12782
rect 30104 12718 30156 12724
rect 30116 11762 30144 12718
rect 30104 11756 30156 11762
rect 30104 11698 30156 11704
rect 30208 11200 30236 14214
rect 30288 12980 30340 12986
rect 30288 12922 30340 12928
rect 30300 12170 30328 12922
rect 30392 12889 30420 14350
rect 30484 14074 30512 17462
rect 30668 14618 30696 18022
rect 31036 17762 31064 19910
rect 31116 19304 31168 19310
rect 31114 19272 31116 19281
rect 31168 19272 31170 19281
rect 31114 19207 31170 19216
rect 31128 18086 31156 19207
rect 31116 18080 31168 18086
rect 31116 18022 31168 18028
rect 30944 17734 31064 17762
rect 30944 16114 30972 17734
rect 31024 17672 31076 17678
rect 31024 17614 31076 17620
rect 30932 16108 30984 16114
rect 30932 16050 30984 16056
rect 30840 15496 30892 15502
rect 30840 15438 30892 15444
rect 30656 14612 30708 14618
rect 30656 14554 30708 14560
rect 30852 14414 30880 15438
rect 30932 14952 30984 14958
rect 30932 14894 30984 14900
rect 30944 14414 30972 14894
rect 31036 14414 31064 17614
rect 31220 16522 31248 20878
rect 31404 20806 31432 21100
rect 31574 20904 31630 20913
rect 31574 20839 31576 20848
rect 31628 20839 31630 20848
rect 31576 20810 31628 20816
rect 31392 20800 31444 20806
rect 31392 20742 31444 20748
rect 31574 20768 31630 20777
rect 31574 20703 31630 20712
rect 31588 20466 31616 20703
rect 31576 20460 31628 20466
rect 31576 20402 31628 20408
rect 31300 20392 31352 20398
rect 31300 20334 31352 20340
rect 31392 20392 31444 20398
rect 31680 20346 31708 21927
rect 31772 21486 31800 22714
rect 31864 22642 31892 22918
rect 31852 22636 31904 22642
rect 31852 22578 31904 22584
rect 31956 22094 31984 24704
rect 32036 24686 32088 24692
rect 32036 24608 32088 24614
rect 32036 24550 32088 24556
rect 32128 24608 32180 24614
rect 32128 24550 32180 24556
rect 32048 23118 32076 24550
rect 32140 23168 32168 24550
rect 32232 24342 32260 29990
rect 32324 29782 32352 30495
rect 32312 29776 32364 29782
rect 32312 29718 32364 29724
rect 32312 28960 32364 28966
rect 32312 28902 32364 28908
rect 32324 28218 32352 28902
rect 32312 28212 32364 28218
rect 32312 28154 32364 28160
rect 32220 24336 32272 24342
rect 32220 24278 32272 24284
rect 32324 23633 32352 28154
rect 32416 27606 32444 30534
rect 32508 30258 32536 30654
rect 32496 30252 32548 30258
rect 32496 30194 32548 30200
rect 32588 30184 32640 30190
rect 32588 30126 32640 30132
rect 32496 29164 32548 29170
rect 32496 29106 32548 29112
rect 32404 27600 32456 27606
rect 32404 27542 32456 27548
rect 32508 27470 32536 29106
rect 32600 28966 32628 30126
rect 32588 28960 32640 28966
rect 32588 28902 32640 28908
rect 32588 28416 32640 28422
rect 32588 28358 32640 28364
rect 32600 28218 32628 28358
rect 32588 28212 32640 28218
rect 32588 28154 32640 28160
rect 32588 27872 32640 27878
rect 32588 27814 32640 27820
rect 32496 27464 32548 27470
rect 32496 27406 32548 27412
rect 32404 26988 32456 26994
rect 32404 26930 32456 26936
rect 32416 25294 32444 26930
rect 32508 25430 32536 27406
rect 32600 27402 32628 27814
rect 32588 27396 32640 27402
rect 32588 27338 32640 27344
rect 32588 26920 32640 26926
rect 32588 26862 32640 26868
rect 32600 26382 32628 26862
rect 32588 26376 32640 26382
rect 32588 26318 32640 26324
rect 32496 25424 32548 25430
rect 32496 25366 32548 25372
rect 32586 25392 32642 25401
rect 32692 25378 32720 30738
rect 32864 30252 32916 30258
rect 32864 30194 32916 30200
rect 32772 30048 32824 30054
rect 32772 29990 32824 29996
rect 32784 29714 32812 29990
rect 32772 29708 32824 29714
rect 32772 29650 32824 29656
rect 32876 29646 32904 30194
rect 32864 29640 32916 29646
rect 32864 29582 32916 29588
rect 32772 29504 32824 29510
rect 32772 29446 32824 29452
rect 32784 28558 32812 29446
rect 32876 29102 32904 29582
rect 32968 29306 32996 31470
rect 33060 30002 33088 32370
rect 33140 32224 33192 32230
rect 33140 32166 33192 32172
rect 33152 30870 33180 32166
rect 33244 31822 33272 33594
rect 33612 33590 33640 33934
rect 33600 33584 33652 33590
rect 33600 33526 33652 33532
rect 33612 33454 33640 33526
rect 33600 33448 33652 33454
rect 33600 33390 33652 33396
rect 33324 32224 33376 32230
rect 33324 32166 33376 32172
rect 33336 32026 33364 32166
rect 33324 32020 33376 32026
rect 33324 31962 33376 31968
rect 33600 31884 33652 31890
rect 33600 31826 33652 31832
rect 33232 31816 33284 31822
rect 33612 31793 33640 31826
rect 33232 31758 33284 31764
rect 33598 31784 33654 31793
rect 33598 31719 33654 31728
rect 33508 31680 33560 31686
rect 33508 31622 33560 31628
rect 33520 31482 33548 31622
rect 33508 31476 33560 31482
rect 33508 31418 33560 31424
rect 33416 31340 33468 31346
rect 33416 31282 33468 31288
rect 33140 30864 33192 30870
rect 33140 30806 33192 30812
rect 33428 30598 33456 31282
rect 33600 31272 33652 31278
rect 33600 31214 33652 31220
rect 33612 31142 33640 31214
rect 33600 31136 33652 31142
rect 33600 31078 33652 31084
rect 33416 30592 33468 30598
rect 33416 30534 33468 30540
rect 33414 30424 33470 30433
rect 33470 30382 33548 30410
rect 33414 30359 33470 30368
rect 33416 30116 33468 30122
rect 33416 30058 33468 30064
rect 33060 29974 33272 30002
rect 32956 29300 33008 29306
rect 32956 29242 33008 29248
rect 33060 29170 33088 29974
rect 33140 29844 33192 29850
rect 33140 29786 33192 29792
rect 33152 29238 33180 29786
rect 33244 29578 33272 29974
rect 33232 29572 33284 29578
rect 33232 29514 33284 29520
rect 33428 29306 33456 30058
rect 33520 29782 33548 30382
rect 33508 29776 33560 29782
rect 33508 29718 33560 29724
rect 33508 29640 33560 29646
rect 33612 29628 33640 31078
rect 33560 29600 33640 29628
rect 33508 29582 33560 29588
rect 33416 29300 33468 29306
rect 33416 29242 33468 29248
rect 33140 29232 33192 29238
rect 33140 29174 33192 29180
rect 33048 29164 33100 29170
rect 33048 29106 33100 29112
rect 32864 29096 32916 29102
rect 32864 29038 32916 29044
rect 32772 28552 32824 28558
rect 32772 28494 32824 28500
rect 32784 28150 32812 28494
rect 32772 28144 32824 28150
rect 32772 28086 32824 28092
rect 32772 27600 32824 27606
rect 32772 27542 32824 27548
rect 32784 27441 32812 27542
rect 32770 27432 32826 27441
rect 32770 27367 32826 27376
rect 32772 26376 32824 26382
rect 32772 26318 32824 26324
rect 32784 25498 32812 26318
rect 32772 25492 32824 25498
rect 32772 25434 32824 25440
rect 32692 25350 32812 25378
rect 32586 25327 32642 25336
rect 32404 25288 32456 25294
rect 32404 25230 32456 25236
rect 32416 24886 32444 25230
rect 32496 25152 32548 25158
rect 32496 25094 32548 25100
rect 32404 24880 32456 24886
rect 32404 24822 32456 24828
rect 32508 24410 32536 25094
rect 32600 24614 32628 25327
rect 32680 25288 32732 25294
rect 32680 25230 32732 25236
rect 32588 24608 32640 24614
rect 32588 24550 32640 24556
rect 32496 24404 32548 24410
rect 32496 24346 32548 24352
rect 32496 24064 32548 24070
rect 32496 24006 32548 24012
rect 32404 23656 32456 23662
rect 32310 23624 32366 23633
rect 32404 23598 32456 23604
rect 32310 23559 32366 23568
rect 32140 23140 32352 23168
rect 32036 23112 32088 23118
rect 32036 23054 32088 23060
rect 32220 23044 32272 23050
rect 32220 22986 32272 22992
rect 32232 22710 32260 22986
rect 32220 22704 32272 22710
rect 32220 22646 32272 22652
rect 32128 22636 32180 22642
rect 32128 22578 32180 22584
rect 32036 22160 32088 22166
rect 32036 22102 32088 22108
rect 31864 22066 31984 22094
rect 31760 21480 31812 21486
rect 31760 21422 31812 21428
rect 31760 21140 31812 21146
rect 31760 21082 31812 21088
rect 31392 20334 31444 20340
rect 31312 19922 31340 20334
rect 31404 20233 31432 20334
rect 31496 20318 31708 20346
rect 31496 20262 31524 20318
rect 31484 20256 31536 20262
rect 31390 20224 31446 20233
rect 31484 20198 31536 20204
rect 31576 20256 31628 20262
rect 31576 20198 31628 20204
rect 31390 20159 31446 20168
rect 31390 19952 31446 19961
rect 31300 19916 31352 19922
rect 31390 19887 31392 19896
rect 31300 19858 31352 19864
rect 31444 19887 31446 19896
rect 31392 19858 31444 19864
rect 31484 19848 31536 19854
rect 31484 19790 31536 19796
rect 31390 18728 31446 18737
rect 31390 18663 31446 18672
rect 31404 18630 31432 18663
rect 31392 18624 31444 18630
rect 31496 18601 31524 19790
rect 31588 19786 31616 20198
rect 31576 19780 31628 19786
rect 31576 19722 31628 19728
rect 31576 19236 31628 19242
rect 31576 19178 31628 19184
rect 31588 18970 31616 19178
rect 31576 18964 31628 18970
rect 31576 18906 31628 18912
rect 31668 18964 31720 18970
rect 31668 18906 31720 18912
rect 31680 18630 31708 18906
rect 31772 18766 31800 21082
rect 31760 18760 31812 18766
rect 31760 18702 31812 18708
rect 31668 18624 31720 18630
rect 31392 18566 31444 18572
rect 31482 18592 31538 18601
rect 31668 18566 31720 18572
rect 31758 18592 31814 18601
rect 31482 18527 31538 18536
rect 31392 18284 31444 18290
rect 31392 18226 31444 18232
rect 31404 18034 31432 18226
rect 31312 18006 31432 18034
rect 31312 17785 31340 18006
rect 31576 17808 31628 17814
rect 31298 17776 31354 17785
rect 31576 17750 31628 17756
rect 31298 17711 31354 17720
rect 31588 16590 31616 17750
rect 31576 16584 31628 16590
rect 31576 16526 31628 16532
rect 31208 16516 31260 16522
rect 31208 16458 31260 16464
rect 31116 16448 31168 16454
rect 31116 16390 31168 16396
rect 31128 16182 31156 16390
rect 31116 16176 31168 16182
rect 31116 16118 31168 16124
rect 31220 15434 31248 16458
rect 31680 16436 31708 18566
rect 31758 18527 31814 18536
rect 31772 17678 31800 18527
rect 31864 18426 31892 22066
rect 32048 22012 32076 22102
rect 32048 21984 32077 22012
rect 31944 21888 31996 21894
rect 32049 21842 32077 21984
rect 31944 21830 31996 21836
rect 31956 20874 31984 21830
rect 32048 21814 32077 21842
rect 31944 20868 31996 20874
rect 31944 20810 31996 20816
rect 31852 18420 31904 18426
rect 31852 18362 31904 18368
rect 31956 18306 31984 20810
rect 32048 20534 32076 21814
rect 32036 20528 32088 20534
rect 32036 20470 32088 20476
rect 32036 19848 32088 19854
rect 32036 19790 32088 19796
rect 31864 18278 31984 18306
rect 31760 17672 31812 17678
rect 31760 17614 31812 17620
rect 31760 16992 31812 16998
rect 31760 16934 31812 16940
rect 31588 16408 31708 16436
rect 31484 16176 31536 16182
rect 31588 16153 31616 16408
rect 31484 16118 31536 16124
rect 31574 16144 31630 16153
rect 31392 16108 31444 16114
rect 31392 16050 31444 16056
rect 31208 15428 31260 15434
rect 31208 15370 31260 15376
rect 30840 14408 30892 14414
rect 30840 14350 30892 14356
rect 30932 14408 30984 14414
rect 30932 14350 30984 14356
rect 31024 14408 31076 14414
rect 31024 14350 31076 14356
rect 31300 14408 31352 14414
rect 31300 14350 31352 14356
rect 30564 14340 30616 14346
rect 30564 14282 30616 14288
rect 30472 14068 30524 14074
rect 30472 14010 30524 14016
rect 30378 12880 30434 12889
rect 30378 12815 30434 12824
rect 30392 12306 30420 12815
rect 30380 12300 30432 12306
rect 30380 12242 30432 12248
rect 30472 12232 30524 12238
rect 30472 12174 30524 12180
rect 30288 12164 30340 12170
rect 30288 12106 30340 12112
rect 30300 11830 30328 12106
rect 30380 12096 30432 12102
rect 30380 12038 30432 12044
rect 30288 11824 30340 11830
rect 30288 11766 30340 11772
rect 30392 11558 30420 12038
rect 30380 11552 30432 11558
rect 30380 11494 30432 11500
rect 30208 11172 30328 11200
rect 30300 11121 30328 11172
rect 30286 11112 30342 11121
rect 30196 11076 30248 11082
rect 30286 11047 30342 11056
rect 30196 11018 30248 11024
rect 30208 10674 30236 11018
rect 30484 10810 30512 12174
rect 30576 11898 30604 14282
rect 30852 13433 30880 14350
rect 31036 13938 31064 14350
rect 31312 14278 31340 14350
rect 31300 14272 31352 14278
rect 31300 14214 31352 14220
rect 31404 14074 31432 16050
rect 31496 14550 31524 16118
rect 31574 16079 31630 16088
rect 31588 15026 31616 16079
rect 31772 15502 31800 16934
rect 31864 16590 31892 18278
rect 31852 16584 31904 16590
rect 31852 16526 31904 16532
rect 31944 16516 31996 16522
rect 31944 16458 31996 16464
rect 31760 15496 31812 15502
rect 31760 15438 31812 15444
rect 31668 15360 31720 15366
rect 31956 15348 31984 16458
rect 31668 15302 31720 15308
rect 31772 15320 31984 15348
rect 31576 15020 31628 15026
rect 31576 14962 31628 14968
rect 31680 14890 31708 15302
rect 31772 14890 31800 15320
rect 31852 15020 31904 15026
rect 32048 15008 32076 19790
rect 31852 14962 31904 14968
rect 31956 14980 32076 15008
rect 31668 14884 31720 14890
rect 31668 14826 31720 14832
rect 31760 14884 31812 14890
rect 31760 14826 31812 14832
rect 31484 14544 31536 14550
rect 31484 14486 31536 14492
rect 31680 14414 31708 14826
rect 31484 14408 31536 14414
rect 31484 14350 31536 14356
rect 31576 14408 31628 14414
rect 31576 14350 31628 14356
rect 31668 14408 31720 14414
rect 31864 14396 31892 14962
rect 31956 14634 31984 14980
rect 32140 14906 32168 22578
rect 32220 20868 32272 20874
rect 32220 20810 32272 20816
rect 32232 19854 32260 20810
rect 32220 19848 32272 19854
rect 32220 19790 32272 19796
rect 32220 19712 32272 19718
rect 32220 19654 32272 19660
rect 32232 16998 32260 19654
rect 32220 16992 32272 16998
rect 32220 16934 32272 16940
rect 32218 16824 32274 16833
rect 32218 16759 32220 16768
rect 32272 16759 32274 16768
rect 32220 16730 32272 16736
rect 32220 16448 32272 16454
rect 32220 16390 32272 16396
rect 32232 15706 32260 16390
rect 32220 15700 32272 15706
rect 32220 15642 32272 15648
rect 32232 15162 32260 15642
rect 32324 15366 32352 23140
rect 32312 15360 32364 15366
rect 32312 15302 32364 15308
rect 32416 15162 32444 23598
rect 32508 22778 32536 24006
rect 32600 23866 32628 24550
rect 32692 23866 32720 25230
rect 32588 23860 32640 23866
rect 32588 23802 32640 23808
rect 32680 23860 32732 23866
rect 32680 23802 32732 23808
rect 32600 23730 32628 23802
rect 32588 23724 32640 23730
rect 32588 23666 32640 23672
rect 32588 23588 32640 23594
rect 32588 23530 32640 23536
rect 32680 23588 32732 23594
rect 32680 23530 32732 23536
rect 32600 23186 32628 23530
rect 32692 23254 32720 23530
rect 32680 23248 32732 23254
rect 32680 23190 32732 23196
rect 32588 23180 32640 23186
rect 32588 23122 32640 23128
rect 32680 22976 32732 22982
rect 32680 22918 32732 22924
rect 32496 22772 32548 22778
rect 32496 22714 32548 22720
rect 32692 22642 32720 22918
rect 32680 22636 32732 22642
rect 32680 22578 32732 22584
rect 32496 22432 32548 22438
rect 32496 22374 32548 22380
rect 32508 22094 32536 22374
rect 32508 22066 32628 22094
rect 32496 21140 32548 21146
rect 32496 21082 32548 21088
rect 32508 20942 32536 21082
rect 32496 20936 32548 20942
rect 32496 20878 32548 20884
rect 32508 18970 32536 20878
rect 32600 20806 32628 22066
rect 32692 22030 32720 22578
rect 32680 22024 32732 22030
rect 32680 21966 32732 21972
rect 32588 20800 32640 20806
rect 32588 20742 32640 20748
rect 32784 19854 32812 25350
rect 32876 24818 32904 29038
rect 32956 28960 33008 28966
rect 32956 28902 33008 28908
rect 32968 25401 32996 28902
rect 33060 26586 33088 29106
rect 33324 27464 33376 27470
rect 33416 27464 33468 27470
rect 33324 27406 33376 27412
rect 33414 27432 33416 27441
rect 33468 27432 33470 27441
rect 33232 27328 33284 27334
rect 33232 27270 33284 27276
rect 33048 26580 33100 26586
rect 33100 26540 33180 26568
rect 33048 26522 33100 26528
rect 32954 25392 33010 25401
rect 32954 25327 33010 25336
rect 32956 25288 33008 25294
rect 33008 25236 33088 25242
rect 32956 25230 33088 25236
rect 32968 25214 33088 25230
rect 32956 25152 33008 25158
rect 32956 25094 33008 25100
rect 32864 24812 32916 24818
rect 32864 24754 32916 24760
rect 32968 24698 32996 25094
rect 32876 24670 32996 24698
rect 32876 24614 32904 24670
rect 32864 24608 32916 24614
rect 32864 24550 32916 24556
rect 32954 24576 33010 24585
rect 32954 24511 33010 24520
rect 32864 24200 32916 24206
rect 32864 24142 32916 24148
rect 32876 23905 32904 24142
rect 32862 23896 32918 23905
rect 32862 23831 32918 23840
rect 32968 23730 32996 24511
rect 32956 23724 33008 23730
rect 32956 23666 33008 23672
rect 32864 23180 32916 23186
rect 32864 23122 32916 23128
rect 32876 21146 32904 23122
rect 32968 23050 32996 23666
rect 32956 23044 33008 23050
rect 32956 22986 33008 22992
rect 32864 21140 32916 21146
rect 32864 21082 32916 21088
rect 32864 20800 32916 20806
rect 32864 20742 32916 20748
rect 32772 19848 32824 19854
rect 32772 19790 32824 19796
rect 32496 18964 32548 18970
rect 32496 18906 32548 18912
rect 32680 18896 32732 18902
rect 32680 18838 32732 18844
rect 32588 18828 32640 18834
rect 32588 18770 32640 18776
rect 32496 18624 32548 18630
rect 32496 18566 32548 18572
rect 32220 15156 32272 15162
rect 32220 15098 32272 15104
rect 32404 15156 32456 15162
rect 32404 15098 32456 15104
rect 32048 14878 32168 14906
rect 32220 14884 32272 14890
rect 32048 14822 32076 14878
rect 32220 14826 32272 14832
rect 32036 14816 32088 14822
rect 32036 14758 32088 14764
rect 31956 14606 32076 14634
rect 31944 14544 31996 14550
rect 31942 14512 31944 14521
rect 31996 14512 31998 14521
rect 31942 14447 31998 14456
rect 31864 14368 31984 14396
rect 31668 14350 31720 14356
rect 31392 14068 31444 14074
rect 31392 14010 31444 14016
rect 31024 13932 31076 13938
rect 31024 13874 31076 13880
rect 30838 13424 30894 13433
rect 30838 13359 30894 13368
rect 30656 12096 30708 12102
rect 30656 12038 30708 12044
rect 30668 11898 30696 12038
rect 30564 11892 30616 11898
rect 30564 11834 30616 11840
rect 30656 11892 30708 11898
rect 30656 11834 30708 11840
rect 30564 11756 30616 11762
rect 30748 11756 30800 11762
rect 30616 11716 30748 11744
rect 30564 11698 30616 11704
rect 30748 11698 30800 11704
rect 30852 11676 30880 13359
rect 31036 12374 31064 13874
rect 31496 13462 31524 14350
rect 31484 13456 31536 13462
rect 31484 13398 31536 13404
rect 31300 12776 31352 12782
rect 31300 12718 31352 12724
rect 31024 12368 31076 12374
rect 31024 12310 31076 12316
rect 30930 12200 30986 12209
rect 30930 12135 30986 12144
rect 31208 12164 31260 12170
rect 30944 12102 30972 12135
rect 31208 12106 31260 12112
rect 30932 12096 30984 12102
rect 30932 12038 30984 12044
rect 31220 11898 31248 12106
rect 31312 11898 31340 12718
rect 31588 12442 31616 14350
rect 31760 13932 31812 13938
rect 31760 13874 31812 13880
rect 31772 12986 31800 13874
rect 31852 13184 31904 13190
rect 31852 13126 31904 13132
rect 31760 12980 31812 12986
rect 31760 12922 31812 12928
rect 31668 12912 31720 12918
rect 31668 12854 31720 12860
rect 31576 12436 31628 12442
rect 31576 12378 31628 12384
rect 31576 12232 31628 12238
rect 31680 12220 31708 12854
rect 31628 12192 31708 12220
rect 31576 12174 31628 12180
rect 31392 12164 31444 12170
rect 31392 12106 31444 12112
rect 31404 11898 31432 12106
rect 31208 11892 31260 11898
rect 31208 11834 31260 11840
rect 31300 11892 31352 11898
rect 31300 11834 31352 11840
rect 31392 11892 31444 11898
rect 31392 11834 31444 11840
rect 31404 11676 31432 11834
rect 31588 11694 31616 12174
rect 31576 11688 31628 11694
rect 30852 11648 31064 11676
rect 31404 11648 31524 11676
rect 30656 11552 30708 11558
rect 30656 11494 30708 11500
rect 30564 11076 30616 11082
rect 30564 11018 30616 11024
rect 30472 10804 30524 10810
rect 30472 10746 30524 10752
rect 30104 10668 30156 10674
rect 30104 10610 30156 10616
rect 30196 10668 30248 10674
rect 30196 10610 30248 10616
rect 30116 9586 30144 10610
rect 30196 10260 30248 10266
rect 30196 10202 30248 10208
rect 30104 9580 30156 9586
rect 30104 9522 30156 9528
rect 30208 9042 30236 10202
rect 30484 10130 30512 10746
rect 30576 10470 30604 11018
rect 30564 10464 30616 10470
rect 30564 10406 30616 10412
rect 30472 10124 30524 10130
rect 30472 10066 30524 10072
rect 30288 9920 30340 9926
rect 30288 9862 30340 9868
rect 30300 9178 30328 9862
rect 30380 9648 30432 9654
rect 30380 9590 30432 9596
rect 30288 9172 30340 9178
rect 30288 9114 30340 9120
rect 30104 9036 30156 9042
rect 30024 8996 30104 9024
rect 30104 8978 30156 8984
rect 30196 9036 30248 9042
rect 30196 8978 30248 8984
rect 29920 8968 29972 8974
rect 29920 8910 29972 8916
rect 30300 8906 30328 9114
rect 30196 8900 30248 8906
rect 30196 8842 30248 8848
rect 30288 8900 30340 8906
rect 30288 8842 30340 8848
rect 30012 8356 30064 8362
rect 29932 8316 30012 8344
rect 29828 8084 29880 8090
rect 29828 8026 29880 8032
rect 29736 7948 29788 7954
rect 29656 7908 29736 7936
rect 29460 7812 29512 7818
rect 29460 7754 29512 7760
rect 29552 7812 29604 7818
rect 29552 7754 29604 7760
rect 29472 7410 29500 7754
rect 29552 7472 29604 7478
rect 29552 7414 29604 7420
rect 29460 7404 29512 7410
rect 29460 7346 29512 7352
rect 29472 6798 29500 7346
rect 29460 6792 29512 6798
rect 29460 6734 29512 6740
rect 29564 6390 29592 7414
rect 29656 7274 29684 7908
rect 29736 7890 29788 7896
rect 29736 7812 29788 7818
rect 29736 7754 29788 7760
rect 29748 7449 29776 7754
rect 29734 7440 29790 7449
rect 29840 7410 29868 8026
rect 29932 7410 29960 8316
rect 30012 8298 30064 8304
rect 30102 7984 30158 7993
rect 30102 7919 30158 7928
rect 30116 7886 30144 7919
rect 30104 7880 30156 7886
rect 30104 7822 30156 7828
rect 30208 7750 30236 8842
rect 30288 8288 30340 8294
rect 30288 8230 30340 8236
rect 30196 7744 30248 7750
rect 30196 7686 30248 7692
rect 30300 7410 30328 8230
rect 30392 7585 30420 9590
rect 30562 9208 30618 9217
rect 30562 9143 30564 9152
rect 30616 9143 30618 9152
rect 30564 9114 30616 9120
rect 30472 9036 30524 9042
rect 30472 8978 30524 8984
rect 30484 8906 30512 8978
rect 30472 8900 30524 8906
rect 30472 8842 30524 8848
rect 30484 8634 30512 8842
rect 30472 8628 30524 8634
rect 30524 8588 30604 8616
rect 30472 8570 30524 8576
rect 30472 7812 30524 7818
rect 30472 7754 30524 7760
rect 30378 7576 30434 7585
rect 30378 7511 30434 7520
rect 29734 7375 29790 7384
rect 29828 7404 29880 7410
rect 29828 7346 29880 7352
rect 29920 7404 29972 7410
rect 29920 7346 29972 7352
rect 30288 7404 30340 7410
rect 30288 7346 30340 7352
rect 29644 7268 29696 7274
rect 29644 7210 29696 7216
rect 29932 7018 29960 7346
rect 29840 6990 29960 7018
rect 29644 6928 29696 6934
rect 29644 6870 29696 6876
rect 29656 6730 29684 6870
rect 29644 6724 29696 6730
rect 29644 6666 29696 6672
rect 29552 6384 29604 6390
rect 29552 6326 29604 6332
rect 29656 6322 29684 6666
rect 29644 6316 29696 6322
rect 29644 6258 29696 6264
rect 29368 5704 29420 5710
rect 29368 5646 29420 5652
rect 29104 5358 29224 5386
rect 29092 5296 29144 5302
rect 29092 5238 29144 5244
rect 28172 5228 28224 5234
rect 28172 5170 28224 5176
rect 28264 5228 28316 5234
rect 28264 5170 28316 5176
rect 27712 5024 27764 5030
rect 27712 4966 27764 4972
rect 28184 4826 28212 5170
rect 29000 5024 29052 5030
rect 29000 4966 29052 4972
rect 27528 4820 27580 4826
rect 27528 4762 27580 4768
rect 28172 4820 28224 4826
rect 28172 4762 28224 4768
rect 29012 4690 29040 4966
rect 29104 4826 29132 5238
rect 29092 4820 29144 4826
rect 29092 4762 29144 4768
rect 29000 4684 29052 4690
rect 29000 4626 29052 4632
rect 29196 4622 29224 5358
rect 29380 5030 29408 5646
rect 29368 5024 29420 5030
rect 29368 4966 29420 4972
rect 27436 4616 27488 4622
rect 27436 4558 27488 4564
rect 29184 4616 29236 4622
rect 29184 4558 29236 4564
rect 29840 2514 29868 6990
rect 30300 6798 30328 7346
rect 30392 7274 30420 7511
rect 30484 7410 30512 7754
rect 30472 7404 30524 7410
rect 30576 7392 30604 8588
rect 30668 7750 30696 11494
rect 31036 11354 31064 11648
rect 31024 11348 31076 11354
rect 31024 11290 31076 11296
rect 30840 11280 30892 11286
rect 30840 11222 30892 11228
rect 30852 10674 30880 11222
rect 31496 11150 31524 11648
rect 31576 11630 31628 11636
rect 31484 11144 31536 11150
rect 31484 11086 31536 11092
rect 31208 11008 31260 11014
rect 31208 10950 31260 10956
rect 30840 10668 30892 10674
rect 30840 10610 30892 10616
rect 31220 10606 31248 10950
rect 31496 10674 31524 11086
rect 31588 10962 31616 11630
rect 31668 11076 31720 11082
rect 31720 11036 31800 11064
rect 31668 11018 31720 11024
rect 31588 10934 31708 10962
rect 31484 10668 31536 10674
rect 31484 10610 31536 10616
rect 31208 10600 31260 10606
rect 31208 10542 31260 10548
rect 31024 10532 31076 10538
rect 31024 10474 31076 10480
rect 31036 10130 31064 10474
rect 31024 10124 31076 10130
rect 31024 10066 31076 10072
rect 31220 10044 31248 10542
rect 31496 10266 31524 10610
rect 31484 10260 31536 10266
rect 31484 10202 31536 10208
rect 31300 10056 31352 10062
rect 31220 10016 31300 10044
rect 31300 9998 31352 10004
rect 31576 10056 31628 10062
rect 31576 9998 31628 10004
rect 31312 8537 31340 9998
rect 31484 9716 31536 9722
rect 31484 9658 31536 9664
rect 31392 9512 31444 9518
rect 31392 9454 31444 9460
rect 31298 8528 31354 8537
rect 31404 8498 31432 9454
rect 31298 8463 31354 8472
rect 31392 8492 31444 8498
rect 31392 8434 31444 8440
rect 31208 8424 31260 8430
rect 31208 8366 31260 8372
rect 30932 8084 30984 8090
rect 30932 8026 30984 8032
rect 30656 7744 30708 7750
rect 30656 7686 30708 7692
rect 30944 7410 30972 8026
rect 31022 7848 31078 7857
rect 31022 7783 31078 7792
rect 30656 7404 30708 7410
rect 30576 7364 30656 7392
rect 30472 7346 30524 7352
rect 30656 7346 30708 7352
rect 30932 7404 30984 7410
rect 30932 7346 30984 7352
rect 30380 7268 30432 7274
rect 30380 7210 30432 7216
rect 30380 6860 30432 6866
rect 30380 6802 30432 6808
rect 30288 6792 30340 6798
rect 30288 6734 30340 6740
rect 30392 6633 30420 6802
rect 30668 6798 30696 7346
rect 30748 7200 30800 7206
rect 30748 7142 30800 7148
rect 30656 6792 30708 6798
rect 30656 6734 30708 6740
rect 30378 6624 30434 6633
rect 30378 6559 30434 6568
rect 30760 5710 30788 7142
rect 30840 6112 30892 6118
rect 30840 6054 30892 6060
rect 30852 5778 30880 6054
rect 30840 5772 30892 5778
rect 30840 5714 30892 5720
rect 30748 5704 30800 5710
rect 30748 5646 30800 5652
rect 30012 5636 30064 5642
rect 30012 5578 30064 5584
rect 29920 5568 29972 5574
rect 29920 5510 29972 5516
rect 29932 5234 29960 5510
rect 29920 5228 29972 5234
rect 29920 5170 29972 5176
rect 30024 4690 30052 5578
rect 31036 5234 31064 7783
rect 31220 7410 31248 8366
rect 31208 7404 31260 7410
rect 31208 7346 31260 7352
rect 31496 7290 31524 9658
rect 31588 9654 31616 9998
rect 31576 9648 31628 9654
rect 31576 9590 31628 9596
rect 31680 9500 31708 10934
rect 31772 10810 31800 11036
rect 31760 10804 31812 10810
rect 31760 10746 31812 10752
rect 31588 9472 31708 9500
rect 31588 7886 31616 9472
rect 31668 9104 31720 9110
rect 31772 9058 31800 10746
rect 31864 10198 31892 13126
rect 31852 10192 31904 10198
rect 31852 10134 31904 10140
rect 31852 9920 31904 9926
rect 31852 9862 31904 9868
rect 31864 9586 31892 9862
rect 31852 9580 31904 9586
rect 31852 9522 31904 9528
rect 31956 9058 31984 14368
rect 32048 14006 32076 14606
rect 32128 14272 32180 14278
rect 32128 14214 32180 14220
rect 32036 14000 32088 14006
rect 32036 13942 32088 13948
rect 32048 11830 32076 13942
rect 32140 13734 32168 14214
rect 32128 13728 32180 13734
rect 32128 13670 32180 13676
rect 32232 13190 32260 14826
rect 32508 14414 32536 18566
rect 32600 17814 32628 18770
rect 32692 18426 32720 18838
rect 32772 18760 32824 18766
rect 32772 18702 32824 18708
rect 32680 18420 32732 18426
rect 32680 18362 32732 18368
rect 32784 18290 32812 18702
rect 32772 18284 32824 18290
rect 32772 18226 32824 18232
rect 32588 17808 32640 17814
rect 32588 17750 32640 17756
rect 32588 17060 32640 17066
rect 32588 17002 32640 17008
rect 32600 15502 32628 17002
rect 32680 16516 32732 16522
rect 32680 16458 32732 16464
rect 32588 15496 32640 15502
rect 32588 15438 32640 15444
rect 32404 14408 32456 14414
rect 32404 14350 32456 14356
rect 32496 14408 32548 14414
rect 32496 14350 32548 14356
rect 32312 13252 32364 13258
rect 32312 13194 32364 13200
rect 32220 13184 32272 13190
rect 32220 13126 32272 13132
rect 32128 12980 32180 12986
rect 32128 12922 32180 12928
rect 32036 11824 32088 11830
rect 32036 11766 32088 11772
rect 32036 11144 32088 11150
rect 32036 11086 32088 11092
rect 32048 10674 32076 11086
rect 32036 10668 32088 10674
rect 32036 10610 32088 10616
rect 32048 9926 32076 10610
rect 32140 10538 32168 12922
rect 32324 12646 32352 13194
rect 32312 12640 32364 12646
rect 32312 12582 32364 12588
rect 32324 12442 32352 12582
rect 32312 12436 32364 12442
rect 32312 12378 32364 12384
rect 32416 12345 32444 14350
rect 32600 14226 32628 15438
rect 32692 14890 32720 16458
rect 32876 16182 32904 20742
rect 32956 19304 33008 19310
rect 32956 19246 33008 19252
rect 32968 19174 32996 19246
rect 32956 19168 33008 19174
rect 32956 19110 33008 19116
rect 32968 18204 32996 19110
rect 33060 18358 33088 25214
rect 33152 24818 33180 26540
rect 33244 26382 33272 27270
rect 33336 26994 33364 27406
rect 33414 27367 33470 27376
rect 33520 27334 33548 29582
rect 33704 29238 33732 34546
rect 33888 34406 33916 35974
rect 33980 35086 34008 35974
rect 34164 35494 34192 36110
rect 34520 35692 34572 35698
rect 34520 35634 34572 35640
rect 34244 35624 34296 35630
rect 34244 35566 34296 35572
rect 34152 35488 34204 35494
rect 34152 35430 34204 35436
rect 33968 35080 34020 35086
rect 33968 35022 34020 35028
rect 34060 34944 34112 34950
rect 34060 34886 34112 34892
rect 34072 34785 34100 34886
rect 34058 34776 34114 34785
rect 33968 34740 34020 34746
rect 34058 34711 34114 34720
rect 33968 34682 34020 34688
rect 33876 34400 33928 34406
rect 33876 34342 33928 34348
rect 33782 34232 33838 34241
rect 33782 34167 33784 34176
rect 33836 34167 33838 34176
rect 33784 34138 33836 34144
rect 33784 33856 33836 33862
rect 33784 33798 33836 33804
rect 33796 33590 33824 33798
rect 33784 33584 33836 33590
rect 33784 33526 33836 33532
rect 33888 32570 33916 34342
rect 33980 33522 34008 34682
rect 33968 33516 34020 33522
rect 33968 33458 34020 33464
rect 34072 32774 34100 34711
rect 34164 34610 34192 35430
rect 34256 35222 34284 35566
rect 34336 35488 34388 35494
rect 34336 35430 34388 35436
rect 34244 35216 34296 35222
rect 34244 35158 34296 35164
rect 34348 35086 34376 35430
rect 34336 35080 34388 35086
rect 34336 35022 34388 35028
rect 34152 34604 34204 34610
rect 34152 34546 34204 34552
rect 34164 32910 34192 34546
rect 34532 33998 34560 35634
rect 34704 35488 34756 35494
rect 34704 35430 34756 35436
rect 34716 35290 34744 35430
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34704 35284 34756 35290
rect 34704 35226 34756 35232
rect 34520 33992 34572 33998
rect 34520 33934 34572 33940
rect 34336 33380 34388 33386
rect 34336 33322 34388 33328
rect 34152 32904 34204 32910
rect 34152 32846 34204 32852
rect 34060 32768 34112 32774
rect 34060 32710 34112 32716
rect 33876 32564 33928 32570
rect 33876 32506 33928 32512
rect 33968 31816 34020 31822
rect 33968 31758 34020 31764
rect 33784 31680 33836 31686
rect 33876 31680 33928 31686
rect 33784 31622 33836 31628
rect 33874 31648 33876 31657
rect 33928 31648 33930 31657
rect 33796 31414 33824 31622
rect 33874 31583 33930 31592
rect 33876 31476 33928 31482
rect 33876 31418 33928 31424
rect 33784 31408 33836 31414
rect 33784 31350 33836 31356
rect 33782 31104 33838 31113
rect 33888 31090 33916 31418
rect 33980 31278 34008 31758
rect 34072 31346 34100 32710
rect 34060 31340 34112 31346
rect 34060 31282 34112 31288
rect 33968 31272 34020 31278
rect 34164 31226 34192 32846
rect 34244 32360 34296 32366
rect 34244 32302 34296 32308
rect 34256 31822 34284 32302
rect 34244 31816 34296 31822
rect 34244 31758 34296 31764
rect 34348 31657 34376 33322
rect 34428 32496 34480 32502
rect 34428 32438 34480 32444
rect 34440 31958 34468 32438
rect 34428 31952 34480 31958
rect 34428 31894 34480 31900
rect 34334 31648 34390 31657
rect 34334 31583 34390 31592
rect 34242 31376 34298 31385
rect 34242 31311 34298 31320
rect 34256 31278 34284 31311
rect 34348 31278 34376 31583
rect 34440 31278 34468 31894
rect 34532 31686 34560 33934
rect 34612 33856 34664 33862
rect 34612 33798 34664 33804
rect 34624 32745 34652 33798
rect 34610 32736 34666 32745
rect 34610 32671 34666 32680
rect 34612 32224 34664 32230
rect 34612 32166 34664 32172
rect 34624 32026 34652 32166
rect 34612 32020 34664 32026
rect 34612 31962 34664 31968
rect 34612 31816 34664 31822
rect 34610 31784 34612 31793
rect 34664 31784 34666 31793
rect 34610 31719 34666 31728
rect 34520 31680 34572 31686
rect 34520 31622 34572 31628
rect 34716 31498 34744 35226
rect 35348 34740 35400 34746
rect 35348 34682 35400 34688
rect 34796 34468 34848 34474
rect 34796 34410 34848 34416
rect 34808 34066 34836 34410
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34796 34060 34848 34066
rect 34796 34002 34848 34008
rect 34888 33992 34940 33998
rect 34888 33934 34940 33940
rect 34900 33658 34928 33934
rect 35360 33862 35388 34682
rect 35532 34536 35584 34542
rect 35532 34478 35584 34484
rect 35440 34468 35492 34474
rect 35440 34410 35492 34416
rect 35452 34134 35480 34410
rect 35440 34128 35492 34134
rect 35440 34070 35492 34076
rect 35348 33856 35400 33862
rect 35348 33798 35400 33804
rect 35440 33856 35492 33862
rect 35440 33798 35492 33804
rect 35360 33658 35388 33798
rect 34888 33652 34940 33658
rect 34888 33594 34940 33600
rect 35348 33652 35400 33658
rect 35348 33594 35400 33600
rect 34900 33402 34928 33594
rect 34808 33374 34928 33402
rect 34808 32910 34836 33374
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34796 32904 34848 32910
rect 34796 32846 34848 32852
rect 35348 32768 35400 32774
rect 35348 32710 35400 32716
rect 34796 32564 34848 32570
rect 34796 32506 34848 32512
rect 34624 31470 34744 31498
rect 33968 31214 34020 31220
rect 33838 31062 33916 31090
rect 33782 31039 33838 31048
rect 33876 30592 33928 30598
rect 33876 30534 33928 30540
rect 33888 30433 33916 30534
rect 33874 30424 33930 30433
rect 33874 30359 33930 30368
rect 33876 30048 33928 30054
rect 33876 29990 33928 29996
rect 33692 29232 33744 29238
rect 33692 29174 33744 29180
rect 33600 28960 33652 28966
rect 33600 28902 33652 28908
rect 33508 27328 33560 27334
rect 33414 27296 33470 27305
rect 33508 27270 33560 27276
rect 33414 27231 33470 27240
rect 33428 27130 33456 27231
rect 33416 27124 33468 27130
rect 33416 27066 33468 27072
rect 33324 26988 33376 26994
rect 33376 26948 33456 26976
rect 33324 26930 33376 26936
rect 33232 26376 33284 26382
rect 33232 26318 33284 26324
rect 33428 25906 33456 26948
rect 33506 26888 33562 26897
rect 33506 26823 33562 26832
rect 33520 26518 33548 26823
rect 33508 26512 33560 26518
rect 33508 26454 33560 26460
rect 33508 26376 33560 26382
rect 33508 26318 33560 26324
rect 33416 25900 33468 25906
rect 33416 25842 33468 25848
rect 33232 25832 33284 25838
rect 33232 25774 33284 25780
rect 33140 24812 33192 24818
rect 33140 24754 33192 24760
rect 33152 23746 33180 24754
rect 33244 24070 33272 25774
rect 33324 25288 33376 25294
rect 33324 25230 33376 25236
rect 33336 25106 33364 25230
rect 33414 25120 33470 25129
rect 33336 25078 33414 25106
rect 33414 25055 33470 25064
rect 33416 24744 33468 24750
rect 33322 24712 33378 24721
rect 33416 24686 33468 24692
rect 33322 24647 33378 24656
rect 33336 24274 33364 24647
rect 33324 24268 33376 24274
rect 33324 24210 33376 24216
rect 33322 24168 33378 24177
rect 33322 24103 33378 24112
rect 33232 24064 33284 24070
rect 33232 24006 33284 24012
rect 33152 23718 33272 23746
rect 33244 23118 33272 23718
rect 33232 23112 33284 23118
rect 33232 23054 33284 23060
rect 33244 22642 33272 23054
rect 33232 22636 33284 22642
rect 33232 22578 33284 22584
rect 33232 22500 33284 22506
rect 33232 22442 33284 22448
rect 33140 21548 33192 21554
rect 33140 21490 33192 21496
rect 33152 20942 33180 21490
rect 33140 20936 33192 20942
rect 33140 20878 33192 20884
rect 33140 19712 33192 19718
rect 33140 19654 33192 19660
rect 33152 19514 33180 19654
rect 33140 19508 33192 19514
rect 33140 19450 33192 19456
rect 33140 19168 33192 19174
rect 33140 19110 33192 19116
rect 33152 18766 33180 19110
rect 33140 18760 33192 18766
rect 33140 18702 33192 18708
rect 33140 18624 33192 18630
rect 33138 18592 33140 18601
rect 33192 18592 33194 18601
rect 33138 18527 33194 18536
rect 33048 18352 33100 18358
rect 33048 18294 33100 18300
rect 32968 18176 33180 18204
rect 33048 18080 33100 18086
rect 33048 18022 33100 18028
rect 32956 17332 33008 17338
rect 32956 17274 33008 17280
rect 32864 16176 32916 16182
rect 32864 16118 32916 16124
rect 32864 15020 32916 15026
rect 32864 14962 32916 14968
rect 32772 14952 32824 14958
rect 32772 14894 32824 14900
rect 32680 14884 32732 14890
rect 32680 14826 32732 14832
rect 32784 14793 32812 14894
rect 32770 14784 32826 14793
rect 32770 14719 32826 14728
rect 32508 14198 32628 14226
rect 32772 14272 32824 14278
rect 32772 14214 32824 14220
rect 32508 13802 32536 14198
rect 32588 14068 32640 14074
rect 32588 14010 32640 14016
rect 32600 13841 32628 14010
rect 32680 13932 32732 13938
rect 32680 13874 32732 13880
rect 32586 13832 32642 13841
rect 32496 13796 32548 13802
rect 32586 13767 32642 13776
rect 32496 13738 32548 13744
rect 32508 12918 32536 13738
rect 32692 13394 32720 13874
rect 32680 13388 32732 13394
rect 32680 13330 32732 13336
rect 32586 13016 32642 13025
rect 32586 12951 32588 12960
rect 32640 12951 32642 12960
rect 32588 12922 32640 12928
rect 32692 12918 32720 13330
rect 32496 12912 32548 12918
rect 32496 12854 32548 12860
rect 32680 12912 32732 12918
rect 32680 12854 32732 12860
rect 32402 12336 32458 12345
rect 32312 12300 32364 12306
rect 32402 12271 32458 12280
rect 32312 12242 32364 12248
rect 32324 11898 32352 12242
rect 32312 11892 32364 11898
rect 32312 11834 32364 11840
rect 32416 11778 32444 12271
rect 32508 12170 32536 12854
rect 32680 12776 32732 12782
rect 32680 12718 32732 12724
rect 32588 12232 32640 12238
rect 32588 12174 32640 12180
rect 32496 12164 32548 12170
rect 32496 12106 32548 12112
rect 32232 11750 32444 11778
rect 32128 10532 32180 10538
rect 32128 10474 32180 10480
rect 32140 10062 32168 10474
rect 32128 10056 32180 10062
rect 32128 9998 32180 10004
rect 32036 9920 32088 9926
rect 32036 9862 32088 9868
rect 32036 9376 32088 9382
rect 32036 9318 32088 9324
rect 31720 9052 31800 9058
rect 31668 9046 31800 9052
rect 31680 9030 31800 9046
rect 31666 8528 31722 8537
rect 31666 8463 31668 8472
rect 31720 8463 31722 8472
rect 31668 8434 31720 8440
rect 31680 8362 31708 8434
rect 31772 8412 31800 9030
rect 31864 9030 31984 9058
rect 31864 8974 31892 9030
rect 32048 8974 32076 9318
rect 31852 8968 31904 8974
rect 31852 8910 31904 8916
rect 32036 8968 32088 8974
rect 32232 8922 32260 11750
rect 32404 11620 32456 11626
rect 32324 11580 32404 11608
rect 32324 10010 32352 11580
rect 32404 11562 32456 11568
rect 32404 10736 32456 10742
rect 32404 10678 32456 10684
rect 32416 10130 32444 10678
rect 32496 10192 32548 10198
rect 32496 10134 32548 10140
rect 32404 10124 32456 10130
rect 32404 10066 32456 10072
rect 32324 9982 32444 10010
rect 32312 9920 32364 9926
rect 32312 9862 32364 9868
rect 32324 9450 32352 9862
rect 32312 9444 32364 9450
rect 32312 9386 32364 9392
rect 32324 8974 32352 9386
rect 32036 8910 32088 8916
rect 32048 8566 32076 8910
rect 32140 8894 32260 8922
rect 32312 8968 32364 8974
rect 32312 8910 32364 8916
rect 32036 8560 32088 8566
rect 32036 8502 32088 8508
rect 32036 8424 32088 8430
rect 31772 8384 32036 8412
rect 32036 8366 32088 8372
rect 31668 8356 31720 8362
rect 31668 8298 31720 8304
rect 32036 8016 32088 8022
rect 32036 7958 32088 7964
rect 31576 7880 31628 7886
rect 31576 7822 31628 7828
rect 31588 7478 31616 7822
rect 32048 7478 32076 7958
rect 32140 7834 32168 8894
rect 32220 8832 32272 8838
rect 32220 8774 32272 8780
rect 32232 8498 32260 8774
rect 32220 8492 32272 8498
rect 32220 8434 32272 8440
rect 32416 8090 32444 9982
rect 32508 8401 32536 10134
rect 32494 8392 32550 8401
rect 32494 8327 32550 8336
rect 32404 8084 32456 8090
rect 32404 8026 32456 8032
rect 32140 7806 32260 7834
rect 32128 7744 32180 7750
rect 32128 7686 32180 7692
rect 32140 7478 32168 7686
rect 31576 7472 31628 7478
rect 31576 7414 31628 7420
rect 32036 7472 32088 7478
rect 32036 7414 32088 7420
rect 32128 7472 32180 7478
rect 32128 7414 32180 7420
rect 31668 7404 31720 7410
rect 31668 7346 31720 7352
rect 31220 7262 31524 7290
rect 31220 7206 31248 7262
rect 31208 7200 31260 7206
rect 31208 7142 31260 7148
rect 31300 7200 31352 7206
rect 31300 7142 31352 7148
rect 31312 6798 31340 7142
rect 31496 6866 31524 7262
rect 31680 6934 31708 7346
rect 32036 7336 32088 7342
rect 32036 7278 32088 7284
rect 32048 7002 32076 7278
rect 32128 7200 32180 7206
rect 32128 7142 32180 7148
rect 32036 6996 32088 7002
rect 32036 6938 32088 6944
rect 31668 6928 31720 6934
rect 31668 6870 31720 6876
rect 32140 6866 32168 7142
rect 32232 7002 32260 7806
rect 32416 7290 32444 8026
rect 32508 7478 32536 8327
rect 32600 8276 32628 12174
rect 32692 10470 32720 12718
rect 32784 12170 32812 14214
rect 32876 13870 32904 14962
rect 32864 13864 32916 13870
rect 32864 13806 32916 13812
rect 32864 13524 32916 13530
rect 32864 13466 32916 13472
rect 32876 12850 32904 13466
rect 32968 12986 32996 17274
rect 33060 16658 33088 18022
rect 33048 16652 33100 16658
rect 33048 16594 33100 16600
rect 33152 14906 33180 18176
rect 33244 15094 33272 22442
rect 33336 22166 33364 24103
rect 33324 22160 33376 22166
rect 33324 22102 33376 22108
rect 33324 21956 33376 21962
rect 33324 21898 33376 21904
rect 33336 19718 33364 21898
rect 33428 20806 33456 24686
rect 33520 24342 33548 26318
rect 33612 25809 33640 28902
rect 33704 28626 33732 29174
rect 33692 28620 33744 28626
rect 33692 28562 33744 28568
rect 33784 27872 33836 27878
rect 33784 27814 33836 27820
rect 33796 27713 33824 27814
rect 33782 27704 33838 27713
rect 33782 27639 33838 27648
rect 33692 27328 33744 27334
rect 33692 27270 33744 27276
rect 33704 26926 33732 27270
rect 33796 27130 33824 27639
rect 33784 27124 33836 27130
rect 33784 27066 33836 27072
rect 33692 26920 33744 26926
rect 33692 26862 33744 26868
rect 33692 26240 33744 26246
rect 33692 26182 33744 26188
rect 33598 25800 33654 25809
rect 33598 25735 33654 25744
rect 33612 25362 33640 25735
rect 33600 25356 33652 25362
rect 33600 25298 33652 25304
rect 33598 25256 33654 25265
rect 33598 25191 33600 25200
rect 33652 25191 33654 25200
rect 33600 25162 33652 25168
rect 33600 24608 33652 24614
rect 33600 24550 33652 24556
rect 33612 24410 33640 24550
rect 33600 24404 33652 24410
rect 33600 24346 33652 24352
rect 33508 24336 33560 24342
rect 33508 24278 33560 24284
rect 33612 23474 33640 24346
rect 33704 23730 33732 26182
rect 33692 23724 33744 23730
rect 33692 23666 33744 23672
rect 33612 23446 33732 23474
rect 33508 22976 33560 22982
rect 33508 22918 33560 22924
rect 33416 20800 33468 20806
rect 33416 20742 33468 20748
rect 33428 20534 33456 20742
rect 33416 20528 33468 20534
rect 33416 20470 33468 20476
rect 33416 20256 33468 20262
rect 33416 20198 33468 20204
rect 33428 19922 33456 20198
rect 33416 19916 33468 19922
rect 33416 19858 33468 19864
rect 33520 19802 33548 22918
rect 33416 19780 33468 19786
rect 33520 19774 33640 19802
rect 33416 19722 33468 19728
rect 33324 19712 33376 19718
rect 33324 19654 33376 19660
rect 33232 15088 33284 15094
rect 33232 15030 33284 15036
rect 33152 14878 33272 14906
rect 33140 14816 33192 14822
rect 33140 14758 33192 14764
rect 33152 13938 33180 14758
rect 33140 13932 33192 13938
rect 33140 13874 33192 13880
rect 32956 12980 33008 12986
rect 32956 12922 33008 12928
rect 33048 12980 33100 12986
rect 33048 12922 33100 12928
rect 32864 12844 32916 12850
rect 32864 12786 32916 12792
rect 32956 12708 33008 12714
rect 32956 12650 33008 12656
rect 32772 12164 32824 12170
rect 32772 12106 32824 12112
rect 32968 11218 32996 12650
rect 33060 12442 33088 12922
rect 33152 12850 33180 13874
rect 33244 13802 33272 14878
rect 33232 13796 33284 13802
rect 33232 13738 33284 13744
rect 33232 13456 33284 13462
rect 33232 13398 33284 13404
rect 33140 12844 33192 12850
rect 33140 12786 33192 12792
rect 33244 12730 33272 13398
rect 33336 13258 33364 19654
rect 33428 19378 33456 19722
rect 33612 19446 33640 19774
rect 33600 19440 33652 19446
rect 33598 19408 33600 19417
rect 33652 19408 33654 19417
rect 33416 19372 33468 19378
rect 33598 19343 33654 19352
rect 33416 19314 33468 19320
rect 33428 18698 33456 19314
rect 33508 19304 33560 19310
rect 33704 19292 33732 23446
rect 33796 22506 33824 27066
rect 33888 26994 33916 29990
rect 33980 28422 34008 31214
rect 34072 31198 34192 31226
rect 34244 31272 34296 31278
rect 34244 31214 34296 31220
rect 34336 31272 34388 31278
rect 34336 31214 34388 31220
rect 34428 31272 34480 31278
rect 34428 31214 34480 31220
rect 34072 30734 34100 31198
rect 34348 31124 34376 31214
rect 34256 31096 34376 31124
rect 34060 30728 34112 30734
rect 34060 30670 34112 30676
rect 34060 29504 34112 29510
rect 34060 29446 34112 29452
rect 34072 29073 34100 29446
rect 34058 29064 34114 29073
rect 34058 28999 34114 29008
rect 34152 28552 34204 28558
rect 34152 28494 34204 28500
rect 33968 28416 34020 28422
rect 33968 28358 34020 28364
rect 33968 28008 34020 28014
rect 33968 27950 34020 27956
rect 33980 27334 34008 27950
rect 34060 27464 34112 27470
rect 34060 27406 34112 27412
rect 33968 27328 34020 27334
rect 33968 27270 34020 27276
rect 33876 26988 33928 26994
rect 33876 26930 33928 26936
rect 33888 24585 33916 26930
rect 34072 26382 34100 27406
rect 34060 26376 34112 26382
rect 34060 26318 34112 26324
rect 34164 26194 34192 28494
rect 34256 26994 34284 31096
rect 34336 29776 34388 29782
rect 34336 29718 34388 29724
rect 34348 29646 34376 29718
rect 34336 29640 34388 29646
rect 34336 29582 34388 29588
rect 34348 28694 34376 29582
rect 34440 29170 34468 31214
rect 34520 30592 34572 30598
rect 34520 30534 34572 30540
rect 34428 29164 34480 29170
rect 34428 29106 34480 29112
rect 34336 28688 34388 28694
rect 34336 28630 34388 28636
rect 34532 28626 34560 30534
rect 34624 30274 34652 31470
rect 34704 31408 34756 31414
rect 34704 31350 34756 31356
rect 34716 30666 34744 31350
rect 34808 31278 34836 32506
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35360 32026 35388 32710
rect 35452 32337 35480 33798
rect 35438 32328 35494 32337
rect 35438 32263 35494 32272
rect 35348 32020 35400 32026
rect 35348 31962 35400 31968
rect 34888 31816 34940 31822
rect 35348 31816 35400 31822
rect 34888 31758 34940 31764
rect 35346 31784 35348 31793
rect 35400 31784 35402 31793
rect 34900 31482 34928 31758
rect 34980 31748 35032 31754
rect 35346 31719 35402 31728
rect 34980 31690 35032 31696
rect 34888 31476 34940 31482
rect 34888 31418 34940 31424
rect 34992 31346 35020 31690
rect 35348 31680 35400 31686
rect 35348 31622 35400 31628
rect 34980 31340 35032 31346
rect 34980 31282 35032 31288
rect 34796 31272 34848 31278
rect 34796 31214 34848 31220
rect 34808 30802 34836 31214
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34796 30796 34848 30802
rect 34796 30738 34848 30744
rect 34704 30660 34756 30666
rect 34704 30602 34756 30608
rect 34794 30560 34850 30569
rect 34794 30495 34850 30504
rect 34624 30246 34744 30274
rect 34612 30116 34664 30122
rect 34612 30058 34664 30064
rect 34520 28620 34572 28626
rect 34520 28562 34572 28568
rect 34624 28393 34652 30058
rect 34716 30054 34744 30246
rect 34808 30190 34836 30495
rect 34796 30184 34848 30190
rect 34796 30126 34848 30132
rect 34704 30048 34756 30054
rect 34704 29990 34756 29996
rect 34716 29646 34744 29990
rect 34704 29640 34756 29646
rect 34704 29582 34756 29588
rect 34704 28688 34756 28694
rect 34704 28630 34756 28636
rect 34610 28384 34666 28393
rect 34610 28319 34666 28328
rect 34336 28212 34388 28218
rect 34336 28154 34388 28160
rect 34348 27010 34376 28154
rect 34520 28076 34572 28082
rect 34520 28018 34572 28024
rect 34428 27396 34480 27402
rect 34428 27338 34480 27344
rect 34440 27305 34468 27338
rect 34426 27296 34482 27305
rect 34426 27231 34482 27240
rect 34244 26988 34296 26994
rect 34348 26982 34468 27010
rect 34244 26930 34296 26936
rect 34256 26450 34284 26930
rect 34440 26790 34468 26982
rect 34428 26784 34480 26790
rect 34428 26726 34480 26732
rect 34244 26444 34296 26450
rect 34244 26386 34296 26392
rect 34440 26353 34468 26726
rect 34426 26344 34482 26353
rect 34426 26279 34482 26288
rect 34072 26166 34192 26194
rect 33968 25424 34020 25430
rect 33968 25366 34020 25372
rect 33980 24886 34008 25366
rect 33968 24880 34020 24886
rect 33968 24822 34020 24828
rect 33874 24576 33930 24585
rect 33874 24511 33930 24520
rect 33876 24336 33928 24342
rect 33876 24278 33928 24284
rect 33888 23730 33916 24278
rect 33980 24206 34008 24822
rect 34072 24818 34100 26166
rect 34244 26036 34296 26042
rect 34244 25978 34296 25984
rect 34336 26036 34388 26042
rect 34336 25978 34388 25984
rect 34256 25362 34284 25978
rect 34244 25356 34296 25362
rect 34244 25298 34296 25304
rect 34152 25288 34204 25294
rect 34152 25230 34204 25236
rect 34242 25256 34298 25265
rect 34060 24812 34112 24818
rect 34060 24754 34112 24760
rect 34164 24721 34192 25230
rect 34348 25242 34376 25978
rect 34426 25392 34482 25401
rect 34426 25327 34482 25336
rect 34298 25214 34376 25242
rect 34242 25191 34298 25200
rect 34336 24880 34388 24886
rect 34336 24822 34388 24828
rect 34244 24744 34296 24750
rect 34150 24712 34206 24721
rect 34244 24686 34296 24692
rect 34150 24647 34206 24656
rect 34152 24336 34204 24342
rect 34152 24278 34204 24284
rect 33968 24200 34020 24206
rect 33968 24142 34020 24148
rect 34060 23860 34112 23866
rect 34060 23802 34112 23808
rect 33876 23724 33928 23730
rect 33876 23666 33928 23672
rect 34072 23526 34100 23802
rect 34060 23520 34112 23526
rect 34060 23462 34112 23468
rect 34060 22704 34112 22710
rect 34060 22646 34112 22652
rect 33876 22568 33928 22574
rect 33876 22510 33928 22516
rect 33784 22500 33836 22506
rect 33784 22442 33836 22448
rect 33888 22030 33916 22510
rect 33876 22024 33928 22030
rect 33796 21984 33876 22012
rect 33796 20262 33824 21984
rect 33876 21966 33928 21972
rect 33968 21956 34020 21962
rect 33968 21898 34020 21904
rect 33876 20800 33928 20806
rect 33876 20742 33928 20748
rect 33784 20256 33836 20262
rect 33784 20198 33836 20204
rect 33784 19984 33836 19990
rect 33784 19926 33836 19932
rect 33796 19854 33824 19926
rect 33888 19854 33916 20742
rect 33784 19848 33836 19854
rect 33784 19790 33836 19796
rect 33876 19848 33928 19854
rect 33876 19790 33928 19796
rect 33784 19372 33836 19378
rect 33784 19314 33836 19320
rect 33560 19264 33732 19292
rect 33508 19246 33560 19252
rect 33796 19224 33824 19314
rect 33704 19196 33824 19224
rect 33704 18698 33732 19196
rect 33416 18692 33468 18698
rect 33416 18634 33468 18640
rect 33692 18692 33744 18698
rect 33692 18634 33744 18640
rect 33428 18290 33456 18634
rect 33508 18624 33560 18630
rect 33508 18566 33560 18572
rect 33520 18358 33548 18566
rect 33508 18352 33560 18358
rect 33508 18294 33560 18300
rect 33416 18284 33468 18290
rect 33416 18226 33468 18232
rect 33414 18184 33470 18193
rect 33414 18119 33470 18128
rect 33428 17134 33456 18119
rect 33704 17762 33732 18634
rect 33782 18456 33838 18465
rect 33782 18391 33838 18400
rect 33796 17814 33824 18391
rect 33980 18358 34008 21898
rect 34072 21690 34100 22646
rect 34060 21684 34112 21690
rect 34060 21626 34112 21632
rect 34060 20392 34112 20398
rect 34060 20334 34112 20340
rect 34072 20058 34100 20334
rect 34164 20330 34192 24278
rect 34152 20324 34204 20330
rect 34152 20266 34204 20272
rect 34060 20052 34112 20058
rect 34060 19994 34112 20000
rect 34164 19922 34192 20266
rect 34060 19916 34112 19922
rect 34060 19858 34112 19864
rect 34152 19916 34204 19922
rect 34152 19858 34204 19864
rect 34072 19786 34100 19858
rect 34060 19780 34112 19786
rect 34060 19722 34112 19728
rect 34152 19780 34204 19786
rect 34152 19722 34204 19728
rect 34072 19145 34100 19722
rect 34164 19446 34192 19722
rect 34152 19440 34204 19446
rect 34152 19382 34204 19388
rect 34058 19136 34114 19145
rect 34058 19071 34114 19080
rect 34060 18964 34112 18970
rect 34060 18906 34112 18912
rect 34072 18766 34100 18906
rect 34060 18760 34112 18766
rect 34060 18702 34112 18708
rect 33968 18352 34020 18358
rect 33968 18294 34020 18300
rect 33876 18080 33928 18086
rect 33876 18022 33928 18028
rect 33612 17734 33732 17762
rect 33784 17808 33836 17814
rect 33784 17750 33836 17756
rect 33612 17610 33640 17734
rect 33692 17672 33744 17678
rect 33692 17614 33744 17620
rect 33784 17672 33836 17678
rect 33784 17614 33836 17620
rect 33600 17604 33652 17610
rect 33600 17546 33652 17552
rect 33508 17536 33560 17542
rect 33508 17478 33560 17484
rect 33520 17241 33548 17478
rect 33506 17232 33562 17241
rect 33506 17167 33562 17176
rect 33416 17128 33468 17134
rect 33416 17070 33468 17076
rect 33506 17096 33562 17105
rect 33506 17031 33562 17040
rect 33520 16998 33548 17031
rect 33508 16992 33560 16998
rect 33508 16934 33560 16940
rect 33414 16688 33470 16697
rect 33414 16623 33416 16632
rect 33468 16623 33470 16632
rect 33508 16652 33560 16658
rect 33416 16594 33468 16600
rect 33508 16594 33560 16600
rect 33416 16516 33468 16522
rect 33416 16458 33468 16464
rect 33428 16250 33456 16458
rect 33416 16244 33468 16250
rect 33416 16186 33468 16192
rect 33416 14408 33468 14414
rect 33416 14350 33468 14356
rect 33324 13252 33376 13258
rect 33324 13194 33376 13200
rect 33152 12702 33272 12730
rect 33048 12436 33100 12442
rect 33048 12378 33100 12384
rect 33152 12374 33180 12702
rect 33140 12368 33192 12374
rect 33140 12310 33192 12316
rect 33152 12170 33180 12310
rect 33140 12164 33192 12170
rect 33140 12106 33192 12112
rect 33152 11626 33180 12106
rect 33140 11620 33192 11626
rect 33140 11562 33192 11568
rect 32956 11212 33008 11218
rect 32956 11154 33008 11160
rect 33336 11098 33364 13194
rect 32876 11082 33364 11098
rect 32876 11076 33376 11082
rect 32876 11070 33324 11076
rect 32876 10826 32904 11070
rect 33324 11018 33376 11024
rect 32956 11008 33008 11014
rect 32956 10950 33008 10956
rect 33140 11008 33192 11014
rect 33140 10950 33192 10956
rect 32784 10798 32904 10826
rect 32784 10742 32812 10798
rect 32772 10736 32824 10742
rect 32772 10678 32824 10684
rect 32968 10674 32996 10950
rect 33046 10840 33102 10849
rect 33046 10775 33048 10784
rect 33100 10775 33102 10784
rect 33048 10746 33100 10752
rect 32956 10668 33008 10674
rect 32956 10610 33008 10616
rect 32680 10464 32732 10470
rect 32680 10406 32732 10412
rect 32692 10266 32720 10406
rect 32680 10260 32732 10266
rect 32680 10202 32732 10208
rect 32692 9178 32720 10202
rect 33152 9926 33180 10950
rect 33140 9920 33192 9926
rect 33140 9862 33192 9868
rect 33152 9722 33180 9862
rect 33140 9716 33192 9722
rect 33140 9658 33192 9664
rect 33428 9586 33456 14350
rect 33520 12442 33548 16594
rect 33612 15502 33640 17546
rect 33600 15496 33652 15502
rect 33600 15438 33652 15444
rect 33600 15020 33652 15026
rect 33600 14962 33652 14968
rect 33612 14278 33640 14962
rect 33704 14618 33732 17614
rect 33796 17134 33824 17614
rect 33888 17542 33916 18022
rect 33876 17536 33928 17542
rect 33876 17478 33928 17484
rect 33784 17128 33836 17134
rect 33784 17070 33836 17076
rect 33796 16658 33824 17070
rect 33784 16652 33836 16658
rect 33784 16594 33836 16600
rect 33888 15026 33916 17478
rect 33980 16998 34008 18294
rect 34060 18216 34112 18222
rect 34060 18158 34112 18164
rect 34072 17202 34100 18158
rect 34256 17814 34284 24686
rect 34348 22094 34376 24822
rect 34440 24138 34468 25327
rect 34428 24132 34480 24138
rect 34428 24074 34480 24080
rect 34532 23798 34560 28018
rect 34624 27962 34652 28319
rect 34716 28218 34744 28630
rect 34808 28558 34836 30126
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34980 29844 35032 29850
rect 34980 29786 35032 29792
rect 34992 29646 35020 29786
rect 35254 29744 35310 29753
rect 35254 29679 35310 29688
rect 34888 29640 34940 29646
rect 34888 29582 34940 29588
rect 34980 29640 35032 29646
rect 34980 29582 35032 29588
rect 34900 29102 34928 29582
rect 34980 29504 35032 29510
rect 34980 29446 35032 29452
rect 34888 29096 34940 29102
rect 34888 29038 34940 29044
rect 34992 29034 35020 29446
rect 35164 29300 35216 29306
rect 35164 29242 35216 29248
rect 35176 29102 35204 29242
rect 35164 29096 35216 29102
rect 35164 29038 35216 29044
rect 34980 29028 35032 29034
rect 34980 28970 35032 28976
rect 35268 28966 35296 29679
rect 35256 28960 35308 28966
rect 35256 28902 35308 28908
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35360 28626 35388 31622
rect 35348 28620 35400 28626
rect 35348 28562 35400 28568
rect 34796 28552 34848 28558
rect 34796 28494 34848 28500
rect 34980 28552 35032 28558
rect 34980 28494 35032 28500
rect 34992 28422 35020 28494
rect 34980 28416 35032 28422
rect 34808 28376 34980 28404
rect 34704 28212 34756 28218
rect 34704 28154 34756 28160
rect 34702 27976 34758 27985
rect 34624 27934 34702 27962
rect 34702 27911 34758 27920
rect 34704 27872 34756 27878
rect 34704 27814 34756 27820
rect 34610 27704 34666 27713
rect 34610 27639 34666 27648
rect 34520 23792 34572 23798
rect 34518 23760 34520 23769
rect 34572 23760 34574 23769
rect 34518 23695 34574 23704
rect 34428 23520 34480 23526
rect 34428 23462 34480 23468
rect 34440 23118 34468 23462
rect 34428 23112 34480 23118
rect 34428 23054 34480 23060
rect 34520 23044 34572 23050
rect 34520 22986 34572 22992
rect 34532 22642 34560 22986
rect 34520 22636 34572 22642
rect 34520 22578 34572 22584
rect 34428 22500 34480 22506
rect 34428 22442 34480 22448
rect 34440 22216 34468 22442
rect 34440 22188 34560 22216
rect 34348 22066 34468 22094
rect 34336 22024 34388 22030
rect 34336 21966 34388 21972
rect 34348 21729 34376 21966
rect 34334 21720 34390 21729
rect 34334 21655 34390 21664
rect 34336 21616 34388 21622
rect 34336 21558 34388 21564
rect 34348 20058 34376 21558
rect 34336 20052 34388 20058
rect 34336 19994 34388 20000
rect 34336 19848 34388 19854
rect 34336 19790 34388 19796
rect 34348 18057 34376 19790
rect 34440 18834 34468 22066
rect 34532 21894 34560 22188
rect 34520 21888 34572 21894
rect 34520 21830 34572 21836
rect 34520 20800 34572 20806
rect 34520 20742 34572 20748
rect 34532 19854 34560 20742
rect 34624 20618 34652 27639
rect 34716 27470 34744 27814
rect 34808 27554 34836 28376
rect 34980 28358 35032 28364
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34808 27526 34928 27554
rect 34704 27464 34756 27470
rect 34704 27406 34756 27412
rect 34704 27328 34756 27334
rect 34704 27270 34756 27276
rect 34796 27328 34848 27334
rect 34796 27270 34848 27276
rect 34716 26858 34744 27270
rect 34704 26852 34756 26858
rect 34704 26794 34756 26800
rect 34716 24721 34744 26794
rect 34808 25838 34836 27270
rect 34900 27130 34928 27526
rect 34980 27464 35032 27470
rect 34980 27406 35032 27412
rect 35070 27432 35126 27441
rect 34888 27124 34940 27130
rect 34888 27066 34940 27072
rect 34992 27062 35020 27406
rect 35070 27367 35072 27376
rect 35124 27367 35126 27376
rect 35072 27338 35124 27344
rect 34980 27056 35032 27062
rect 34980 26998 35032 27004
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35070 26208 35126 26217
rect 35070 26143 35126 26152
rect 35084 25974 35112 26143
rect 35072 25968 35124 25974
rect 35072 25910 35124 25916
rect 35360 25838 35388 28562
rect 35452 27614 35480 32263
rect 35544 31414 35572 34478
rect 35532 31408 35584 31414
rect 35532 31350 35584 31356
rect 35532 30728 35584 30734
rect 35532 30670 35584 30676
rect 35544 29646 35572 30670
rect 35636 30172 35664 37130
rect 36084 35284 36136 35290
rect 36084 35226 36136 35232
rect 35716 34604 35768 34610
rect 35716 34546 35768 34552
rect 35728 33862 35756 34546
rect 35716 33856 35768 33862
rect 35716 33798 35768 33804
rect 35728 33522 35756 33798
rect 35716 33516 35768 33522
rect 35716 33458 35768 33464
rect 35728 33318 35756 33458
rect 35992 33448 36044 33454
rect 35992 33390 36044 33396
rect 35716 33312 35768 33318
rect 35716 33254 35768 33260
rect 36004 33114 36032 33390
rect 35992 33108 36044 33114
rect 35992 33050 36044 33056
rect 35992 32564 36044 32570
rect 35992 32506 36044 32512
rect 36004 31929 36032 32506
rect 35990 31920 36046 31929
rect 35716 31884 35768 31890
rect 35990 31855 36046 31864
rect 35716 31826 35768 31832
rect 35728 31754 35756 31826
rect 36096 31793 36124 35226
rect 36360 34944 36412 34950
rect 36360 34886 36412 34892
rect 36820 34944 36872 34950
rect 36820 34886 36872 34892
rect 36372 34610 36400 34886
rect 36360 34604 36412 34610
rect 36360 34546 36412 34552
rect 36452 34536 36504 34542
rect 36452 34478 36504 34484
rect 36360 34468 36412 34474
rect 36360 34410 36412 34416
rect 36176 34060 36228 34066
rect 36176 34002 36228 34008
rect 36188 33590 36216 34002
rect 36372 33930 36400 34410
rect 36360 33924 36412 33930
rect 36360 33866 36412 33872
rect 36176 33584 36228 33590
rect 36176 33526 36228 33532
rect 36372 33386 36400 33866
rect 36360 33380 36412 33386
rect 36360 33322 36412 33328
rect 36372 33046 36400 33322
rect 36360 33040 36412 33046
rect 36360 32982 36412 32988
rect 36464 32434 36492 34478
rect 36636 33448 36688 33454
rect 36556 33396 36636 33402
rect 36556 33390 36688 33396
rect 36556 33374 36676 33390
rect 36268 32428 36320 32434
rect 36268 32370 36320 32376
rect 36452 32428 36504 32434
rect 36452 32370 36504 32376
rect 36082 31784 36138 31793
rect 35728 31726 35940 31754
rect 35716 31680 35768 31686
rect 35716 31622 35768 31628
rect 35728 30734 35756 31622
rect 35808 31476 35860 31482
rect 35808 31418 35860 31424
rect 35716 30728 35768 30734
rect 35716 30670 35768 30676
rect 35636 30144 35756 30172
rect 35820 30161 35848 31418
rect 35912 30274 35940 31726
rect 36082 31719 36138 31728
rect 35912 30246 36216 30274
rect 36280 30258 36308 32370
rect 36556 32178 36584 33374
rect 36372 32150 36584 32178
rect 36372 31521 36400 32150
rect 36636 32020 36688 32026
rect 36636 31962 36688 31968
rect 36728 32020 36780 32026
rect 36728 31962 36780 31968
rect 36648 31754 36676 31962
rect 36464 31726 36676 31754
rect 36358 31512 36414 31521
rect 36358 31447 36414 31456
rect 36372 30258 36400 31447
rect 35900 30184 35952 30190
rect 35532 29640 35584 29646
rect 35532 29582 35584 29588
rect 35544 28994 35572 29582
rect 35544 28966 35664 28994
rect 35532 28552 35584 28558
rect 35532 28494 35584 28500
rect 35544 28014 35572 28494
rect 35636 28422 35664 28966
rect 35624 28416 35676 28422
rect 35624 28358 35676 28364
rect 35728 28150 35756 30144
rect 35806 30152 35862 30161
rect 35952 30144 36124 30172
rect 35900 30126 35952 30132
rect 35806 30087 35862 30096
rect 35808 30048 35860 30054
rect 35808 29990 35860 29996
rect 35992 30048 36044 30054
rect 35992 29990 36044 29996
rect 35820 29850 35848 29990
rect 35808 29844 35860 29850
rect 35808 29786 35860 29792
rect 35820 29594 35848 29786
rect 36004 29714 36032 29990
rect 35992 29708 36044 29714
rect 35992 29650 36044 29656
rect 35820 29566 35940 29594
rect 35808 29504 35860 29510
rect 35808 29446 35860 29452
rect 35820 28558 35848 29446
rect 35912 29238 35940 29566
rect 35900 29232 35952 29238
rect 35900 29174 35952 29180
rect 36004 29170 36032 29650
rect 35992 29164 36044 29170
rect 35992 29106 36044 29112
rect 35900 29096 35952 29102
rect 35900 29038 35952 29044
rect 35808 28552 35860 28558
rect 35808 28494 35860 28500
rect 35716 28144 35768 28150
rect 35716 28086 35768 28092
rect 35532 28008 35584 28014
rect 35532 27950 35584 27956
rect 35452 27586 35664 27614
rect 35532 27328 35584 27334
rect 35532 27270 35584 27276
rect 35544 26353 35572 27270
rect 35530 26344 35586 26353
rect 35530 26279 35586 26288
rect 35532 26036 35584 26042
rect 35532 25978 35584 25984
rect 34796 25832 34848 25838
rect 34796 25774 34848 25780
rect 35348 25832 35400 25838
rect 35544 25786 35572 25978
rect 35348 25774 35400 25780
rect 34796 25696 34848 25702
rect 34796 25638 34848 25644
rect 34808 25498 34836 25638
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34796 25492 34848 25498
rect 34796 25434 34848 25440
rect 35360 24954 35388 25774
rect 35452 25758 35572 25786
rect 35348 24948 35400 24954
rect 35348 24890 35400 24896
rect 35348 24812 35400 24818
rect 35348 24754 35400 24760
rect 34702 24712 34758 24721
rect 34702 24647 34758 24656
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34794 24440 34850 24449
rect 34934 24443 35242 24452
rect 35360 24410 35388 24754
rect 34794 24375 34850 24384
rect 35348 24404 35400 24410
rect 34704 21616 34756 21622
rect 34704 21558 34756 21564
rect 34716 20874 34744 21558
rect 34704 20868 34756 20874
rect 34704 20810 34756 20816
rect 34624 20590 34744 20618
rect 34610 20496 34666 20505
rect 34610 20431 34666 20440
rect 34624 20058 34652 20431
rect 34612 20052 34664 20058
rect 34612 19994 34664 20000
rect 34520 19848 34572 19854
rect 34520 19790 34572 19796
rect 34428 18828 34480 18834
rect 34428 18770 34480 18776
rect 34532 18290 34560 19790
rect 34612 19440 34664 19446
rect 34612 19382 34664 19388
rect 34520 18284 34572 18290
rect 34520 18226 34572 18232
rect 34334 18048 34390 18057
rect 34334 17983 34390 17992
rect 34244 17808 34296 17814
rect 34244 17750 34296 17756
rect 34256 17626 34284 17750
rect 34164 17598 34284 17626
rect 34336 17672 34388 17678
rect 34336 17614 34388 17620
rect 34060 17196 34112 17202
rect 34060 17138 34112 17144
rect 33968 16992 34020 16998
rect 33968 16934 34020 16940
rect 33876 15020 33928 15026
rect 33876 14962 33928 14968
rect 33692 14612 33744 14618
rect 33744 14572 33824 14600
rect 33692 14554 33744 14560
rect 33692 14340 33744 14346
rect 33692 14282 33744 14288
rect 33600 14272 33652 14278
rect 33600 14214 33652 14220
rect 33508 12436 33560 12442
rect 33508 12378 33560 12384
rect 33704 12306 33732 14282
rect 33796 14006 33824 14572
rect 33784 14000 33836 14006
rect 33784 13942 33836 13948
rect 33782 13832 33838 13841
rect 33782 13767 33838 13776
rect 33796 13190 33824 13767
rect 33888 13394 33916 14962
rect 33980 14278 34008 16934
rect 34072 16697 34100 17138
rect 34058 16688 34114 16697
rect 34164 16658 34192 17598
rect 34348 17524 34376 17614
rect 34256 17496 34376 17524
rect 34058 16623 34114 16632
rect 34152 16652 34204 16658
rect 34152 16594 34204 16600
rect 34256 16538 34284 17496
rect 34532 16794 34560 18226
rect 34336 16788 34388 16794
rect 34336 16730 34388 16736
rect 34520 16788 34572 16794
rect 34520 16730 34572 16736
rect 34072 16510 34284 16538
rect 34072 16454 34100 16510
rect 34060 16448 34112 16454
rect 34060 16390 34112 16396
rect 34348 16096 34376 16730
rect 34426 16552 34482 16561
rect 34426 16487 34428 16496
rect 34480 16487 34482 16496
rect 34520 16516 34572 16522
rect 34428 16458 34480 16464
rect 34520 16458 34572 16464
rect 34532 16425 34560 16458
rect 34518 16416 34574 16425
rect 34518 16351 34574 16360
rect 34624 16250 34652 19382
rect 34716 18873 34744 20590
rect 34808 18952 34836 24375
rect 35348 24346 35400 24352
rect 35164 24132 35216 24138
rect 35164 24074 35216 24080
rect 35176 23730 35204 24074
rect 35164 23724 35216 23730
rect 35216 23684 35388 23712
rect 35164 23666 35216 23672
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34888 22772 34940 22778
rect 34888 22714 34940 22720
rect 34900 22545 34928 22714
rect 35360 22642 35388 23684
rect 35348 22636 35400 22642
rect 35348 22578 35400 22584
rect 34886 22536 34942 22545
rect 34886 22471 34942 22480
rect 35360 22438 35388 22578
rect 35348 22432 35400 22438
rect 35348 22374 35400 22380
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35452 22094 35480 25758
rect 35636 25684 35664 27586
rect 35820 26994 35848 28494
rect 35912 28082 35940 29038
rect 35900 28076 35952 28082
rect 35900 28018 35952 28024
rect 35898 27976 35954 27985
rect 36004 27946 36032 29106
rect 35898 27911 35954 27920
rect 35992 27940 36044 27946
rect 35808 26988 35860 26994
rect 35808 26930 35860 26936
rect 35820 25906 35848 26930
rect 35808 25900 35860 25906
rect 35808 25842 35860 25848
rect 35808 25764 35860 25770
rect 35808 25706 35860 25712
rect 35544 25656 35664 25684
rect 35544 24410 35572 25656
rect 35820 25362 35848 25706
rect 35808 25356 35860 25362
rect 35808 25298 35860 25304
rect 35624 24812 35676 24818
rect 35624 24754 35676 24760
rect 35532 24404 35584 24410
rect 35532 24346 35584 24352
rect 35532 23656 35584 23662
rect 35532 23598 35584 23604
rect 35544 22681 35572 23598
rect 35530 22672 35586 22681
rect 35530 22607 35586 22616
rect 35532 22568 35584 22574
rect 35532 22510 35584 22516
rect 35544 22234 35572 22510
rect 35532 22228 35584 22234
rect 35532 22170 35584 22176
rect 35360 22066 35480 22094
rect 35360 21622 35388 22066
rect 35348 21616 35400 21622
rect 35348 21558 35400 21564
rect 35636 21486 35664 24754
rect 35808 23044 35860 23050
rect 35808 22986 35860 22992
rect 35820 22642 35848 22986
rect 35808 22636 35860 22642
rect 35808 22578 35860 22584
rect 35808 22228 35860 22234
rect 35808 22170 35860 22176
rect 35348 21480 35400 21486
rect 35348 21422 35400 21428
rect 35624 21480 35676 21486
rect 35624 21422 35676 21428
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34808 18924 35020 18952
rect 34702 18864 34758 18873
rect 34702 18799 34758 18808
rect 34888 18828 34940 18834
rect 34888 18770 34940 18776
rect 34704 18760 34756 18766
rect 34704 18702 34756 18708
rect 34612 16244 34664 16250
rect 34612 16186 34664 16192
rect 34520 16176 34572 16182
rect 34520 16118 34572 16124
rect 34428 16108 34480 16114
rect 34348 16068 34428 16096
rect 34428 16050 34480 16056
rect 34440 15484 34468 16050
rect 34532 15638 34560 16118
rect 34520 15632 34572 15638
rect 34520 15574 34572 15580
rect 34440 15456 34560 15484
rect 34060 15428 34112 15434
rect 34060 15370 34112 15376
rect 33968 14272 34020 14278
rect 33968 14214 34020 14220
rect 33876 13388 33928 13394
rect 33876 13330 33928 13336
rect 34072 13326 34100 15370
rect 34244 15360 34296 15366
rect 34244 15302 34296 15308
rect 34256 15026 34284 15302
rect 34244 15020 34296 15026
rect 34244 14962 34296 14968
rect 34256 14414 34284 14962
rect 34428 14952 34480 14958
rect 34428 14894 34480 14900
rect 34440 14822 34468 14894
rect 34428 14816 34480 14822
rect 34428 14758 34480 14764
rect 34336 14476 34388 14482
rect 34440 14464 34468 14758
rect 34388 14436 34468 14464
rect 34336 14418 34388 14424
rect 34244 14408 34296 14414
rect 34244 14350 34296 14356
rect 34152 13796 34204 13802
rect 34152 13738 34204 13744
rect 33968 13320 34020 13326
rect 33968 13262 34020 13268
rect 34060 13320 34112 13326
rect 34060 13262 34112 13268
rect 33784 13184 33836 13190
rect 33784 13126 33836 13132
rect 33784 12844 33836 12850
rect 33784 12786 33836 12792
rect 33692 12300 33744 12306
rect 33692 12242 33744 12248
rect 33600 12164 33652 12170
rect 33600 12106 33652 12112
rect 33508 11280 33560 11286
rect 33612 11268 33640 12106
rect 33796 11694 33824 12786
rect 33876 12640 33928 12646
rect 33876 12582 33928 12588
rect 33888 11762 33916 12582
rect 33876 11756 33928 11762
rect 33876 11698 33928 11704
rect 33784 11688 33836 11694
rect 33784 11630 33836 11636
rect 33560 11240 33640 11268
rect 33508 11222 33560 11228
rect 33876 11212 33928 11218
rect 33876 11154 33928 11160
rect 33600 11144 33652 11150
rect 33598 11112 33600 11121
rect 33652 11112 33654 11121
rect 33598 11047 33654 11056
rect 33888 10962 33916 11154
rect 33704 10934 33916 10962
rect 33508 10668 33560 10674
rect 33704 10656 33732 10934
rect 33560 10628 33732 10656
rect 33784 10668 33836 10674
rect 33508 10610 33560 10616
rect 33784 10610 33836 10616
rect 33520 10062 33548 10610
rect 33508 10056 33560 10062
rect 33508 9998 33560 10004
rect 33520 9654 33548 9998
rect 33692 9920 33744 9926
rect 33692 9862 33744 9868
rect 33600 9716 33652 9722
rect 33600 9658 33652 9664
rect 33508 9648 33560 9654
rect 33508 9590 33560 9596
rect 33416 9580 33468 9586
rect 33416 9522 33468 9528
rect 32772 9512 32824 9518
rect 32772 9454 32824 9460
rect 32784 9217 32812 9454
rect 32770 9208 32826 9217
rect 32680 9172 32732 9178
rect 33428 9178 33456 9522
rect 33508 9444 33560 9450
rect 33612 9432 33640 9658
rect 33560 9404 33640 9432
rect 33508 9386 33560 9392
rect 33520 9178 33548 9386
rect 32770 9143 32826 9152
rect 33416 9172 33468 9178
rect 32680 9114 32732 9120
rect 33416 9114 33468 9120
rect 33508 9172 33560 9178
rect 33508 9114 33560 9120
rect 33048 8968 33100 8974
rect 33048 8910 33100 8916
rect 33060 8430 33088 8910
rect 33520 8634 33548 9114
rect 33704 8974 33732 9862
rect 33692 8968 33744 8974
rect 33692 8910 33744 8916
rect 33796 8906 33824 10610
rect 33980 9654 34008 13262
rect 34058 12880 34114 12889
rect 34164 12850 34192 13738
rect 34058 12815 34060 12824
rect 34112 12815 34114 12824
rect 34152 12844 34204 12850
rect 34060 12786 34112 12792
rect 34152 12786 34204 12792
rect 34072 12238 34100 12786
rect 34152 12708 34204 12714
rect 34256 12696 34284 14350
rect 34348 13682 34376 14418
rect 34428 14340 34480 14346
rect 34428 14282 34480 14288
rect 34440 13802 34468 14282
rect 34532 13841 34560 15456
rect 34624 15366 34652 16186
rect 34612 15360 34664 15366
rect 34612 15302 34664 15308
rect 34612 14476 34664 14482
rect 34716 14464 34744 18702
rect 34900 18290 34928 18770
rect 34888 18284 34940 18290
rect 34888 18226 34940 18232
rect 34900 18170 34928 18226
rect 34992 18193 35020 18924
rect 35070 18864 35126 18873
rect 35070 18799 35126 18808
rect 35084 18306 35112 18799
rect 35164 18692 35216 18698
rect 35164 18634 35216 18640
rect 35176 18426 35204 18634
rect 35164 18420 35216 18426
rect 35164 18362 35216 18368
rect 35084 18290 35296 18306
rect 35084 18284 35308 18290
rect 35084 18278 35256 18284
rect 35256 18226 35308 18232
rect 34808 18142 34928 18170
rect 34978 18184 35034 18193
rect 34808 16794 34836 18142
rect 34978 18119 35034 18128
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35360 17610 35388 21422
rect 35440 21344 35492 21350
rect 35440 21286 35492 21292
rect 35532 21344 35584 21350
rect 35532 21286 35584 21292
rect 35452 20942 35480 21286
rect 35544 20942 35572 21286
rect 35440 20936 35492 20942
rect 35440 20878 35492 20884
rect 35532 20936 35584 20942
rect 35532 20878 35584 20884
rect 35452 19854 35480 20878
rect 35440 19848 35492 19854
rect 35440 19790 35492 19796
rect 35452 18970 35480 19790
rect 35440 18964 35492 18970
rect 35440 18906 35492 18912
rect 35452 17678 35480 18906
rect 35440 17672 35492 17678
rect 35440 17614 35492 17620
rect 35348 17604 35400 17610
rect 35348 17546 35400 17552
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35452 16794 35480 17614
rect 34796 16788 34848 16794
rect 34796 16730 34848 16736
rect 35440 16788 35492 16794
rect 35440 16730 35492 16736
rect 34978 16552 35034 16561
rect 34978 16487 35034 16496
rect 35164 16516 35216 16522
rect 34992 16250 35020 16487
rect 35164 16458 35216 16464
rect 35256 16516 35308 16522
rect 35256 16458 35308 16464
rect 35348 16516 35400 16522
rect 35544 16504 35572 20878
rect 35716 20868 35768 20874
rect 35820 20856 35848 22170
rect 35912 20942 35940 27911
rect 35992 27882 36044 27888
rect 36004 26382 36032 27882
rect 36096 27674 36124 30144
rect 36188 30122 36216 30246
rect 36268 30252 36320 30258
rect 36268 30194 36320 30200
rect 36360 30252 36412 30258
rect 36360 30194 36412 30200
rect 36176 30116 36228 30122
rect 36176 30058 36228 30064
rect 36188 29073 36216 30058
rect 36280 29578 36308 30194
rect 36268 29572 36320 29578
rect 36268 29514 36320 29520
rect 36266 29472 36322 29481
rect 36266 29407 36322 29416
rect 36174 29064 36230 29073
rect 36174 28999 36230 29008
rect 36280 28762 36308 29407
rect 36268 28756 36320 28762
rect 36268 28698 36320 28704
rect 36372 27878 36400 30194
rect 36464 28014 36492 31726
rect 36740 30802 36768 31962
rect 36832 31890 36860 34886
rect 36820 31884 36872 31890
rect 36820 31826 36872 31832
rect 36728 30796 36780 30802
rect 36728 30738 36780 30744
rect 36636 30048 36688 30054
rect 36636 29990 36688 29996
rect 36648 29850 36676 29990
rect 36636 29844 36688 29850
rect 36636 29786 36688 29792
rect 36636 29504 36688 29510
rect 36636 29446 36688 29452
rect 36452 28008 36504 28014
rect 36452 27950 36504 27956
rect 36544 28008 36596 28014
rect 36544 27950 36596 27956
rect 36360 27872 36412 27878
rect 36360 27814 36412 27820
rect 36084 27668 36136 27674
rect 36084 27610 36136 27616
rect 36096 27316 36124 27610
rect 36372 27470 36400 27814
rect 36360 27464 36412 27470
rect 36360 27406 36412 27412
rect 36096 27288 36400 27316
rect 36084 27056 36136 27062
rect 36084 26998 36136 27004
rect 36096 26382 36124 26998
rect 35992 26376 36044 26382
rect 35992 26318 36044 26324
rect 36084 26376 36136 26382
rect 36084 26318 36136 26324
rect 36084 25832 36136 25838
rect 36082 25800 36084 25809
rect 36136 25800 36138 25809
rect 36082 25735 36138 25744
rect 36084 25696 36136 25702
rect 36084 25638 36136 25644
rect 36096 25294 36124 25638
rect 36084 25288 36136 25294
rect 36084 25230 36136 25236
rect 36176 25152 36228 25158
rect 36176 25094 36228 25100
rect 36188 24614 36216 25094
rect 36176 24608 36228 24614
rect 36176 24550 36228 24556
rect 35992 24064 36044 24070
rect 35992 24006 36044 24012
rect 35900 20936 35952 20942
rect 35900 20878 35952 20884
rect 35768 20828 35848 20856
rect 35716 20810 35768 20816
rect 35624 20596 35676 20602
rect 35624 20538 35676 20544
rect 35636 19446 35664 20538
rect 35624 19440 35676 19446
rect 35624 19382 35676 19388
rect 35728 19378 35756 20810
rect 35900 19848 35952 19854
rect 35898 19816 35900 19825
rect 35952 19816 35954 19825
rect 35898 19751 35954 19760
rect 35716 19372 35768 19378
rect 35716 19314 35768 19320
rect 35716 18760 35768 18766
rect 35636 18737 35716 18748
rect 35622 18728 35716 18737
rect 35678 18720 35716 18728
rect 35716 18702 35768 18708
rect 35808 18760 35860 18766
rect 35808 18702 35860 18708
rect 35622 18663 35678 18672
rect 35820 18601 35848 18702
rect 35806 18592 35862 18601
rect 35806 18527 35862 18536
rect 35820 17626 35848 18527
rect 35912 18465 35940 19751
rect 35898 18456 35954 18465
rect 35898 18391 35954 18400
rect 35900 18284 35952 18290
rect 35900 18226 35952 18232
rect 35636 17598 35848 17626
rect 35636 17202 35664 17598
rect 35716 17536 35768 17542
rect 35716 17478 35768 17484
rect 35808 17536 35860 17542
rect 35808 17478 35860 17484
rect 35728 17377 35756 17478
rect 35714 17368 35770 17377
rect 35714 17303 35770 17312
rect 35624 17196 35676 17202
rect 35624 17138 35676 17144
rect 35624 16788 35676 16794
rect 35624 16730 35676 16736
rect 35348 16458 35400 16464
rect 35452 16476 35572 16504
rect 34980 16244 35032 16250
rect 34980 16186 35032 16192
rect 35176 16114 35204 16458
rect 35268 16182 35296 16458
rect 35256 16176 35308 16182
rect 35256 16118 35308 16124
rect 35164 16108 35216 16114
rect 35164 16050 35216 16056
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35360 15722 35388 16458
rect 35452 16289 35480 16476
rect 35438 16280 35494 16289
rect 35438 16215 35440 16224
rect 35492 16215 35494 16224
rect 35440 16186 35492 16192
rect 35636 16182 35664 16730
rect 35624 16176 35676 16182
rect 35438 16144 35494 16153
rect 35624 16118 35676 16124
rect 35438 16079 35440 16088
rect 35492 16079 35494 16088
rect 35440 16050 35492 16056
rect 35624 16040 35676 16046
rect 35268 15694 35388 15722
rect 35544 16000 35624 16028
rect 34794 15328 34850 15337
rect 34794 15263 34850 15272
rect 34664 14436 34744 14464
rect 34808 14464 34836 15263
rect 35268 15026 35296 15694
rect 35348 15428 35400 15434
rect 35348 15370 35400 15376
rect 35256 15020 35308 15026
rect 35256 14962 35308 14968
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34808 14436 35204 14464
rect 34612 14418 34664 14424
rect 34518 13832 34574 13841
rect 34428 13796 34480 13802
rect 34518 13767 34574 13776
rect 34428 13738 34480 13744
rect 34520 13728 34572 13734
rect 34348 13654 34468 13682
rect 34520 13670 34572 13676
rect 34204 12668 34284 12696
rect 34152 12650 34204 12656
rect 34060 12232 34112 12238
rect 34060 12174 34112 12180
rect 34152 11688 34204 11694
rect 34152 11630 34204 11636
rect 34060 11552 34112 11558
rect 34060 11494 34112 11500
rect 34072 11150 34100 11494
rect 34060 11144 34112 11150
rect 34060 11086 34112 11092
rect 34060 10600 34112 10606
rect 34060 10542 34112 10548
rect 33968 9648 34020 9654
rect 33968 9590 34020 9596
rect 33876 9580 33928 9586
rect 33876 9522 33928 9528
rect 33784 8900 33836 8906
rect 33784 8842 33836 8848
rect 33692 8832 33744 8838
rect 33692 8774 33744 8780
rect 33704 8634 33732 8774
rect 33508 8628 33560 8634
rect 33508 8570 33560 8576
rect 33692 8628 33744 8634
rect 33692 8570 33744 8576
rect 33048 8424 33100 8430
rect 33888 8378 33916 9522
rect 33966 9480 34022 9489
rect 33966 9415 33968 9424
rect 34020 9415 34022 9424
rect 33968 9386 34020 9392
rect 34072 9194 34100 10542
rect 33980 9166 34100 9194
rect 33980 8430 34008 9166
rect 34060 9104 34112 9110
rect 34060 9046 34112 9052
rect 33048 8366 33100 8372
rect 33232 8356 33284 8362
rect 33232 8298 33284 8304
rect 33796 8350 33916 8378
rect 33968 8424 34020 8430
rect 33968 8366 34020 8372
rect 32772 8288 32824 8294
rect 32600 8248 32772 8276
rect 32772 8230 32824 8236
rect 32496 7472 32548 7478
rect 32496 7414 32548 7420
rect 32784 7410 32812 8230
rect 33244 7410 33272 8298
rect 33796 7818 33824 8350
rect 33876 8288 33928 8294
rect 33876 8230 33928 8236
rect 33784 7812 33836 7818
rect 33784 7754 33836 7760
rect 33692 7472 33744 7478
rect 33690 7440 33692 7449
rect 33744 7440 33746 7449
rect 32772 7404 32824 7410
rect 32772 7346 32824 7352
rect 33140 7404 33192 7410
rect 33140 7346 33192 7352
rect 33232 7404 33284 7410
rect 33416 7404 33468 7410
rect 33232 7346 33284 7352
rect 33336 7364 33416 7392
rect 33152 7290 33180 7346
rect 33336 7290 33364 7364
rect 33690 7375 33746 7384
rect 33416 7346 33468 7352
rect 32416 7262 32536 7290
rect 33152 7262 33364 7290
rect 32312 7200 32364 7206
rect 32312 7142 32364 7148
rect 32404 7200 32456 7206
rect 32404 7142 32456 7148
rect 32324 7002 32352 7142
rect 32220 6996 32272 7002
rect 32220 6938 32272 6944
rect 32312 6996 32364 7002
rect 32312 6938 32364 6944
rect 31484 6860 31536 6866
rect 31484 6802 31536 6808
rect 32128 6860 32180 6866
rect 32128 6802 32180 6808
rect 31300 6792 31352 6798
rect 31300 6734 31352 6740
rect 31312 6322 31340 6734
rect 31576 6656 31628 6662
rect 31576 6598 31628 6604
rect 31300 6316 31352 6322
rect 31300 6258 31352 6264
rect 31588 5370 31616 6598
rect 32232 6322 32260 6938
rect 32416 6798 32444 7142
rect 32508 6934 32536 7262
rect 32496 6928 32548 6934
rect 33336 6905 33364 7262
rect 33796 7206 33824 7754
rect 33888 7410 33916 8230
rect 34072 8090 34100 9046
rect 34060 8084 34112 8090
rect 34060 8026 34112 8032
rect 33876 7404 33928 7410
rect 33876 7346 33928 7352
rect 33784 7200 33836 7206
rect 33784 7142 33836 7148
rect 33508 6928 33560 6934
rect 32496 6870 32548 6876
rect 33322 6896 33378 6905
rect 33508 6870 33560 6876
rect 33322 6831 33378 6840
rect 32404 6792 32456 6798
rect 32404 6734 32456 6740
rect 32496 6792 32548 6798
rect 33324 6792 33376 6798
rect 32496 6734 32548 6740
rect 33322 6760 33324 6769
rect 33376 6760 33378 6769
rect 32508 6662 32536 6734
rect 33048 6724 33100 6730
rect 33232 6724 33284 6730
rect 33100 6684 33232 6712
rect 33048 6666 33100 6672
rect 33322 6695 33378 6704
rect 33232 6666 33284 6672
rect 32496 6656 32548 6662
rect 32496 6598 32548 6604
rect 32680 6656 32732 6662
rect 32680 6598 32732 6604
rect 32220 6316 32272 6322
rect 32220 6258 32272 6264
rect 32588 5704 32640 5710
rect 32586 5672 32588 5681
rect 32640 5672 32642 5681
rect 32586 5607 32642 5616
rect 31666 5400 31722 5409
rect 31576 5364 31628 5370
rect 31666 5335 31668 5344
rect 31576 5306 31628 5312
rect 31720 5335 31722 5344
rect 31668 5306 31720 5312
rect 32600 5234 32628 5607
rect 32692 5370 32720 6598
rect 32772 5636 32824 5642
rect 32772 5578 32824 5584
rect 32784 5370 32812 5578
rect 33232 5568 33284 5574
rect 33232 5510 33284 5516
rect 32680 5364 32732 5370
rect 32680 5306 32732 5312
rect 32772 5364 32824 5370
rect 32772 5306 32824 5312
rect 33244 5234 33272 5510
rect 33520 5302 33548 6870
rect 33888 6730 33916 7346
rect 34164 7002 34192 11630
rect 34256 9654 34284 12668
rect 34336 12232 34388 12238
rect 34336 12174 34388 12180
rect 34244 9648 34296 9654
rect 34244 9590 34296 9596
rect 34244 9444 34296 9450
rect 34244 9386 34296 9392
rect 34256 9042 34284 9386
rect 34348 9110 34376 12174
rect 34440 11914 34468 13654
rect 34532 13297 34560 13670
rect 34624 13530 34652 14418
rect 35176 14346 35204 14436
rect 35072 14340 35124 14346
rect 35072 14282 35124 14288
rect 35164 14340 35216 14346
rect 35164 14282 35216 14288
rect 34704 14272 34756 14278
rect 34704 14214 34756 14220
rect 34716 14074 34744 14214
rect 34794 14104 34850 14113
rect 34704 14068 34756 14074
rect 34794 14039 34850 14048
rect 34704 14010 34756 14016
rect 34612 13524 34664 13530
rect 34612 13466 34664 13472
rect 34518 13288 34574 13297
rect 34518 13223 34574 13232
rect 34532 13190 34560 13223
rect 34520 13184 34572 13190
rect 34520 13126 34572 13132
rect 34520 12776 34572 12782
rect 34520 12718 34572 12724
rect 34532 12102 34560 12718
rect 34520 12096 34572 12102
rect 34520 12038 34572 12044
rect 34440 11886 34560 11914
rect 34426 11792 34482 11801
rect 34426 11727 34482 11736
rect 34440 11694 34468 11727
rect 34428 11688 34480 11694
rect 34428 11630 34480 11636
rect 34440 10810 34468 11630
rect 34532 11558 34560 11886
rect 34808 11812 34836 14039
rect 35084 13841 35112 14282
rect 35176 13938 35204 14282
rect 35164 13932 35216 13938
rect 35164 13874 35216 13880
rect 35070 13832 35126 13841
rect 35070 13767 35126 13776
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35256 13388 35308 13394
rect 35256 13330 35308 13336
rect 34888 13252 34940 13258
rect 34888 13194 34940 13200
rect 34900 12986 34928 13194
rect 34888 12980 34940 12986
rect 34888 12922 34940 12928
rect 35268 12714 35296 13330
rect 35256 12708 35308 12714
rect 35256 12650 35308 12656
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35256 12300 35308 12306
rect 35256 12242 35308 12248
rect 35268 11830 35296 12242
rect 34888 11824 34940 11830
rect 34808 11784 34888 11812
rect 35072 11824 35124 11830
rect 34888 11766 34940 11772
rect 35070 11792 35072 11801
rect 35256 11824 35308 11830
rect 35124 11792 35126 11801
rect 35256 11766 35308 11772
rect 35070 11727 35126 11736
rect 34520 11552 34572 11558
rect 34520 11494 34572 11500
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35164 11144 35216 11150
rect 35164 11086 35216 11092
rect 35360 11098 35388 15370
rect 35438 14784 35494 14793
rect 35438 14719 35494 14728
rect 35452 14414 35480 14719
rect 35440 14408 35492 14414
rect 35440 14350 35492 14356
rect 35544 14346 35572 16000
rect 35624 15982 35676 15988
rect 35624 15496 35676 15502
rect 35676 15456 35756 15484
rect 35624 15438 35676 15444
rect 35624 15360 35676 15366
rect 35624 15302 35676 15308
rect 35636 14346 35664 15302
rect 35728 14958 35756 15456
rect 35716 14952 35768 14958
rect 35716 14894 35768 14900
rect 35532 14340 35584 14346
rect 35532 14282 35584 14288
rect 35624 14340 35676 14346
rect 35624 14282 35676 14288
rect 35440 13320 35492 13326
rect 35440 13262 35492 13268
rect 35452 11218 35480 13262
rect 35440 11212 35492 11218
rect 35440 11154 35492 11160
rect 34428 10804 34480 10810
rect 34428 10746 34480 10752
rect 35176 10520 35204 11086
rect 35360 11070 35480 11098
rect 35452 10606 35480 11070
rect 35440 10600 35492 10606
rect 35440 10542 35492 10548
rect 35176 10492 35388 10520
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35360 9674 35388 10492
rect 34520 9648 34572 9654
rect 35268 9646 35388 9674
rect 34520 9590 34572 9596
rect 34610 9616 34666 9625
rect 34428 9580 34480 9586
rect 34428 9522 34480 9528
rect 34440 9178 34468 9522
rect 34428 9172 34480 9178
rect 34428 9114 34480 9120
rect 34336 9104 34388 9110
rect 34532 9058 34560 9590
rect 34610 9551 34666 9560
rect 34624 9450 34652 9551
rect 35268 9518 35296 9646
rect 35256 9512 35308 9518
rect 35254 9480 35256 9489
rect 35348 9512 35400 9518
rect 35308 9480 35310 9489
rect 34612 9444 34664 9450
rect 35348 9454 35400 9460
rect 35254 9415 35310 9424
rect 34612 9386 34664 9392
rect 34336 9046 34388 9052
rect 34244 9036 34296 9042
rect 34244 8978 34296 8984
rect 34440 9030 34560 9058
rect 34256 8498 34284 8978
rect 34440 8838 34468 9030
rect 34624 8974 34652 9386
rect 34796 9376 34848 9382
rect 34716 9336 34796 9364
rect 34612 8968 34664 8974
rect 34612 8910 34664 8916
rect 34336 8832 34388 8838
rect 34336 8774 34388 8780
rect 34428 8832 34480 8838
rect 34428 8774 34480 8780
rect 34244 8492 34296 8498
rect 34244 8434 34296 8440
rect 34348 8294 34376 8774
rect 34440 8566 34468 8774
rect 34428 8560 34480 8566
rect 34428 8502 34480 8508
rect 34520 8560 34572 8566
rect 34520 8502 34572 8508
rect 34532 8412 34560 8502
rect 34440 8384 34560 8412
rect 34336 8288 34388 8294
rect 34336 8230 34388 8236
rect 34440 8106 34468 8384
rect 34256 8078 34468 8106
rect 34152 6996 34204 7002
rect 34152 6938 34204 6944
rect 33968 6792 34020 6798
rect 33968 6734 34020 6740
rect 34152 6792 34204 6798
rect 34256 6780 34284 8078
rect 34336 7540 34388 7546
rect 34336 7482 34388 7488
rect 34348 7002 34376 7482
rect 34336 6996 34388 7002
rect 34336 6938 34388 6944
rect 34624 6866 34652 8910
rect 34716 7750 34744 9336
rect 34796 9318 34848 9324
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 35360 8498 35388 9454
rect 35348 8492 35400 8498
rect 35348 8434 35400 8440
rect 34796 8424 34848 8430
rect 34796 8366 34848 8372
rect 34808 8072 34836 8366
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34808 8044 35020 8072
rect 34992 7886 35020 8044
rect 34888 7880 34940 7886
rect 34888 7822 34940 7828
rect 34980 7880 35032 7886
rect 34980 7822 35032 7828
rect 34704 7744 34756 7750
rect 34704 7686 34756 7692
rect 34716 7002 34744 7686
rect 34900 7410 34928 7822
rect 35072 7812 35124 7818
rect 35072 7754 35124 7760
rect 34980 7744 35032 7750
rect 34980 7686 35032 7692
rect 34992 7478 35020 7686
rect 35084 7546 35112 7754
rect 35348 7744 35400 7750
rect 35268 7704 35348 7732
rect 35072 7540 35124 7546
rect 35072 7482 35124 7488
rect 34980 7472 35032 7478
rect 34980 7414 35032 7420
rect 35162 7440 35218 7449
rect 34888 7404 34940 7410
rect 34888 7346 34940 7352
rect 34900 7274 34928 7346
rect 34992 7274 35020 7414
rect 35268 7410 35296 7704
rect 35348 7686 35400 7692
rect 35348 7472 35400 7478
rect 35348 7414 35400 7420
rect 35162 7375 35164 7384
rect 35216 7375 35218 7384
rect 35256 7404 35308 7410
rect 35164 7346 35216 7352
rect 35256 7346 35308 7352
rect 34888 7268 34940 7274
rect 34888 7210 34940 7216
rect 34980 7268 35032 7274
rect 34980 7210 35032 7216
rect 34796 7200 34848 7206
rect 34796 7142 34848 7148
rect 34704 6996 34756 7002
rect 34704 6938 34756 6944
rect 34612 6860 34664 6866
rect 34612 6802 34664 6808
rect 34204 6752 34284 6780
rect 34428 6792 34480 6798
rect 34152 6734 34204 6740
rect 34808 6780 34836 7142
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35360 6798 35388 7414
rect 34980 6792 35032 6798
rect 34808 6752 34980 6780
rect 34428 6734 34480 6740
rect 34980 6734 35032 6740
rect 35348 6792 35400 6798
rect 35452 6769 35480 10542
rect 35544 7290 35572 14282
rect 35728 13870 35756 14894
rect 35716 13864 35768 13870
rect 35716 13806 35768 13812
rect 35624 13728 35676 13734
rect 35624 13670 35676 13676
rect 35636 12986 35664 13670
rect 35728 13308 35756 13806
rect 35820 13530 35848 17478
rect 35912 17270 35940 18226
rect 35900 17264 35952 17270
rect 35900 17206 35952 17212
rect 35900 17060 35952 17066
rect 35900 17002 35952 17008
rect 35912 15434 35940 17002
rect 35900 15428 35952 15434
rect 35900 15370 35952 15376
rect 36004 14618 36032 24006
rect 36188 23186 36216 24550
rect 36176 23180 36228 23186
rect 36176 23122 36228 23128
rect 36268 23112 36320 23118
rect 36268 23054 36320 23060
rect 36174 22944 36230 22953
rect 36280 22930 36308 23054
rect 36230 22902 36308 22930
rect 36174 22879 36230 22888
rect 36372 22642 36400 27288
rect 36464 26994 36492 27950
rect 36452 26988 36504 26994
rect 36452 26930 36504 26936
rect 36556 26790 36584 27950
rect 36648 27470 36676 29446
rect 36726 28792 36782 28801
rect 36726 28727 36728 28736
rect 36780 28727 36782 28736
rect 36728 28698 36780 28704
rect 36832 28642 36860 31826
rect 36924 31482 36952 41386
rect 41892 41274 41920 43893
rect 41880 41268 41932 41274
rect 41880 41210 41932 41216
rect 40776 41132 40828 41138
rect 40776 41074 40828 41080
rect 40788 40186 40816 41074
rect 40960 40928 41012 40934
rect 40958 40896 40960 40905
rect 41012 40896 41014 40905
rect 40958 40831 41014 40840
rect 40776 40180 40828 40186
rect 40776 40122 40828 40128
rect 40776 37256 40828 37262
rect 40776 37198 40828 37204
rect 40040 36916 40092 36922
rect 40040 36858 40092 36864
rect 37740 34536 37792 34542
rect 37740 34478 37792 34484
rect 37464 34400 37516 34406
rect 37464 34342 37516 34348
rect 37476 34202 37504 34342
rect 37464 34196 37516 34202
rect 37464 34138 37516 34144
rect 37372 33924 37424 33930
rect 37372 33866 37424 33872
rect 37280 33516 37332 33522
rect 37280 33458 37332 33464
rect 37292 32978 37320 33458
rect 37384 33114 37412 33866
rect 37372 33108 37424 33114
rect 37372 33050 37424 33056
rect 37096 32972 37148 32978
rect 37096 32914 37148 32920
rect 37280 32972 37332 32978
rect 37280 32914 37332 32920
rect 37004 32768 37056 32774
rect 37004 32710 37056 32716
rect 37016 31890 37044 32710
rect 37108 32570 37136 32914
rect 37292 32774 37320 32914
rect 37280 32768 37332 32774
rect 37280 32710 37332 32716
rect 37556 32768 37608 32774
rect 37556 32710 37608 32716
rect 37648 32768 37700 32774
rect 37648 32710 37700 32716
rect 37096 32564 37148 32570
rect 37096 32506 37148 32512
rect 37108 32026 37136 32506
rect 37292 32366 37320 32710
rect 37464 32428 37516 32434
rect 37464 32370 37516 32376
rect 37280 32360 37332 32366
rect 37280 32302 37332 32308
rect 37096 32020 37148 32026
rect 37096 31962 37148 31968
rect 37004 31884 37056 31890
rect 37004 31826 37056 31832
rect 37292 31754 37320 32302
rect 37476 32026 37504 32370
rect 37568 32230 37596 32710
rect 37556 32224 37608 32230
rect 37556 32166 37608 32172
rect 37464 32020 37516 32026
rect 37464 31962 37516 31968
rect 37280 31748 37332 31754
rect 37280 31690 37332 31696
rect 36912 31476 36964 31482
rect 36912 31418 36964 31424
rect 37292 31142 37320 31690
rect 37280 31136 37332 31142
rect 37280 31078 37332 31084
rect 37292 30802 37320 31078
rect 37280 30796 37332 30802
rect 37280 30738 37332 30744
rect 36912 30592 36964 30598
rect 36912 30534 36964 30540
rect 36924 29646 36952 30534
rect 37370 30288 37426 30297
rect 37370 30223 37426 30232
rect 36912 29640 36964 29646
rect 36912 29582 36964 29588
rect 36740 28614 36860 28642
rect 36636 27464 36688 27470
rect 36636 27406 36688 27412
rect 36648 27062 36676 27406
rect 36636 27056 36688 27062
rect 36636 26998 36688 27004
rect 36544 26784 36596 26790
rect 36544 26726 36596 26732
rect 36544 26512 36596 26518
rect 36544 26454 36596 26460
rect 36556 24818 36584 26454
rect 36740 25498 36768 28614
rect 36820 28484 36872 28490
rect 36820 28426 36872 28432
rect 36728 25492 36780 25498
rect 36728 25434 36780 25440
rect 36544 24812 36596 24818
rect 36544 24754 36596 24760
rect 36452 24744 36504 24750
rect 36452 24686 36504 24692
rect 36464 23662 36492 24686
rect 36728 24132 36780 24138
rect 36728 24074 36780 24080
rect 36452 23656 36504 23662
rect 36452 23598 36504 23604
rect 36360 22636 36412 22642
rect 36360 22578 36412 22584
rect 36360 21888 36412 21894
rect 36360 21830 36412 21836
rect 36372 21690 36400 21830
rect 36360 21684 36412 21690
rect 36360 21626 36412 21632
rect 36084 21140 36136 21146
rect 36084 21082 36136 21088
rect 36268 21140 36320 21146
rect 36268 21082 36320 21088
rect 36096 20262 36124 21082
rect 36084 20256 36136 20262
rect 36084 20198 36136 20204
rect 36174 19544 36230 19553
rect 36174 19479 36230 19488
rect 36188 18358 36216 19479
rect 36176 18352 36228 18358
rect 36176 18294 36228 18300
rect 36174 17776 36230 17785
rect 36174 17711 36230 17720
rect 36084 17332 36136 17338
rect 36084 17274 36136 17280
rect 36096 16658 36124 17274
rect 36084 16652 36136 16658
rect 36084 16594 36136 16600
rect 36082 16552 36138 16561
rect 36082 16487 36138 16496
rect 36096 16114 36124 16487
rect 36084 16108 36136 16114
rect 36084 16050 36136 16056
rect 36084 15428 36136 15434
rect 36084 15370 36136 15376
rect 35992 14612 36044 14618
rect 35992 14554 36044 14560
rect 35992 14340 36044 14346
rect 35992 14282 36044 14288
rect 36004 13938 36032 14282
rect 36096 13938 36124 15370
rect 35992 13932 36044 13938
rect 35992 13874 36044 13880
rect 36084 13932 36136 13938
rect 36084 13874 36136 13880
rect 35808 13524 35860 13530
rect 35808 13466 35860 13472
rect 35808 13320 35860 13326
rect 35728 13280 35808 13308
rect 35808 13262 35860 13268
rect 35624 12980 35676 12986
rect 35624 12922 35676 12928
rect 35820 12238 35848 13262
rect 36004 13190 36032 13874
rect 35992 13184 36044 13190
rect 35992 13126 36044 13132
rect 35900 12980 35952 12986
rect 35900 12922 35952 12928
rect 35808 12232 35860 12238
rect 35808 12174 35860 12180
rect 35716 11756 35768 11762
rect 35716 11698 35768 11704
rect 35728 9654 35756 11698
rect 35912 10742 35940 12922
rect 35990 12064 36046 12073
rect 35990 11999 36046 12008
rect 36004 11830 36032 11999
rect 35992 11824 36044 11830
rect 35992 11766 36044 11772
rect 36096 11762 36124 13874
rect 36188 12986 36216 17711
rect 36280 16697 36308 21082
rect 36372 20942 36400 21626
rect 36360 20936 36412 20942
rect 36360 20878 36412 20884
rect 36464 20641 36492 23598
rect 36544 23520 36596 23526
rect 36544 23462 36596 23468
rect 36556 20777 36584 23462
rect 36636 23044 36688 23050
rect 36636 22986 36688 22992
rect 36648 22710 36676 22986
rect 36636 22704 36688 22710
rect 36636 22646 36688 22652
rect 36648 21622 36676 22646
rect 36636 21616 36688 21622
rect 36636 21558 36688 21564
rect 36648 20924 36676 21558
rect 36740 21146 36768 24074
rect 36728 21140 36780 21146
rect 36728 21082 36780 21088
rect 36728 20936 36780 20942
rect 36648 20896 36728 20924
rect 36728 20878 36780 20884
rect 36636 20800 36688 20806
rect 36542 20768 36598 20777
rect 36636 20742 36688 20748
rect 36542 20703 36598 20712
rect 36450 20632 36506 20641
rect 36450 20567 36506 20576
rect 36544 20256 36596 20262
rect 36544 20198 36596 20204
rect 36360 18692 36412 18698
rect 36360 18634 36412 18640
rect 36372 17814 36400 18634
rect 36452 18624 36504 18630
rect 36452 18566 36504 18572
rect 36464 18154 36492 18566
rect 36556 18290 36584 20198
rect 36648 18902 36676 20742
rect 36636 18896 36688 18902
rect 36636 18838 36688 18844
rect 36544 18284 36596 18290
rect 36544 18226 36596 18232
rect 36452 18148 36504 18154
rect 36452 18090 36504 18096
rect 36636 18080 36688 18086
rect 36636 18022 36688 18028
rect 36648 17882 36676 18022
rect 36636 17876 36688 17882
rect 36636 17818 36688 17824
rect 36360 17808 36412 17814
rect 36360 17750 36412 17756
rect 36544 17536 36596 17542
rect 36544 17478 36596 17484
rect 36556 17241 36584 17478
rect 36542 17232 36598 17241
rect 36542 17167 36598 17176
rect 36266 16688 36322 16697
rect 36266 16623 36322 16632
rect 36360 16448 36412 16454
rect 36360 16390 36412 16396
rect 36266 16280 36322 16289
rect 36266 16215 36322 16224
rect 36280 16114 36308 16215
rect 36268 16108 36320 16114
rect 36268 16050 36320 16056
rect 36268 14612 36320 14618
rect 36268 14554 36320 14560
rect 36280 13938 36308 14554
rect 36268 13932 36320 13938
rect 36268 13874 36320 13880
rect 36372 13818 36400 16390
rect 36544 16108 36596 16114
rect 36544 16050 36596 16056
rect 36280 13790 36400 13818
rect 36452 13796 36504 13802
rect 36176 12980 36228 12986
rect 36176 12922 36228 12928
rect 36280 12238 36308 13790
rect 36452 13738 36504 13744
rect 36360 13456 36412 13462
rect 36360 13398 36412 13404
rect 36372 13297 36400 13398
rect 36464 13326 36492 13738
rect 36452 13320 36504 13326
rect 36358 13288 36414 13297
rect 36452 13262 36504 13268
rect 36358 13223 36414 13232
rect 36464 12458 36492 13262
rect 36556 12850 36584 16050
rect 36740 13802 36768 20878
rect 36728 13796 36780 13802
rect 36728 13738 36780 13744
rect 36636 13184 36688 13190
rect 36636 13126 36688 13132
rect 36544 12844 36596 12850
rect 36648 12832 36676 13126
rect 36648 12804 36768 12832
rect 36544 12786 36596 12792
rect 36556 12594 36584 12786
rect 36556 12566 36676 12594
rect 36464 12430 36584 12458
rect 36452 12300 36504 12306
rect 36452 12242 36504 12248
rect 36268 12232 36320 12238
rect 36268 12174 36320 12180
rect 36268 12096 36320 12102
rect 36268 12038 36320 12044
rect 36084 11756 36136 11762
rect 36084 11698 36136 11704
rect 36084 11348 36136 11354
rect 36084 11290 36136 11296
rect 36176 11348 36228 11354
rect 36176 11290 36228 11296
rect 36096 11150 36124 11290
rect 36188 11150 36216 11290
rect 36084 11144 36136 11150
rect 36084 11086 36136 11092
rect 36176 11144 36228 11150
rect 36176 11086 36228 11092
rect 35992 11076 36044 11082
rect 35992 11018 36044 11024
rect 35900 10736 35952 10742
rect 35900 10678 35952 10684
rect 36004 10146 36032 11018
rect 36096 10996 36124 11086
rect 36280 10996 36308 12038
rect 36360 11552 36412 11558
rect 36360 11494 36412 11500
rect 36372 11286 36400 11494
rect 36360 11280 36412 11286
rect 36360 11222 36412 11228
rect 36360 11144 36412 11150
rect 36360 11086 36412 11092
rect 36096 10968 36308 10996
rect 36084 10668 36136 10674
rect 36084 10610 36136 10616
rect 35912 10118 36032 10146
rect 35716 9648 35768 9654
rect 35716 9590 35768 9596
rect 35808 8968 35860 8974
rect 35808 8910 35860 8916
rect 35820 8634 35848 8910
rect 35808 8628 35860 8634
rect 35808 8570 35860 8576
rect 35912 8566 35940 10118
rect 35992 9376 36044 9382
rect 35992 9318 36044 9324
rect 36004 9178 36032 9318
rect 35992 9172 36044 9178
rect 35992 9114 36044 9120
rect 36096 9058 36124 10610
rect 36372 10606 36400 11086
rect 36360 10600 36412 10606
rect 36360 10542 36412 10548
rect 36004 9030 36124 9058
rect 36004 8906 36032 9030
rect 35992 8900 36044 8906
rect 35992 8842 36044 8848
rect 35900 8560 35952 8566
rect 35900 8502 35952 8508
rect 35898 8392 35954 8401
rect 35898 8327 35954 8336
rect 35716 8288 35768 8294
rect 35622 8256 35678 8265
rect 35716 8230 35768 8236
rect 35622 8191 35678 8200
rect 35636 7449 35664 8191
rect 35728 7818 35756 8230
rect 35716 7812 35768 7818
rect 35716 7754 35768 7760
rect 35808 7812 35860 7818
rect 35808 7754 35860 7760
rect 35728 7546 35756 7754
rect 35716 7540 35768 7546
rect 35716 7482 35768 7488
rect 35622 7440 35678 7449
rect 35716 7404 35768 7410
rect 35678 7384 35716 7392
rect 35622 7375 35716 7384
rect 35636 7364 35716 7375
rect 35716 7346 35768 7352
rect 35544 7274 35756 7290
rect 35544 7268 35768 7274
rect 35544 7262 35716 7268
rect 35716 7210 35768 7216
rect 35624 7200 35676 7206
rect 35624 7142 35676 7148
rect 35636 6866 35664 7142
rect 35820 6905 35848 7754
rect 35912 7206 35940 8327
rect 36004 7886 36032 8842
rect 36082 7984 36138 7993
rect 36082 7919 36138 7928
rect 35992 7880 36044 7886
rect 35992 7822 36044 7828
rect 36096 7750 36124 7919
rect 36084 7744 36136 7750
rect 36084 7686 36136 7692
rect 36464 7546 36492 12242
rect 36176 7540 36228 7546
rect 36176 7482 36228 7488
rect 36452 7540 36504 7546
rect 36452 7482 36504 7488
rect 35992 7472 36044 7478
rect 35992 7414 36044 7420
rect 36004 7313 36032 7414
rect 35990 7304 36046 7313
rect 35990 7239 36046 7248
rect 35900 7200 35952 7206
rect 35900 7142 35952 7148
rect 35806 6896 35862 6905
rect 35624 6860 35676 6866
rect 35806 6831 35862 6840
rect 35624 6802 35676 6808
rect 35820 6798 35848 6831
rect 35808 6792 35860 6798
rect 35348 6734 35400 6740
rect 35438 6760 35494 6769
rect 33876 6724 33928 6730
rect 33876 6666 33928 6672
rect 33980 6633 34008 6734
rect 34336 6724 34388 6730
rect 34336 6666 34388 6672
rect 33966 6624 34022 6633
rect 33966 6559 34022 6568
rect 33692 6384 33744 6390
rect 33692 6326 33744 6332
rect 33600 6112 33652 6118
rect 33600 6054 33652 6060
rect 33612 5914 33640 6054
rect 33600 5908 33652 5914
rect 33600 5850 33652 5856
rect 33612 5710 33640 5850
rect 33704 5710 33732 6326
rect 34348 6254 34376 6666
rect 34440 6458 34468 6734
rect 35808 6734 35860 6740
rect 35438 6695 35494 6704
rect 35452 6644 35480 6695
rect 35532 6656 35584 6662
rect 35452 6616 35532 6644
rect 35532 6598 35584 6604
rect 34428 6452 34480 6458
rect 34428 6394 34480 6400
rect 34336 6248 34388 6254
rect 34336 6190 34388 6196
rect 34796 6248 34848 6254
rect 34796 6190 34848 6196
rect 34152 6180 34204 6186
rect 34152 6122 34204 6128
rect 34164 5710 34192 6122
rect 34612 6112 34664 6118
rect 34808 6066 34836 6190
rect 34664 6060 34836 6066
rect 34612 6054 34836 6060
rect 35716 6112 35768 6118
rect 35716 6054 35768 6060
rect 34624 6038 34836 6054
rect 34808 5778 34836 6038
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34796 5772 34848 5778
rect 34796 5714 34848 5720
rect 33600 5704 33652 5710
rect 33600 5646 33652 5652
rect 33692 5704 33744 5710
rect 33692 5646 33744 5652
rect 34152 5704 34204 5710
rect 34152 5646 34204 5652
rect 33508 5296 33560 5302
rect 33508 5238 33560 5244
rect 31024 5228 31076 5234
rect 31024 5170 31076 5176
rect 31760 5228 31812 5234
rect 31760 5170 31812 5176
rect 32588 5228 32640 5234
rect 32588 5170 32640 5176
rect 33232 5228 33284 5234
rect 33232 5170 33284 5176
rect 30932 5024 30984 5030
rect 30932 4966 30984 4972
rect 31668 5024 31720 5030
rect 31668 4966 31720 4972
rect 30012 4684 30064 4690
rect 30012 4626 30064 4632
rect 30564 4548 30616 4554
rect 30564 4490 30616 4496
rect 30576 4282 30604 4490
rect 30944 4282 30972 4966
rect 31680 4690 31708 4966
rect 31772 4826 31800 5170
rect 32956 5024 33008 5030
rect 32956 4966 33008 4972
rect 31760 4820 31812 4826
rect 31760 4762 31812 4768
rect 32968 4690 32996 4966
rect 33612 4826 33640 5646
rect 34336 5568 34388 5574
rect 34336 5510 34388 5516
rect 34348 5409 34376 5510
rect 34334 5400 34390 5409
rect 34334 5335 34390 5344
rect 34060 5296 34112 5302
rect 34060 5238 34112 5244
rect 33600 4820 33652 4826
rect 33600 4762 33652 4768
rect 31668 4684 31720 4690
rect 31668 4626 31720 4632
rect 32956 4684 33008 4690
rect 32956 4626 33008 4632
rect 34072 4486 34100 5238
rect 34808 5166 34836 5714
rect 35728 5710 35756 6054
rect 36188 5914 36216 7482
rect 36452 7404 36504 7410
rect 36452 7346 36504 7352
rect 36464 7002 36492 7346
rect 36556 7206 36584 12430
rect 36648 11898 36676 12566
rect 36636 11892 36688 11898
rect 36636 11834 36688 11840
rect 36636 11756 36688 11762
rect 36636 11698 36688 11704
rect 36648 11286 36676 11698
rect 36636 11280 36688 11286
rect 36636 11222 36688 11228
rect 36636 11008 36688 11014
rect 36740 10996 36768 12804
rect 36832 12102 36860 28426
rect 36924 28082 36952 29582
rect 37004 29504 37056 29510
rect 37004 29446 37056 29452
rect 37016 29345 37044 29446
rect 37002 29336 37058 29345
rect 37002 29271 37058 29280
rect 37384 29073 37412 30223
rect 37476 29850 37504 31962
rect 37568 31822 37596 32166
rect 37660 31822 37688 32710
rect 37556 31816 37608 31822
rect 37556 31758 37608 31764
rect 37648 31816 37700 31822
rect 37648 31758 37700 31764
rect 37568 30938 37596 31758
rect 37556 30932 37608 30938
rect 37556 30874 37608 30880
rect 37660 30870 37688 31758
rect 37648 30864 37700 30870
rect 37648 30806 37700 30812
rect 37556 30116 37608 30122
rect 37556 30058 37608 30064
rect 37464 29844 37516 29850
rect 37464 29786 37516 29792
rect 37464 29164 37516 29170
rect 37464 29106 37516 29112
rect 37370 29064 37426 29073
rect 37370 28999 37372 29008
rect 37424 28999 37426 29008
rect 37372 28970 37424 28976
rect 37476 28218 37504 29106
rect 37568 28558 37596 30058
rect 37648 29572 37700 29578
rect 37648 29514 37700 29520
rect 37660 29170 37688 29514
rect 37648 29164 37700 29170
rect 37648 29106 37700 29112
rect 37648 28960 37700 28966
rect 37648 28902 37700 28908
rect 37556 28552 37608 28558
rect 37556 28494 37608 28500
rect 37464 28212 37516 28218
rect 37464 28154 37516 28160
rect 36912 28076 36964 28082
rect 36912 28018 36964 28024
rect 37372 28008 37424 28014
rect 37372 27950 37424 27956
rect 37280 27872 37332 27878
rect 37280 27814 37332 27820
rect 37292 27470 37320 27814
rect 37384 27538 37412 27950
rect 37372 27532 37424 27538
rect 37372 27474 37424 27480
rect 37280 27464 37332 27470
rect 37280 27406 37332 27412
rect 37384 26994 37412 27474
rect 37004 26988 37056 26994
rect 37004 26930 37056 26936
rect 37372 26988 37424 26994
rect 37372 26930 37424 26936
rect 37016 25294 37044 26930
rect 37372 26580 37424 26586
rect 37372 26522 37424 26528
rect 37096 26308 37148 26314
rect 37096 26250 37148 26256
rect 37108 25294 37136 26250
rect 37384 25294 37412 26522
rect 37476 26042 37504 28154
rect 37556 27872 37608 27878
rect 37660 27860 37688 28902
rect 37608 27832 37688 27860
rect 37556 27814 37608 27820
rect 37568 26586 37596 27814
rect 37648 27668 37700 27674
rect 37648 27610 37700 27616
rect 37660 26790 37688 27610
rect 37752 26874 37780 34478
rect 37832 33924 37884 33930
rect 37832 33866 37884 33872
rect 37844 33522 37872 33866
rect 37832 33516 37884 33522
rect 37832 33458 37884 33464
rect 38016 33516 38068 33522
rect 38016 33458 38068 33464
rect 37844 32842 37872 33458
rect 38028 33114 38056 33458
rect 39212 33448 39264 33454
rect 39212 33390 39264 33396
rect 38384 33380 38436 33386
rect 38384 33322 38436 33328
rect 38396 33114 38424 33322
rect 38016 33108 38068 33114
rect 38016 33050 38068 33056
rect 38384 33108 38436 33114
rect 38384 33050 38436 33056
rect 37832 32836 37884 32842
rect 37832 32778 37884 32784
rect 38028 32570 38056 33050
rect 38108 32904 38160 32910
rect 38108 32846 38160 32852
rect 38016 32564 38068 32570
rect 38016 32506 38068 32512
rect 37832 32496 37884 32502
rect 37832 32438 37884 32444
rect 37844 28694 37872 32438
rect 38028 32434 38056 32506
rect 38016 32428 38068 32434
rect 38016 32370 38068 32376
rect 38028 31346 38056 32370
rect 38120 32298 38148 32846
rect 38396 32434 38424 33050
rect 38476 32972 38528 32978
rect 38476 32914 38528 32920
rect 38488 32434 38516 32914
rect 38660 32904 38712 32910
rect 38660 32846 38712 32852
rect 38568 32768 38620 32774
rect 38568 32710 38620 32716
rect 38384 32428 38436 32434
rect 38384 32370 38436 32376
rect 38476 32428 38528 32434
rect 38476 32370 38528 32376
rect 38108 32292 38160 32298
rect 38108 32234 38160 32240
rect 38580 31958 38608 32710
rect 38672 32570 38700 32846
rect 38660 32564 38712 32570
rect 38660 32506 38712 32512
rect 39224 32502 39252 33390
rect 39856 32904 39908 32910
rect 39856 32846 39908 32852
rect 39580 32768 39632 32774
rect 39580 32710 39632 32716
rect 39212 32496 39264 32502
rect 39212 32438 39264 32444
rect 38568 31952 38620 31958
rect 38568 31894 38620 31900
rect 39224 31754 39252 32438
rect 39592 32366 39620 32710
rect 39580 32360 39632 32366
rect 39580 32302 39632 32308
rect 38200 31748 38252 31754
rect 38200 31690 38252 31696
rect 39040 31726 39252 31754
rect 38212 31385 38240 31690
rect 38198 31376 38254 31385
rect 38016 31340 38068 31346
rect 38198 31311 38254 31320
rect 38568 31340 38620 31346
rect 38016 31282 38068 31288
rect 38568 31282 38620 31288
rect 38936 31340 38988 31346
rect 38936 31282 38988 31288
rect 38028 30734 38056 31282
rect 38200 31272 38252 31278
rect 38200 31214 38252 31220
rect 38212 30938 38240 31214
rect 38384 31136 38436 31142
rect 38384 31078 38436 31084
rect 38200 30932 38252 30938
rect 38200 30874 38252 30880
rect 38396 30734 38424 31078
rect 38580 30802 38608 31282
rect 38660 31136 38712 31142
rect 38660 31078 38712 31084
rect 38752 31136 38804 31142
rect 38752 31078 38804 31084
rect 38568 30796 38620 30802
rect 38568 30738 38620 30744
rect 38016 30728 38068 30734
rect 38016 30670 38068 30676
rect 38384 30728 38436 30734
rect 38384 30670 38436 30676
rect 38016 30048 38068 30054
rect 38016 29990 38068 29996
rect 38028 28994 38056 29990
rect 38200 29844 38252 29850
rect 38200 29786 38252 29792
rect 38028 28966 38148 28994
rect 37832 28688 37884 28694
rect 37884 28636 38056 28642
rect 37832 28630 38056 28636
rect 37844 28614 38056 28630
rect 37832 28552 37884 28558
rect 37832 28494 37884 28500
rect 37844 26994 37872 28494
rect 38028 28082 38056 28614
rect 38016 28076 38068 28082
rect 38016 28018 38068 28024
rect 38120 26994 38148 28966
rect 38212 28529 38240 29786
rect 38396 29628 38424 30670
rect 38476 30592 38528 30598
rect 38476 30534 38528 30540
rect 38488 30326 38516 30534
rect 38580 30394 38608 30738
rect 38568 30388 38620 30394
rect 38568 30330 38620 30336
rect 38476 30320 38528 30326
rect 38476 30262 38528 30268
rect 38672 30122 38700 31078
rect 38764 30938 38792 31078
rect 38752 30932 38804 30938
rect 38752 30874 38804 30880
rect 38764 30258 38792 30874
rect 38844 30728 38896 30734
rect 38844 30670 38896 30676
rect 38856 30598 38884 30670
rect 38948 30666 38976 31282
rect 39040 31278 39068 31726
rect 39028 31272 39080 31278
rect 39028 31214 39080 31220
rect 39580 31272 39632 31278
rect 39580 31214 39632 31220
rect 38936 30660 38988 30666
rect 38936 30602 38988 30608
rect 38844 30592 38896 30598
rect 38844 30534 38896 30540
rect 38752 30252 38804 30258
rect 38752 30194 38804 30200
rect 38660 30116 38712 30122
rect 38660 30058 38712 30064
rect 38568 29776 38620 29782
rect 38568 29718 38620 29724
rect 38476 29640 38528 29646
rect 38396 29600 38476 29628
rect 38476 29582 38528 29588
rect 38580 28994 38608 29718
rect 38764 29646 38792 30194
rect 38856 30054 38884 30534
rect 38948 30122 38976 30602
rect 39040 30190 39068 31214
rect 39592 30938 39620 31214
rect 39580 30932 39632 30938
rect 39580 30874 39632 30880
rect 39212 30592 39264 30598
rect 39212 30534 39264 30540
rect 39028 30184 39080 30190
rect 39028 30126 39080 30132
rect 38936 30116 38988 30122
rect 38936 30058 38988 30064
rect 38844 30048 38896 30054
rect 38844 29990 38896 29996
rect 38752 29640 38804 29646
rect 38752 29582 38804 29588
rect 38856 29510 38884 29990
rect 38948 29850 38976 30058
rect 38936 29844 38988 29850
rect 38936 29786 38988 29792
rect 38752 29504 38804 29510
rect 38752 29446 38804 29452
rect 38844 29504 38896 29510
rect 38844 29446 38896 29452
rect 38488 28966 38608 28994
rect 38382 28656 38438 28665
rect 38382 28591 38438 28600
rect 38198 28520 38254 28529
rect 38198 28455 38254 28464
rect 38212 27470 38240 28455
rect 38396 28218 38424 28591
rect 38384 28212 38436 28218
rect 38384 28154 38436 28160
rect 38292 28076 38344 28082
rect 38292 28018 38344 28024
rect 38200 27464 38252 27470
rect 38200 27406 38252 27412
rect 38304 27402 38332 28018
rect 38396 27713 38424 28154
rect 38382 27704 38438 27713
rect 38382 27639 38438 27648
rect 38488 27470 38516 28966
rect 38764 27656 38792 29446
rect 38856 29034 38884 29446
rect 38844 29028 38896 29034
rect 38844 28970 38896 28976
rect 39040 28082 39068 30126
rect 39120 30048 39172 30054
rect 39120 29990 39172 29996
rect 39132 29306 39160 29990
rect 39224 29714 39252 30534
rect 39580 30184 39632 30190
rect 39580 30126 39632 30132
rect 39592 29850 39620 30126
rect 39580 29844 39632 29850
rect 39580 29786 39632 29792
rect 39212 29708 39264 29714
rect 39212 29650 39264 29656
rect 39868 29345 39896 32846
rect 40052 31414 40080 36858
rect 40788 36378 40816 37198
rect 40960 37120 41012 37126
rect 40960 37062 41012 37068
rect 40972 36825 41000 37062
rect 40958 36816 41014 36825
rect 40958 36751 41014 36760
rect 40776 36372 40828 36378
rect 40776 36314 40828 36320
rect 40592 33516 40644 33522
rect 40592 33458 40644 33464
rect 40500 32904 40552 32910
rect 40500 32846 40552 32852
rect 40512 32570 40540 32846
rect 40500 32564 40552 32570
rect 40500 32506 40552 32512
rect 40604 32434 40632 33458
rect 41052 33448 41104 33454
rect 41052 33390 41104 33396
rect 40960 33312 41012 33318
rect 40960 33254 41012 33260
rect 40972 32858 41000 33254
rect 41064 33114 41092 33390
rect 41052 33108 41104 33114
rect 41052 33050 41104 33056
rect 40972 32830 41092 32858
rect 40958 32736 41014 32745
rect 40958 32671 41014 32680
rect 40972 32570 41000 32671
rect 40960 32564 41012 32570
rect 40960 32506 41012 32512
rect 40774 32464 40830 32473
rect 40592 32428 40644 32434
rect 40774 32399 40776 32408
rect 40592 32370 40644 32376
rect 40828 32399 40830 32408
rect 40776 32370 40828 32376
rect 40040 31408 40092 31414
rect 40040 31350 40092 31356
rect 40052 30326 40080 31350
rect 40040 30320 40092 30326
rect 40040 30262 40092 30268
rect 39854 29336 39910 29345
rect 39120 29300 39172 29306
rect 39854 29271 39910 29280
rect 39120 29242 39172 29248
rect 39488 29028 39540 29034
rect 39488 28970 39540 28976
rect 39028 28076 39080 28082
rect 39028 28018 39080 28024
rect 39304 28008 39356 28014
rect 39304 27950 39356 27956
rect 39316 27674 39344 27950
rect 39304 27668 39356 27674
rect 38764 27628 39160 27656
rect 38476 27464 38528 27470
rect 38396 27424 38476 27452
rect 38292 27396 38344 27402
rect 38292 27338 38344 27344
rect 38304 27062 38332 27338
rect 38292 27056 38344 27062
rect 38292 26998 38344 27004
rect 37832 26988 37884 26994
rect 38108 26988 38160 26994
rect 37832 26930 37884 26936
rect 38028 26948 38108 26976
rect 37752 26846 37964 26874
rect 37648 26784 37700 26790
rect 37648 26726 37700 26732
rect 37556 26580 37608 26586
rect 37556 26522 37608 26528
rect 37464 26036 37516 26042
rect 37464 25978 37516 25984
rect 37464 25900 37516 25906
rect 37464 25842 37516 25848
rect 37004 25288 37056 25294
rect 37004 25230 37056 25236
rect 37096 25288 37148 25294
rect 37096 25230 37148 25236
rect 37372 25288 37424 25294
rect 37372 25230 37424 25236
rect 37016 23526 37044 25230
rect 37096 25152 37148 25158
rect 37096 25094 37148 25100
rect 37108 24993 37136 25094
rect 37094 24984 37150 24993
rect 37094 24919 37150 24928
rect 37280 24200 37332 24206
rect 37280 24142 37332 24148
rect 37004 23520 37056 23526
rect 37292 23474 37320 24142
rect 37372 24064 37424 24070
rect 37372 24006 37424 24012
rect 37004 23462 37056 23468
rect 37200 23446 37320 23474
rect 37200 23118 37228 23446
rect 37188 23112 37240 23118
rect 37188 23054 37240 23060
rect 37280 22976 37332 22982
rect 37280 22918 37332 22924
rect 37292 21622 37320 22918
rect 37280 21616 37332 21622
rect 37280 21558 37332 21564
rect 37384 21486 37412 24006
rect 37476 23730 37504 25842
rect 37556 25424 37608 25430
rect 37556 25366 37608 25372
rect 37568 24274 37596 25366
rect 37556 24268 37608 24274
rect 37556 24210 37608 24216
rect 37464 23724 37516 23730
rect 37464 23666 37516 23672
rect 37556 23588 37608 23594
rect 37556 23530 37608 23536
rect 37568 23497 37596 23530
rect 37554 23488 37610 23497
rect 37554 23423 37610 23432
rect 37464 22976 37516 22982
rect 37464 22918 37516 22924
rect 37476 22778 37504 22918
rect 37464 22772 37516 22778
rect 37464 22714 37516 22720
rect 37660 22094 37688 26726
rect 37740 26036 37792 26042
rect 37740 25978 37792 25984
rect 37752 25401 37780 25978
rect 37832 25900 37884 25906
rect 37832 25842 37884 25848
rect 37844 25498 37872 25842
rect 37832 25492 37884 25498
rect 37832 25434 37884 25440
rect 37738 25392 37794 25401
rect 37738 25327 37794 25336
rect 37740 25152 37792 25158
rect 37740 25094 37792 25100
rect 37752 24206 37780 25094
rect 37740 24200 37792 24206
rect 37740 24142 37792 24148
rect 37832 24200 37884 24206
rect 37832 24142 37884 24148
rect 37844 23866 37872 24142
rect 37832 23860 37884 23866
rect 37832 23802 37884 23808
rect 37740 23520 37792 23526
rect 37738 23488 37740 23497
rect 37792 23488 37794 23497
rect 37738 23423 37794 23432
rect 37832 22432 37884 22438
rect 37832 22374 37884 22380
rect 37660 22066 37780 22094
rect 37464 21548 37516 21554
rect 37464 21490 37516 21496
rect 37372 21480 37424 21486
rect 37372 21422 37424 21428
rect 36912 21140 36964 21146
rect 36912 21082 36964 21088
rect 36924 17678 36952 21082
rect 37476 21078 37504 21490
rect 37648 21344 37700 21350
rect 37648 21286 37700 21292
rect 37280 21072 37332 21078
rect 37464 21072 37516 21078
rect 37332 21020 37412 21026
rect 37280 21014 37412 21020
rect 37464 21014 37516 21020
rect 37292 20998 37412 21014
rect 37188 20868 37240 20874
rect 37240 20828 37320 20856
rect 37188 20810 37240 20816
rect 37186 20768 37242 20777
rect 37186 20703 37242 20712
rect 37096 18080 37148 18086
rect 37096 18022 37148 18028
rect 36912 17672 36964 17678
rect 36912 17614 36964 17620
rect 37004 15496 37056 15502
rect 37004 15438 37056 15444
rect 37016 14822 37044 15438
rect 37004 14816 37056 14822
rect 37004 14758 37056 14764
rect 37016 14414 37044 14758
rect 37108 14618 37136 18022
rect 37200 15570 37228 20703
rect 37292 18970 37320 20828
rect 37384 20466 37412 20998
rect 37464 20936 37516 20942
rect 37464 20878 37516 20884
rect 37476 20602 37504 20878
rect 37464 20596 37516 20602
rect 37464 20538 37516 20544
rect 37372 20460 37424 20466
rect 37556 20460 37608 20466
rect 37372 20402 37424 20408
rect 37476 20420 37556 20448
rect 37372 20256 37424 20262
rect 37372 20198 37424 20204
rect 37384 19242 37412 20198
rect 37372 19236 37424 19242
rect 37372 19178 37424 19184
rect 37280 18964 37332 18970
rect 37280 18906 37332 18912
rect 37384 18766 37412 19178
rect 37372 18760 37424 18766
rect 37372 18702 37424 18708
rect 37280 18692 37332 18698
rect 37280 18634 37332 18640
rect 37292 16250 37320 18634
rect 37372 16992 37424 16998
rect 37372 16934 37424 16940
rect 37384 16794 37412 16934
rect 37372 16788 37424 16794
rect 37372 16730 37424 16736
rect 37476 16674 37504 20420
rect 37556 20402 37608 20408
rect 37556 18828 37608 18834
rect 37556 18770 37608 18776
rect 37568 17746 37596 18770
rect 37660 18358 37688 21286
rect 37752 20942 37780 22066
rect 37844 21350 37872 22374
rect 37832 21344 37884 21350
rect 37832 21286 37884 21292
rect 37740 20936 37792 20942
rect 37740 20878 37792 20884
rect 37936 20346 37964 26846
rect 38028 23866 38056 26948
rect 38108 26930 38160 26936
rect 38304 26586 38332 26998
rect 38292 26580 38344 26586
rect 38292 26522 38344 26528
rect 38304 25906 38332 26522
rect 38292 25900 38344 25906
rect 38292 25842 38344 25848
rect 38292 25696 38344 25702
rect 38292 25638 38344 25644
rect 38304 25362 38332 25638
rect 38292 25356 38344 25362
rect 38292 25298 38344 25304
rect 38108 25152 38160 25158
rect 38108 25094 38160 25100
rect 38016 23860 38068 23866
rect 38016 23802 38068 23808
rect 38016 21684 38068 21690
rect 38016 21626 38068 21632
rect 38028 20942 38056 21626
rect 38016 20936 38068 20942
rect 38016 20878 38068 20884
rect 38016 20800 38068 20806
rect 38016 20742 38068 20748
rect 37752 20318 37964 20346
rect 37752 19174 37780 20318
rect 37924 19712 37976 19718
rect 37924 19654 37976 19660
rect 37740 19168 37792 19174
rect 37740 19110 37792 19116
rect 37832 18964 37884 18970
rect 37832 18906 37884 18912
rect 37648 18352 37700 18358
rect 37648 18294 37700 18300
rect 37648 18216 37700 18222
rect 37648 18158 37700 18164
rect 37556 17740 37608 17746
rect 37556 17682 37608 17688
rect 37384 16646 37504 16674
rect 37384 16590 37412 16646
rect 37372 16584 37424 16590
rect 37372 16526 37424 16532
rect 37464 16584 37516 16590
rect 37464 16526 37516 16532
rect 37280 16244 37332 16250
rect 37280 16186 37332 16192
rect 37278 16144 37334 16153
rect 37334 16102 37412 16130
rect 37476 16114 37504 16526
rect 37556 16244 37608 16250
rect 37556 16186 37608 16192
rect 37278 16079 37334 16088
rect 37384 15910 37412 16102
rect 37464 16108 37516 16114
rect 37464 16050 37516 16056
rect 37372 15904 37424 15910
rect 37372 15846 37424 15852
rect 37188 15564 37240 15570
rect 37188 15506 37240 15512
rect 37188 15360 37240 15366
rect 37188 15302 37240 15308
rect 37096 14612 37148 14618
rect 37096 14554 37148 14560
rect 36912 14408 36964 14414
rect 36912 14350 36964 14356
rect 37004 14408 37056 14414
rect 37004 14350 37056 14356
rect 36924 13938 36952 14350
rect 37094 14240 37150 14249
rect 37094 14175 37150 14184
rect 36912 13932 36964 13938
rect 36912 13874 36964 13880
rect 36820 12096 36872 12102
rect 36820 12038 36872 12044
rect 36820 11892 36872 11898
rect 36820 11834 36872 11840
rect 36832 11801 36860 11834
rect 36818 11792 36874 11801
rect 36818 11727 36874 11736
rect 36832 11150 36860 11727
rect 36820 11144 36872 11150
rect 36820 11086 36872 11092
rect 36832 11014 36860 11086
rect 36688 10968 36768 10996
rect 36820 11008 36872 11014
rect 36636 10950 36688 10956
rect 36820 10950 36872 10956
rect 36924 7546 36952 13874
rect 37004 13796 37056 13802
rect 37004 13738 37056 13744
rect 37016 12306 37044 13738
rect 37004 12300 37056 12306
rect 37004 12242 37056 12248
rect 37108 11014 37136 14175
rect 37200 14074 37228 15302
rect 37188 14068 37240 14074
rect 37188 14010 37240 14016
rect 37280 13932 37332 13938
rect 37280 13874 37332 13880
rect 37292 13433 37320 13874
rect 37278 13424 37334 13433
rect 37278 13359 37334 13368
rect 37280 13320 37332 13326
rect 37280 13262 37332 13268
rect 37188 13252 37240 13258
rect 37188 13194 37240 13200
rect 37200 12442 37228 13194
rect 37292 13025 37320 13262
rect 37278 13016 37334 13025
rect 37278 12951 37334 12960
rect 37188 12436 37240 12442
rect 37188 12378 37240 12384
rect 37188 12164 37240 12170
rect 37188 12106 37240 12112
rect 37200 11082 37228 12106
rect 37188 11076 37240 11082
rect 37188 11018 37240 11024
rect 37096 11008 37148 11014
rect 37096 10950 37148 10956
rect 37384 9042 37412 15846
rect 37476 15706 37504 16050
rect 37568 15910 37596 16186
rect 37556 15904 37608 15910
rect 37556 15846 37608 15852
rect 37464 15700 37516 15706
rect 37464 15642 37516 15648
rect 37464 15496 37516 15502
rect 37464 15438 37516 15444
rect 37476 11898 37504 15438
rect 37554 15192 37610 15201
rect 37554 15127 37610 15136
rect 37660 15144 37688 18158
rect 37740 17672 37792 17678
rect 37740 17614 37792 17620
rect 37752 16794 37780 17614
rect 37740 16788 37792 16794
rect 37740 16730 37792 16736
rect 37568 14006 37596 15127
rect 37660 15116 37780 15144
rect 37648 15020 37700 15026
rect 37648 14962 37700 14968
rect 37556 14000 37608 14006
rect 37556 13942 37608 13948
rect 37660 13326 37688 14962
rect 37648 13320 37700 13326
rect 37648 13262 37700 13268
rect 37464 11892 37516 11898
rect 37464 11834 37516 11840
rect 37660 11286 37688 13262
rect 37752 11694 37780 15116
rect 37844 14906 37872 18906
rect 37936 18766 37964 19654
rect 38028 18970 38056 20742
rect 38016 18964 38068 18970
rect 38016 18906 38068 18912
rect 37924 18760 37976 18766
rect 37924 18702 37976 18708
rect 37936 18442 37964 18702
rect 38120 18698 38148 25094
rect 38304 24410 38332 25298
rect 38292 24404 38344 24410
rect 38292 24346 38344 24352
rect 38304 23730 38332 24346
rect 38396 24206 38424 27424
rect 38476 27406 38528 27412
rect 38844 27464 38896 27470
rect 38844 27406 38896 27412
rect 38856 26790 38884 27406
rect 38844 26784 38896 26790
rect 38844 26726 38896 26732
rect 38384 24200 38436 24206
rect 38384 24142 38436 24148
rect 38660 24132 38712 24138
rect 38660 24074 38712 24080
rect 38476 24064 38528 24070
rect 38476 24006 38528 24012
rect 38292 23724 38344 23730
rect 38292 23666 38344 23672
rect 38384 23724 38436 23730
rect 38384 23666 38436 23672
rect 38292 21072 38344 21078
rect 38292 21014 38344 21020
rect 38304 18902 38332 21014
rect 38292 18896 38344 18902
rect 38292 18838 38344 18844
rect 38108 18692 38160 18698
rect 38108 18634 38160 18640
rect 38200 18624 38252 18630
rect 38200 18566 38252 18572
rect 37936 18414 38056 18442
rect 38212 18426 38240 18566
rect 37924 18284 37976 18290
rect 37924 18226 37976 18232
rect 37936 17882 37964 18226
rect 37924 17876 37976 17882
rect 37924 17818 37976 17824
rect 38028 17746 38056 18414
rect 38200 18420 38252 18426
rect 38200 18362 38252 18368
rect 38108 18284 38160 18290
rect 38108 18226 38160 18232
rect 38120 18086 38148 18226
rect 38108 18080 38160 18086
rect 38108 18022 38160 18028
rect 38016 17740 38068 17746
rect 38016 17682 38068 17688
rect 38200 17604 38252 17610
rect 38200 17546 38252 17552
rect 38108 15020 38160 15026
rect 38108 14962 38160 14968
rect 37844 14878 37964 14906
rect 37832 14408 37884 14414
rect 37832 14350 37884 14356
rect 37844 14074 37872 14350
rect 37832 14068 37884 14074
rect 37832 14010 37884 14016
rect 37830 13696 37886 13705
rect 37830 13631 37886 13640
rect 37844 13326 37872 13631
rect 37936 13530 37964 14878
rect 37924 13524 37976 13530
rect 37924 13466 37976 13472
rect 37936 13410 37964 13466
rect 37936 13382 38056 13410
rect 37832 13320 37884 13326
rect 37832 13262 37884 13268
rect 37740 11688 37792 11694
rect 37740 11630 37792 11636
rect 37648 11280 37700 11286
rect 37648 11222 37700 11228
rect 37556 11144 37608 11150
rect 37556 11086 37608 11092
rect 37568 10606 37596 11086
rect 37660 10674 37688 11222
rect 37648 10668 37700 10674
rect 37648 10610 37700 10616
rect 37556 10600 37608 10606
rect 37556 10542 37608 10548
rect 37832 10464 37884 10470
rect 37832 10406 37884 10412
rect 37844 10266 37872 10406
rect 37832 10260 37884 10266
rect 37832 10202 37884 10208
rect 37462 9616 37518 9625
rect 37462 9551 37518 9560
rect 37476 9178 37504 9551
rect 37464 9172 37516 9178
rect 37464 9114 37516 9120
rect 37372 9036 37424 9042
rect 37372 8978 37424 8984
rect 37844 8974 37872 10202
rect 37832 8968 37884 8974
rect 37832 8910 37884 8916
rect 37924 8968 37976 8974
rect 37924 8910 37976 8916
rect 37936 8634 37964 8910
rect 37924 8628 37976 8634
rect 37924 8570 37976 8576
rect 37464 8492 37516 8498
rect 37464 8434 37516 8440
rect 37556 8492 37608 8498
rect 38028 8480 38056 13382
rect 38120 13326 38148 14962
rect 38212 14618 38240 17546
rect 38396 16454 38424 23666
rect 38488 23662 38516 24006
rect 38672 23780 38700 24074
rect 38752 23792 38804 23798
rect 38672 23752 38752 23780
rect 38476 23656 38528 23662
rect 38476 23598 38528 23604
rect 38568 23112 38620 23118
rect 38568 23054 38620 23060
rect 38580 22642 38608 23054
rect 38672 22710 38700 23752
rect 38752 23734 38804 23740
rect 38752 23520 38804 23526
rect 38752 23462 38804 23468
rect 38764 23050 38792 23462
rect 38752 23044 38804 23050
rect 38752 22986 38804 22992
rect 38660 22704 38712 22710
rect 38660 22646 38712 22652
rect 38568 22636 38620 22642
rect 38568 22578 38620 22584
rect 38660 21480 38712 21486
rect 38660 21422 38712 21428
rect 38476 21412 38528 21418
rect 38476 21354 38528 21360
rect 38488 17105 38516 21354
rect 38568 21344 38620 21350
rect 38568 21286 38620 21292
rect 38580 21146 38608 21286
rect 38568 21140 38620 21146
rect 38568 21082 38620 21088
rect 38566 18592 38622 18601
rect 38566 18527 38622 18536
rect 38474 17096 38530 17105
rect 38474 17031 38530 17040
rect 38384 16448 38436 16454
rect 38384 16390 38436 16396
rect 38384 15428 38436 15434
rect 38384 15370 38436 15376
rect 38396 15094 38424 15370
rect 38384 15088 38436 15094
rect 38384 15030 38436 15036
rect 38488 14958 38516 17031
rect 38580 15094 38608 18527
rect 38672 16794 38700 21422
rect 38764 19310 38792 22986
rect 38856 22710 38884 26726
rect 39028 24812 39080 24818
rect 39028 24754 39080 24760
rect 38936 23724 38988 23730
rect 38936 23666 38988 23672
rect 38844 22704 38896 22710
rect 38844 22646 38896 22652
rect 38844 22500 38896 22506
rect 38844 22442 38896 22448
rect 38856 21554 38884 22442
rect 38844 21548 38896 21554
rect 38948 21536 38976 23666
rect 39040 23254 39068 24754
rect 39132 23866 39160 27628
rect 39304 27610 39356 27616
rect 39396 27328 39448 27334
rect 39396 27270 39448 27276
rect 39408 27130 39436 27270
rect 39500 27130 39528 28970
rect 40052 28150 40080 30262
rect 40040 28144 40092 28150
rect 40040 28086 40092 28092
rect 39856 27464 39908 27470
rect 39856 27406 39908 27412
rect 39396 27124 39448 27130
rect 39396 27066 39448 27072
rect 39488 27124 39540 27130
rect 39488 27066 39540 27072
rect 39304 26784 39356 26790
rect 39304 26726 39356 26732
rect 39212 26240 39264 26246
rect 39212 26182 39264 26188
rect 39224 25974 39252 26182
rect 39212 25968 39264 25974
rect 39212 25910 39264 25916
rect 39316 25838 39344 26726
rect 39764 26308 39816 26314
rect 39764 26250 39816 26256
rect 39776 26042 39804 26250
rect 39764 26036 39816 26042
rect 39764 25978 39816 25984
rect 39304 25832 39356 25838
rect 39304 25774 39356 25780
rect 39580 25832 39632 25838
rect 39580 25774 39632 25780
rect 39316 24750 39344 25774
rect 39592 25498 39620 25774
rect 39580 25492 39632 25498
rect 39580 25434 39632 25440
rect 39776 25294 39804 25978
rect 39764 25288 39816 25294
rect 39764 25230 39816 25236
rect 39304 24744 39356 24750
rect 39304 24686 39356 24692
rect 39580 24744 39632 24750
rect 39580 24686 39632 24692
rect 39592 24410 39620 24686
rect 39580 24404 39632 24410
rect 39580 24346 39632 24352
rect 39120 23860 39172 23866
rect 39120 23802 39172 23808
rect 39580 23724 39632 23730
rect 39580 23666 39632 23672
rect 39120 23588 39172 23594
rect 39120 23530 39172 23536
rect 39028 23248 39080 23254
rect 39028 23190 39080 23196
rect 39028 22636 39080 22642
rect 39028 22578 39080 22584
rect 39040 21690 39068 22578
rect 39132 22574 39160 23530
rect 39592 23118 39620 23666
rect 39764 23520 39816 23526
rect 39764 23462 39816 23468
rect 39580 23112 39632 23118
rect 39580 23054 39632 23060
rect 39212 22976 39264 22982
rect 39212 22918 39264 22924
rect 39120 22568 39172 22574
rect 39120 22510 39172 22516
rect 39224 22438 39252 22918
rect 39396 22636 39448 22642
rect 39396 22578 39448 22584
rect 39120 22432 39172 22438
rect 39120 22374 39172 22380
rect 39212 22432 39264 22438
rect 39212 22374 39264 22380
rect 39028 21684 39080 21690
rect 39028 21626 39080 21632
rect 38948 21508 39068 21536
rect 38844 21490 38896 21496
rect 38856 20777 38884 21490
rect 38936 21004 38988 21010
rect 38936 20946 38988 20952
rect 38842 20768 38898 20777
rect 38842 20703 38898 20712
rect 38948 20602 38976 20946
rect 38936 20596 38988 20602
rect 38936 20538 38988 20544
rect 38844 20392 38896 20398
rect 38844 20334 38896 20340
rect 38856 19786 38884 20334
rect 38844 19780 38896 19786
rect 38844 19722 38896 19728
rect 39040 19334 39068 21508
rect 39132 19446 39160 22374
rect 39408 22234 39436 22578
rect 39488 22568 39540 22574
rect 39488 22510 39540 22516
rect 39396 22228 39448 22234
rect 39396 22170 39448 22176
rect 39212 21344 39264 21350
rect 39212 21286 39264 21292
rect 39304 21344 39356 21350
rect 39304 21286 39356 21292
rect 39224 21146 39252 21286
rect 39212 21140 39264 21146
rect 39212 21082 39264 21088
rect 39212 20800 39264 20806
rect 39212 20742 39264 20748
rect 39224 20602 39252 20742
rect 39212 20596 39264 20602
rect 39212 20538 39264 20544
rect 39120 19440 39172 19446
rect 39120 19382 39172 19388
rect 38752 19304 38804 19310
rect 38752 19246 38804 19252
rect 38948 19306 39068 19334
rect 38752 18760 38804 18766
rect 38752 18702 38804 18708
rect 38660 16788 38712 16794
rect 38660 16730 38712 16736
rect 38660 15904 38712 15910
rect 38660 15846 38712 15852
rect 38672 15162 38700 15846
rect 38764 15162 38792 18702
rect 38844 17876 38896 17882
rect 38844 17818 38896 17824
rect 38660 15156 38712 15162
rect 38660 15098 38712 15104
rect 38752 15156 38804 15162
rect 38752 15098 38804 15104
rect 38568 15088 38620 15094
rect 38568 15030 38620 15036
rect 38476 14952 38528 14958
rect 38476 14894 38528 14900
rect 38200 14612 38252 14618
rect 38200 14554 38252 14560
rect 38660 14612 38712 14618
rect 38660 14554 38712 14560
rect 38108 13320 38160 13326
rect 38108 13262 38160 13268
rect 38120 12442 38148 13262
rect 38212 12986 38240 14554
rect 38566 13424 38622 13433
rect 38566 13359 38622 13368
rect 38200 12980 38252 12986
rect 38200 12922 38252 12928
rect 38108 12436 38160 12442
rect 38108 12378 38160 12384
rect 38580 11937 38608 13359
rect 38672 13258 38700 14554
rect 38764 14482 38792 15098
rect 38752 14476 38804 14482
rect 38752 14418 38804 14424
rect 38856 14414 38884 17818
rect 38948 15502 38976 19306
rect 39120 19304 39172 19310
rect 39120 19246 39172 19252
rect 39028 18692 39080 18698
rect 39028 18634 39080 18640
rect 39040 18154 39068 18634
rect 39028 18148 39080 18154
rect 39028 18090 39080 18096
rect 39040 17678 39068 18090
rect 39028 17672 39080 17678
rect 39028 17614 39080 17620
rect 39028 16108 39080 16114
rect 39028 16050 39080 16056
rect 39040 15706 39068 16050
rect 39028 15700 39080 15706
rect 39028 15642 39080 15648
rect 38936 15496 38988 15502
rect 38936 15438 38988 15444
rect 38948 15026 38976 15438
rect 38936 15020 38988 15026
rect 38936 14962 38988 14968
rect 38844 14408 38896 14414
rect 38844 14350 38896 14356
rect 39132 13870 39160 19246
rect 39316 19174 39344 21286
rect 39500 21010 39528 22510
rect 39776 21010 39804 23462
rect 39868 23322 39896 27406
rect 40052 27062 40080 28086
rect 40406 27976 40462 27985
rect 40406 27911 40462 27920
rect 40040 27056 40092 27062
rect 40040 26998 40092 27004
rect 39948 26308 40000 26314
rect 39948 26250 40000 26256
rect 39960 24750 39988 26250
rect 40052 25974 40080 26998
rect 40040 25968 40092 25974
rect 40092 25916 40172 25922
rect 40040 25910 40172 25916
rect 40052 25894 40172 25910
rect 40144 25498 40172 25894
rect 40132 25492 40184 25498
rect 40132 25434 40184 25440
rect 40040 25288 40092 25294
rect 40040 25230 40092 25236
rect 39948 24744 40000 24750
rect 39948 24686 40000 24692
rect 39856 23316 39908 23322
rect 39856 23258 39908 23264
rect 39948 23044 40000 23050
rect 39948 22986 40000 22992
rect 39960 22778 39988 22986
rect 39948 22772 40000 22778
rect 39948 22714 40000 22720
rect 39856 22432 39908 22438
rect 39856 22374 39908 22380
rect 39488 21004 39540 21010
rect 39488 20946 39540 20952
rect 39764 21004 39816 21010
rect 39764 20946 39816 20952
rect 39672 20936 39724 20942
rect 39672 20878 39724 20884
rect 39580 20256 39632 20262
rect 39580 20198 39632 20204
rect 39488 19780 39540 19786
rect 39488 19722 39540 19728
rect 39304 19168 39356 19174
rect 39304 19110 39356 19116
rect 39396 17536 39448 17542
rect 39396 17478 39448 17484
rect 39212 16584 39264 16590
rect 39212 16526 39264 16532
rect 39224 15910 39252 16526
rect 39304 16516 39356 16522
rect 39304 16458 39356 16464
rect 39212 15904 39264 15910
rect 39212 15846 39264 15852
rect 39212 14408 39264 14414
rect 39212 14350 39264 14356
rect 38936 13864 38988 13870
rect 38936 13806 38988 13812
rect 39120 13864 39172 13870
rect 39120 13806 39172 13812
rect 38764 13394 38884 13410
rect 38764 13388 38896 13394
rect 38764 13382 38844 13388
rect 38660 13252 38712 13258
rect 38660 13194 38712 13200
rect 38660 12776 38712 12782
rect 38660 12718 38712 12724
rect 38566 11928 38622 11937
rect 38566 11863 38622 11872
rect 38672 11354 38700 12718
rect 38660 11348 38712 11354
rect 38660 11290 38712 11296
rect 38764 11150 38792 13382
rect 38844 13330 38896 13336
rect 38844 13252 38896 13258
rect 38844 13194 38896 13200
rect 38856 12850 38884 13194
rect 38948 12918 38976 13806
rect 39026 13696 39082 13705
rect 39026 13631 39082 13640
rect 39040 13326 39068 13631
rect 39118 13560 39174 13569
rect 39118 13495 39174 13504
rect 39028 13320 39080 13326
rect 39028 13262 39080 13268
rect 39132 12918 39160 13495
rect 38936 12912 38988 12918
rect 39120 12912 39172 12918
rect 38988 12872 39068 12900
rect 38936 12854 38988 12860
rect 38844 12844 38896 12850
rect 38844 12786 38896 12792
rect 38856 11626 38884 12786
rect 38936 12708 38988 12714
rect 38936 12650 38988 12656
rect 38844 11620 38896 11626
rect 38844 11562 38896 11568
rect 38384 11144 38436 11150
rect 38384 11086 38436 11092
rect 38752 11144 38804 11150
rect 38752 11086 38804 11092
rect 38106 10976 38162 10985
rect 38106 10911 38162 10920
rect 38120 10062 38148 10911
rect 38200 10124 38252 10130
rect 38200 10066 38252 10072
rect 38108 10056 38160 10062
rect 38108 9998 38160 10004
rect 38108 8492 38160 8498
rect 38028 8452 38108 8480
rect 37556 8434 37608 8440
rect 38108 8434 38160 8440
rect 37476 7954 37504 8434
rect 37568 7954 37596 8434
rect 38212 8430 38240 10066
rect 38396 10062 38424 11086
rect 38384 10056 38436 10062
rect 38384 9998 38436 10004
rect 38948 9654 38976 12650
rect 39040 12374 39068 12872
rect 39120 12854 39172 12860
rect 39028 12368 39080 12374
rect 39028 12310 39080 12316
rect 39040 11014 39068 12310
rect 39120 11688 39172 11694
rect 39118 11656 39120 11665
rect 39172 11656 39174 11665
rect 39118 11591 39174 11600
rect 39224 11558 39252 14350
rect 39212 11552 39264 11558
rect 39212 11494 39264 11500
rect 39316 11354 39344 16458
rect 39408 16114 39436 17478
rect 39500 16250 39528 19722
rect 39592 19378 39620 20198
rect 39684 19514 39712 20878
rect 39776 20466 39804 20946
rect 39868 20942 39896 22374
rect 39948 21684 40000 21690
rect 39948 21626 40000 21632
rect 39856 20936 39908 20942
rect 39856 20878 39908 20884
rect 39764 20460 39816 20466
rect 39764 20402 39816 20408
rect 39672 19508 39724 19514
rect 39672 19450 39724 19456
rect 39580 19372 39632 19378
rect 39580 19314 39632 19320
rect 39672 19372 39724 19378
rect 39672 19314 39724 19320
rect 39592 18290 39620 19314
rect 39580 18284 39632 18290
rect 39580 18226 39632 18232
rect 39580 18148 39632 18154
rect 39580 18090 39632 18096
rect 39592 17678 39620 18090
rect 39684 17882 39712 19314
rect 39856 19168 39908 19174
rect 39856 19110 39908 19116
rect 39868 18970 39896 19110
rect 39856 18964 39908 18970
rect 39856 18906 39908 18912
rect 39764 18080 39816 18086
rect 39764 18022 39816 18028
rect 39672 17876 39724 17882
rect 39672 17818 39724 17824
rect 39580 17672 39632 17678
rect 39580 17614 39632 17620
rect 39684 16998 39712 17818
rect 39776 17270 39804 18022
rect 39960 17626 39988 21626
rect 40052 20602 40080 25230
rect 40144 24886 40172 25434
rect 40132 24880 40184 24886
rect 40132 24822 40184 24828
rect 40316 24200 40368 24206
rect 40316 24142 40368 24148
rect 40328 23322 40356 24142
rect 40224 23316 40276 23322
rect 40224 23258 40276 23264
rect 40316 23316 40368 23322
rect 40316 23258 40368 23264
rect 40040 20596 40092 20602
rect 40040 20538 40092 20544
rect 40132 19508 40184 19514
rect 40132 19450 40184 19456
rect 40040 18624 40092 18630
rect 40040 18566 40092 18572
rect 40052 18086 40080 18566
rect 40144 18306 40172 19450
rect 40236 18970 40264 23258
rect 40224 18964 40276 18970
rect 40224 18906 40276 18912
rect 40144 18278 40264 18306
rect 40132 18216 40184 18222
rect 40132 18158 40184 18164
rect 40040 18080 40092 18086
rect 40040 18022 40092 18028
rect 40144 17814 40172 18158
rect 40132 17808 40184 17814
rect 40132 17750 40184 17756
rect 39960 17598 40172 17626
rect 40040 17536 40092 17542
rect 40040 17478 40092 17484
rect 40052 17354 40080 17478
rect 39960 17338 40080 17354
rect 39948 17332 40080 17338
rect 40000 17326 40080 17332
rect 39948 17274 40000 17280
rect 39764 17264 39816 17270
rect 39764 17206 39816 17212
rect 40040 17196 40092 17202
rect 40040 17138 40092 17144
rect 39948 17128 40000 17134
rect 39948 17070 40000 17076
rect 39580 16992 39632 16998
rect 39580 16934 39632 16940
rect 39672 16992 39724 16998
rect 39672 16934 39724 16940
rect 39488 16244 39540 16250
rect 39488 16186 39540 16192
rect 39396 16108 39448 16114
rect 39396 16050 39448 16056
rect 39592 16046 39620 16934
rect 39960 16794 39988 17070
rect 39948 16788 40000 16794
rect 39948 16730 40000 16736
rect 39580 16040 39632 16046
rect 39580 15982 39632 15988
rect 39856 15972 39908 15978
rect 39856 15914 39908 15920
rect 39672 15904 39724 15910
rect 39672 15846 39724 15852
rect 39684 15706 39712 15846
rect 39868 15706 39896 15914
rect 39672 15700 39724 15706
rect 39672 15642 39724 15648
rect 39856 15700 39908 15706
rect 39856 15642 39908 15648
rect 39764 15564 39816 15570
rect 39764 15506 39816 15512
rect 39396 15020 39448 15026
rect 39396 14962 39448 14968
rect 39408 12850 39436 14962
rect 39776 14618 39804 15506
rect 39764 14612 39816 14618
rect 39764 14554 39816 14560
rect 39946 14512 40002 14521
rect 39946 14447 39948 14456
rect 40000 14447 40002 14456
rect 39948 14418 40000 14424
rect 40052 14414 40080 17138
rect 40144 16810 40172 17598
rect 40236 17202 40264 18278
rect 40316 18284 40368 18290
rect 40316 18226 40368 18232
rect 40224 17196 40276 17202
rect 40224 17138 40276 17144
rect 40144 16782 40264 16810
rect 40132 16720 40184 16726
rect 40132 16662 40184 16668
rect 40040 14408 40092 14414
rect 39762 14376 39818 14385
rect 39818 14334 39988 14362
rect 40040 14350 40092 14356
rect 39762 14311 39818 14320
rect 39488 13932 39540 13938
rect 39488 13874 39540 13880
rect 39500 13394 39528 13874
rect 39856 13524 39908 13530
rect 39856 13466 39908 13472
rect 39488 13388 39540 13394
rect 39488 13330 39540 13336
rect 39396 12844 39448 12850
rect 39396 12786 39448 12792
rect 39500 12714 39528 13330
rect 39868 12986 39896 13466
rect 39856 12980 39908 12986
rect 39856 12922 39908 12928
rect 39868 12866 39896 12922
rect 39684 12838 39896 12866
rect 39488 12708 39540 12714
rect 39488 12650 39540 12656
rect 39394 12336 39450 12345
rect 39394 12271 39450 12280
rect 39408 11830 39436 12271
rect 39396 11824 39448 11830
rect 39396 11766 39448 11772
rect 39120 11348 39172 11354
rect 39120 11290 39172 11296
rect 39304 11348 39356 11354
rect 39304 11290 39356 11296
rect 39132 11150 39160 11290
rect 39120 11144 39172 11150
rect 39120 11086 39172 11092
rect 39028 11008 39080 11014
rect 39028 10950 39080 10956
rect 39408 9674 39436 11766
rect 39684 11762 39712 12838
rect 39672 11756 39724 11762
rect 39672 11698 39724 11704
rect 39856 11756 39908 11762
rect 39856 11698 39908 11704
rect 39868 10266 39896 11698
rect 39960 11286 39988 14334
rect 40052 13530 40080 14350
rect 40040 13524 40092 13530
rect 40040 13466 40092 13472
rect 40144 11762 40172 16662
rect 40236 12345 40264 16782
rect 40328 14618 40356 18226
rect 40420 17746 40448 27911
rect 40500 26240 40552 26246
rect 40604 26228 40632 32370
rect 41064 31754 41092 32830
rect 41604 31816 41656 31822
rect 41604 31758 41656 31764
rect 40972 31726 41092 31754
rect 40684 29572 40736 29578
rect 40684 29514 40736 29520
rect 40696 28150 40724 29514
rect 40684 28144 40736 28150
rect 40684 28086 40736 28092
rect 40684 26308 40736 26314
rect 40736 26268 40908 26296
rect 40684 26250 40736 26256
rect 40552 26200 40632 26228
rect 40500 26182 40552 26188
rect 40512 25226 40540 26182
rect 40500 25220 40552 25226
rect 40500 25162 40552 25168
rect 40512 19854 40540 25162
rect 40592 23044 40644 23050
rect 40592 22986 40644 22992
rect 40500 19848 40552 19854
rect 40500 19790 40552 19796
rect 40500 18284 40552 18290
rect 40500 18226 40552 18232
rect 40408 17740 40460 17746
rect 40408 17682 40460 17688
rect 40512 17338 40540 18226
rect 40500 17332 40552 17338
rect 40500 17274 40552 17280
rect 40604 15706 40632 22986
rect 40684 22568 40736 22574
rect 40684 22510 40736 22516
rect 40696 16590 40724 22510
rect 40880 21690 40908 26268
rect 40868 21684 40920 21690
rect 40868 21626 40920 21632
rect 40776 20800 40828 20806
rect 40776 20742 40828 20748
rect 40788 20262 40816 20742
rect 40776 20256 40828 20262
rect 40776 20198 40828 20204
rect 40684 16584 40736 16590
rect 40684 16526 40736 16532
rect 40592 15700 40644 15706
rect 40592 15642 40644 15648
rect 40316 14612 40368 14618
rect 40316 14554 40368 14560
rect 40222 12336 40278 12345
rect 40222 12271 40278 12280
rect 40132 11756 40184 11762
rect 40132 11698 40184 11704
rect 40040 11688 40092 11694
rect 40038 11656 40040 11665
rect 40092 11656 40094 11665
rect 40038 11591 40094 11600
rect 39948 11280 40000 11286
rect 39948 11222 40000 11228
rect 40972 10810 41000 31726
rect 41052 31476 41104 31482
rect 41052 31418 41104 31424
rect 40960 10804 41012 10810
rect 40960 10746 41012 10752
rect 39856 10260 39908 10266
rect 39856 10202 39908 10208
rect 39408 9654 39620 9674
rect 38936 9648 38988 9654
rect 39408 9648 39632 9654
rect 39408 9646 39580 9648
rect 38936 9590 38988 9596
rect 39580 9590 39632 9596
rect 38948 8974 38976 9590
rect 38936 8968 38988 8974
rect 38936 8910 38988 8916
rect 38384 8492 38436 8498
rect 38384 8434 38436 8440
rect 38200 8424 38252 8430
rect 38200 8366 38252 8372
rect 38396 8090 38424 8434
rect 41064 8294 41092 31418
rect 41328 30728 41380 30734
rect 41328 30670 41380 30676
rect 41142 28248 41198 28257
rect 41142 28183 41198 28192
rect 41156 8362 41184 28183
rect 41236 20460 41288 20466
rect 41236 20402 41288 20408
rect 41248 11898 41276 20402
rect 41340 18426 41368 30670
rect 41512 29640 41564 29646
rect 41512 29582 41564 29588
rect 41420 21548 41472 21554
rect 41420 21490 41472 21496
rect 41432 21185 41460 21490
rect 41418 21176 41474 21185
rect 41418 21111 41474 21120
rect 41524 18426 41552 29582
rect 41328 18420 41380 18426
rect 41328 18362 41380 18368
rect 41512 18420 41564 18426
rect 41512 18362 41564 18368
rect 41616 17542 41644 31758
rect 41696 27464 41748 27470
rect 41696 27406 41748 27412
rect 41708 18222 41736 27406
rect 41878 23080 41934 23089
rect 41878 23015 41934 23024
rect 41696 18216 41748 18222
rect 41696 18158 41748 18164
rect 41604 17536 41656 17542
rect 41604 17478 41656 17484
rect 41892 12434 41920 23015
rect 41616 12406 41920 12434
rect 41236 11892 41288 11898
rect 41236 11834 41288 11840
rect 41616 9625 41644 12406
rect 41602 9616 41658 9625
rect 41602 9551 41658 9560
rect 41144 8356 41196 8362
rect 41144 8298 41196 8304
rect 41052 8288 41104 8294
rect 41052 8230 41104 8236
rect 38384 8084 38436 8090
rect 38384 8026 38436 8032
rect 37464 7948 37516 7954
rect 37464 7890 37516 7896
rect 37556 7948 37608 7954
rect 37556 7890 37608 7896
rect 40776 7744 40828 7750
rect 40776 7686 40828 7692
rect 36912 7540 36964 7546
rect 36912 7482 36964 7488
rect 36544 7200 36596 7206
rect 36544 7142 36596 7148
rect 36452 6996 36504 7002
rect 36452 6938 36504 6944
rect 36556 6934 36584 7142
rect 36544 6928 36596 6934
rect 36544 6870 36596 6876
rect 36176 5908 36228 5914
rect 36176 5850 36228 5856
rect 35716 5704 35768 5710
rect 35714 5672 35716 5681
rect 36912 5704 36964 5710
rect 35768 5672 35770 5681
rect 36912 5646 36964 5652
rect 35714 5607 35770 5616
rect 35348 5568 35400 5574
rect 35348 5510 35400 5516
rect 35990 5536 36046 5545
rect 35360 5302 35388 5510
rect 35990 5471 36046 5480
rect 35348 5296 35400 5302
rect 35348 5238 35400 5244
rect 34796 5160 34848 5166
rect 34796 5102 34848 5108
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 36004 4622 36032 5471
rect 36924 5370 36952 5646
rect 36912 5364 36964 5370
rect 36912 5306 36964 5312
rect 36176 5160 36228 5166
rect 36176 5102 36228 5108
rect 35992 4616 36044 4622
rect 35992 4558 36044 4564
rect 36188 4486 36216 5102
rect 34060 4480 34112 4486
rect 34060 4422 34112 4428
rect 36176 4480 36228 4486
rect 36176 4422 36228 4428
rect 30564 4276 30616 4282
rect 30564 4218 30616 4224
rect 30932 4276 30984 4282
rect 30932 4218 30984 4224
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 36728 3460 36780 3466
rect 36728 3402 36780 3408
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 29828 2508 29880 2514
rect 29828 2450 29880 2456
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 29012 800 29040 2382
rect 33140 2304 33192 2310
rect 33140 2246 33192 2252
rect 33152 1442 33180 2246
rect 32876 1414 33180 1442
rect 32876 800 32904 1414
rect 36740 800 36768 3402
rect 40788 2650 40816 7686
rect 40960 6384 41012 6390
rect 40960 6326 41012 6332
rect 40972 5914 41000 6326
rect 40960 5908 41012 5914
rect 40960 5850 41012 5856
rect 41328 5568 41380 5574
rect 41326 5536 41328 5545
rect 41380 5536 41382 5545
rect 41326 5471 41382 5480
rect 40776 2644 40828 2650
rect 40776 2586 40828 2592
rect 40684 2372 40736 2378
rect 40684 2314 40736 2320
rect 40696 1170 40724 2314
rect 40604 1142 40724 1170
rect 40604 800 40632 1142
rect 18 0 74 800
rect 3238 0 3294 800
rect 7102 0 7158 800
rect 10966 0 11022 800
rect 14186 0 14242 800
rect 18050 0 18106 800
rect 21914 0 21970 800
rect 25778 0 25834 800
rect 28998 0 29054 800
rect 32862 0 32918 800
rect 36726 0 36782 800
rect 40590 0 40646 800
<< via2 >>
rect 3422 42880 3478 42936
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 3790 38800 3846 38856
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 1030 34740 1086 34776
rect 1030 34720 1032 34740
rect 1032 34720 1084 34740
rect 1084 34720 1086 34740
rect 1858 34604 1914 34640
rect 1858 34584 1860 34604
rect 1860 34584 1912 34604
rect 1912 34584 1914 34604
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 2778 30640 2834 30696
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 3422 29164 3478 29200
rect 3422 29144 3424 29164
rect 3424 29144 3476 29164
rect 3476 29144 3478 29164
rect 3606 23160 3662 23216
rect 3330 19080 3386 19136
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4526 29688 4582 29744
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4066 27240 4122 27296
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 5170 28872 5226 28928
rect 7102 29588 7104 29608
rect 7104 29588 7156 29608
rect 7156 29588 7158 29608
rect 7102 29552 7158 29588
rect 6274 28872 6330 28928
rect 5078 24812 5134 24848
rect 5078 24792 5080 24812
rect 5080 24792 5132 24812
rect 5132 24792 5134 24812
rect 4986 24656 5042 24712
rect 5262 24692 5264 24712
rect 5264 24692 5316 24712
rect 5316 24692 5318 24712
rect 5262 24656 5318 24692
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 5078 22888 5134 22944
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 1582 15136 1638 15192
rect 938 11600 994 11656
rect 938 7520 994 7576
rect 5538 24812 5594 24848
rect 5538 24792 5540 24812
rect 5540 24792 5592 24812
rect 5592 24792 5594 24812
rect 5906 24692 5908 24712
rect 5908 24692 5960 24712
rect 5960 24692 5962 24712
rect 5906 24656 5962 24692
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4710 19372 4766 19408
rect 4710 19352 4712 19372
rect 4712 19352 4764 19372
rect 4764 19352 4766 19372
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4894 12688 4950 12744
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 5354 15136 5410 15192
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 7194 29008 7250 29064
rect 6458 24148 6460 24168
rect 6460 24148 6512 24168
rect 6512 24148 6514 24168
rect 6458 24112 6514 24148
rect 7746 29588 7748 29608
rect 7748 29588 7800 29608
rect 7800 29588 7802 29608
rect 7746 29552 7802 29588
rect 6826 20168 6882 20224
rect 7286 19352 7342 19408
rect 5998 12688 6054 12744
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 7378 12960 7434 13016
rect 7930 26832 7986 26888
rect 8298 29824 8354 29880
rect 8390 27512 8446 27568
rect 8206 24812 8262 24848
rect 8206 24792 8208 24812
rect 8208 24792 8260 24812
rect 8260 24792 8262 24812
rect 7746 19352 7802 19408
rect 8574 27240 8630 27296
rect 8850 29824 8906 29880
rect 8758 27512 8814 27568
rect 8850 27376 8906 27432
rect 9034 29044 9036 29064
rect 9036 29044 9088 29064
rect 9088 29044 9090 29064
rect 9034 29008 9090 29044
rect 9862 40180 9918 40216
rect 9862 40160 9864 40180
rect 9864 40160 9916 40180
rect 9916 40160 9918 40180
rect 10598 40180 10654 40216
rect 10598 40160 10600 40180
rect 10600 40160 10652 40180
rect 10652 40160 10654 40180
rect 10046 40044 10102 40080
rect 10046 40024 10048 40044
rect 10048 40024 10100 40044
rect 10100 40024 10102 40044
rect 10782 40044 10838 40080
rect 10782 40024 10784 40044
rect 10784 40024 10836 40044
rect 10836 40024 10838 40044
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 9862 29688 9918 29744
rect 10138 29552 10194 29608
rect 9954 29416 10010 29472
rect 10322 29144 10378 29200
rect 9218 27512 9274 27568
rect 9126 26696 9182 26752
rect 9494 26968 9550 27024
rect 9126 25744 9182 25800
rect 7838 12960 7894 13016
rect 8022 12824 8078 12880
rect 9218 24928 9274 24984
rect 9218 24676 9274 24712
rect 9218 24656 9220 24676
rect 9220 24656 9272 24676
rect 9272 24656 9274 24676
rect 9770 27124 9826 27160
rect 9770 27104 9772 27124
rect 9772 27104 9824 27124
rect 9824 27104 9826 27124
rect 10046 26988 10102 27024
rect 10046 26968 10048 26988
rect 10048 26968 10100 26988
rect 10100 26968 10102 26988
rect 9494 24112 9550 24168
rect 10322 27240 10378 27296
rect 10322 26288 10378 26344
rect 10046 21972 10048 21992
rect 10048 21972 10100 21992
rect 10100 21972 10102 21992
rect 10046 21936 10102 21972
rect 9126 19760 9182 19816
rect 9034 16224 9090 16280
rect 9586 16244 9642 16280
rect 9586 16224 9588 16244
rect 9588 16224 9640 16244
rect 9640 16224 9642 16244
rect 9218 12960 9274 13016
rect 9126 12824 9182 12880
rect 10138 20168 10194 20224
rect 10690 27512 10746 27568
rect 10690 25200 10746 25256
rect 11610 34992 11666 35048
rect 11610 32852 11612 32872
rect 11612 32852 11664 32872
rect 11664 32852 11666 32872
rect 11610 32816 11666 32852
rect 10966 28464 11022 28520
rect 10966 28056 11022 28112
rect 11978 30540 11980 30560
rect 11980 30540 12032 30560
rect 12032 30540 12034 30560
rect 11978 30504 12034 30540
rect 11610 30368 11666 30424
rect 10230 19352 10286 19408
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 938 3440 994 3496
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 10046 12844 10102 12880
rect 10046 12824 10048 12844
rect 10048 12824 10100 12844
rect 10100 12824 10102 12844
rect 10506 19352 10562 19408
rect 10598 13232 10654 13288
rect 11150 19488 11206 19544
rect 11426 26324 11428 26344
rect 11428 26324 11480 26344
rect 11480 26324 11482 26344
rect 11426 26288 11482 26324
rect 11610 24928 11666 24984
rect 11978 28872 12034 28928
rect 12162 28500 12164 28520
rect 12164 28500 12216 28520
rect 12216 28500 12218 28520
rect 12162 28464 12218 28500
rect 12070 27004 12072 27024
rect 12072 27004 12124 27024
rect 12124 27004 12126 27024
rect 12070 26968 12126 27004
rect 12714 30368 12770 30424
rect 12530 29688 12586 29744
rect 13266 29416 13322 29472
rect 12622 28464 12678 28520
rect 13450 29008 13506 29064
rect 12530 27124 12586 27160
rect 12530 27104 12532 27124
rect 12532 27104 12584 27124
rect 12584 27104 12586 27124
rect 11702 23432 11758 23488
rect 11150 16496 11206 16552
rect 12070 22636 12126 22672
rect 12070 22616 12072 22636
rect 12072 22616 12124 22636
rect 12124 22616 12126 22636
rect 12530 24284 12532 24304
rect 12532 24284 12584 24304
rect 12584 24284 12586 24304
rect 12530 24248 12586 24284
rect 12530 23432 12586 23488
rect 11794 20576 11850 20632
rect 11058 12008 11114 12064
rect 11610 12708 11666 12744
rect 11610 12688 11612 12708
rect 11612 12688 11664 12708
rect 11664 12688 11666 12708
rect 11242 9036 11298 9072
rect 11242 9016 11244 9036
rect 11244 9016 11296 9036
rect 11296 9016 11298 9036
rect 11610 9424 11666 9480
rect 11518 8744 11574 8800
rect 12806 24384 12862 24440
rect 13174 26988 13230 27024
rect 13174 26968 13176 26988
rect 13176 26968 13228 26988
rect 13228 26968 13230 26988
rect 15106 35536 15162 35592
rect 14002 29416 14058 29472
rect 13726 26732 13728 26752
rect 13728 26732 13780 26752
rect 13780 26732 13782 26752
rect 13726 26696 13782 26732
rect 12990 24520 13046 24576
rect 12714 19352 12770 19408
rect 12898 21936 12954 21992
rect 12070 13504 12126 13560
rect 11794 12960 11850 13016
rect 11978 10920 12034 10976
rect 12622 12824 12678 12880
rect 12530 12280 12586 12336
rect 13818 22616 13874 22672
rect 14186 28076 14242 28112
rect 14186 28056 14188 28076
rect 14188 28056 14240 28076
rect 14240 28056 14242 28076
rect 16486 35028 16488 35048
rect 16488 35028 16540 35048
rect 16540 35028 16542 35048
rect 16486 34992 16542 35028
rect 14462 24656 14518 24712
rect 14462 24404 14518 24440
rect 14186 24248 14242 24304
rect 13818 19760 13874 19816
rect 13542 13676 13544 13696
rect 13544 13676 13596 13696
rect 13596 13676 13598 13696
rect 13542 13640 13598 13676
rect 13450 10784 13506 10840
rect 13082 10648 13138 10704
rect 12530 9424 12586 9480
rect 11978 9016 12034 9072
rect 11518 8492 11574 8528
rect 11518 8472 11520 8492
rect 11520 8472 11572 8492
rect 11572 8472 11574 8492
rect 11978 8744 12034 8800
rect 12714 7248 12770 7304
rect 12622 6840 12678 6896
rect 14462 24384 14464 24404
rect 14464 24384 14516 24404
rect 14516 24384 14518 24404
rect 14830 28464 14886 28520
rect 14922 27124 14978 27160
rect 14922 27104 14924 27124
rect 14924 27104 14976 27124
rect 14976 27104 14978 27124
rect 14278 21956 14334 21992
rect 14278 21936 14280 21956
rect 14280 21936 14332 21956
rect 14332 21936 14334 21956
rect 15750 29144 15806 29200
rect 15934 29044 15936 29064
rect 15936 29044 15988 29064
rect 15988 29044 15990 29064
rect 15934 29008 15990 29044
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 16394 30912 16450 30968
rect 15382 26988 15438 27024
rect 15934 27124 15990 27160
rect 15934 27104 15936 27124
rect 15936 27104 15988 27124
rect 15988 27104 15990 27124
rect 15382 26968 15384 26988
rect 15384 26968 15436 26988
rect 15436 26968 15438 26988
rect 14738 20032 14794 20088
rect 13910 12144 13966 12200
rect 14462 12280 14518 12336
rect 13634 6740 13636 6760
rect 13636 6740 13688 6760
rect 13688 6740 13690 6760
rect 13634 6704 13690 6740
rect 15842 24012 15844 24032
rect 15844 24012 15896 24032
rect 15896 24012 15898 24032
rect 15842 23976 15898 24012
rect 16486 29164 16542 29200
rect 16486 29144 16488 29164
rect 16488 29144 16540 29164
rect 16540 29144 16542 29164
rect 16946 30640 17002 30696
rect 16302 27104 16358 27160
rect 16946 28056 17002 28112
rect 16486 27512 16542 27568
rect 16670 26832 16726 26888
rect 16302 26288 16358 26344
rect 16026 22888 16082 22944
rect 16486 24656 16542 24712
rect 16486 24148 16488 24168
rect 16488 24148 16540 24168
rect 16540 24148 16542 24168
rect 16486 24112 16542 24148
rect 17682 30504 17738 30560
rect 16394 22888 16450 22944
rect 16210 20868 16266 20904
rect 16210 20848 16212 20868
rect 16212 20848 16264 20868
rect 16264 20848 16266 20868
rect 16210 20712 16266 20768
rect 16118 19216 16174 19272
rect 15290 15444 15292 15464
rect 15292 15444 15344 15464
rect 15344 15444 15346 15464
rect 15290 15408 15346 15444
rect 15750 18128 15806 18184
rect 15658 14728 15714 14784
rect 14646 12144 14702 12200
rect 15106 11756 15162 11792
rect 15106 11736 15108 11756
rect 15108 11736 15160 11756
rect 15160 11736 15162 11756
rect 14646 8472 14702 8528
rect 15474 12960 15530 13016
rect 16118 17720 16174 17776
rect 15750 13504 15806 13560
rect 14462 7248 14518 7304
rect 15014 6860 15070 6896
rect 15014 6840 15016 6860
rect 15016 6840 15068 6860
rect 15068 6840 15070 6860
rect 15566 12844 15622 12880
rect 15566 12824 15568 12844
rect 15568 12824 15620 12844
rect 15620 12824 15622 12844
rect 16118 13096 16174 13152
rect 16394 13524 16450 13560
rect 16394 13504 16396 13524
rect 16396 13504 16448 13524
rect 16448 13504 16450 13524
rect 17406 23976 17462 24032
rect 17406 23160 17462 23216
rect 16854 20576 16910 20632
rect 16762 13776 16818 13832
rect 16670 13232 16726 13288
rect 17406 21956 17462 21992
rect 17406 21936 17408 21956
rect 17408 21936 17460 21956
rect 17460 21936 17462 21956
rect 17314 21120 17370 21176
rect 17130 20848 17186 20904
rect 17498 20168 17554 20224
rect 18786 35128 18842 35184
rect 17958 29688 18014 29744
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19614 34040 19670 34096
rect 20074 33904 20130 33960
rect 19982 33768 20038 33824
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 20258 34584 20314 34640
rect 20166 32816 20222 32872
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19982 32272 20038 32328
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 18694 29144 18750 29200
rect 18326 28600 18382 28656
rect 17958 23160 18014 23216
rect 18418 23976 18474 24032
rect 17498 19352 17554 19408
rect 17590 17448 17646 17504
rect 17222 17176 17278 17232
rect 18234 19760 18290 19816
rect 17774 17856 17830 17912
rect 17130 15408 17186 15464
rect 16854 10784 16910 10840
rect 16946 9444 17002 9480
rect 17590 13640 17646 13696
rect 17682 12960 17738 13016
rect 18234 17584 18290 17640
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19890 29688 19946 29744
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19798 28756 19854 28792
rect 19798 28736 19800 28756
rect 19800 28736 19852 28756
rect 19852 28736 19854 28756
rect 19798 28484 19854 28520
rect 19798 28464 19800 28484
rect 19800 28464 19852 28484
rect 19852 28464 19854 28484
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19982 27648 20038 27704
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 20534 34060 20590 34096
rect 20534 34040 20536 34060
rect 20536 34040 20588 34060
rect 20588 34040 20590 34060
rect 20534 33768 20590 33824
rect 22006 37304 22062 37360
rect 21454 34060 21510 34096
rect 21454 34040 21456 34060
rect 21456 34040 21508 34060
rect 21508 34040 21510 34060
rect 21362 33940 21364 33960
rect 21364 33940 21416 33960
rect 21416 33940 21418 33960
rect 21362 33904 21418 33940
rect 21362 32408 21418 32464
rect 20442 30116 20498 30152
rect 20442 30096 20444 30116
rect 20444 30096 20496 30116
rect 20496 30096 20498 30116
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 18510 17620 18512 17640
rect 18512 17620 18564 17640
rect 18564 17620 18566 17640
rect 18510 17584 18566 17620
rect 18418 13096 18474 13152
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19706 24404 19762 24440
rect 19706 24384 19708 24404
rect 19708 24384 19760 24404
rect 19760 24384 19762 24404
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19522 21392 19578 21448
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 20258 23568 20314 23624
rect 19706 20304 19762 20360
rect 19614 20032 19670 20088
rect 19246 18944 19302 19000
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 18970 17856 19026 17912
rect 19338 17720 19394 17776
rect 19062 17584 19118 17640
rect 18878 17448 18934 17504
rect 19246 16108 19302 16144
rect 19246 16088 19248 16108
rect 19248 16088 19300 16108
rect 19300 16088 19302 16108
rect 19154 15408 19210 15464
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19890 16768 19946 16824
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19430 14864 19486 14920
rect 20074 19080 20130 19136
rect 20166 18400 20222 18456
rect 20166 15156 20222 15192
rect 20166 15136 20168 15156
rect 20168 15136 20220 15156
rect 20220 15136 20222 15156
rect 19890 14320 19946 14376
rect 16946 9424 16948 9444
rect 16948 9424 17000 9444
rect 17000 9424 17002 9444
rect 15842 7284 15844 7304
rect 15844 7284 15896 7304
rect 15896 7284 15898 7304
rect 15842 7248 15898 7284
rect 15382 6704 15438 6760
rect 17130 5616 17186 5672
rect 16946 5480 17002 5536
rect 18418 9152 18474 9208
rect 18418 8472 18474 8528
rect 18786 12688 18842 12744
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19522 13912 19578 13968
rect 19798 13932 19854 13968
rect 19798 13912 19800 13932
rect 19800 13912 19852 13932
rect 19852 13912 19854 13932
rect 19062 10684 19064 10704
rect 19064 10684 19116 10704
rect 19116 10684 19118 10704
rect 19062 10648 19118 10684
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19430 9968 19486 10024
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19062 8064 19118 8120
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 20718 28736 20774 28792
rect 21086 30776 21142 30832
rect 21178 30132 21180 30152
rect 21180 30132 21232 30152
rect 21232 30132 21234 30152
rect 21178 30096 21234 30132
rect 20994 28600 21050 28656
rect 20994 28500 20996 28520
rect 20996 28500 21048 28520
rect 21048 28500 21050 28520
rect 20994 28464 21050 28500
rect 20810 27648 20866 27704
rect 20994 25880 21050 25936
rect 20718 23604 20720 23624
rect 20720 23604 20772 23624
rect 20772 23604 20774 23624
rect 20718 23568 20774 23604
rect 20626 21972 20628 21992
rect 20628 21972 20680 21992
rect 20680 21972 20682 21992
rect 20626 21936 20682 21972
rect 20718 21120 20774 21176
rect 20994 22888 21050 22944
rect 21178 25064 21234 25120
rect 21730 31084 21732 31104
rect 21732 31084 21784 31104
rect 21784 31084 21786 31104
rect 21730 31048 21786 31084
rect 22098 31728 22154 31784
rect 22558 34720 22614 34776
rect 22834 34992 22890 35048
rect 22834 33904 22890 33960
rect 22558 31728 22614 31784
rect 22282 31184 22338 31240
rect 22190 30776 22246 30832
rect 21546 28328 21602 28384
rect 21454 28192 21510 28248
rect 21454 27648 21510 27704
rect 21546 26324 21548 26344
rect 21548 26324 21600 26344
rect 21600 26324 21602 26344
rect 21546 26288 21602 26324
rect 21546 25644 21548 25664
rect 21548 25644 21600 25664
rect 21600 25644 21602 25664
rect 21546 25608 21602 25644
rect 21546 25472 21602 25528
rect 21086 22208 21142 22264
rect 21086 21936 21142 21992
rect 21270 23044 21326 23080
rect 21270 23024 21272 23044
rect 21272 23024 21324 23044
rect 21324 23024 21326 23044
rect 21270 22636 21326 22672
rect 21270 22616 21272 22636
rect 21272 22616 21324 22636
rect 21324 22616 21326 22636
rect 22006 29280 22062 29336
rect 22006 29180 22008 29200
rect 22008 29180 22060 29200
rect 22060 29180 22062 29200
rect 22006 29144 22062 29180
rect 21822 28872 21878 28928
rect 21730 28192 21786 28248
rect 21730 26696 21786 26752
rect 21914 27240 21970 27296
rect 22466 29452 22468 29472
rect 22468 29452 22520 29472
rect 22520 29452 22522 29472
rect 22466 29416 22522 29452
rect 22098 28620 22154 28656
rect 22098 28600 22100 28620
rect 22100 28600 22152 28620
rect 22152 28600 22154 28620
rect 22558 28736 22614 28792
rect 22190 27920 22246 27976
rect 21822 25472 21878 25528
rect 22190 26832 22246 26888
rect 22006 25064 22062 25120
rect 21362 22208 21418 22264
rect 21638 22228 21694 22264
rect 21638 22208 21640 22228
rect 21640 22208 21692 22228
rect 21692 22208 21694 22228
rect 20350 14456 20406 14512
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 15014 3984 15070 4040
rect 14738 3576 14794 3632
rect 20994 18672 21050 18728
rect 21086 18264 21142 18320
rect 20718 17992 20774 18048
rect 20718 16904 20774 16960
rect 20902 15036 20904 15056
rect 20904 15036 20956 15056
rect 20956 15036 20958 15056
rect 20902 15000 20958 15036
rect 21730 21936 21786 21992
rect 21454 21664 21510 21720
rect 22190 23316 22246 23352
rect 22190 23296 22192 23316
rect 22192 23296 22244 23316
rect 22244 23296 22246 23316
rect 22190 22752 22246 22808
rect 22190 22616 22246 22672
rect 22466 23704 22522 23760
rect 22282 22228 22338 22264
rect 22282 22208 22284 22228
rect 22284 22208 22336 22228
rect 22336 22208 22338 22228
rect 22466 22344 22522 22400
rect 22558 22208 22614 22264
rect 22466 21972 22468 21992
rect 22468 21972 22520 21992
rect 22520 21972 22522 21992
rect 22466 21936 22522 21972
rect 22374 21800 22430 21856
rect 22190 21256 22246 21312
rect 22006 20712 22062 20768
rect 22374 20304 22430 20360
rect 22006 18828 22062 18864
rect 22006 18808 22008 18828
rect 22008 18808 22060 18828
rect 22060 18808 22062 18828
rect 21914 17040 21970 17096
rect 21270 15000 21326 15056
rect 21638 15952 21694 16008
rect 22190 15680 22246 15736
rect 21914 15000 21970 15056
rect 21638 14884 21694 14920
rect 21638 14864 21640 14884
rect 21640 14864 21692 14884
rect 21692 14864 21694 14884
rect 21638 10920 21694 10976
rect 24122 35264 24178 35320
rect 23938 35128 23994 35184
rect 23294 31592 23350 31648
rect 23018 28500 23020 28520
rect 23020 28500 23072 28520
rect 23072 28500 23074 28520
rect 23018 28464 23074 28500
rect 23110 26832 23166 26888
rect 22742 24148 22744 24168
rect 22744 24148 22796 24168
rect 22796 24148 22798 24168
rect 22742 24112 22798 24148
rect 22834 23704 22890 23760
rect 22926 22888 22982 22944
rect 22926 22772 22982 22808
rect 22926 22752 22928 22772
rect 22928 22752 22980 22772
rect 22980 22752 22982 22772
rect 23846 31864 23902 31920
rect 24306 31456 24362 31512
rect 24030 31320 24086 31376
rect 23570 28464 23626 28520
rect 23754 28500 23756 28520
rect 23756 28500 23808 28520
rect 23808 28500 23810 28520
rect 23754 28464 23810 28500
rect 23386 26288 23442 26344
rect 23294 24268 23350 24304
rect 23294 24248 23296 24268
rect 23296 24248 23348 24268
rect 23348 24248 23350 24268
rect 23202 22888 23258 22944
rect 23202 22108 23204 22128
rect 23204 22108 23256 22128
rect 23256 22108 23258 22128
rect 23202 22072 23258 22108
rect 23938 29144 23994 29200
rect 23662 26324 23664 26344
rect 23664 26324 23716 26344
rect 23716 26324 23718 26344
rect 23662 26288 23718 26324
rect 23478 23588 23534 23624
rect 23478 23568 23480 23588
rect 23480 23568 23532 23588
rect 23532 23568 23534 23588
rect 24030 27920 24086 27976
rect 23662 24384 23718 24440
rect 23846 23840 23902 23896
rect 23662 23568 23718 23624
rect 23570 23432 23626 23488
rect 23662 23160 23718 23216
rect 23386 22752 23442 22808
rect 23570 22344 23626 22400
rect 23202 21020 23204 21040
rect 23204 21020 23256 21040
rect 23256 21020 23258 21040
rect 23202 20984 23258 21020
rect 23110 20884 23112 20904
rect 23112 20884 23164 20904
rect 23164 20884 23166 20904
rect 23110 20848 23166 20884
rect 23478 21800 23534 21856
rect 22926 19488 22982 19544
rect 22650 17196 22706 17232
rect 22650 17176 22652 17196
rect 22652 17176 22704 17196
rect 22704 17176 22706 17196
rect 22650 14592 22706 14648
rect 22742 14456 22798 14512
rect 23018 17448 23074 17504
rect 23294 20576 23350 20632
rect 23202 19624 23258 19680
rect 24582 35164 24584 35184
rect 24584 35164 24636 35184
rect 24636 35164 24638 35184
rect 24582 35128 24638 35164
rect 24582 34584 24638 34640
rect 25042 35808 25098 35864
rect 24950 35264 25006 35320
rect 34518 42220 34574 42256
rect 34518 42200 34520 42220
rect 34520 42200 34572 42220
rect 34572 42200 34574 42220
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 31298 41384 31354 41440
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 25410 35028 25412 35048
rect 25412 35028 25464 35048
rect 25464 35028 25466 35048
rect 24766 33768 24822 33824
rect 24858 31728 24914 31784
rect 25410 34992 25466 35028
rect 26238 35828 26294 35864
rect 26238 35808 26240 35828
rect 26240 35808 26292 35828
rect 26292 35808 26294 35828
rect 25410 33904 25466 33960
rect 24398 30096 24454 30152
rect 24766 31220 24768 31240
rect 24768 31220 24820 31240
rect 24820 31220 24822 31240
rect 24766 31184 24822 31220
rect 24490 29044 24492 29064
rect 24492 29044 24544 29064
rect 24544 29044 24546 29064
rect 24490 29008 24546 29044
rect 24490 28872 24546 28928
rect 24306 28464 24362 28520
rect 23478 19216 23534 19272
rect 23570 17856 23626 17912
rect 23754 16768 23810 16824
rect 23570 16632 23626 16688
rect 23938 17448 23994 17504
rect 24582 26732 24584 26752
rect 24584 26732 24636 26752
rect 24636 26732 24638 26752
rect 24582 26696 24638 26732
rect 24950 31048 25006 31104
rect 25042 30504 25098 30560
rect 24766 27512 24822 27568
rect 25226 29008 25282 29064
rect 26330 35536 26386 35592
rect 26146 34856 26202 34912
rect 26698 35128 26754 35184
rect 26606 34720 26662 34776
rect 26422 33088 26478 33144
rect 25410 29280 25466 29336
rect 25318 28872 25374 28928
rect 25318 27648 25374 27704
rect 25042 26424 25098 26480
rect 25502 28600 25558 28656
rect 25134 24928 25190 24984
rect 24674 23704 24730 23760
rect 24582 23568 24638 23624
rect 24398 21972 24400 21992
rect 24400 21972 24452 21992
rect 24452 21972 24454 21992
rect 24398 21936 24454 21972
rect 24398 21428 24400 21448
rect 24400 21428 24452 21448
rect 24452 21428 24454 21448
rect 24398 21392 24454 21428
rect 23386 12824 23442 12880
rect 24858 22616 24914 22672
rect 25042 23976 25098 24032
rect 25042 23180 25098 23216
rect 25042 23160 25044 23180
rect 25044 23160 25096 23180
rect 25096 23160 25098 23180
rect 25042 21800 25098 21856
rect 25594 26308 25650 26344
rect 25594 26288 25596 26308
rect 25596 26288 25648 26308
rect 25648 26288 25650 26308
rect 25870 30368 25926 30424
rect 26146 32272 26202 32328
rect 25870 29416 25926 29472
rect 26330 31900 26332 31920
rect 26332 31900 26384 31920
rect 26384 31900 26386 31920
rect 26330 31864 26386 31900
rect 27066 33768 27122 33824
rect 26698 33224 26754 33280
rect 25962 28600 26018 28656
rect 26146 28328 26202 28384
rect 27618 34740 27674 34776
rect 27618 34720 27620 34740
rect 27620 34720 27672 34740
rect 27672 34720 27674 34740
rect 26974 32272 27030 32328
rect 27342 31184 27398 31240
rect 26698 28328 26754 28384
rect 26606 27920 26662 27976
rect 26238 24248 26294 24304
rect 25962 23976 26018 24032
rect 25410 22480 25466 22536
rect 24950 20984 25006 21040
rect 24766 20168 24822 20224
rect 24582 19352 24638 19408
rect 24766 18400 24822 18456
rect 24582 15136 24638 15192
rect 23478 12300 23534 12336
rect 23478 12280 23480 12300
rect 23480 12280 23532 12300
rect 23532 12280 23534 12300
rect 22742 11736 22798 11792
rect 24306 13640 24362 13696
rect 24398 12416 24454 12472
rect 25134 18944 25190 19000
rect 25594 19508 25650 19544
rect 25594 19488 25596 19508
rect 25596 19488 25648 19508
rect 25648 19488 25650 19508
rect 26054 23568 26110 23624
rect 26054 22616 26110 22672
rect 26698 23432 26754 23488
rect 25778 20712 25834 20768
rect 25962 21972 25964 21992
rect 25964 21972 26016 21992
rect 26016 21972 26018 21992
rect 25962 21936 26018 21972
rect 25962 21800 26018 21856
rect 26882 28192 26938 28248
rect 26882 27648 26938 27704
rect 27158 28500 27160 28520
rect 27160 28500 27212 28520
rect 27212 28500 27214 28520
rect 27158 28464 27214 28500
rect 27434 28736 27490 28792
rect 26974 25880 27030 25936
rect 26974 24148 26976 24168
rect 26976 24148 27028 24168
rect 27028 24148 27030 24168
rect 26974 24112 27030 24148
rect 25502 14356 25504 14376
rect 25504 14356 25556 14376
rect 25556 14356 25558 14376
rect 25502 14320 25558 14356
rect 25226 14048 25282 14104
rect 26238 19352 26294 19408
rect 25870 17992 25926 18048
rect 25870 16632 25926 16688
rect 26330 18944 26386 19000
rect 26330 17076 26332 17096
rect 26332 17076 26384 17096
rect 26384 17076 26386 17096
rect 26330 17040 26386 17076
rect 26054 16904 26110 16960
rect 26330 16632 26386 16688
rect 26146 16496 26202 16552
rect 25594 12280 25650 12336
rect 25778 15136 25834 15192
rect 26238 15272 26294 15328
rect 26606 21392 26662 21448
rect 26606 19236 26662 19272
rect 26606 19216 26608 19236
rect 26608 19216 26660 19236
rect 26660 19216 26662 19236
rect 26606 18672 26662 18728
rect 26514 17856 26570 17912
rect 26698 17332 26754 17368
rect 26698 17312 26700 17332
rect 26700 17312 26752 17332
rect 26752 17312 26754 17332
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 28262 36116 28264 36136
rect 28264 36116 28316 36136
rect 28316 36116 28318 36136
rect 28262 36080 28318 36116
rect 27986 32544 28042 32600
rect 27894 31628 27896 31648
rect 27896 31628 27948 31648
rect 27948 31628 27950 31648
rect 27894 31592 27950 31628
rect 27710 28192 27766 28248
rect 27894 29280 27950 29336
rect 27986 28192 28042 28248
rect 28170 31456 28226 31512
rect 28262 30232 28318 30288
rect 28170 29416 28226 29472
rect 28262 29008 28318 29064
rect 28630 35944 28686 36000
rect 28446 31320 28502 31376
rect 28814 33088 28870 33144
rect 28814 32680 28870 32736
rect 28354 28736 28410 28792
rect 30010 34720 30066 34776
rect 29918 34584 29974 34640
rect 29734 34468 29790 34504
rect 29734 34448 29736 34468
rect 29736 34448 29788 34468
rect 29788 34448 29790 34468
rect 29550 34176 29606 34232
rect 28906 30504 28962 30560
rect 28814 29280 28870 29336
rect 28814 29008 28870 29064
rect 28630 28872 28686 28928
rect 28446 28600 28502 28656
rect 28630 28600 28686 28656
rect 28262 28192 28318 28248
rect 28538 28056 28594 28112
rect 27986 27512 28042 27568
rect 28170 27648 28226 27704
rect 27986 26188 27988 26208
rect 27988 26188 28040 26208
rect 28040 26188 28042 26208
rect 27986 26152 28042 26188
rect 26882 19080 26938 19136
rect 26882 15308 26884 15328
rect 26884 15308 26936 15328
rect 26936 15308 26938 15328
rect 26882 15272 26938 15308
rect 26882 15136 26938 15192
rect 26882 14184 26938 14240
rect 28814 28192 28870 28248
rect 29182 28500 29184 28520
rect 29184 28500 29236 28520
rect 29236 28500 29238 28520
rect 29182 28464 29238 28500
rect 29090 28056 29146 28112
rect 29458 31084 29460 31104
rect 29460 31084 29512 31104
rect 29512 31084 29514 31104
rect 29458 31048 29514 31084
rect 29458 30368 29514 30424
rect 29366 29280 29422 29336
rect 29458 28192 29514 28248
rect 28998 27648 29054 27704
rect 28814 25608 28870 25664
rect 28078 23840 28134 23896
rect 28446 24248 28502 24304
rect 27618 21120 27674 21176
rect 27342 19896 27398 19952
rect 28538 23432 28594 23488
rect 28446 23296 28502 23352
rect 28538 22888 28594 22944
rect 28630 22344 28686 22400
rect 28354 20984 28410 21040
rect 27894 20324 27950 20360
rect 27894 20304 27896 20324
rect 27896 20304 27948 20324
rect 27948 20304 27950 20324
rect 27526 19216 27582 19272
rect 27710 19660 27712 19680
rect 27712 19660 27764 19680
rect 27764 19660 27766 19680
rect 27710 19624 27766 19660
rect 27710 19508 27766 19544
rect 27710 19488 27712 19508
rect 27712 19488 27764 19508
rect 27764 19488 27766 19508
rect 27710 19372 27766 19408
rect 27710 19352 27712 19372
rect 27712 19352 27764 19372
rect 27764 19352 27766 19372
rect 27894 20032 27950 20088
rect 26514 12280 26570 12336
rect 22558 10004 22560 10024
rect 22560 10004 22612 10024
rect 22612 10004 22614 10024
rect 22558 9968 22614 10004
rect 20810 7248 20866 7304
rect 24490 10376 24546 10432
rect 27066 13932 27122 13968
rect 27066 13912 27068 13932
rect 27068 13912 27120 13932
rect 27120 13912 27122 13932
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 27434 14612 27490 14648
rect 27434 14592 27436 14612
rect 27436 14592 27488 14612
rect 27488 14592 27490 14612
rect 27250 13776 27306 13832
rect 27250 13640 27306 13696
rect 27894 15136 27950 15192
rect 27802 14340 27858 14376
rect 27802 14320 27804 14340
rect 27804 14320 27856 14340
rect 27856 14320 27858 14340
rect 27802 14184 27858 14240
rect 27618 13812 27620 13832
rect 27620 13812 27672 13832
rect 27672 13812 27674 13832
rect 27618 13776 27674 13812
rect 27434 13504 27490 13560
rect 27526 12280 27582 12336
rect 27434 10920 27490 10976
rect 27618 10104 27674 10160
rect 27434 8236 27436 8256
rect 27436 8236 27488 8256
rect 27488 8236 27490 8256
rect 27434 8200 27490 8236
rect 28262 17720 28318 17776
rect 28078 17040 28134 17096
rect 28998 22480 29054 22536
rect 29458 27376 29514 27432
rect 29458 26288 29514 26344
rect 29274 24112 29330 24168
rect 29458 24148 29460 24168
rect 29460 24148 29512 24168
rect 29512 24148 29514 24168
rect 29458 24112 29514 24148
rect 28998 19932 29000 19952
rect 29000 19932 29052 19952
rect 29052 19932 29054 19952
rect 28998 19896 29054 19932
rect 28538 19352 28594 19408
rect 31390 35128 31446 35184
rect 30654 34040 30710 34096
rect 29826 29280 29882 29336
rect 29826 29008 29882 29064
rect 30010 26580 30066 26616
rect 30010 26560 30012 26580
rect 30012 26560 30064 26580
rect 30064 26560 30066 26580
rect 30010 25064 30066 25120
rect 30010 24248 30066 24304
rect 30654 32136 30710 32192
rect 30286 30912 30342 30968
rect 30470 31728 30526 31784
rect 30286 29280 30342 29336
rect 30378 25780 30380 25800
rect 30380 25780 30432 25800
rect 30432 25780 30434 25800
rect 30378 25744 30434 25780
rect 30378 24384 30434 24440
rect 28630 17196 28686 17232
rect 28630 17176 28632 17196
rect 28632 17176 28684 17196
rect 28684 17176 28686 17196
rect 29182 19488 29238 19544
rect 28906 17060 28962 17096
rect 28906 17040 28908 17060
rect 28908 17040 28960 17060
rect 28960 17040 28962 17060
rect 28446 15156 28502 15192
rect 28446 15136 28448 15156
rect 28448 15136 28500 15156
rect 28500 15136 28502 15156
rect 28170 13932 28226 13968
rect 28170 13912 28172 13932
rect 28172 13912 28224 13932
rect 28224 13912 28226 13932
rect 28354 14456 28410 14512
rect 28354 14048 28410 14104
rect 30102 22616 30158 22672
rect 30010 20032 30066 20088
rect 29642 17604 29698 17640
rect 29642 17584 29644 17604
rect 29644 17584 29696 17604
rect 29696 17584 29698 17604
rect 29458 15136 29514 15192
rect 28630 12416 28686 12472
rect 30838 29280 30894 29336
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 31666 34856 31722 34912
rect 33506 35536 33562 35592
rect 32310 35264 32366 35320
rect 31666 33224 31722 33280
rect 30930 27648 30986 27704
rect 30838 27412 30840 27432
rect 30840 27412 30892 27432
rect 30892 27412 30894 27432
rect 30838 27376 30894 27412
rect 30562 24384 30618 24440
rect 30470 22228 30526 22264
rect 30470 22208 30472 22228
rect 30472 22208 30524 22228
rect 30524 22208 30526 22228
rect 30010 17332 30066 17368
rect 30010 17312 30012 17332
rect 30012 17312 30064 17332
rect 30064 17312 30066 17332
rect 29734 14320 29790 14376
rect 30378 20032 30434 20088
rect 31022 27104 31078 27160
rect 31206 26152 31262 26208
rect 30746 22480 30802 22536
rect 30654 19488 30710 19544
rect 30838 22072 30894 22128
rect 31390 27784 31446 27840
rect 31206 23588 31262 23624
rect 31206 23568 31208 23588
rect 31208 23568 31260 23588
rect 31260 23568 31262 23588
rect 31666 27784 31722 27840
rect 31390 22480 31446 22536
rect 31298 21936 31354 21992
rect 33414 34992 33470 35048
rect 32862 31456 32918 31512
rect 32310 30504 32366 30560
rect 32126 28484 32182 28520
rect 32126 28464 32128 28484
rect 32128 28464 32180 28484
rect 32180 28464 32182 28484
rect 32126 27512 32182 27568
rect 32034 26696 32090 26752
rect 31666 21936 31722 21992
rect 29274 11872 29330 11928
rect 28998 10240 29054 10296
rect 28538 10124 28594 10160
rect 28538 10104 28540 10124
rect 28540 10104 28592 10124
rect 28592 10104 28594 10124
rect 28354 8200 28410 8256
rect 28170 7792 28226 7848
rect 28630 7384 28686 7440
rect 27710 5480 27766 5536
rect 29642 10784 29698 10840
rect 30194 14728 30250 14784
rect 31114 19252 31116 19272
rect 31116 19252 31168 19272
rect 31168 19252 31170 19272
rect 31114 19216 31170 19252
rect 31574 20868 31630 20904
rect 31574 20848 31576 20868
rect 31576 20848 31628 20868
rect 31628 20848 31630 20868
rect 31574 20712 31630 20768
rect 32586 25336 32642 25392
rect 33598 31728 33654 31784
rect 33414 30368 33470 30424
rect 32770 27376 32826 27432
rect 32310 23568 32366 23624
rect 31390 20168 31446 20224
rect 31390 19916 31446 19952
rect 31390 19896 31392 19916
rect 31392 19896 31444 19916
rect 31444 19896 31446 19916
rect 31390 18672 31446 18728
rect 31482 18536 31538 18592
rect 31298 17720 31354 17776
rect 31758 18536 31814 18592
rect 30378 12824 30434 12880
rect 30286 11056 30342 11112
rect 31574 16088 31630 16144
rect 32218 16788 32274 16824
rect 32218 16768 32220 16788
rect 32220 16768 32272 16788
rect 32272 16768 32274 16788
rect 33414 27412 33416 27432
rect 33416 27412 33468 27432
rect 33468 27412 33470 27432
rect 32954 25336 33010 25392
rect 32954 24520 33010 24576
rect 32862 23840 32918 23896
rect 31942 14492 31944 14512
rect 31944 14492 31996 14512
rect 31996 14492 31998 14512
rect 31942 14456 31998 14492
rect 30838 13368 30894 13424
rect 30930 12144 30986 12200
rect 29734 7384 29790 7440
rect 30102 7928 30158 7984
rect 30562 9172 30618 9208
rect 30562 9152 30564 9172
rect 30564 9152 30616 9172
rect 30616 9152 30618 9172
rect 30378 7520 30434 7576
rect 31298 8472 31354 8528
rect 31022 7792 31078 7848
rect 30378 6568 30434 6624
rect 33414 27376 33470 27412
rect 34058 34720 34114 34776
rect 33782 34196 33838 34232
rect 33782 34176 33784 34196
rect 33784 34176 33836 34196
rect 33836 34176 33838 34196
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 33874 31628 33876 31648
rect 33876 31628 33928 31648
rect 33928 31628 33930 31648
rect 33874 31592 33930 31628
rect 33782 31048 33838 31104
rect 34334 31592 34390 31648
rect 34242 31320 34298 31376
rect 34610 32680 34666 32736
rect 34610 31764 34612 31784
rect 34612 31764 34664 31784
rect 34664 31764 34666 31784
rect 34610 31728 34666 31764
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 33874 30368 33930 30424
rect 33414 27240 33470 27296
rect 33506 26832 33562 26888
rect 33414 25064 33470 25120
rect 33322 24656 33378 24712
rect 33322 24112 33378 24168
rect 33138 18572 33140 18592
rect 33140 18572 33192 18592
rect 33192 18572 33194 18592
rect 33138 18536 33194 18572
rect 32770 14728 32826 14784
rect 32586 13776 32642 13832
rect 32586 12980 32642 13016
rect 32586 12960 32588 12980
rect 32588 12960 32640 12980
rect 32640 12960 32642 12980
rect 32402 12280 32458 12336
rect 31666 8492 31722 8528
rect 31666 8472 31668 8492
rect 31668 8472 31720 8492
rect 31720 8472 31722 8492
rect 32494 8336 32550 8392
rect 33782 27648 33838 27704
rect 33598 25744 33654 25800
rect 33598 25220 33654 25256
rect 33598 25200 33600 25220
rect 33600 25200 33652 25220
rect 33652 25200 33654 25220
rect 33598 19388 33600 19408
rect 33600 19388 33652 19408
rect 33652 19388 33654 19408
rect 33598 19352 33654 19388
rect 34058 29008 34114 29064
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35438 32272 35494 32328
rect 35346 31764 35348 31784
rect 35348 31764 35400 31784
rect 35400 31764 35402 31784
rect 35346 31728 35402 31764
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34794 30504 34850 30560
rect 34610 28328 34666 28384
rect 34426 27240 34482 27296
rect 34426 26288 34482 26344
rect 33874 24520 33930 24576
rect 34242 25200 34298 25256
rect 34426 25336 34482 25392
rect 34150 24656 34206 24712
rect 33414 18128 33470 18184
rect 33782 18400 33838 18456
rect 34058 19080 34114 19136
rect 33506 17176 33562 17232
rect 33506 17040 33562 17096
rect 33414 16652 33470 16688
rect 33414 16632 33416 16652
rect 33416 16632 33468 16652
rect 33468 16632 33470 16652
rect 33046 10804 33102 10840
rect 33046 10784 33048 10804
rect 33048 10784 33100 10804
rect 33100 10784 33102 10804
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 35254 29688 35310 29744
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34702 27920 34758 27976
rect 34610 27648 34666 27704
rect 34518 23740 34520 23760
rect 34520 23740 34572 23760
rect 34572 23740 34574 23760
rect 34518 23704 34574 23740
rect 34334 21664 34390 21720
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 35070 27396 35126 27432
rect 35070 27376 35072 27396
rect 35072 27376 35124 27396
rect 35124 27376 35126 27396
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35070 26152 35126 26208
rect 35990 31864 36046 31920
rect 36082 31728 36138 31784
rect 36358 31456 36414 31512
rect 35806 30096 35862 30152
rect 35530 26288 35586 26344
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34702 24656 34758 24712
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34794 24384 34850 24440
rect 34610 20440 34666 20496
rect 34334 17992 34390 18048
rect 33782 13776 33838 13832
rect 34058 16632 34114 16688
rect 34426 16516 34482 16552
rect 34426 16496 34428 16516
rect 34428 16496 34480 16516
rect 34480 16496 34482 16516
rect 34518 16360 34574 16416
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34886 22480 34942 22536
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 35898 27920 35954 27976
rect 35530 22616 35586 22672
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34702 18808 34758 18864
rect 33598 11092 33600 11112
rect 33600 11092 33652 11112
rect 33652 11092 33654 11112
rect 33598 11056 33654 11092
rect 32770 9152 32826 9208
rect 34058 12844 34114 12880
rect 34058 12824 34060 12844
rect 34060 12824 34112 12844
rect 34112 12824 34114 12844
rect 35070 18808 35126 18864
rect 34978 18128 35034 18184
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34978 16496 35034 16552
rect 36266 29416 36322 29472
rect 36174 29008 36230 29064
rect 36082 25780 36084 25800
rect 36084 25780 36136 25800
rect 36136 25780 36138 25800
rect 36082 25744 36138 25780
rect 35898 19796 35900 19816
rect 35900 19796 35952 19816
rect 35952 19796 35954 19816
rect 35898 19760 35954 19796
rect 35622 18672 35678 18728
rect 35806 18536 35862 18592
rect 35898 18400 35954 18456
rect 35714 17312 35770 17368
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 35438 16244 35494 16280
rect 35438 16224 35440 16244
rect 35440 16224 35492 16244
rect 35492 16224 35494 16244
rect 35438 16108 35494 16144
rect 35438 16088 35440 16108
rect 35440 16088 35492 16108
rect 35492 16088 35494 16108
rect 34794 15272 34850 15328
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34518 13776 34574 13832
rect 33966 9444 34022 9480
rect 33966 9424 33968 9444
rect 33968 9424 34020 9444
rect 34020 9424 34022 9444
rect 33690 7420 33692 7440
rect 33692 7420 33744 7440
rect 33744 7420 33746 7440
rect 33690 7384 33746 7420
rect 33322 6840 33378 6896
rect 33322 6740 33324 6760
rect 33324 6740 33376 6760
rect 33376 6740 33378 6760
rect 33322 6704 33378 6740
rect 32586 5652 32588 5672
rect 32588 5652 32640 5672
rect 32640 5652 32642 5672
rect 32586 5616 32642 5652
rect 31666 5364 31722 5400
rect 31666 5344 31668 5364
rect 31668 5344 31720 5364
rect 31720 5344 31722 5364
rect 34794 14048 34850 14104
rect 34518 13232 34574 13288
rect 34426 11736 34482 11792
rect 35070 13776 35126 13832
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 35070 11772 35072 11792
rect 35072 11772 35124 11792
rect 35124 11772 35126 11792
rect 35070 11736 35126 11772
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35438 14728 35494 14784
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34610 9560 34666 9616
rect 35254 9460 35256 9480
rect 35256 9460 35308 9480
rect 35308 9460 35310 9480
rect 35254 9424 35310 9460
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 35162 7404 35218 7440
rect 35162 7384 35164 7404
rect 35164 7384 35216 7404
rect 35216 7384 35218 7404
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 36174 22888 36230 22944
rect 36726 28756 36782 28792
rect 36726 28736 36728 28756
rect 36728 28736 36780 28756
rect 36780 28736 36782 28756
rect 40958 40876 40960 40896
rect 40960 40876 41012 40896
rect 41012 40876 41014 40896
rect 40958 40840 41014 40876
rect 37370 30232 37426 30288
rect 36174 19488 36230 19544
rect 36174 17720 36230 17776
rect 36082 16496 36138 16552
rect 35990 12008 36046 12064
rect 36542 20712 36598 20768
rect 36450 20576 36506 20632
rect 36542 17176 36598 17232
rect 36266 16632 36322 16688
rect 36266 16224 36322 16280
rect 36358 13232 36414 13288
rect 35898 8336 35954 8392
rect 35622 8200 35678 8256
rect 35622 7384 35678 7440
rect 36082 7928 36138 7984
rect 35990 7248 36046 7304
rect 35806 6840 35862 6896
rect 33966 6568 34022 6624
rect 35438 6704 35494 6760
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34334 5344 34390 5400
rect 37002 29280 37058 29336
rect 37370 29028 37426 29064
rect 37370 29008 37372 29028
rect 37372 29008 37424 29028
rect 37424 29008 37426 29028
rect 38198 31320 38254 31376
rect 38382 28600 38438 28656
rect 38198 28464 38254 28520
rect 38382 27648 38438 27704
rect 40958 36760 41014 36816
rect 40958 32680 41014 32736
rect 40774 32428 40830 32464
rect 40774 32408 40776 32428
rect 40776 32408 40828 32428
rect 40828 32408 40830 32428
rect 39854 29280 39910 29336
rect 37094 24928 37150 24984
rect 37554 23432 37610 23488
rect 37738 25336 37794 25392
rect 37738 23468 37740 23488
rect 37740 23468 37792 23488
rect 37792 23468 37794 23488
rect 37738 23432 37794 23468
rect 37186 20712 37242 20768
rect 37278 16088 37334 16144
rect 37094 14184 37150 14240
rect 36818 11736 36874 11792
rect 37278 13368 37334 13424
rect 37278 12960 37334 13016
rect 37554 15136 37610 15192
rect 37830 13640 37886 13696
rect 37462 9560 37518 9616
rect 38566 18536 38622 18592
rect 38474 17040 38530 17096
rect 38842 20712 38898 20768
rect 38566 13368 38622 13424
rect 40406 27920 40462 27976
rect 38566 11872 38622 11928
rect 39026 13640 39082 13696
rect 39118 13504 39174 13560
rect 38106 10920 38162 10976
rect 39118 11636 39120 11656
rect 39120 11636 39172 11656
rect 39172 11636 39174 11656
rect 39118 11600 39174 11636
rect 39946 14476 40002 14512
rect 39946 14456 39948 14476
rect 39948 14456 40000 14476
rect 40000 14456 40002 14476
rect 39762 14320 39818 14376
rect 39394 12280 39450 12336
rect 40222 12280 40278 12336
rect 40038 11636 40040 11656
rect 40040 11636 40092 11656
rect 40092 11636 40094 11656
rect 40038 11600 40094 11636
rect 41142 28192 41198 28248
rect 41418 21120 41474 21176
rect 41878 23024 41934 23080
rect 41602 9560 41658 9616
rect 35714 5652 35716 5672
rect 35716 5652 35768 5672
rect 35768 5652 35770 5672
rect 35714 5616 35770 5652
rect 35990 5480 36046 5536
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 41326 5516 41328 5536
rect 41328 5516 41380 5536
rect 41380 5516 41382 5536
rect 41326 5480 41382 5516
<< metal3 >>
rect 0 42938 800 42968
rect 3417 42938 3483 42941
rect 0 42936 3483 42938
rect 0 42880 3422 42936
rect 3478 42880 3483 42936
rect 0 42878 3483 42880
rect 0 42848 800 42878
rect 3417 42875 3483 42878
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 17718 42196 17724 42260
rect 17788 42258 17794 42260
rect 34513 42258 34579 42261
rect 17788 42256 34579 42258
rect 17788 42200 34518 42256
rect 34574 42200 34579 42256
rect 17788 42198 34579 42200
rect 17788 42196 17794 42198
rect 34513 42195 34579 42198
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 31293 41444 31359 41445
rect 31293 41440 31340 41444
rect 31404 41442 31410 41444
rect 31293 41384 31298 41440
rect 31293 41380 31340 41384
rect 31404 41382 31450 41442
rect 31404 41380 31410 41382
rect 31293 41379 31359 41380
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 40953 40898 41019 40901
rect 41749 40898 42549 40928
rect 40953 40896 42549 40898
rect 40953 40840 40958 40896
rect 41014 40840 42549 40896
rect 40953 40838 42549 40840
rect 40953 40835 41019 40838
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 41749 40808 42549 40838
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 9857 40218 9923 40221
rect 10593 40218 10659 40221
rect 9857 40216 10659 40218
rect 9857 40160 9862 40216
rect 9918 40160 10598 40216
rect 10654 40160 10659 40216
rect 9857 40158 10659 40160
rect 9857 40155 9923 40158
rect 10593 40155 10659 40158
rect 10041 40082 10107 40085
rect 10777 40082 10843 40085
rect 10041 40080 10843 40082
rect 10041 40024 10046 40080
rect 10102 40024 10782 40080
rect 10838 40024 10843 40080
rect 10041 40022 10843 40024
rect 10041 40019 10107 40022
rect 10777 40019 10843 40022
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 0 38858 800 38888
rect 3785 38858 3851 38861
rect 0 38856 3851 38858
rect 0 38800 3790 38856
rect 3846 38800 3851 38856
rect 0 38798 3851 38800
rect 0 38768 800 38798
rect 3785 38795 3851 38798
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 17350 37300 17356 37364
rect 17420 37362 17426 37364
rect 22001 37362 22067 37365
rect 17420 37360 22067 37362
rect 17420 37304 22006 37360
rect 22062 37304 22067 37360
rect 17420 37302 22067 37304
rect 17420 37300 17426 37302
rect 22001 37299 22067 37302
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 40953 36818 41019 36821
rect 41749 36818 42549 36848
rect 40953 36816 42549 36818
rect 40953 36760 40958 36816
rect 41014 36760 42549 36816
rect 40953 36758 42549 36760
rect 40953 36755 41019 36758
rect 41749 36728 42549 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 28257 36138 28323 36141
rect 31886 36138 31892 36140
rect 28257 36136 31892 36138
rect 28257 36080 28262 36136
rect 28318 36080 31892 36136
rect 28257 36078 31892 36080
rect 28257 36075 28323 36078
rect 31886 36076 31892 36078
rect 31956 36076 31962 36140
rect 28625 36002 28691 36005
rect 28758 36002 28764 36004
rect 28625 36000 28764 36002
rect 28625 35944 28630 36000
rect 28686 35944 28764 36000
rect 28625 35942 28764 35944
rect 28625 35939 28691 35942
rect 28758 35940 28764 35942
rect 28828 35940 28834 36004
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 25037 35866 25103 35869
rect 26233 35866 26299 35869
rect 25037 35864 26299 35866
rect 25037 35808 25042 35864
rect 25098 35808 26238 35864
rect 26294 35808 26299 35864
rect 25037 35806 26299 35808
rect 25037 35803 25103 35806
rect 26233 35803 26299 35806
rect 10910 35532 10916 35596
rect 10980 35594 10986 35596
rect 15101 35594 15167 35597
rect 10980 35592 15167 35594
rect 10980 35536 15106 35592
rect 15162 35536 15167 35592
rect 10980 35534 15167 35536
rect 10980 35532 10986 35534
rect 15101 35531 15167 35534
rect 26325 35594 26391 35597
rect 29126 35594 29132 35596
rect 26325 35592 29132 35594
rect 26325 35536 26330 35592
rect 26386 35536 29132 35592
rect 26325 35534 29132 35536
rect 26325 35531 26391 35534
rect 29126 35532 29132 35534
rect 29196 35594 29202 35596
rect 33501 35594 33567 35597
rect 29196 35592 33567 35594
rect 29196 35536 33506 35592
rect 33562 35536 33567 35592
rect 29196 35534 33567 35536
rect 29196 35532 29202 35534
rect 33501 35531 33567 35534
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 24117 35322 24183 35325
rect 24945 35322 25011 35325
rect 32305 35322 32371 35325
rect 24117 35320 32371 35322
rect 24117 35264 24122 35320
rect 24178 35264 24950 35320
rect 25006 35264 32310 35320
rect 32366 35264 32371 35320
rect 24117 35262 32371 35264
rect 24117 35259 24183 35262
rect 24945 35259 25011 35262
rect 32305 35259 32371 35262
rect 18781 35186 18847 35189
rect 23933 35186 23999 35189
rect 18781 35184 23999 35186
rect 18781 35128 18786 35184
rect 18842 35128 23938 35184
rect 23994 35128 23999 35184
rect 18781 35126 23999 35128
rect 18781 35123 18847 35126
rect 23933 35123 23999 35126
rect 24577 35186 24643 35189
rect 26693 35186 26759 35189
rect 31385 35186 31451 35189
rect 24577 35184 31451 35186
rect 24577 35128 24582 35184
rect 24638 35128 26698 35184
rect 26754 35128 31390 35184
rect 31446 35128 31451 35184
rect 24577 35126 31451 35128
rect 24577 35123 24643 35126
rect 26693 35123 26759 35126
rect 31385 35123 31451 35126
rect 11605 35050 11671 35053
rect 16481 35050 16547 35053
rect 11605 35048 16547 35050
rect 11605 34992 11610 35048
rect 11666 34992 16486 35048
rect 16542 34992 16547 35048
rect 11605 34990 16547 34992
rect 11605 34987 11671 34990
rect 16481 34987 16547 34990
rect 22686 34988 22692 35052
rect 22756 35050 22762 35052
rect 22829 35050 22895 35053
rect 25405 35050 25471 35053
rect 33409 35050 33475 35053
rect 22756 35048 33475 35050
rect 22756 34992 22834 35048
rect 22890 34992 25410 35048
rect 25466 34992 33414 35048
rect 33470 34992 33475 35048
rect 22756 34990 33475 34992
rect 22756 34988 22762 34990
rect 22829 34987 22895 34990
rect 25405 34987 25471 34990
rect 33409 34987 33475 34990
rect 26141 34914 26207 34917
rect 31661 34914 31727 34917
rect 26141 34912 31727 34914
rect 26141 34856 26146 34912
rect 26202 34856 31666 34912
rect 31722 34856 31727 34912
rect 26141 34854 31727 34856
rect 26141 34851 26207 34854
rect 31661 34851 31727 34854
rect 19570 34848 19886 34849
rect 0 34778 800 34808
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 1025 34778 1091 34781
rect 0 34776 1091 34778
rect 0 34720 1030 34776
rect 1086 34720 1091 34776
rect 0 34718 1091 34720
rect 0 34688 800 34718
rect 1025 34715 1091 34718
rect 20110 34716 20116 34780
rect 20180 34778 20186 34780
rect 22553 34778 22619 34781
rect 20180 34776 22619 34778
rect 20180 34720 22558 34776
rect 22614 34720 22619 34776
rect 20180 34718 22619 34720
rect 20180 34716 20186 34718
rect 22553 34715 22619 34718
rect 26601 34778 26667 34781
rect 27613 34778 27679 34781
rect 26601 34776 27679 34778
rect 26601 34720 26606 34776
rect 26662 34720 27618 34776
rect 27674 34720 27679 34776
rect 26601 34718 27679 34720
rect 26601 34715 26667 34718
rect 27613 34715 27679 34718
rect 30005 34778 30071 34781
rect 34053 34778 34119 34781
rect 30005 34776 34119 34778
rect 30005 34720 30010 34776
rect 30066 34720 34058 34776
rect 34114 34720 34119 34776
rect 30005 34718 34119 34720
rect 30005 34715 30071 34718
rect 34053 34715 34119 34718
rect 1853 34642 1919 34645
rect 20253 34642 20319 34645
rect 24577 34644 24643 34645
rect 29913 34644 29979 34645
rect 1853 34640 20319 34642
rect 1853 34584 1858 34640
rect 1914 34584 20258 34640
rect 20314 34584 20319 34640
rect 1853 34582 20319 34584
rect 1853 34579 1919 34582
rect 20253 34579 20319 34582
rect 24526 34580 24532 34644
rect 24596 34642 24643 34644
rect 24596 34640 24688 34642
rect 24638 34584 24688 34640
rect 24596 34582 24688 34584
rect 24596 34580 24643 34582
rect 28942 34580 28948 34644
rect 29012 34642 29018 34644
rect 29012 34582 29746 34642
rect 29012 34580 29018 34582
rect 24577 34579 24643 34580
rect 29686 34509 29746 34582
rect 29862 34580 29868 34644
rect 29932 34642 29979 34644
rect 29932 34640 30024 34642
rect 29974 34584 30024 34640
rect 29932 34582 30024 34584
rect 29932 34580 29979 34582
rect 29913 34579 29979 34580
rect 29686 34504 29795 34509
rect 29686 34448 29734 34504
rect 29790 34448 29795 34504
rect 29686 34446 29795 34448
rect 29729 34443 29795 34446
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 29545 34234 29611 34237
rect 33777 34234 33843 34237
rect 34646 34234 34652 34236
rect 29545 34232 34652 34234
rect 29545 34176 29550 34232
rect 29606 34176 33782 34232
rect 33838 34176 34652 34232
rect 29545 34174 34652 34176
rect 29545 34171 29611 34174
rect 33777 34171 33843 34174
rect 34646 34172 34652 34174
rect 34716 34172 34722 34236
rect 19609 34098 19675 34101
rect 20529 34098 20595 34101
rect 19609 34096 20595 34098
rect 19609 34040 19614 34096
rect 19670 34040 20534 34096
rect 20590 34040 20595 34096
rect 19609 34038 20595 34040
rect 19609 34035 19675 34038
rect 20529 34035 20595 34038
rect 21449 34098 21515 34101
rect 30649 34098 30715 34101
rect 21449 34096 30715 34098
rect 21449 34040 21454 34096
rect 21510 34040 30654 34096
rect 30710 34040 30715 34096
rect 21449 34038 30715 34040
rect 21449 34035 21515 34038
rect 30649 34035 30715 34038
rect 20069 33962 20135 33965
rect 21357 33962 21423 33965
rect 20069 33960 21423 33962
rect 20069 33904 20074 33960
rect 20130 33904 21362 33960
rect 21418 33904 21423 33960
rect 20069 33902 21423 33904
rect 20069 33899 20135 33902
rect 21357 33899 21423 33902
rect 22829 33962 22895 33965
rect 25405 33962 25471 33965
rect 22829 33960 25471 33962
rect 22829 33904 22834 33960
rect 22890 33904 25410 33960
rect 25466 33904 25471 33960
rect 22829 33902 25471 33904
rect 22829 33899 22895 33902
rect 25405 33899 25471 33902
rect 19977 33826 20043 33829
rect 20529 33826 20595 33829
rect 19977 33824 20595 33826
rect 19977 33768 19982 33824
rect 20038 33768 20534 33824
rect 20590 33768 20595 33824
rect 19977 33766 20595 33768
rect 19977 33763 20043 33766
rect 20529 33763 20595 33766
rect 24761 33826 24827 33829
rect 27061 33826 27127 33829
rect 24761 33824 27127 33826
rect 24761 33768 24766 33824
rect 24822 33768 27066 33824
rect 27122 33768 27127 33824
rect 24761 33766 27127 33768
rect 24761 33763 24827 33766
rect 27061 33763 27127 33766
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 26693 33284 26759 33285
rect 26693 33282 26740 33284
rect 26648 33280 26740 33282
rect 26648 33224 26698 33280
rect 26648 33222 26740 33224
rect 26693 33220 26740 33222
rect 26804 33220 26810 33284
rect 31661 33282 31727 33285
rect 32438 33282 32444 33284
rect 31661 33280 32444 33282
rect 31661 33224 31666 33280
rect 31722 33224 32444 33280
rect 31661 33222 32444 33224
rect 26693 33219 26759 33220
rect 31661 33219 31727 33222
rect 32438 33220 32444 33222
rect 32508 33220 32514 33284
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 26417 33146 26483 33149
rect 28809 33146 28875 33149
rect 26417 33144 28875 33146
rect 26417 33088 26422 33144
rect 26478 33088 28814 33144
rect 28870 33088 28875 33144
rect 26417 33086 28875 33088
rect 26417 33083 26483 33086
rect 28809 33083 28875 33086
rect 11605 32874 11671 32877
rect 11830 32874 11836 32876
rect 11605 32872 11836 32874
rect 11605 32816 11610 32872
rect 11666 32816 11836 32872
rect 11605 32814 11836 32816
rect 11605 32811 11671 32814
rect 11830 32812 11836 32814
rect 11900 32812 11906 32876
rect 20161 32874 20227 32877
rect 20478 32874 20484 32876
rect 20161 32872 20484 32874
rect 20161 32816 20166 32872
rect 20222 32816 20484 32872
rect 20161 32814 20484 32816
rect 20161 32811 20227 32814
rect 20478 32812 20484 32814
rect 20548 32812 20554 32876
rect 28809 32738 28875 32741
rect 34462 32738 34468 32740
rect 28809 32736 34468 32738
rect 28809 32680 28814 32736
rect 28870 32680 34468 32736
rect 28809 32678 34468 32680
rect 28809 32675 28875 32678
rect 34462 32676 34468 32678
rect 34532 32738 34538 32740
rect 34605 32738 34671 32741
rect 34532 32736 34671 32738
rect 34532 32680 34610 32736
rect 34666 32680 34671 32736
rect 34532 32678 34671 32680
rect 34532 32676 34538 32678
rect 34605 32675 34671 32678
rect 40953 32738 41019 32741
rect 41749 32738 42549 32768
rect 40953 32736 42549 32738
rect 40953 32680 40958 32736
rect 41014 32680 42549 32736
rect 40953 32678 42549 32680
rect 40953 32675 41019 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 41749 32648 42549 32678
rect 19570 32607 19886 32608
rect 27981 32604 28047 32605
rect 27981 32602 28028 32604
rect 27936 32600 28028 32602
rect 27936 32544 27986 32600
rect 27936 32542 28028 32544
rect 27981 32540 28028 32542
rect 28092 32540 28098 32604
rect 27981 32539 28047 32540
rect 21357 32466 21423 32469
rect 40769 32466 40835 32469
rect 21357 32464 40835 32466
rect 21357 32408 21362 32464
rect 21418 32408 40774 32464
rect 40830 32408 40835 32464
rect 21357 32406 40835 32408
rect 21357 32403 21423 32406
rect 40769 32403 40835 32406
rect 15878 32268 15884 32332
rect 15948 32330 15954 32332
rect 19977 32330 20043 32333
rect 15948 32328 20043 32330
rect 15948 32272 19982 32328
rect 20038 32272 20043 32328
rect 15948 32270 20043 32272
rect 15948 32268 15954 32270
rect 19977 32267 20043 32270
rect 26141 32330 26207 32333
rect 26969 32330 27035 32333
rect 35433 32330 35499 32333
rect 26141 32328 35499 32330
rect 26141 32272 26146 32328
rect 26202 32272 26974 32328
rect 27030 32272 35438 32328
rect 35494 32272 35499 32328
rect 26141 32270 35499 32272
rect 26141 32267 26207 32270
rect 26969 32267 27035 32270
rect 35433 32267 35499 32270
rect 30649 32196 30715 32197
rect 30598 32132 30604 32196
rect 30668 32194 30715 32196
rect 30668 32192 30760 32194
rect 30710 32136 30760 32192
rect 30668 32134 30760 32136
rect 30668 32132 30715 32134
rect 30649 32131 30715 32132
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 23841 31922 23907 31925
rect 26325 31922 26391 31925
rect 35985 31924 36051 31925
rect 35934 31922 35940 31924
rect 23841 31920 26391 31922
rect 23841 31864 23846 31920
rect 23902 31864 26330 31920
rect 26386 31864 26391 31920
rect 23841 31862 26391 31864
rect 23841 31859 23907 31862
rect 26325 31859 26391 31862
rect 31894 31862 35940 31922
rect 36004 31920 36051 31924
rect 36046 31864 36051 31920
rect 22093 31786 22159 31789
rect 22553 31786 22619 31789
rect 22093 31784 22619 31786
rect 22093 31728 22098 31784
rect 22154 31728 22558 31784
rect 22614 31728 22619 31784
rect 22093 31726 22619 31728
rect 22093 31723 22159 31726
rect 22553 31723 22619 31726
rect 24853 31786 24919 31789
rect 30465 31786 30531 31789
rect 31894 31786 31954 31862
rect 35934 31860 35940 31862
rect 36004 31860 36051 31864
rect 35985 31859 36051 31860
rect 24853 31784 25468 31786
rect 24853 31728 24858 31784
rect 24914 31728 25468 31784
rect 24853 31726 25468 31728
rect 24853 31723 24919 31726
rect 23289 31652 23355 31653
rect 23238 31650 23244 31652
rect 23198 31590 23244 31650
rect 23308 31648 23355 31652
rect 23350 31592 23355 31648
rect 23238 31588 23244 31590
rect 23308 31588 23355 31592
rect 25408 31650 25468 31726
rect 30465 31784 31954 31786
rect 30465 31728 30470 31784
rect 30526 31728 31954 31784
rect 30465 31726 31954 31728
rect 33593 31786 33659 31789
rect 34605 31786 34671 31789
rect 35341 31788 35407 31789
rect 35341 31786 35388 31788
rect 33593 31784 34671 31786
rect 33593 31728 33598 31784
rect 33654 31728 34610 31784
rect 34666 31728 34671 31784
rect 33593 31726 34671 31728
rect 35296 31784 35388 31786
rect 35452 31786 35458 31788
rect 36077 31786 36143 31789
rect 35452 31784 36143 31786
rect 35296 31728 35346 31784
rect 35452 31728 36082 31784
rect 36138 31728 36143 31784
rect 35296 31726 35388 31728
rect 30465 31723 30531 31726
rect 33593 31723 33659 31726
rect 34605 31723 34671 31726
rect 35341 31724 35388 31726
rect 35452 31726 36143 31728
rect 35452 31724 35458 31726
rect 35341 31723 35407 31724
rect 36077 31723 36143 31726
rect 27889 31650 27955 31653
rect 25408 31648 27955 31650
rect 25408 31592 27894 31648
rect 27950 31592 27955 31648
rect 25408 31590 27955 31592
rect 23289 31587 23355 31588
rect 27889 31587 27955 31590
rect 33869 31650 33935 31653
rect 34329 31650 34395 31653
rect 33869 31648 34395 31650
rect 33869 31592 33874 31648
rect 33930 31592 34334 31648
rect 34390 31592 34395 31648
rect 33869 31590 34395 31592
rect 33869 31587 33935 31590
rect 34329 31587 34395 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 24301 31514 24367 31517
rect 28165 31514 28231 31517
rect 24301 31512 28231 31514
rect 24301 31456 24306 31512
rect 24362 31456 28170 31512
rect 28226 31456 28231 31512
rect 24301 31454 28231 31456
rect 24301 31451 24367 31454
rect 28165 31451 28231 31454
rect 32857 31514 32923 31517
rect 36353 31514 36419 31517
rect 32857 31512 36419 31514
rect 32857 31456 32862 31512
rect 32918 31456 36358 31512
rect 36414 31456 36419 31512
rect 32857 31454 36419 31456
rect 32857 31451 32923 31454
rect 36353 31451 36419 31454
rect 24025 31378 24091 31381
rect 28441 31378 28507 31381
rect 24025 31376 28507 31378
rect 24025 31320 24030 31376
rect 24086 31320 28446 31376
rect 28502 31320 28507 31376
rect 24025 31318 28507 31320
rect 24025 31315 24091 31318
rect 28441 31315 28507 31318
rect 34237 31378 34303 31381
rect 38193 31378 38259 31381
rect 34237 31376 38259 31378
rect 34237 31320 34242 31376
rect 34298 31320 38198 31376
rect 38254 31320 38259 31376
rect 34237 31318 38259 31320
rect 34237 31315 34303 31318
rect 38193 31315 38259 31318
rect 22277 31244 22343 31245
rect 22277 31242 22324 31244
rect 22232 31240 22324 31242
rect 22232 31184 22282 31240
rect 22232 31182 22324 31184
rect 22277 31180 22324 31182
rect 22388 31180 22394 31244
rect 24761 31242 24827 31245
rect 27337 31242 27403 31245
rect 24761 31240 27403 31242
rect 24761 31184 24766 31240
rect 24822 31184 27342 31240
rect 27398 31184 27403 31240
rect 24761 31182 27403 31184
rect 22277 31179 22343 31180
rect 24761 31179 24827 31182
rect 27337 31179 27403 31182
rect 21725 31106 21791 31109
rect 24945 31106 25011 31109
rect 21725 31104 25011 31106
rect 21725 31048 21730 31104
rect 21786 31048 24950 31104
rect 25006 31048 25011 31104
rect 21725 31046 25011 31048
rect 21725 31043 21791 31046
rect 24945 31043 25011 31046
rect 29453 31106 29519 31109
rect 32254 31106 32260 31108
rect 29453 31104 32260 31106
rect 29453 31048 29458 31104
rect 29514 31048 32260 31104
rect 29453 31046 32260 31048
rect 29453 31043 29519 31046
rect 32254 31044 32260 31046
rect 32324 31106 32330 31108
rect 33777 31106 33843 31109
rect 32324 31104 33843 31106
rect 32324 31048 33782 31104
rect 33838 31048 33843 31104
rect 32324 31046 33843 31048
rect 32324 31044 32330 31046
rect 33777 31043 33843 31046
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 16389 30970 16455 30973
rect 16982 30970 16988 30972
rect 16389 30968 16988 30970
rect 16389 30912 16394 30968
rect 16450 30912 16988 30968
rect 16389 30910 16988 30912
rect 16389 30907 16455 30910
rect 16982 30908 16988 30910
rect 17052 30908 17058 30972
rect 24894 30908 24900 30972
rect 24964 30970 24970 30972
rect 30281 30970 30347 30973
rect 24964 30968 30347 30970
rect 24964 30912 30286 30968
rect 30342 30912 30347 30968
rect 24964 30910 30347 30912
rect 24964 30908 24970 30910
rect 30281 30907 30347 30910
rect 21081 30834 21147 30837
rect 22185 30834 22251 30837
rect 21081 30832 22251 30834
rect 21081 30776 21086 30832
rect 21142 30776 22190 30832
rect 22246 30776 22251 30832
rect 21081 30774 22251 30776
rect 21081 30771 21147 30774
rect 22185 30771 22251 30774
rect 0 30698 800 30728
rect 2773 30698 2839 30701
rect 0 30696 2839 30698
rect 0 30640 2778 30696
rect 2834 30640 2839 30696
rect 0 30638 2839 30640
rect 0 30608 800 30638
rect 2773 30635 2839 30638
rect 16941 30698 17007 30701
rect 17534 30698 17540 30700
rect 16941 30696 17540 30698
rect 16941 30640 16946 30696
rect 17002 30640 17540 30696
rect 16941 30638 17540 30640
rect 16941 30635 17007 30638
rect 17534 30636 17540 30638
rect 17604 30636 17610 30700
rect 11973 30564 12039 30565
rect 11973 30562 12020 30564
rect 11928 30560 12020 30562
rect 11928 30504 11978 30560
rect 11928 30502 12020 30504
rect 11973 30500 12020 30502
rect 12084 30500 12090 30564
rect 13670 30500 13676 30564
rect 13740 30562 13746 30564
rect 17677 30562 17743 30565
rect 13740 30560 17743 30562
rect 13740 30504 17682 30560
rect 17738 30504 17743 30560
rect 13740 30502 17743 30504
rect 13740 30500 13746 30502
rect 11973 30499 12039 30500
rect 17677 30499 17743 30502
rect 25037 30562 25103 30565
rect 26182 30562 26188 30564
rect 25037 30560 26188 30562
rect 25037 30504 25042 30560
rect 25098 30504 26188 30560
rect 25037 30502 26188 30504
rect 25037 30499 25103 30502
rect 26182 30500 26188 30502
rect 26252 30500 26258 30564
rect 28574 30500 28580 30564
rect 28644 30562 28650 30564
rect 28901 30562 28967 30565
rect 28644 30560 28967 30562
rect 28644 30504 28906 30560
rect 28962 30504 28967 30560
rect 28644 30502 28967 30504
rect 28644 30500 28650 30502
rect 28901 30499 28967 30502
rect 32305 30562 32371 30565
rect 34789 30562 34855 30565
rect 32305 30560 34855 30562
rect 32305 30504 32310 30560
rect 32366 30504 34794 30560
rect 34850 30504 34855 30560
rect 32305 30502 34855 30504
rect 32305 30499 32371 30502
rect 34789 30499 34855 30502
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 11094 30364 11100 30428
rect 11164 30426 11170 30428
rect 11605 30426 11671 30429
rect 12709 30428 12775 30429
rect 25865 30428 25931 30429
rect 12709 30426 12756 30428
rect 11164 30424 11671 30426
rect 11164 30368 11610 30424
rect 11666 30368 11671 30424
rect 11164 30366 11671 30368
rect 12664 30424 12756 30426
rect 12664 30368 12714 30424
rect 12664 30366 12756 30368
rect 11164 30364 11170 30366
rect 11605 30363 11671 30366
rect 12709 30364 12756 30366
rect 12820 30364 12826 30428
rect 25814 30364 25820 30428
rect 25884 30426 25931 30428
rect 29453 30426 29519 30429
rect 33409 30426 33475 30429
rect 25884 30424 25976 30426
rect 25926 30368 25976 30424
rect 25884 30366 25976 30368
rect 29453 30424 33475 30426
rect 29453 30368 29458 30424
rect 29514 30368 33414 30424
rect 33470 30368 33475 30424
rect 29453 30366 33475 30368
rect 25884 30364 25931 30366
rect 12709 30363 12775 30364
rect 25865 30363 25931 30364
rect 29453 30363 29519 30366
rect 33409 30363 33475 30366
rect 33542 30364 33548 30428
rect 33612 30426 33618 30428
rect 33869 30426 33935 30429
rect 33612 30424 33935 30426
rect 33612 30368 33874 30424
rect 33930 30368 33935 30424
rect 33612 30366 33935 30368
rect 33612 30364 33618 30366
rect 33869 30363 33935 30366
rect 28257 30290 28323 30293
rect 37365 30290 37431 30293
rect 28257 30288 37431 30290
rect 28257 30232 28262 30288
rect 28318 30232 37370 30288
rect 37426 30232 37431 30288
rect 28257 30230 37431 30232
rect 28257 30227 28323 30230
rect 37365 30227 37431 30230
rect 20437 30154 20503 30157
rect 21173 30154 21239 30157
rect 24393 30156 24459 30157
rect 20437 30152 21239 30154
rect 20437 30096 20442 30152
rect 20498 30096 21178 30152
rect 21234 30096 21239 30152
rect 20437 30094 21239 30096
rect 20437 30091 20503 30094
rect 21173 30091 21239 30094
rect 24342 30092 24348 30156
rect 24412 30154 24459 30156
rect 35801 30154 35867 30157
rect 24412 30152 24504 30154
rect 24454 30096 24504 30152
rect 24412 30094 24504 30096
rect 31710 30152 35867 30154
rect 31710 30096 35806 30152
rect 35862 30096 35867 30152
rect 31710 30094 35867 30096
rect 24412 30092 24459 30094
rect 24393 30091 24459 30092
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 8293 29882 8359 29885
rect 8845 29882 8911 29885
rect 8293 29880 8911 29882
rect 8293 29824 8298 29880
rect 8354 29824 8850 29880
rect 8906 29824 8911 29880
rect 8293 29822 8911 29824
rect 8293 29819 8359 29822
rect 8845 29819 8911 29822
rect 4521 29746 4587 29749
rect 9857 29746 9923 29749
rect 12525 29746 12591 29749
rect 4521 29744 12591 29746
rect 4521 29688 4526 29744
rect 4582 29688 9862 29744
rect 9918 29688 12530 29744
rect 12586 29688 12591 29744
rect 4521 29686 12591 29688
rect 4521 29683 4587 29686
rect 9857 29683 9923 29686
rect 12525 29683 12591 29686
rect 17953 29746 18019 29749
rect 18086 29746 18092 29748
rect 17953 29744 18092 29746
rect 17953 29688 17958 29744
rect 18014 29688 18092 29744
rect 17953 29686 18092 29688
rect 17953 29683 18019 29686
rect 18086 29684 18092 29686
rect 18156 29684 18162 29748
rect 19885 29746 19951 29749
rect 29862 29746 29868 29748
rect 19885 29744 29868 29746
rect 19885 29688 19890 29744
rect 19946 29688 29868 29744
rect 19885 29686 29868 29688
rect 19885 29683 19951 29686
rect 29862 29684 29868 29686
rect 29932 29684 29938 29748
rect 7097 29610 7163 29613
rect 7741 29610 7807 29613
rect 10133 29610 10199 29613
rect 31710 29610 31770 30094
rect 35801 30091 35867 30094
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 35249 29746 35315 29749
rect 35382 29746 35388 29748
rect 35249 29744 35388 29746
rect 35249 29688 35254 29744
rect 35310 29688 35388 29744
rect 35249 29686 35388 29688
rect 35249 29683 35315 29686
rect 35382 29684 35388 29686
rect 35452 29684 35458 29748
rect 7097 29608 10199 29610
rect 7097 29552 7102 29608
rect 7158 29552 7746 29608
rect 7802 29552 10138 29608
rect 10194 29552 10199 29608
rect 7097 29550 10199 29552
rect 7097 29547 7163 29550
rect 7741 29547 7807 29550
rect 10133 29547 10199 29550
rect 10320 29550 31770 29610
rect 9806 29412 9812 29476
rect 9876 29474 9882 29476
rect 9949 29474 10015 29477
rect 10320 29474 10380 29550
rect 9876 29472 10380 29474
rect 9876 29416 9954 29472
rect 10010 29416 10380 29472
rect 9876 29414 10380 29416
rect 13261 29474 13327 29477
rect 13997 29474 14063 29477
rect 13261 29472 14063 29474
rect 13261 29416 13266 29472
rect 13322 29416 14002 29472
rect 14058 29416 14063 29472
rect 13261 29414 14063 29416
rect 9876 29412 9882 29414
rect 9949 29411 10015 29414
rect 13261 29411 13327 29414
rect 13997 29411 14063 29414
rect 22461 29474 22527 29477
rect 25865 29474 25931 29477
rect 22461 29472 25931 29474
rect 22461 29416 22466 29472
rect 22522 29416 25870 29472
rect 25926 29416 25931 29472
rect 22461 29414 25931 29416
rect 22461 29411 22527 29414
rect 25865 29411 25931 29414
rect 28165 29474 28231 29477
rect 36261 29474 36327 29477
rect 28165 29472 36327 29474
rect 28165 29416 28170 29472
rect 28226 29416 36266 29472
rect 36322 29416 36327 29472
rect 28165 29414 36327 29416
rect 28165 29411 28231 29414
rect 36261 29411 36327 29414
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 22001 29338 22067 29341
rect 25405 29338 25471 29341
rect 22001 29336 25471 29338
rect 22001 29280 22006 29336
rect 22062 29280 25410 29336
rect 25466 29280 25471 29336
rect 22001 29278 25471 29280
rect 22001 29275 22067 29278
rect 25405 29275 25471 29278
rect 27889 29338 27955 29341
rect 28809 29338 28875 29341
rect 27889 29336 28875 29338
rect 27889 29280 27894 29336
rect 27950 29280 28814 29336
rect 28870 29280 28875 29336
rect 27889 29278 28875 29280
rect 27889 29275 27955 29278
rect 28809 29275 28875 29278
rect 29361 29338 29427 29341
rect 29821 29338 29887 29341
rect 30281 29338 30347 29341
rect 29361 29336 30347 29338
rect 29361 29280 29366 29336
rect 29422 29280 29826 29336
rect 29882 29280 30286 29336
rect 30342 29280 30347 29336
rect 29361 29278 30347 29280
rect 29361 29275 29427 29278
rect 29821 29275 29887 29278
rect 30281 29275 30347 29278
rect 30833 29338 30899 29341
rect 31518 29338 31524 29340
rect 30833 29336 31524 29338
rect 30833 29280 30838 29336
rect 30894 29280 31524 29336
rect 30833 29278 31524 29280
rect 30833 29275 30899 29278
rect 31518 29276 31524 29278
rect 31588 29338 31594 29340
rect 36997 29338 37063 29341
rect 31588 29336 37063 29338
rect 31588 29280 37002 29336
rect 37058 29280 37063 29336
rect 31588 29278 37063 29280
rect 31588 29276 31594 29278
rect 36997 29275 37063 29278
rect 39849 29338 39915 29341
rect 41749 29338 42549 29368
rect 39849 29336 42549 29338
rect 39849 29280 39854 29336
rect 39910 29280 42549 29336
rect 39849 29278 42549 29280
rect 39849 29275 39915 29278
rect 41749 29248 42549 29278
rect 3417 29202 3483 29205
rect 10317 29202 10383 29205
rect 3417 29200 10383 29202
rect 3417 29144 3422 29200
rect 3478 29144 10322 29200
rect 10378 29144 10383 29200
rect 3417 29142 10383 29144
rect 3417 29139 3483 29142
rect 10317 29139 10383 29142
rect 15745 29202 15811 29205
rect 16481 29202 16547 29205
rect 18689 29202 18755 29205
rect 15745 29200 18755 29202
rect 15745 29144 15750 29200
rect 15806 29144 16486 29200
rect 16542 29144 18694 29200
rect 18750 29144 18755 29200
rect 15745 29142 18755 29144
rect 15745 29139 15811 29142
rect 16481 29139 16547 29142
rect 18689 29139 18755 29142
rect 22001 29202 22067 29205
rect 23933 29202 23999 29205
rect 22001 29200 23999 29202
rect 22001 29144 22006 29200
rect 22062 29144 23938 29200
rect 23994 29144 23999 29200
rect 22001 29142 23999 29144
rect 22001 29139 22067 29142
rect 23933 29139 23999 29142
rect 29686 29142 31770 29202
rect 7189 29066 7255 29069
rect 9029 29066 9095 29069
rect 7189 29064 9095 29066
rect 7189 29008 7194 29064
rect 7250 29008 9034 29064
rect 9090 29008 9095 29064
rect 7189 29006 9095 29008
rect 7189 29003 7255 29006
rect 9029 29003 9095 29006
rect 13445 29066 13511 29069
rect 15929 29066 15995 29069
rect 13445 29064 15995 29066
rect 13445 29008 13450 29064
rect 13506 29008 15934 29064
rect 15990 29008 15995 29064
rect 13445 29006 15995 29008
rect 13445 29003 13511 29006
rect 15929 29003 15995 29006
rect 22134 29004 22140 29068
rect 22204 29066 22210 29068
rect 24485 29066 24551 29069
rect 22204 29064 24551 29066
rect 22204 29008 24490 29064
rect 24546 29008 24551 29064
rect 22204 29006 24551 29008
rect 22204 29004 22210 29006
rect 24485 29003 24551 29006
rect 25078 29004 25084 29068
rect 25148 29066 25154 29068
rect 25221 29066 25287 29069
rect 25148 29064 25287 29066
rect 25148 29008 25226 29064
rect 25282 29008 25287 29064
rect 25148 29006 25287 29008
rect 25148 29004 25154 29006
rect 25221 29003 25287 29006
rect 28257 29066 28323 29069
rect 28390 29066 28396 29068
rect 28257 29064 28396 29066
rect 28257 29008 28262 29064
rect 28318 29008 28396 29064
rect 28257 29006 28396 29008
rect 28257 29003 28323 29006
rect 28390 29004 28396 29006
rect 28460 29004 28466 29068
rect 28809 29066 28875 29069
rect 29686 29066 29746 29142
rect 28809 29064 29746 29066
rect 28809 29008 28814 29064
rect 28870 29008 29746 29064
rect 28809 29006 29746 29008
rect 29821 29066 29887 29069
rect 30230 29066 30236 29068
rect 29821 29064 30236 29066
rect 29821 29008 29826 29064
rect 29882 29008 30236 29064
rect 29821 29006 30236 29008
rect 28809 29003 28875 29006
rect 29821 29003 29887 29006
rect 30230 29004 30236 29006
rect 30300 29004 30306 29068
rect 31710 29066 31770 29142
rect 34053 29068 34119 29069
rect 34053 29066 34100 29068
rect 31710 29064 34100 29066
rect 31710 29008 34058 29064
rect 31710 29006 34100 29008
rect 34053 29004 34100 29006
rect 34164 29004 34170 29068
rect 35382 29004 35388 29068
rect 35452 29066 35458 29068
rect 36169 29066 36235 29069
rect 37365 29068 37431 29069
rect 37365 29066 37412 29068
rect 35452 29064 36235 29066
rect 35452 29008 36174 29064
rect 36230 29008 36235 29064
rect 35452 29006 36235 29008
rect 37320 29064 37412 29066
rect 37320 29008 37370 29064
rect 37320 29006 37412 29008
rect 35452 29004 35458 29006
rect 5165 28930 5231 28933
rect 6269 28930 6335 28933
rect 5165 28928 6335 28930
rect 5165 28872 5170 28928
rect 5226 28872 6274 28928
rect 6330 28872 6335 28928
rect 5165 28870 6335 28872
rect 5165 28867 5231 28870
rect 6269 28867 6335 28870
rect 11973 28930 12039 28933
rect 13448 28930 13508 29003
rect 11973 28928 13508 28930
rect 11973 28872 11978 28928
rect 12034 28872 13508 28928
rect 11973 28870 13508 28872
rect 21817 28930 21883 28933
rect 24485 28930 24551 28933
rect 21817 28928 24551 28930
rect 21817 28872 21822 28928
rect 21878 28872 24490 28928
rect 24546 28872 24551 28928
rect 21817 28870 24551 28872
rect 11973 28867 12039 28870
rect 21817 28867 21883 28870
rect 24485 28867 24551 28870
rect 25313 28930 25379 28933
rect 27286 28930 27292 28932
rect 25313 28928 27292 28930
rect 25313 28872 25318 28928
rect 25374 28872 27292 28928
rect 25313 28870 27292 28872
rect 25313 28867 25379 28870
rect 27286 28868 27292 28870
rect 27356 28868 27362 28932
rect 28625 28930 28691 28933
rect 28582 28928 28691 28930
rect 28582 28872 28630 28928
rect 28686 28872 28691 28928
rect 28582 28867 28691 28872
rect 30238 28930 30298 29004
rect 34053 29003 34119 29004
rect 36169 29003 36235 29006
rect 37365 29004 37412 29006
rect 37476 29004 37482 29068
rect 37365 29003 37431 29004
rect 30238 28870 34714 28930
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 19793 28794 19859 28797
rect 20713 28794 20779 28797
rect 19793 28792 20779 28794
rect 19793 28736 19798 28792
rect 19854 28736 20718 28792
rect 20774 28736 20779 28792
rect 19793 28734 20779 28736
rect 19793 28731 19859 28734
rect 20713 28731 20779 28734
rect 22553 28794 22619 28797
rect 22686 28794 22692 28796
rect 22553 28792 22692 28794
rect 22553 28736 22558 28792
rect 22614 28736 22692 28792
rect 22553 28734 22692 28736
rect 22553 28731 22619 28734
rect 22686 28732 22692 28734
rect 22756 28732 22762 28796
rect 27429 28794 27495 28797
rect 25960 28792 27495 28794
rect 25960 28736 27434 28792
rect 27490 28736 27495 28792
rect 25960 28734 27495 28736
rect 25960 28661 26020 28734
rect 27429 28731 27495 28734
rect 27838 28732 27844 28796
rect 27908 28794 27914 28796
rect 28349 28794 28415 28797
rect 27908 28792 28415 28794
rect 27908 28736 28354 28792
rect 28410 28736 28415 28792
rect 27908 28734 28415 28736
rect 27908 28732 27914 28734
rect 28349 28731 28415 28734
rect 28582 28661 28642 28867
rect 18321 28658 18387 28661
rect 20989 28658 21055 28661
rect 22093 28658 22159 28661
rect 18321 28656 22159 28658
rect 18321 28600 18326 28656
rect 18382 28600 20994 28656
rect 21050 28600 22098 28656
rect 22154 28600 22159 28656
rect 18321 28598 22159 28600
rect 18321 28595 18387 28598
rect 20989 28595 21055 28598
rect 22093 28595 22159 28598
rect 23422 28596 23428 28660
rect 23492 28658 23498 28660
rect 25497 28658 25563 28661
rect 23492 28656 25563 28658
rect 23492 28600 25502 28656
rect 25558 28600 25563 28656
rect 23492 28598 25563 28600
rect 23492 28596 23498 28598
rect 25497 28595 25563 28598
rect 25957 28656 26023 28661
rect 25957 28600 25962 28656
rect 26018 28600 26023 28656
rect 25957 28595 26023 28600
rect 28206 28596 28212 28660
rect 28276 28658 28282 28660
rect 28441 28658 28507 28661
rect 28276 28656 28507 28658
rect 28276 28600 28446 28656
rect 28502 28600 28507 28656
rect 28276 28598 28507 28600
rect 28582 28656 28691 28661
rect 28582 28600 28630 28656
rect 28686 28600 28691 28656
rect 28582 28598 28691 28600
rect 34654 28658 34714 28870
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 36721 28794 36787 28797
rect 36854 28794 36860 28796
rect 36721 28792 36860 28794
rect 36721 28736 36726 28792
rect 36782 28736 36860 28792
rect 36721 28734 36860 28736
rect 36721 28731 36787 28734
rect 36854 28732 36860 28734
rect 36924 28732 36930 28796
rect 38377 28658 38443 28661
rect 34654 28656 38443 28658
rect 34654 28600 38382 28656
rect 38438 28600 38443 28656
rect 34654 28598 38443 28600
rect 28276 28596 28282 28598
rect 28441 28595 28507 28598
rect 28625 28595 28691 28598
rect 38377 28595 38443 28598
rect 10961 28522 11027 28525
rect 12157 28522 12223 28525
rect 10961 28520 12223 28522
rect 10961 28464 10966 28520
rect 11022 28464 12162 28520
rect 12218 28464 12223 28520
rect 10961 28462 12223 28464
rect 10961 28459 11027 28462
rect 12157 28459 12223 28462
rect 12617 28522 12683 28525
rect 14825 28522 14891 28525
rect 12617 28520 14891 28522
rect 12617 28464 12622 28520
rect 12678 28464 14830 28520
rect 14886 28464 14891 28520
rect 12617 28462 14891 28464
rect 12617 28459 12683 28462
rect 14825 28459 14891 28462
rect 19793 28522 19859 28525
rect 20846 28522 20852 28524
rect 19793 28520 20852 28522
rect 19793 28464 19798 28520
rect 19854 28464 20852 28520
rect 19793 28462 20852 28464
rect 19793 28459 19859 28462
rect 20846 28460 20852 28462
rect 20916 28460 20922 28524
rect 20989 28522 21055 28525
rect 23013 28522 23079 28525
rect 23565 28522 23631 28525
rect 20989 28520 21098 28522
rect 20989 28464 20994 28520
rect 21050 28464 21098 28520
rect 20989 28459 21098 28464
rect 23013 28520 23631 28522
rect 23013 28464 23018 28520
rect 23074 28464 23570 28520
rect 23626 28464 23631 28520
rect 23013 28462 23631 28464
rect 23013 28459 23079 28462
rect 23565 28459 23631 28462
rect 23749 28522 23815 28525
rect 24301 28522 24367 28525
rect 27153 28522 27219 28525
rect 29177 28522 29243 28525
rect 23749 28520 24367 28522
rect 23749 28464 23754 28520
rect 23810 28464 24306 28520
rect 24362 28464 24367 28520
rect 23749 28462 24367 28464
rect 23749 28459 23815 28462
rect 24301 28459 24367 28462
rect 26420 28520 29243 28522
rect 26420 28464 27158 28520
rect 27214 28464 29182 28520
rect 29238 28464 29243 28520
rect 26420 28462 29243 28464
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 21038 28250 21098 28459
rect 21541 28386 21607 28389
rect 26141 28386 26207 28389
rect 26420 28386 26480 28462
rect 27153 28459 27219 28462
rect 29177 28459 29243 28462
rect 32121 28522 32187 28525
rect 34278 28522 34284 28524
rect 32121 28520 34284 28522
rect 32121 28464 32126 28520
rect 32182 28464 34284 28520
rect 32121 28462 34284 28464
rect 32121 28459 32187 28462
rect 34278 28460 34284 28462
rect 34348 28522 34354 28524
rect 38193 28522 38259 28525
rect 34348 28520 38259 28522
rect 34348 28464 38198 28520
rect 38254 28464 38259 28520
rect 34348 28462 38259 28464
rect 34348 28460 34354 28462
rect 38193 28459 38259 28462
rect 26693 28388 26759 28389
rect 26693 28386 26740 28388
rect 21541 28384 26480 28386
rect 21541 28328 21546 28384
rect 21602 28328 26146 28384
rect 26202 28328 26480 28384
rect 21541 28326 26480 28328
rect 26652 28384 26740 28386
rect 26804 28386 26810 28388
rect 34605 28386 34671 28389
rect 26804 28384 34671 28386
rect 26652 28328 26698 28384
rect 26804 28328 34610 28384
rect 34666 28328 34671 28384
rect 26652 28326 26740 28328
rect 21541 28323 21607 28326
rect 26141 28323 26207 28326
rect 26693 28324 26740 28326
rect 26804 28326 34671 28328
rect 26804 28324 26810 28326
rect 26693 28323 26759 28324
rect 34605 28323 34671 28326
rect 21449 28250 21515 28253
rect 21038 28248 21515 28250
rect 21038 28192 21454 28248
rect 21510 28192 21515 28248
rect 21038 28190 21515 28192
rect 21449 28187 21515 28190
rect 21725 28250 21791 28253
rect 26877 28250 26943 28253
rect 21725 28248 26943 28250
rect 21725 28192 21730 28248
rect 21786 28192 26882 28248
rect 26938 28192 26943 28248
rect 21725 28190 26943 28192
rect 21725 28187 21791 28190
rect 26877 28187 26943 28190
rect 27705 28250 27771 28253
rect 27981 28250 28047 28253
rect 27705 28248 28047 28250
rect 27705 28192 27710 28248
rect 27766 28192 27986 28248
rect 28042 28192 28047 28248
rect 27705 28190 28047 28192
rect 27705 28187 27771 28190
rect 27981 28187 28047 28190
rect 28257 28248 28323 28253
rect 28257 28192 28262 28248
rect 28318 28192 28323 28248
rect 28257 28187 28323 28192
rect 28809 28250 28875 28253
rect 28942 28250 28948 28252
rect 28809 28248 28948 28250
rect 28809 28192 28814 28248
rect 28870 28192 28948 28248
rect 28809 28190 28948 28192
rect 28809 28187 28875 28190
rect 28942 28188 28948 28190
rect 29012 28188 29018 28252
rect 29453 28250 29519 28253
rect 31334 28250 31340 28252
rect 29453 28248 31340 28250
rect 29453 28192 29458 28248
rect 29514 28192 31340 28248
rect 29453 28190 31340 28192
rect 29453 28187 29519 28190
rect 31334 28188 31340 28190
rect 31404 28250 31410 28252
rect 41137 28250 41203 28253
rect 31404 28248 41203 28250
rect 31404 28192 41142 28248
rect 41198 28192 41203 28248
rect 31404 28190 41203 28192
rect 31404 28188 31410 28190
rect 41137 28187 41203 28190
rect 10961 28114 11027 28117
rect 14181 28114 14247 28117
rect 10961 28112 14247 28114
rect 10961 28056 10966 28112
rect 11022 28056 14186 28112
rect 14242 28056 14247 28112
rect 10961 28054 14247 28056
rect 10961 28051 11027 28054
rect 14181 28051 14247 28054
rect 16941 28114 17007 28117
rect 28260 28114 28320 28187
rect 16941 28112 28320 28114
rect 16941 28056 16946 28112
rect 17002 28056 28320 28112
rect 16941 28054 28320 28056
rect 28533 28114 28599 28117
rect 29085 28114 29151 28117
rect 28533 28112 29151 28114
rect 28533 28056 28538 28112
rect 28594 28056 29090 28112
rect 29146 28056 29151 28112
rect 28533 28054 29151 28056
rect 16941 28051 17007 28054
rect 28533 28051 28599 28054
rect 29085 28051 29151 28054
rect 31710 28054 36186 28114
rect 22185 27978 22251 27981
rect 22318 27978 22324 27980
rect 22185 27976 22324 27978
rect 22185 27920 22190 27976
rect 22246 27920 22324 27976
rect 22185 27918 22324 27920
rect 22185 27915 22251 27918
rect 22318 27916 22324 27918
rect 22388 27916 22394 27980
rect 24025 27978 24091 27981
rect 24894 27978 24900 27980
rect 24025 27976 24900 27978
rect 24025 27920 24030 27976
rect 24086 27920 24900 27976
rect 24025 27918 24900 27920
rect 24025 27915 24091 27918
rect 24894 27916 24900 27918
rect 24964 27916 24970 27980
rect 26601 27978 26667 27981
rect 31710 27978 31770 28054
rect 26601 27976 31770 27978
rect 26601 27920 26606 27976
rect 26662 27920 31770 27976
rect 26601 27918 31770 27920
rect 34697 27978 34763 27981
rect 35893 27978 35959 27981
rect 34697 27976 35959 27978
rect 34697 27920 34702 27976
rect 34758 27920 35898 27976
rect 35954 27920 35959 27976
rect 34697 27918 35959 27920
rect 36126 27978 36186 28054
rect 40401 27978 40467 27981
rect 36126 27976 40467 27978
rect 36126 27920 40406 27976
rect 40462 27920 40467 27976
rect 36126 27918 40467 27920
rect 26601 27915 26667 27918
rect 34697 27915 34763 27918
rect 35893 27915 35959 27918
rect 40401 27915 40467 27918
rect 20846 27780 20852 27844
rect 20916 27842 20922 27844
rect 24710 27842 24716 27844
rect 20916 27782 24716 27842
rect 20916 27780 20922 27782
rect 24710 27780 24716 27782
rect 24780 27780 24786 27844
rect 31385 27842 31451 27845
rect 31661 27842 31727 27845
rect 25316 27840 31727 27842
rect 25316 27784 31390 27840
rect 31446 27784 31666 27840
rect 31722 27784 31727 27840
rect 25316 27782 31727 27784
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 25316 27709 25376 27782
rect 31385 27779 31451 27782
rect 31661 27779 31727 27782
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19374 27644 19380 27708
rect 19444 27706 19450 27708
rect 19977 27706 20043 27709
rect 20805 27708 20871 27709
rect 20805 27706 20852 27708
rect 19444 27704 20043 27706
rect 19444 27648 19982 27704
rect 20038 27648 20043 27704
rect 19444 27646 20043 27648
rect 20760 27704 20852 27706
rect 20760 27648 20810 27704
rect 20760 27646 20852 27648
rect 19444 27644 19450 27646
rect 19977 27643 20043 27646
rect 20805 27644 20852 27646
rect 20916 27644 20922 27708
rect 21449 27706 21515 27709
rect 25313 27706 25379 27709
rect 21449 27704 25379 27706
rect 21449 27648 21454 27704
rect 21510 27648 25318 27704
rect 25374 27648 25379 27704
rect 21449 27646 25379 27648
rect 20805 27643 20871 27644
rect 21449 27643 21515 27646
rect 25313 27643 25379 27646
rect 26366 27644 26372 27708
rect 26436 27706 26442 27708
rect 26877 27706 26943 27709
rect 26436 27704 26943 27706
rect 26436 27648 26882 27704
rect 26938 27648 26943 27704
rect 26436 27646 26943 27648
rect 26436 27644 26442 27646
rect 26877 27643 26943 27646
rect 28022 27644 28028 27708
rect 28092 27706 28098 27708
rect 28165 27706 28231 27709
rect 28092 27704 28231 27706
rect 28092 27648 28170 27704
rect 28226 27648 28231 27704
rect 28092 27646 28231 27648
rect 28092 27644 28098 27646
rect 28165 27643 28231 27646
rect 28993 27706 29059 27709
rect 29126 27706 29132 27708
rect 28993 27704 29132 27706
rect 28993 27648 28998 27704
rect 29054 27648 29132 27704
rect 28993 27646 29132 27648
rect 28993 27643 29059 27646
rect 29126 27644 29132 27646
rect 29196 27644 29202 27708
rect 30925 27706 30991 27709
rect 33777 27706 33843 27709
rect 30925 27704 33843 27706
rect 30925 27648 30930 27704
rect 30986 27648 33782 27704
rect 33838 27648 33843 27704
rect 30925 27646 33843 27648
rect 30925 27643 30991 27646
rect 33777 27643 33843 27646
rect 34462 27644 34468 27708
rect 34532 27706 34538 27708
rect 34605 27706 34671 27709
rect 34532 27704 34671 27706
rect 34532 27648 34610 27704
rect 34666 27648 34671 27704
rect 34532 27646 34671 27648
rect 34532 27644 34538 27646
rect 34605 27643 34671 27646
rect 38377 27706 38443 27709
rect 39062 27706 39068 27708
rect 38377 27704 39068 27706
rect 38377 27648 38382 27704
rect 38438 27648 39068 27704
rect 38377 27646 39068 27648
rect 38377 27643 38443 27646
rect 39062 27644 39068 27646
rect 39132 27644 39138 27708
rect 8385 27570 8451 27573
rect 8753 27570 8819 27573
rect 8385 27568 8819 27570
rect 8385 27512 8390 27568
rect 8446 27512 8758 27568
rect 8814 27512 8819 27568
rect 8385 27510 8819 27512
rect 8385 27507 8451 27510
rect 8753 27507 8819 27510
rect 9213 27570 9279 27573
rect 10685 27570 10751 27573
rect 16481 27570 16547 27573
rect 9213 27568 22110 27570
rect 9213 27512 9218 27568
rect 9274 27512 10690 27568
rect 10746 27512 16486 27568
rect 16542 27512 22110 27568
rect 9213 27510 22110 27512
rect 9213 27507 9279 27510
rect 10685 27507 10751 27510
rect 16481 27507 16547 27510
rect 8845 27434 8911 27437
rect 10910 27434 10916 27436
rect 8845 27432 10916 27434
rect 8845 27376 8850 27432
rect 8906 27376 10916 27432
rect 8845 27374 10916 27376
rect 8845 27371 8911 27374
rect 10910 27372 10916 27374
rect 10980 27372 10986 27436
rect 22050 27434 22110 27510
rect 24342 27508 24348 27572
rect 24412 27570 24418 27572
rect 24761 27570 24827 27573
rect 24412 27568 24827 27570
rect 24412 27512 24766 27568
rect 24822 27512 24827 27568
rect 24412 27510 24827 27512
rect 24412 27508 24418 27510
rect 24761 27507 24827 27510
rect 27981 27570 28047 27573
rect 30966 27570 30972 27572
rect 27981 27568 30972 27570
rect 27981 27512 27986 27568
rect 28042 27512 30972 27568
rect 27981 27510 30972 27512
rect 27981 27507 28047 27510
rect 30966 27508 30972 27510
rect 31036 27570 31042 27572
rect 32121 27570 32187 27573
rect 31036 27568 32187 27570
rect 31036 27512 32126 27568
rect 32182 27512 32187 27568
rect 31036 27510 32187 27512
rect 31036 27508 31042 27510
rect 32121 27507 32187 27510
rect 29453 27434 29519 27437
rect 22050 27432 29519 27434
rect 22050 27376 29458 27432
rect 29514 27376 29519 27432
rect 22050 27374 29519 27376
rect 29453 27371 29519 27374
rect 30833 27434 30899 27437
rect 32765 27434 32831 27437
rect 30833 27432 32831 27434
rect 30833 27376 30838 27432
rect 30894 27376 32770 27432
rect 32826 27376 32831 27432
rect 30833 27374 32831 27376
rect 30833 27371 30899 27374
rect 32765 27371 32831 27374
rect 33409 27434 33475 27437
rect 35065 27434 35131 27437
rect 33409 27432 35131 27434
rect 33409 27376 33414 27432
rect 33470 27376 35070 27432
rect 35126 27376 35131 27432
rect 33409 27374 35131 27376
rect 33409 27371 33475 27374
rect 35065 27371 35131 27374
rect 0 27298 800 27328
rect 4061 27298 4127 27301
rect 0 27296 4127 27298
rect 0 27240 4066 27296
rect 4122 27240 4127 27296
rect 0 27238 4127 27240
rect 0 27208 800 27238
rect 4061 27235 4127 27238
rect 8569 27298 8635 27301
rect 10317 27298 10383 27301
rect 8569 27296 10383 27298
rect 8569 27240 8574 27296
rect 8630 27240 10322 27296
rect 10378 27240 10383 27296
rect 8569 27238 10383 27240
rect 8569 27235 8635 27238
rect 10317 27235 10383 27238
rect 21909 27300 21975 27301
rect 21909 27296 21956 27300
rect 22020 27298 22026 27300
rect 33409 27298 33475 27301
rect 34421 27298 34487 27301
rect 21909 27240 21914 27296
rect 21909 27236 21956 27240
rect 22020 27238 22066 27298
rect 33409 27296 34487 27298
rect 33409 27240 33414 27296
rect 33470 27240 34426 27296
rect 34482 27240 34487 27296
rect 33409 27238 34487 27240
rect 22020 27236 22026 27238
rect 21909 27235 21975 27236
rect 33409 27235 33475 27238
rect 34421 27235 34487 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 9765 27164 9831 27165
rect 12525 27164 12591 27165
rect 9765 27162 9812 27164
rect 9720 27160 9812 27162
rect 9720 27104 9770 27160
rect 9720 27102 9812 27104
rect 9765 27100 9812 27102
rect 9876 27100 9882 27164
rect 12525 27162 12572 27164
rect 12484 27160 12572 27162
rect 12636 27162 12642 27164
rect 13670 27162 13676 27164
rect 12484 27104 12530 27160
rect 12484 27102 12572 27104
rect 12525 27100 12572 27102
rect 12636 27102 13676 27162
rect 12636 27100 12642 27102
rect 13670 27100 13676 27102
rect 13740 27100 13746 27164
rect 14917 27162 14983 27165
rect 15929 27162 15995 27165
rect 16297 27164 16363 27165
rect 16246 27162 16252 27164
rect 14917 27160 15995 27162
rect 14917 27104 14922 27160
rect 14978 27104 15934 27160
rect 15990 27104 15995 27160
rect 14917 27102 15995 27104
rect 16206 27102 16252 27162
rect 16316 27160 16363 27164
rect 16358 27104 16363 27160
rect 9765 27099 9831 27100
rect 12525 27099 12591 27100
rect 14917 27099 14983 27102
rect 15929 27099 15995 27102
rect 16246 27100 16252 27102
rect 16316 27100 16363 27104
rect 16297 27099 16363 27100
rect 31017 27162 31083 27165
rect 35934 27162 35940 27164
rect 31017 27160 35940 27162
rect 31017 27104 31022 27160
rect 31078 27104 35940 27160
rect 31017 27102 35940 27104
rect 31017 27099 31083 27102
rect 35934 27100 35940 27102
rect 36004 27162 36010 27164
rect 39246 27162 39252 27164
rect 36004 27102 39252 27162
rect 36004 27100 36010 27102
rect 39246 27100 39252 27102
rect 39316 27100 39322 27164
rect 9489 27026 9555 27029
rect 10041 27026 10107 27029
rect 9489 27024 10107 27026
rect 9489 26968 9494 27024
rect 9550 26968 10046 27024
rect 10102 26968 10107 27024
rect 9489 26966 10107 26968
rect 9489 26963 9555 26966
rect 10041 26963 10107 26966
rect 12065 27026 12131 27029
rect 13169 27026 13235 27029
rect 15377 27026 15443 27029
rect 12065 27024 15443 27026
rect 12065 26968 12070 27024
rect 12126 26968 13174 27024
rect 13230 26968 15382 27024
rect 15438 26968 15443 27024
rect 12065 26966 15443 26968
rect 12065 26963 12131 26966
rect 13169 26963 13235 26966
rect 15377 26963 15443 26966
rect 7925 26890 7991 26893
rect 16665 26890 16731 26893
rect 7925 26888 16731 26890
rect 7925 26832 7930 26888
rect 7986 26832 16670 26888
rect 16726 26832 16731 26888
rect 7925 26830 16731 26832
rect 7925 26827 7991 26830
rect 16665 26827 16731 26830
rect 22185 26890 22251 26893
rect 23105 26890 23171 26893
rect 33501 26890 33567 26893
rect 22185 26888 33567 26890
rect 22185 26832 22190 26888
rect 22246 26832 23110 26888
rect 23166 26832 33506 26888
rect 33562 26832 33567 26888
rect 22185 26830 33567 26832
rect 22185 26827 22251 26830
rect 23105 26827 23171 26830
rect 33501 26827 33567 26830
rect 9121 26756 9187 26757
rect 9070 26692 9076 26756
rect 9140 26754 9187 26756
rect 13721 26754 13787 26757
rect 15878 26754 15884 26756
rect 9140 26752 9232 26754
rect 9182 26696 9232 26752
rect 9140 26694 9232 26696
rect 13721 26752 15884 26754
rect 13721 26696 13726 26752
rect 13782 26696 15884 26752
rect 13721 26694 15884 26696
rect 9140 26692 9187 26694
rect 9121 26691 9187 26692
rect 13721 26691 13787 26694
rect 15878 26692 15884 26694
rect 15948 26692 15954 26756
rect 21725 26754 21791 26757
rect 24577 26754 24643 26757
rect 21725 26752 24643 26754
rect 21725 26696 21730 26752
rect 21786 26696 24582 26752
rect 24638 26696 24643 26752
rect 21725 26694 24643 26696
rect 21725 26691 21791 26694
rect 24577 26691 24643 26694
rect 26182 26692 26188 26756
rect 26252 26754 26258 26756
rect 32029 26754 32095 26757
rect 26252 26752 32095 26754
rect 26252 26696 32034 26752
rect 32090 26696 32095 26752
rect 26252 26694 32095 26696
rect 26252 26692 26258 26694
rect 32029 26691 32095 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19190 26556 19196 26620
rect 19260 26618 19266 26620
rect 30005 26618 30071 26621
rect 19260 26616 30071 26618
rect 19260 26560 30010 26616
rect 30066 26560 30071 26616
rect 19260 26558 30071 26560
rect 19260 26556 19266 26558
rect 30005 26555 30071 26558
rect 25037 26482 25103 26485
rect 25262 26482 25268 26484
rect 25037 26480 25268 26482
rect 25037 26424 25042 26480
rect 25098 26424 25268 26480
rect 25037 26422 25268 26424
rect 25037 26419 25103 26422
rect 25262 26420 25268 26422
rect 25332 26420 25338 26484
rect 10317 26348 10383 26349
rect 11421 26348 11487 26349
rect 10317 26344 10364 26348
rect 10428 26346 10434 26348
rect 10317 26288 10322 26344
rect 10317 26284 10364 26288
rect 10428 26286 10474 26346
rect 11421 26344 11468 26348
rect 11532 26346 11538 26348
rect 16297 26346 16363 26349
rect 16430 26346 16436 26348
rect 11421 26288 11426 26344
rect 10428 26284 10434 26286
rect 11421 26284 11468 26288
rect 11532 26286 11578 26346
rect 16297 26344 16436 26346
rect 16297 26288 16302 26344
rect 16358 26288 16436 26344
rect 16297 26286 16436 26288
rect 11532 26284 11538 26286
rect 10317 26283 10383 26284
rect 11421 26283 11487 26284
rect 16297 26283 16363 26286
rect 16430 26284 16436 26286
rect 16500 26284 16506 26348
rect 21541 26346 21607 26349
rect 23381 26346 23447 26349
rect 21541 26344 23447 26346
rect 21541 26288 21546 26344
rect 21602 26288 23386 26344
rect 23442 26288 23447 26344
rect 21541 26286 23447 26288
rect 21541 26283 21607 26286
rect 23381 26283 23447 26286
rect 23657 26346 23723 26349
rect 25589 26346 25655 26349
rect 29453 26348 29519 26349
rect 34421 26348 34487 26349
rect 29453 26346 29500 26348
rect 23657 26344 25655 26346
rect 23657 26288 23662 26344
rect 23718 26288 25594 26344
rect 25650 26288 25655 26344
rect 23657 26286 25655 26288
rect 29408 26344 29500 26346
rect 29408 26288 29458 26344
rect 29408 26286 29500 26288
rect 23657 26283 23723 26286
rect 25589 26283 25655 26286
rect 29453 26284 29500 26286
rect 29564 26284 29570 26348
rect 34421 26346 34468 26348
rect 34376 26344 34468 26346
rect 34376 26288 34426 26344
rect 34376 26286 34468 26288
rect 34421 26284 34468 26286
rect 34532 26284 34538 26348
rect 35525 26346 35591 26349
rect 35750 26346 35756 26348
rect 35525 26344 35756 26346
rect 35525 26288 35530 26344
rect 35586 26288 35756 26344
rect 35525 26286 35756 26288
rect 29453 26283 29519 26284
rect 34421 26283 34487 26284
rect 35525 26283 35591 26286
rect 35750 26284 35756 26286
rect 35820 26284 35826 26348
rect 27981 26212 28047 26213
rect 27981 26208 28028 26212
rect 28092 26210 28098 26212
rect 31201 26210 31267 26213
rect 31518 26210 31524 26212
rect 27981 26152 27986 26208
rect 27981 26148 28028 26152
rect 28092 26150 28138 26210
rect 31201 26208 31524 26210
rect 31201 26152 31206 26208
rect 31262 26152 31524 26208
rect 31201 26150 31524 26152
rect 28092 26148 28098 26150
rect 27981 26147 28047 26148
rect 31201 26147 31267 26150
rect 31518 26148 31524 26150
rect 31588 26148 31594 26212
rect 34646 26148 34652 26212
rect 34716 26210 34722 26212
rect 35065 26210 35131 26213
rect 34716 26208 35131 26210
rect 34716 26152 35070 26208
rect 35126 26152 35131 26208
rect 34716 26150 35131 26152
rect 34716 26148 34722 26150
rect 35065 26147 35131 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 20989 25938 21055 25941
rect 26969 25938 27035 25941
rect 20989 25936 27035 25938
rect 20989 25880 20994 25936
rect 21050 25880 26974 25936
rect 27030 25880 27035 25936
rect 20989 25878 27035 25880
rect 20989 25875 21055 25878
rect 26969 25875 27035 25878
rect 9121 25802 9187 25805
rect 9121 25800 12450 25802
rect 9121 25744 9126 25800
rect 9182 25744 12450 25800
rect 9121 25742 12450 25744
rect 9121 25739 9187 25742
rect 12390 25666 12450 25742
rect 14774 25740 14780 25804
rect 14844 25802 14850 25804
rect 30373 25802 30439 25805
rect 14844 25800 30439 25802
rect 14844 25744 30378 25800
rect 30434 25744 30439 25800
rect 14844 25742 30439 25744
rect 14844 25740 14850 25742
rect 30373 25739 30439 25742
rect 33593 25802 33659 25805
rect 36077 25802 36143 25805
rect 33593 25800 36143 25802
rect 33593 25744 33598 25800
rect 33654 25744 36082 25800
rect 36138 25744 36143 25800
rect 33593 25742 36143 25744
rect 33593 25739 33659 25742
rect 36077 25739 36143 25742
rect 20294 25666 20300 25668
rect 12390 25606 20300 25666
rect 20294 25604 20300 25606
rect 20364 25666 20370 25668
rect 21541 25666 21607 25669
rect 20364 25664 21607 25666
rect 20364 25608 21546 25664
rect 21602 25608 21607 25664
rect 20364 25606 21607 25608
rect 20364 25604 20370 25606
rect 21541 25603 21607 25606
rect 28206 25604 28212 25668
rect 28276 25666 28282 25668
rect 28809 25666 28875 25669
rect 28276 25664 28875 25666
rect 28276 25608 28814 25664
rect 28870 25608 28875 25664
rect 28276 25606 28875 25608
rect 28276 25604 28282 25606
rect 28809 25603 28875 25606
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 21541 25530 21607 25533
rect 21817 25530 21883 25533
rect 21541 25528 21883 25530
rect 21541 25472 21546 25528
rect 21602 25472 21822 25528
rect 21878 25472 21883 25528
rect 21541 25470 21883 25472
rect 21541 25467 21607 25470
rect 21817 25467 21883 25470
rect 32581 25394 32647 25397
rect 32949 25394 33015 25397
rect 32581 25392 33015 25394
rect 32581 25336 32586 25392
rect 32642 25336 32954 25392
rect 33010 25336 33015 25392
rect 32581 25334 33015 25336
rect 32581 25331 32647 25334
rect 32949 25331 33015 25334
rect 34278 25332 34284 25396
rect 34348 25394 34354 25396
rect 34421 25394 34487 25397
rect 34348 25392 34487 25394
rect 34348 25336 34426 25392
rect 34482 25336 34487 25392
rect 34348 25334 34487 25336
rect 34348 25332 34354 25334
rect 34421 25331 34487 25334
rect 37590 25332 37596 25396
rect 37660 25394 37666 25396
rect 37733 25394 37799 25397
rect 37660 25392 37799 25394
rect 37660 25336 37738 25392
rect 37794 25336 37799 25392
rect 37660 25334 37799 25336
rect 37660 25332 37666 25334
rect 37733 25331 37799 25334
rect 9806 25196 9812 25260
rect 9876 25258 9882 25260
rect 10685 25258 10751 25261
rect 9876 25256 10751 25258
rect 9876 25200 10690 25256
rect 10746 25200 10751 25256
rect 9876 25198 10751 25200
rect 9876 25196 9882 25198
rect 10685 25195 10751 25198
rect 18270 25196 18276 25260
rect 18340 25258 18346 25260
rect 33593 25258 33659 25261
rect 18340 25256 33659 25258
rect 18340 25200 33598 25256
rect 33654 25200 33659 25256
rect 18340 25198 33659 25200
rect 18340 25196 18346 25198
rect 33593 25195 33659 25198
rect 34237 25258 34303 25261
rect 41749 25258 42549 25288
rect 34237 25256 42549 25258
rect 34237 25200 34242 25256
rect 34298 25200 42549 25256
rect 34237 25198 42549 25200
rect 34237 25195 34303 25198
rect 41749 25168 42549 25198
rect 21173 25124 21239 25125
rect 22001 25124 22067 25125
rect 21173 25122 21220 25124
rect 21128 25120 21220 25122
rect 21128 25064 21178 25120
rect 21128 25062 21220 25064
rect 21173 25060 21220 25062
rect 21284 25060 21290 25124
rect 21950 25060 21956 25124
rect 22020 25122 22067 25124
rect 22020 25120 22112 25122
rect 22062 25064 22112 25120
rect 22020 25062 22112 25064
rect 22020 25060 22067 25062
rect 24526 25060 24532 25124
rect 24596 25122 24602 25124
rect 29862 25122 29868 25124
rect 24596 25062 29868 25122
rect 24596 25060 24602 25062
rect 29862 25060 29868 25062
rect 29932 25122 29938 25124
rect 30005 25122 30071 25125
rect 33409 25124 33475 25125
rect 29932 25120 30071 25122
rect 29932 25064 30010 25120
rect 30066 25064 30071 25120
rect 29932 25062 30071 25064
rect 29932 25060 29938 25062
rect 21173 25059 21239 25060
rect 22001 25059 22067 25060
rect 30005 25059 30071 25062
rect 33358 25060 33364 25124
rect 33428 25122 33475 25124
rect 33428 25120 33520 25122
rect 33470 25064 33520 25120
rect 33428 25062 33520 25064
rect 33428 25060 33475 25062
rect 33409 25059 33475 25060
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 9213 24988 9279 24989
rect 9213 24986 9260 24988
rect 9168 24984 9260 24986
rect 9168 24928 9218 24984
rect 9168 24926 9260 24928
rect 9213 24924 9260 24926
rect 9324 24924 9330 24988
rect 11605 24986 11671 24989
rect 13854 24986 13860 24988
rect 11605 24984 13860 24986
rect 11605 24928 11610 24984
rect 11666 24928 13860 24984
rect 11605 24926 13860 24928
rect 9213 24923 9279 24924
rect 11605 24923 11671 24926
rect 13854 24924 13860 24926
rect 13924 24924 13930 24988
rect 24894 24924 24900 24988
rect 24964 24986 24970 24988
rect 25129 24986 25195 24989
rect 37089 24988 37155 24989
rect 37038 24986 37044 24988
rect 24964 24984 25195 24986
rect 24964 24928 25134 24984
rect 25190 24928 25195 24984
rect 24964 24926 25195 24928
rect 36998 24926 37044 24986
rect 37108 24984 37155 24988
rect 37150 24928 37155 24984
rect 24964 24924 24970 24926
rect 25129 24923 25195 24926
rect 37038 24924 37044 24926
rect 37108 24924 37155 24928
rect 37089 24923 37155 24924
rect 5073 24850 5139 24853
rect 5533 24850 5599 24853
rect 8201 24850 8267 24853
rect 5073 24848 8267 24850
rect 5073 24792 5078 24848
rect 5134 24792 5538 24848
rect 5594 24792 8206 24848
rect 8262 24792 8267 24848
rect 5073 24790 8267 24792
rect 5073 24787 5139 24790
rect 5533 24787 5599 24790
rect 8201 24787 8267 24790
rect 4981 24714 5047 24717
rect 5257 24714 5323 24717
rect 5901 24714 5967 24717
rect 9213 24714 9279 24717
rect 4981 24712 9279 24714
rect 4981 24656 4986 24712
rect 5042 24656 5262 24712
rect 5318 24656 5906 24712
rect 5962 24656 9218 24712
rect 9274 24656 9279 24712
rect 4981 24654 9279 24656
rect 4981 24651 5047 24654
rect 5257 24651 5323 24654
rect 5901 24651 5967 24654
rect 9213 24651 9279 24654
rect 14457 24714 14523 24717
rect 16481 24714 16547 24717
rect 33317 24714 33383 24717
rect 34145 24714 34211 24717
rect 34697 24714 34763 24717
rect 14457 24712 33383 24714
rect 14457 24656 14462 24712
rect 14518 24656 16486 24712
rect 16542 24656 33322 24712
rect 33378 24656 33383 24712
rect 14457 24654 33383 24656
rect 14457 24651 14523 24654
rect 16481 24651 16547 24654
rect 33317 24651 33383 24654
rect 34102 24712 34211 24714
rect 34102 24656 34150 24712
rect 34206 24656 34211 24712
rect 34102 24651 34211 24656
rect 34654 24712 34763 24714
rect 34654 24656 34702 24712
rect 34758 24656 34763 24712
rect 34654 24651 34763 24656
rect 12985 24580 13051 24581
rect 12934 24516 12940 24580
rect 13004 24578 13051 24580
rect 32949 24578 33015 24581
rect 33869 24578 33935 24581
rect 13004 24576 13096 24578
rect 13046 24520 13096 24576
rect 13004 24518 13096 24520
rect 32949 24576 33935 24578
rect 32949 24520 32954 24576
rect 33010 24520 33874 24576
rect 33930 24520 33935 24576
rect 32949 24518 33935 24520
rect 13004 24516 13051 24518
rect 12985 24515 13051 24516
rect 32949 24515 33015 24518
rect 33869 24515 33935 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 12801 24442 12867 24445
rect 14457 24442 14523 24445
rect 12801 24440 14523 24442
rect 12801 24384 12806 24440
rect 12862 24384 14462 24440
rect 14518 24384 14523 24440
rect 12801 24382 14523 24384
rect 12801 24379 12867 24382
rect 14457 24379 14523 24382
rect 19701 24442 19767 24445
rect 23657 24442 23723 24445
rect 19701 24440 23723 24442
rect 19701 24384 19706 24440
rect 19762 24384 23662 24440
rect 23718 24384 23723 24440
rect 19701 24382 23723 24384
rect 19701 24379 19767 24382
rect 23657 24379 23723 24382
rect 30046 24380 30052 24444
rect 30116 24442 30122 24444
rect 30373 24442 30439 24445
rect 30116 24440 30439 24442
rect 30116 24384 30378 24440
rect 30434 24384 30439 24440
rect 30116 24382 30439 24384
rect 30116 24380 30122 24382
rect 30373 24379 30439 24382
rect 30557 24444 30623 24445
rect 30557 24440 30604 24444
rect 30668 24442 30674 24444
rect 30557 24384 30562 24440
rect 30557 24380 30604 24384
rect 30668 24382 30714 24442
rect 30668 24380 30674 24382
rect 30557 24379 30623 24380
rect 12525 24306 12591 24309
rect 14181 24306 14247 24309
rect 12525 24304 14247 24306
rect 12525 24248 12530 24304
rect 12586 24248 14186 24304
rect 14242 24248 14247 24304
rect 12525 24246 14247 24248
rect 12525 24243 12591 24246
rect 14181 24243 14247 24246
rect 20478 24244 20484 24308
rect 20548 24306 20554 24308
rect 23289 24306 23355 24309
rect 20548 24304 23355 24306
rect 20548 24248 23294 24304
rect 23350 24248 23355 24304
rect 20548 24246 23355 24248
rect 20548 24244 20554 24246
rect 23289 24243 23355 24246
rect 26233 24306 26299 24309
rect 28441 24306 28507 24309
rect 26233 24304 28507 24306
rect 26233 24248 26238 24304
rect 26294 24248 28446 24304
rect 28502 24248 28507 24304
rect 26233 24246 28507 24248
rect 26233 24243 26299 24246
rect 28441 24243 28507 24246
rect 30005 24306 30071 24309
rect 30598 24306 30604 24308
rect 30005 24304 30604 24306
rect 30005 24248 30010 24304
rect 30066 24248 30604 24304
rect 30005 24246 30604 24248
rect 30005 24243 30071 24246
rect 30598 24244 30604 24246
rect 30668 24244 30674 24308
rect 6453 24170 6519 24173
rect 9489 24170 9555 24173
rect 6453 24168 9555 24170
rect 6453 24112 6458 24168
rect 6514 24112 9494 24168
rect 9550 24112 9555 24168
rect 6453 24110 9555 24112
rect 6453 24107 6519 24110
rect 9489 24107 9555 24110
rect 16481 24170 16547 24173
rect 22737 24170 22803 24173
rect 16481 24168 22803 24170
rect 16481 24112 16486 24168
rect 16542 24112 22742 24168
rect 22798 24112 22803 24168
rect 16481 24110 22803 24112
rect 16481 24107 16547 24110
rect 22737 24107 22803 24110
rect 26969 24170 27035 24173
rect 27102 24170 27108 24172
rect 26969 24168 27108 24170
rect 26969 24112 26974 24168
rect 27030 24112 27108 24168
rect 26969 24110 27108 24112
rect 26969 24107 27035 24110
rect 27102 24108 27108 24110
rect 27172 24170 27178 24172
rect 29269 24170 29335 24173
rect 27172 24168 29335 24170
rect 27172 24112 29274 24168
rect 29330 24112 29335 24168
rect 27172 24110 29335 24112
rect 27172 24108 27178 24110
rect 29269 24107 29335 24110
rect 29453 24170 29519 24173
rect 30230 24170 30236 24172
rect 29453 24168 30236 24170
rect 29453 24112 29458 24168
rect 29514 24112 30236 24168
rect 29453 24110 30236 24112
rect 29453 24107 29519 24110
rect 30230 24108 30236 24110
rect 30300 24108 30306 24172
rect 33317 24170 33383 24173
rect 34102 24170 34162 24651
rect 34654 24442 34714 24651
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 34789 24442 34855 24445
rect 34654 24440 34855 24442
rect 34654 24384 34794 24440
rect 34850 24384 34855 24440
rect 34654 24382 34855 24384
rect 34789 24379 34855 24382
rect 33317 24168 34162 24170
rect 33317 24112 33322 24168
rect 33378 24112 34162 24168
rect 33317 24110 34162 24112
rect 33317 24107 33383 24110
rect 15837 24034 15903 24037
rect 17401 24034 17467 24037
rect 18413 24034 18479 24037
rect 15837 24032 18479 24034
rect 15837 23976 15842 24032
rect 15898 23976 17406 24032
rect 17462 23976 18418 24032
rect 18474 23976 18479 24032
rect 15837 23974 18479 23976
rect 15837 23971 15903 23974
rect 17401 23971 17467 23974
rect 18413 23971 18479 23974
rect 25037 24034 25103 24037
rect 25957 24034 26023 24037
rect 26550 24034 26556 24036
rect 25037 24032 26556 24034
rect 25037 23976 25042 24032
rect 25098 23976 25962 24032
rect 26018 23976 26556 24032
rect 25037 23974 26556 23976
rect 25037 23971 25103 23974
rect 25957 23971 26023 23974
rect 26550 23972 26556 23974
rect 26620 23972 26626 24036
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 23841 23898 23907 23901
rect 28073 23898 28139 23901
rect 23841 23896 28139 23898
rect 23841 23840 23846 23896
rect 23902 23840 28078 23896
rect 28134 23840 28139 23896
rect 23841 23838 28139 23840
rect 23841 23835 23907 23838
rect 28073 23835 28139 23838
rect 32857 23898 32923 23901
rect 37590 23898 37596 23900
rect 32857 23896 37596 23898
rect 32857 23840 32862 23896
rect 32918 23840 37596 23896
rect 32857 23838 37596 23840
rect 32857 23835 32923 23838
rect 37590 23836 37596 23838
rect 37660 23836 37666 23900
rect 22461 23762 22527 23765
rect 22829 23762 22895 23765
rect 22461 23760 22895 23762
rect 22461 23704 22466 23760
rect 22522 23704 22834 23760
rect 22890 23704 22895 23760
rect 22461 23702 22895 23704
rect 22461 23699 22527 23702
rect 22829 23699 22895 23702
rect 24669 23762 24735 23765
rect 25814 23762 25820 23764
rect 24669 23760 25820 23762
rect 24669 23704 24674 23760
rect 24730 23704 25820 23760
rect 24669 23702 25820 23704
rect 24669 23699 24735 23702
rect 25814 23700 25820 23702
rect 25884 23762 25890 23764
rect 34513 23762 34579 23765
rect 25884 23760 34579 23762
rect 25884 23704 34518 23760
rect 34574 23704 34579 23760
rect 25884 23702 34579 23704
rect 25884 23700 25890 23702
rect 34513 23699 34579 23702
rect 18638 23564 18644 23628
rect 18708 23626 18714 23628
rect 20253 23626 20319 23629
rect 18708 23624 20319 23626
rect 18708 23568 20258 23624
rect 20314 23568 20319 23624
rect 18708 23566 20319 23568
rect 18708 23564 18714 23566
rect 20253 23563 20319 23566
rect 20713 23626 20779 23629
rect 23473 23626 23539 23629
rect 20713 23624 23539 23626
rect 20713 23568 20718 23624
rect 20774 23568 23478 23624
rect 23534 23568 23539 23624
rect 20713 23566 23539 23568
rect 20713 23563 20779 23566
rect 23473 23563 23539 23566
rect 23657 23626 23723 23629
rect 23790 23626 23796 23628
rect 23657 23624 23796 23626
rect 23657 23568 23662 23624
rect 23718 23568 23796 23624
rect 23657 23566 23796 23568
rect 23657 23563 23723 23566
rect 23790 23564 23796 23566
rect 23860 23564 23866 23628
rect 24577 23626 24643 23629
rect 25078 23626 25084 23628
rect 24577 23624 25084 23626
rect 24577 23568 24582 23624
rect 24638 23568 25084 23624
rect 24577 23566 25084 23568
rect 24577 23563 24643 23566
rect 25078 23564 25084 23566
rect 25148 23564 25154 23628
rect 26049 23626 26115 23629
rect 26734 23626 26740 23628
rect 26049 23624 26740 23626
rect 26049 23568 26054 23624
rect 26110 23568 26740 23624
rect 26049 23566 26740 23568
rect 26049 23563 26115 23566
rect 26734 23564 26740 23566
rect 26804 23564 26810 23628
rect 31201 23626 31267 23629
rect 31518 23626 31524 23628
rect 31201 23624 31524 23626
rect 31201 23568 31206 23624
rect 31262 23568 31524 23624
rect 31201 23566 31524 23568
rect 31201 23563 31267 23566
rect 31518 23564 31524 23566
rect 31588 23626 31594 23628
rect 32305 23626 32371 23629
rect 31588 23624 32371 23626
rect 31588 23568 32310 23624
rect 32366 23568 32371 23624
rect 31588 23566 32371 23568
rect 31588 23564 31594 23566
rect 32305 23563 32371 23566
rect 11697 23490 11763 23493
rect 12525 23492 12591 23493
rect 11830 23490 11836 23492
rect 11697 23488 11836 23490
rect 11697 23432 11702 23488
rect 11758 23432 11836 23488
rect 11697 23430 11836 23432
rect 11697 23427 11763 23430
rect 11830 23428 11836 23430
rect 11900 23428 11906 23492
rect 12525 23490 12572 23492
rect 12480 23488 12572 23490
rect 12480 23432 12530 23488
rect 12480 23430 12572 23432
rect 12525 23428 12572 23430
rect 12636 23428 12642 23492
rect 23565 23490 23631 23493
rect 25630 23490 25636 23492
rect 23565 23488 25636 23490
rect 23565 23432 23570 23488
rect 23626 23432 25636 23488
rect 23565 23430 25636 23432
rect 12525 23427 12591 23428
rect 23565 23427 23631 23430
rect 25630 23428 25636 23430
rect 25700 23428 25706 23492
rect 26693 23490 26759 23493
rect 28533 23492 28599 23493
rect 26918 23490 26924 23492
rect 26693 23488 26924 23490
rect 26693 23432 26698 23488
rect 26754 23432 26924 23488
rect 26693 23430 26924 23432
rect 26693 23427 26759 23430
rect 26918 23428 26924 23430
rect 26988 23428 26994 23492
rect 28533 23490 28580 23492
rect 28488 23488 28580 23490
rect 28488 23432 28538 23488
rect 28488 23430 28580 23432
rect 28533 23428 28580 23430
rect 28644 23428 28650 23492
rect 37222 23428 37228 23492
rect 37292 23490 37298 23492
rect 37549 23490 37615 23493
rect 37292 23488 37615 23490
rect 37292 23432 37554 23488
rect 37610 23432 37615 23488
rect 37292 23430 37615 23432
rect 37292 23428 37298 23430
rect 28533 23427 28599 23428
rect 37549 23427 37615 23430
rect 37733 23492 37799 23493
rect 37733 23488 37780 23492
rect 37844 23490 37850 23492
rect 37733 23432 37738 23488
rect 37733 23428 37780 23432
rect 37844 23430 37890 23490
rect 37844 23428 37850 23430
rect 37733 23427 37799 23428
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 22185 23354 22251 23357
rect 22185 23352 23858 23354
rect 22185 23296 22190 23352
rect 22246 23296 23858 23352
rect 22185 23294 23858 23296
rect 22185 23291 22251 23294
rect 0 23218 800 23248
rect 3601 23218 3667 23221
rect 0 23216 3667 23218
rect 0 23160 3606 23216
rect 3662 23160 3667 23216
rect 0 23158 3667 23160
rect 0 23128 800 23158
rect 3601 23155 3667 23158
rect 17401 23218 17467 23221
rect 17953 23218 18019 23221
rect 17401 23216 18019 23218
rect 17401 23160 17406 23216
rect 17462 23160 17958 23216
rect 18014 23160 18019 23216
rect 17401 23158 18019 23160
rect 17401 23155 17467 23158
rect 17953 23155 18019 23158
rect 23238 23156 23244 23220
rect 23308 23218 23314 23220
rect 23657 23218 23723 23221
rect 23308 23216 23723 23218
rect 23308 23160 23662 23216
rect 23718 23160 23723 23216
rect 23308 23158 23723 23160
rect 23798 23218 23858 23294
rect 24710 23292 24716 23356
rect 24780 23354 24786 23356
rect 28441 23354 28507 23357
rect 24780 23352 28507 23354
rect 24780 23296 28446 23352
rect 28502 23296 28507 23352
rect 24780 23294 28507 23296
rect 24780 23292 24786 23294
rect 28441 23291 28507 23294
rect 25037 23218 25103 23221
rect 23798 23216 25103 23218
rect 23798 23160 25042 23216
rect 25098 23160 25103 23216
rect 23798 23158 25103 23160
rect 23308 23156 23314 23158
rect 23657 23155 23723 23158
rect 25037 23155 25103 23158
rect 21265 23082 21331 23085
rect 41873 23082 41939 23085
rect 21265 23080 41939 23082
rect 21265 23024 21270 23080
rect 21326 23024 41878 23080
rect 41934 23024 41939 23080
rect 21265 23022 41939 23024
rect 21265 23019 21331 23022
rect 41873 23019 41939 23022
rect 5073 22946 5139 22949
rect 5390 22946 5396 22948
rect 5073 22944 5396 22946
rect 5073 22888 5078 22944
rect 5134 22888 5396 22944
rect 5073 22886 5396 22888
rect 5073 22883 5139 22886
rect 5390 22884 5396 22886
rect 5460 22884 5466 22948
rect 16021 22946 16087 22949
rect 16389 22946 16455 22949
rect 16021 22944 16455 22946
rect 16021 22888 16026 22944
rect 16082 22888 16394 22944
rect 16450 22888 16455 22944
rect 16021 22886 16455 22888
rect 16021 22883 16087 22886
rect 16389 22883 16455 22886
rect 20989 22946 21055 22949
rect 22921 22946 22987 22949
rect 20989 22944 22987 22946
rect 20989 22888 20994 22944
rect 21050 22888 22926 22944
rect 22982 22888 22987 22944
rect 20989 22886 22987 22888
rect 20989 22883 21055 22886
rect 22921 22883 22987 22886
rect 23197 22946 23263 22949
rect 26366 22946 26372 22948
rect 23197 22944 26372 22946
rect 23197 22888 23202 22944
rect 23258 22888 26372 22944
rect 23197 22886 26372 22888
rect 23197 22883 23263 22886
rect 26366 22884 26372 22886
rect 26436 22884 26442 22948
rect 28533 22946 28599 22949
rect 36169 22948 36235 22949
rect 29494 22946 29500 22948
rect 28533 22944 29500 22946
rect 28533 22888 28538 22944
rect 28594 22888 29500 22944
rect 28533 22886 29500 22888
rect 28533 22883 28599 22886
rect 29494 22884 29500 22886
rect 29564 22884 29570 22948
rect 36118 22884 36124 22948
rect 36188 22946 36235 22948
rect 36188 22944 36280 22946
rect 36230 22888 36280 22944
rect 36188 22886 36280 22888
rect 36188 22884 36235 22886
rect 36169 22883 36235 22884
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 22185 22810 22251 22813
rect 22921 22810 22987 22813
rect 22185 22808 22987 22810
rect 22185 22752 22190 22808
rect 22246 22752 22926 22808
rect 22982 22752 22987 22808
rect 22185 22750 22987 22752
rect 22185 22747 22251 22750
rect 22921 22747 22987 22750
rect 23381 22810 23447 22813
rect 23606 22810 23612 22812
rect 23381 22808 23612 22810
rect 23381 22752 23386 22808
rect 23442 22752 23612 22808
rect 23381 22750 23612 22752
rect 23381 22747 23447 22750
rect 23606 22748 23612 22750
rect 23676 22748 23682 22812
rect 12065 22674 12131 22677
rect 13813 22674 13879 22677
rect 12065 22672 13879 22674
rect 12065 22616 12070 22672
rect 12126 22616 13818 22672
rect 13874 22616 13879 22672
rect 12065 22614 13879 22616
rect 12065 22611 12131 22614
rect 13813 22611 13879 22614
rect 21265 22674 21331 22677
rect 22185 22674 22251 22677
rect 24853 22674 24919 22677
rect 21265 22672 24919 22674
rect 21265 22616 21270 22672
rect 21326 22616 22190 22672
rect 22246 22616 24858 22672
rect 24914 22616 24919 22672
rect 21265 22614 24919 22616
rect 21265 22611 21331 22614
rect 22185 22611 22251 22614
rect 24853 22611 24919 22614
rect 25814 22612 25820 22676
rect 25884 22674 25890 22676
rect 26049 22674 26115 22677
rect 25884 22672 26115 22674
rect 25884 22616 26054 22672
rect 26110 22616 26115 22672
rect 25884 22614 26115 22616
rect 25884 22612 25890 22614
rect 26049 22611 26115 22614
rect 30097 22674 30163 22677
rect 35525 22674 35591 22677
rect 35934 22674 35940 22676
rect 30097 22672 35940 22674
rect 30097 22616 30102 22672
rect 30158 22616 35530 22672
rect 35586 22616 35940 22672
rect 30097 22614 35940 22616
rect 30097 22611 30163 22614
rect 35525 22611 35591 22614
rect 35934 22612 35940 22614
rect 36004 22612 36010 22676
rect 25405 22538 25471 22541
rect 28993 22538 29059 22541
rect 30741 22538 30807 22541
rect 25405 22536 30807 22538
rect 25405 22480 25410 22536
rect 25466 22480 28998 22536
rect 29054 22480 30746 22536
rect 30802 22480 30807 22536
rect 25405 22478 30807 22480
rect 25405 22475 25471 22478
rect 28993 22475 29059 22478
rect 30741 22475 30807 22478
rect 31385 22538 31451 22541
rect 32254 22538 32260 22540
rect 31385 22536 32260 22538
rect 31385 22480 31390 22536
rect 31446 22480 32260 22536
rect 31385 22478 32260 22480
rect 31385 22475 31451 22478
rect 32254 22476 32260 22478
rect 32324 22476 32330 22540
rect 34646 22476 34652 22540
rect 34716 22538 34722 22540
rect 34881 22538 34947 22541
rect 34716 22536 34947 22538
rect 34716 22480 34886 22536
rect 34942 22480 34947 22536
rect 34716 22478 34947 22480
rect 34716 22476 34722 22478
rect 34881 22475 34947 22478
rect 22461 22402 22527 22405
rect 23565 22402 23631 22405
rect 28625 22402 28691 22405
rect 22461 22400 28691 22402
rect 22461 22344 22466 22400
rect 22522 22344 23570 22400
rect 23626 22344 28630 22400
rect 28686 22344 28691 22400
rect 22461 22342 28691 22344
rect 22461 22339 22527 22342
rect 23565 22339 23631 22342
rect 28625 22339 28691 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 21081 22266 21147 22269
rect 21357 22266 21423 22269
rect 21081 22264 21423 22266
rect 21081 22208 21086 22264
rect 21142 22208 21362 22264
rect 21418 22208 21423 22264
rect 21081 22206 21423 22208
rect 21081 22203 21147 22206
rect 21357 22203 21423 22206
rect 21633 22266 21699 22269
rect 22277 22266 22343 22269
rect 21633 22264 22343 22266
rect 21633 22208 21638 22264
rect 21694 22208 22282 22264
rect 22338 22208 22343 22264
rect 21633 22206 22343 22208
rect 21633 22203 21699 22206
rect 22277 22203 22343 22206
rect 22553 22266 22619 22269
rect 30465 22266 30531 22269
rect 22553 22264 30531 22266
rect 22553 22208 22558 22264
rect 22614 22208 30470 22264
rect 30526 22208 30531 22264
rect 22553 22206 30531 22208
rect 22553 22203 22619 22206
rect 30465 22203 30531 22206
rect 20662 22068 20668 22132
rect 20732 22130 20738 22132
rect 23197 22130 23263 22133
rect 30046 22130 30052 22132
rect 20732 22128 23263 22130
rect 20732 22072 23202 22128
rect 23258 22072 23263 22128
rect 20732 22070 23263 22072
rect 20732 22068 20738 22070
rect 23197 22067 23263 22070
rect 23384 22070 30052 22130
rect 9070 21932 9076 21996
rect 9140 21994 9146 21996
rect 10041 21994 10107 21997
rect 12893 21996 12959 21997
rect 12893 21994 12940 21996
rect 9140 21992 10107 21994
rect 9140 21936 10046 21992
rect 10102 21936 10107 21992
rect 9140 21934 10107 21936
rect 12848 21992 12940 21994
rect 12848 21936 12898 21992
rect 12848 21934 12940 21936
rect 9140 21932 9146 21934
rect 10041 21931 10107 21934
rect 12893 21932 12940 21934
rect 13004 21932 13010 21996
rect 13854 21932 13860 21996
rect 13924 21994 13930 21996
rect 14273 21994 14339 21997
rect 13924 21992 14339 21994
rect 13924 21936 14278 21992
rect 14334 21936 14339 21992
rect 13924 21934 14339 21936
rect 13924 21932 13930 21934
rect 12893 21931 12959 21932
rect 14273 21931 14339 21934
rect 17401 21994 17467 21997
rect 17534 21994 17540 21996
rect 17401 21992 17540 21994
rect 17401 21936 17406 21992
rect 17462 21936 17540 21992
rect 17401 21934 17540 21936
rect 17401 21931 17467 21934
rect 17534 21932 17540 21934
rect 17604 21932 17610 21996
rect 20621 21994 20687 21997
rect 21081 21994 21147 21997
rect 21725 21994 21791 21997
rect 22461 21996 22527 21997
rect 22461 21994 22508 21996
rect 20621 21992 20914 21994
rect 20621 21936 20626 21992
rect 20682 21936 20914 21992
rect 20621 21934 20914 21936
rect 20621 21931 20687 21934
rect 20854 21858 20914 21934
rect 21081 21992 21791 21994
rect 21081 21936 21086 21992
rect 21142 21936 21730 21992
rect 21786 21936 21791 21992
rect 21081 21934 21791 21936
rect 22420 21992 22508 21994
rect 22572 21994 22578 21996
rect 23384 21994 23444 22070
rect 30046 22068 30052 22070
rect 30116 22068 30122 22132
rect 30833 22130 30899 22133
rect 30966 22130 30972 22132
rect 30833 22128 30972 22130
rect 30833 22072 30838 22128
rect 30894 22072 30972 22128
rect 30833 22070 30972 22072
rect 30833 22067 30899 22070
rect 30966 22068 30972 22070
rect 31036 22068 31042 22132
rect 22420 21936 22466 21992
rect 22420 21934 22508 21936
rect 21081 21931 21147 21934
rect 21725 21931 21791 21934
rect 22461 21932 22508 21934
rect 22572 21934 23444 21994
rect 24393 21994 24459 21997
rect 25957 21996 26023 21997
rect 24526 21994 24532 21996
rect 24393 21992 24532 21994
rect 24393 21936 24398 21992
rect 24454 21936 24532 21992
rect 24393 21934 24532 21936
rect 22572 21932 22578 21934
rect 22461 21931 22527 21932
rect 24393 21931 24459 21934
rect 24526 21932 24532 21934
rect 24596 21932 24602 21996
rect 25630 21932 25636 21996
rect 25700 21994 25706 21996
rect 25957 21994 26004 21996
rect 25700 21992 26004 21994
rect 25700 21936 25962 21992
rect 25700 21934 26004 21936
rect 25700 21932 25706 21934
rect 25957 21932 26004 21934
rect 26068 21932 26074 21996
rect 31293 21994 31359 21997
rect 31661 21994 31727 21997
rect 31293 21992 31727 21994
rect 31293 21936 31298 21992
rect 31354 21936 31666 21992
rect 31722 21936 31727 21992
rect 31293 21934 31727 21936
rect 25957 21931 26023 21932
rect 31293 21931 31359 21934
rect 31661 21931 31727 21934
rect 21030 21858 21036 21860
rect 20854 21798 21036 21858
rect 21030 21796 21036 21798
rect 21100 21796 21106 21860
rect 22369 21858 22435 21861
rect 23473 21858 23539 21861
rect 22369 21856 23539 21858
rect 22369 21800 22374 21856
rect 22430 21800 23478 21856
rect 23534 21800 23539 21856
rect 22369 21798 23539 21800
rect 22369 21795 22435 21798
rect 23473 21795 23539 21798
rect 25037 21858 25103 21861
rect 25957 21858 26023 21861
rect 25037 21856 26023 21858
rect 25037 21800 25042 21856
rect 25098 21800 25962 21856
rect 26018 21800 26023 21856
rect 25037 21798 26023 21800
rect 25037 21795 25103 21798
rect 25957 21795 26023 21798
rect 31702 21796 31708 21860
rect 31772 21858 31778 21860
rect 36118 21858 36124 21860
rect 31772 21798 36124 21858
rect 31772 21796 31778 21798
rect 36118 21796 36124 21798
rect 36188 21796 36194 21860
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 21449 21722 21515 21725
rect 34329 21722 34395 21725
rect 34462 21722 34468 21724
rect 21449 21720 34468 21722
rect 21449 21664 21454 21720
rect 21510 21664 34334 21720
rect 34390 21664 34468 21720
rect 21449 21662 34468 21664
rect 21449 21659 21515 21662
rect 34329 21659 34395 21662
rect 34462 21660 34468 21662
rect 34532 21660 34538 21724
rect 19374 21388 19380 21452
rect 19444 21450 19450 21452
rect 19517 21450 19583 21453
rect 19444 21448 19583 21450
rect 19444 21392 19522 21448
rect 19578 21392 19583 21448
rect 19444 21390 19583 21392
rect 19444 21388 19450 21390
rect 19517 21387 19583 21390
rect 24393 21450 24459 21453
rect 26601 21450 26667 21453
rect 24393 21448 26667 21450
rect 24393 21392 24398 21448
rect 24454 21392 26606 21448
rect 26662 21392 26667 21448
rect 24393 21390 26667 21392
rect 24393 21387 24459 21390
rect 26601 21387 26667 21390
rect 21214 21252 21220 21316
rect 21284 21314 21290 21316
rect 22185 21314 22251 21317
rect 21284 21312 22251 21314
rect 21284 21256 22190 21312
rect 22246 21256 22251 21312
rect 21284 21254 22251 21256
rect 21284 21252 21290 21254
rect 22185 21251 22251 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 9254 21116 9260 21180
rect 9324 21178 9330 21180
rect 17309 21178 17375 21181
rect 18270 21178 18276 21180
rect 9324 21176 18276 21178
rect 9324 21120 17314 21176
rect 17370 21120 18276 21176
rect 9324 21118 18276 21120
rect 9324 21116 9330 21118
rect 17309 21115 17375 21118
rect 18270 21116 18276 21118
rect 18340 21116 18346 21180
rect 20713 21178 20779 21181
rect 27613 21178 27679 21181
rect 20713 21176 27679 21178
rect 20713 21120 20718 21176
rect 20774 21120 27618 21176
rect 27674 21120 27679 21176
rect 20713 21118 27679 21120
rect 20713 21115 20779 21118
rect 27613 21115 27679 21118
rect 41413 21178 41479 21181
rect 41749 21178 42549 21208
rect 41413 21176 42549 21178
rect 41413 21120 41418 21176
rect 41474 21120 42549 21176
rect 41413 21118 42549 21120
rect 41413 21115 41479 21118
rect 41749 21088 42549 21118
rect 23197 21042 23263 21045
rect 24945 21042 25011 21045
rect 23197 21040 25011 21042
rect 23197 20984 23202 21040
rect 23258 20984 24950 21040
rect 25006 20984 25011 21040
rect 23197 20982 25011 20984
rect 23197 20979 23263 20982
rect 24945 20979 25011 20982
rect 27286 20980 27292 21044
rect 27356 21042 27362 21044
rect 28349 21042 28415 21045
rect 27356 21040 28415 21042
rect 27356 20984 28354 21040
rect 28410 20984 28415 21040
rect 27356 20982 28415 20984
rect 27356 20980 27362 20982
rect 28349 20979 28415 20982
rect 16205 20906 16271 20909
rect 17125 20906 17191 20909
rect 16205 20904 17191 20906
rect 16205 20848 16210 20904
rect 16266 20848 17130 20904
rect 17186 20848 17191 20904
rect 16205 20846 17191 20848
rect 16205 20843 16271 20846
rect 17125 20843 17191 20846
rect 22870 20844 22876 20908
rect 22940 20906 22946 20908
rect 23105 20906 23171 20909
rect 22940 20904 23171 20906
rect 22940 20848 23110 20904
rect 23166 20848 23171 20904
rect 22940 20846 23171 20848
rect 22940 20844 22946 20846
rect 23105 20843 23171 20846
rect 31569 20906 31635 20909
rect 31569 20904 34898 20906
rect 31569 20848 31574 20904
rect 31630 20848 34898 20904
rect 31569 20846 34898 20848
rect 31569 20843 31635 20846
rect 16205 20772 16271 20773
rect 16205 20770 16252 20772
rect 16160 20768 16252 20770
rect 16160 20712 16210 20768
rect 16160 20710 16252 20712
rect 16205 20708 16252 20710
rect 16316 20708 16322 20772
rect 22001 20770 22067 20773
rect 25773 20770 25839 20773
rect 22001 20768 25839 20770
rect 22001 20712 22006 20768
rect 22062 20712 25778 20768
rect 25834 20712 25839 20768
rect 22001 20710 25839 20712
rect 16205 20707 16271 20708
rect 22001 20707 22067 20710
rect 25773 20707 25839 20710
rect 31569 20770 31635 20773
rect 33358 20770 33364 20772
rect 31569 20768 33364 20770
rect 31569 20712 31574 20768
rect 31630 20712 33364 20768
rect 31569 20710 33364 20712
rect 31569 20707 31635 20710
rect 33358 20708 33364 20710
rect 33428 20708 33434 20772
rect 34838 20770 34898 20846
rect 36537 20770 36603 20773
rect 37181 20770 37247 20773
rect 38837 20772 38903 20773
rect 38837 20770 38884 20772
rect 34838 20768 37247 20770
rect 34838 20712 36542 20768
rect 36598 20712 37186 20768
rect 37242 20712 37247 20768
rect 34838 20710 37247 20712
rect 38792 20768 38884 20770
rect 38792 20712 38842 20768
rect 38792 20710 38884 20712
rect 36537 20707 36603 20710
rect 37181 20707 37247 20710
rect 38837 20708 38884 20710
rect 38948 20708 38954 20772
rect 38837 20707 38903 20708
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 11789 20634 11855 20637
rect 16849 20634 16915 20637
rect 11789 20632 16915 20634
rect 11789 20576 11794 20632
rect 11850 20576 16854 20632
rect 16910 20576 16915 20632
rect 11789 20574 16915 20576
rect 11789 20571 11855 20574
rect 16849 20571 16915 20574
rect 23289 20634 23355 20637
rect 23422 20634 23428 20636
rect 23289 20632 23428 20634
rect 23289 20576 23294 20632
rect 23350 20576 23428 20632
rect 23289 20574 23428 20576
rect 23289 20571 23355 20574
rect 23422 20572 23428 20574
rect 23492 20572 23498 20636
rect 29494 20572 29500 20636
rect 29564 20634 29570 20636
rect 36445 20634 36511 20637
rect 29564 20632 36511 20634
rect 29564 20576 36450 20632
rect 36506 20576 36511 20632
rect 29564 20574 36511 20576
rect 29564 20572 29570 20574
rect 36445 20571 36511 20574
rect 32438 20436 32444 20500
rect 32508 20498 32514 20500
rect 34605 20498 34671 20501
rect 32508 20496 34671 20498
rect 32508 20440 34610 20496
rect 34666 20440 34671 20496
rect 32508 20438 34671 20440
rect 32508 20436 32514 20438
rect 34605 20435 34671 20438
rect 19190 20300 19196 20364
rect 19260 20362 19266 20364
rect 19701 20362 19767 20365
rect 19260 20360 19767 20362
rect 19260 20304 19706 20360
rect 19762 20304 19767 20360
rect 19260 20302 19767 20304
rect 19260 20300 19266 20302
rect 19701 20299 19767 20302
rect 22369 20362 22435 20365
rect 27889 20362 27955 20365
rect 22369 20360 27955 20362
rect 22369 20304 22374 20360
rect 22430 20304 27894 20360
rect 27950 20304 27955 20360
rect 22369 20302 27955 20304
rect 22369 20299 22435 20302
rect 27889 20299 27955 20302
rect 6821 20226 6887 20229
rect 10133 20226 10199 20229
rect 17493 20226 17559 20229
rect 6821 20224 17559 20226
rect 6821 20168 6826 20224
rect 6882 20168 10138 20224
rect 10194 20168 17498 20224
rect 17554 20168 17559 20224
rect 6821 20166 17559 20168
rect 6821 20163 6887 20166
rect 10133 20163 10199 20166
rect 17493 20163 17559 20166
rect 24761 20226 24827 20229
rect 31385 20226 31451 20229
rect 24761 20224 31451 20226
rect 24761 20168 24766 20224
rect 24822 20168 31390 20224
rect 31446 20168 31451 20224
rect 24761 20166 31451 20168
rect 24761 20163 24827 20166
rect 31385 20163 31451 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 14733 20092 14799 20093
rect 14733 20090 14780 20092
rect 14688 20088 14780 20090
rect 14688 20032 14738 20088
rect 14688 20030 14780 20032
rect 14733 20028 14780 20030
rect 14844 20028 14850 20092
rect 19609 20090 19675 20093
rect 27889 20090 27955 20093
rect 19609 20088 27955 20090
rect 19609 20032 19614 20088
rect 19670 20032 27894 20088
rect 27950 20032 27955 20088
rect 19609 20030 27955 20032
rect 14733 20027 14799 20028
rect 19609 20027 19675 20030
rect 27889 20027 27955 20030
rect 30005 20090 30071 20093
rect 30373 20090 30439 20093
rect 30005 20088 30439 20090
rect 30005 20032 30010 20088
rect 30066 20032 30378 20088
rect 30434 20032 30439 20088
rect 30005 20030 30439 20032
rect 30005 20027 30071 20030
rect 30373 20027 30439 20030
rect 23606 19892 23612 19956
rect 23676 19954 23682 19956
rect 27337 19954 27403 19957
rect 23676 19952 27403 19954
rect 23676 19896 27342 19952
rect 27398 19896 27403 19952
rect 23676 19894 27403 19896
rect 23676 19892 23682 19894
rect 27337 19891 27403 19894
rect 28993 19954 29059 19957
rect 31385 19954 31451 19957
rect 28993 19952 31451 19954
rect 28993 19896 28998 19952
rect 29054 19896 31390 19952
rect 31446 19896 31451 19952
rect 28993 19894 31451 19896
rect 28993 19891 29059 19894
rect 31385 19891 31451 19894
rect 9121 19818 9187 19821
rect 13813 19818 13879 19821
rect 9121 19816 13879 19818
rect 9121 19760 9126 19816
rect 9182 19760 13818 19816
rect 13874 19760 13879 19816
rect 9121 19758 13879 19760
rect 9121 19755 9187 19758
rect 13813 19755 13879 19758
rect 18229 19818 18295 19821
rect 35893 19818 35959 19821
rect 18229 19816 35959 19818
rect 18229 19760 18234 19816
rect 18290 19760 35898 19816
rect 35954 19760 35959 19816
rect 18229 19758 35959 19760
rect 18229 19755 18295 19758
rect 35893 19755 35959 19758
rect 23197 19682 23263 19685
rect 27705 19682 27771 19685
rect 28022 19682 28028 19684
rect 23197 19680 28028 19682
rect 23197 19624 23202 19680
rect 23258 19624 27710 19680
rect 27766 19624 28028 19680
rect 23197 19622 28028 19624
rect 23197 19619 23263 19622
rect 27705 19619 27771 19622
rect 28022 19620 28028 19622
rect 28092 19620 28098 19684
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 11145 19546 11211 19549
rect 10366 19544 11211 19546
rect 10366 19488 11150 19544
rect 11206 19488 11211 19544
rect 10366 19486 11211 19488
rect 4705 19410 4771 19413
rect 7281 19410 7347 19413
rect 4705 19408 7347 19410
rect 4705 19352 4710 19408
rect 4766 19352 7286 19408
rect 7342 19352 7347 19408
rect 4705 19350 7347 19352
rect 4705 19347 4771 19350
rect 7281 19347 7347 19350
rect 7741 19410 7807 19413
rect 10225 19410 10291 19413
rect 10366 19410 10426 19486
rect 11145 19483 11211 19486
rect 22921 19546 22987 19549
rect 25589 19546 25655 19549
rect 22921 19544 25655 19546
rect 22921 19488 22926 19544
rect 22982 19488 25594 19544
rect 25650 19488 25655 19544
rect 22921 19486 25655 19488
rect 22921 19483 22987 19486
rect 25589 19483 25655 19486
rect 27705 19546 27771 19549
rect 29177 19548 29243 19549
rect 30649 19548 30715 19549
rect 29126 19546 29132 19548
rect 27705 19544 29132 19546
rect 29196 19546 29243 19548
rect 30598 19546 30604 19548
rect 29196 19544 29324 19546
rect 27705 19488 27710 19544
rect 27766 19488 29132 19544
rect 29238 19488 29324 19544
rect 27705 19486 29132 19488
rect 27705 19483 27771 19486
rect 29126 19484 29132 19486
rect 29196 19486 29324 19488
rect 30522 19486 30604 19546
rect 30668 19546 30715 19548
rect 36169 19546 36235 19549
rect 30668 19544 36235 19546
rect 30710 19488 36174 19544
rect 36230 19488 36235 19544
rect 29196 19484 29243 19486
rect 30598 19484 30604 19486
rect 30668 19486 36235 19488
rect 30668 19484 30715 19486
rect 29177 19483 29243 19484
rect 30649 19483 30715 19484
rect 36169 19483 36235 19486
rect 7741 19408 10426 19410
rect 7741 19352 7746 19408
rect 7802 19352 10230 19408
rect 10286 19352 10426 19408
rect 7741 19350 10426 19352
rect 10501 19410 10567 19413
rect 12709 19410 12775 19413
rect 17493 19412 17559 19413
rect 24577 19412 24643 19413
rect 17493 19410 17540 19412
rect 10501 19408 12775 19410
rect 10501 19352 10506 19408
rect 10562 19352 12714 19408
rect 12770 19352 12775 19408
rect 10501 19350 12775 19352
rect 17448 19408 17540 19410
rect 17448 19352 17498 19408
rect 17448 19350 17540 19352
rect 7741 19347 7807 19350
rect 10225 19347 10291 19350
rect 10501 19347 10567 19350
rect 12709 19347 12775 19350
rect 17493 19348 17540 19350
rect 17604 19348 17610 19412
rect 24526 19348 24532 19412
rect 24596 19410 24643 19412
rect 26233 19410 26299 19413
rect 27705 19410 27771 19413
rect 28533 19410 28599 19413
rect 24596 19408 24688 19410
rect 24638 19352 24688 19408
rect 24596 19350 24688 19352
rect 26233 19408 28599 19410
rect 26233 19352 26238 19408
rect 26294 19352 27710 19408
rect 27766 19352 28538 19408
rect 28594 19352 28599 19408
rect 26233 19350 28599 19352
rect 24596 19348 24643 19350
rect 17493 19347 17559 19348
rect 24577 19347 24643 19348
rect 26233 19347 26299 19350
rect 27705 19347 27771 19350
rect 28533 19347 28599 19350
rect 33593 19410 33659 19413
rect 33726 19410 33732 19412
rect 33593 19408 33732 19410
rect 33593 19352 33598 19408
rect 33654 19352 33732 19408
rect 33593 19350 33732 19352
rect 33593 19347 33659 19350
rect 33726 19348 33732 19350
rect 33796 19348 33802 19412
rect 11462 19212 11468 19276
rect 11532 19274 11538 19276
rect 16113 19274 16179 19277
rect 11532 19272 16179 19274
rect 11532 19216 16118 19272
rect 16174 19216 16179 19272
rect 11532 19214 16179 19216
rect 11532 19212 11538 19214
rect 16113 19211 16179 19214
rect 20846 19212 20852 19276
rect 20916 19274 20922 19276
rect 23473 19274 23539 19277
rect 20916 19272 23539 19274
rect 20916 19216 23478 19272
rect 23534 19216 23539 19272
rect 20916 19214 23539 19216
rect 20916 19212 20922 19214
rect 23473 19211 23539 19214
rect 26601 19274 26667 19277
rect 27521 19274 27587 19277
rect 26601 19272 27587 19274
rect 26601 19216 26606 19272
rect 26662 19216 27526 19272
rect 27582 19216 27587 19272
rect 26601 19214 27587 19216
rect 26601 19211 26667 19214
rect 27521 19211 27587 19214
rect 31109 19274 31175 19277
rect 31518 19274 31524 19276
rect 31109 19272 31524 19274
rect 31109 19216 31114 19272
rect 31170 19216 31524 19272
rect 31109 19214 31524 19216
rect 31109 19211 31175 19214
rect 31518 19212 31524 19214
rect 31588 19212 31594 19276
rect 0 19138 800 19168
rect 3325 19138 3391 19141
rect 0 19136 3391 19138
rect 0 19080 3330 19136
rect 3386 19080 3391 19136
rect 0 19078 3391 19080
rect 0 19048 800 19078
rect 3325 19075 3391 19078
rect 14958 19076 14964 19140
rect 15028 19138 15034 19140
rect 17902 19138 17908 19140
rect 15028 19078 17908 19138
rect 15028 19076 15034 19078
rect 17902 19076 17908 19078
rect 17972 19076 17978 19140
rect 20069 19138 20135 19141
rect 21398 19138 21404 19140
rect 20069 19136 21404 19138
rect 20069 19080 20074 19136
rect 20130 19080 21404 19136
rect 20069 19078 21404 19080
rect 20069 19075 20135 19078
rect 21398 19076 21404 19078
rect 21468 19076 21474 19140
rect 26877 19138 26943 19141
rect 22050 19136 26943 19138
rect 22050 19080 26882 19136
rect 26938 19080 26943 19136
rect 22050 19078 26943 19080
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 19241 19002 19307 19005
rect 22050 19002 22110 19078
rect 26877 19075 26943 19078
rect 33910 19076 33916 19140
rect 33980 19138 33986 19140
rect 34053 19138 34119 19141
rect 33980 19136 34119 19138
rect 33980 19080 34058 19136
rect 34114 19080 34119 19136
rect 33980 19078 34119 19080
rect 33980 19076 33986 19078
rect 34053 19075 34119 19078
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19241 19000 22110 19002
rect 19241 18944 19246 19000
rect 19302 18944 22110 19000
rect 19241 18942 22110 18944
rect 25129 19002 25195 19005
rect 25262 19002 25268 19004
rect 25129 19000 25268 19002
rect 25129 18944 25134 19000
rect 25190 18944 25268 19000
rect 25129 18942 25268 18944
rect 19241 18939 19307 18942
rect 25129 18939 25195 18942
rect 25262 18940 25268 18942
rect 25332 18940 25338 19004
rect 26325 19002 26391 19005
rect 26734 19002 26740 19004
rect 26325 19000 26740 19002
rect 26325 18944 26330 19000
rect 26386 18944 26740 19000
rect 26325 18942 26740 18944
rect 26325 18939 26391 18942
rect 26734 18940 26740 18942
rect 26804 18940 26810 19004
rect 22001 18866 22067 18869
rect 34697 18866 34763 18869
rect 35065 18866 35131 18869
rect 22001 18864 35131 18866
rect 22001 18808 22006 18864
rect 22062 18808 34702 18864
rect 34758 18808 35070 18864
rect 35126 18808 35131 18864
rect 22001 18806 35131 18808
rect 22001 18803 22067 18806
rect 34697 18803 34763 18806
rect 35065 18803 35131 18806
rect 20989 18730 21055 18733
rect 26601 18730 26667 18733
rect 20989 18728 26667 18730
rect 20989 18672 20994 18728
rect 21050 18672 26606 18728
rect 26662 18672 26667 18728
rect 20989 18670 26667 18672
rect 20989 18667 21055 18670
rect 26601 18667 26667 18670
rect 31385 18730 31451 18733
rect 35382 18730 35388 18732
rect 31385 18728 35388 18730
rect 31385 18672 31390 18728
rect 31446 18672 35388 18728
rect 31385 18670 35388 18672
rect 31385 18667 31451 18670
rect 35382 18668 35388 18670
rect 35452 18730 35458 18732
rect 35617 18730 35683 18733
rect 35452 18728 35683 18730
rect 35452 18672 35622 18728
rect 35678 18672 35683 18728
rect 35452 18670 35683 18672
rect 35452 18668 35458 18670
rect 35617 18667 35683 18670
rect 20846 18532 20852 18596
rect 20916 18594 20922 18596
rect 22502 18594 22508 18596
rect 20916 18534 22508 18594
rect 20916 18532 20922 18534
rect 22502 18532 22508 18534
rect 22572 18532 22578 18596
rect 31477 18594 31543 18597
rect 31753 18594 31819 18597
rect 33133 18594 33199 18597
rect 35801 18594 35867 18597
rect 31477 18592 35867 18594
rect 31477 18536 31482 18592
rect 31538 18536 31758 18592
rect 31814 18536 33138 18592
rect 33194 18536 35806 18592
rect 35862 18536 35867 18592
rect 31477 18534 35867 18536
rect 31477 18531 31543 18534
rect 31753 18531 31819 18534
rect 33133 18531 33199 18534
rect 35801 18531 35867 18534
rect 36854 18532 36860 18596
rect 36924 18594 36930 18596
rect 38561 18594 38627 18597
rect 36924 18592 38627 18594
rect 36924 18536 38566 18592
rect 38622 18536 38627 18592
rect 36924 18534 38627 18536
rect 36924 18532 36930 18534
rect 38561 18531 38627 18534
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 20161 18458 20227 18461
rect 24761 18458 24827 18461
rect 20161 18456 24827 18458
rect 20161 18400 20166 18456
rect 20222 18400 24766 18456
rect 24822 18400 24827 18456
rect 20161 18398 24827 18400
rect 20161 18395 20227 18398
rect 24761 18395 24827 18398
rect 33777 18458 33843 18461
rect 34094 18458 34100 18460
rect 33777 18456 34100 18458
rect 33777 18400 33782 18456
rect 33838 18400 34100 18456
rect 33777 18398 34100 18400
rect 33777 18395 33843 18398
rect 34094 18396 34100 18398
rect 34164 18396 34170 18460
rect 35893 18458 35959 18461
rect 36302 18458 36308 18460
rect 35893 18456 36308 18458
rect 35893 18400 35898 18456
rect 35954 18400 36308 18456
rect 35893 18398 36308 18400
rect 35893 18395 35959 18398
rect 36302 18396 36308 18398
rect 36372 18396 36378 18460
rect 17350 18260 17356 18324
rect 17420 18322 17426 18324
rect 21081 18322 21147 18325
rect 17420 18320 21147 18322
rect 17420 18264 21086 18320
rect 21142 18264 21147 18320
rect 17420 18262 21147 18264
rect 17420 18260 17426 18262
rect 21081 18259 21147 18262
rect 15745 18186 15811 18189
rect 15878 18186 15884 18188
rect 15745 18184 15884 18186
rect 15745 18128 15750 18184
rect 15806 18128 15884 18184
rect 15745 18126 15884 18128
rect 15745 18123 15811 18126
rect 15878 18124 15884 18126
rect 15948 18124 15954 18188
rect 33409 18186 33475 18189
rect 33542 18186 33548 18188
rect 33409 18184 33548 18186
rect 33409 18128 33414 18184
rect 33470 18128 33548 18184
rect 33409 18126 33548 18128
rect 33409 18123 33475 18126
rect 33542 18124 33548 18126
rect 33612 18124 33618 18188
rect 34973 18186 35039 18189
rect 35382 18186 35388 18188
rect 34973 18184 35388 18186
rect 34973 18128 34978 18184
rect 35034 18128 35388 18184
rect 34973 18126 35388 18128
rect 34973 18123 35039 18126
rect 35382 18124 35388 18126
rect 35452 18124 35458 18188
rect 20713 18052 20779 18053
rect 20662 17988 20668 18052
rect 20732 18050 20779 18052
rect 20732 18048 20824 18050
rect 20774 17992 20824 18048
rect 20732 17990 20824 17992
rect 20732 17988 20779 17990
rect 24894 17988 24900 18052
rect 24964 18050 24970 18052
rect 25865 18050 25931 18053
rect 24964 18048 25931 18050
rect 24964 17992 25870 18048
rect 25926 17992 25931 18048
rect 24964 17990 25931 17992
rect 24964 17988 24970 17990
rect 20713 17987 20779 17988
rect 25865 17987 25931 17990
rect 33174 17988 33180 18052
rect 33244 18050 33250 18052
rect 34329 18050 34395 18053
rect 33244 18048 34395 18050
rect 33244 17992 34334 18048
rect 34390 17992 34395 18048
rect 33244 17990 34395 17992
rect 33244 17988 33250 17990
rect 34329 17987 34395 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 17769 17914 17835 17917
rect 18965 17914 19031 17917
rect 17769 17912 19031 17914
rect 17769 17856 17774 17912
rect 17830 17856 18970 17912
rect 19026 17856 19031 17912
rect 17769 17854 19031 17856
rect 17769 17851 17835 17854
rect 18965 17851 19031 17854
rect 23565 17914 23631 17917
rect 23790 17914 23796 17916
rect 23565 17912 23796 17914
rect 23565 17856 23570 17912
rect 23626 17856 23796 17912
rect 23565 17854 23796 17856
rect 23565 17851 23631 17854
rect 23790 17852 23796 17854
rect 23860 17852 23866 17916
rect 26509 17914 26575 17917
rect 27102 17914 27108 17916
rect 26509 17912 27108 17914
rect 26509 17856 26514 17912
rect 26570 17856 27108 17912
rect 26509 17854 27108 17856
rect 26509 17851 26575 17854
rect 27102 17852 27108 17854
rect 27172 17852 27178 17916
rect 16113 17778 16179 17781
rect 19333 17778 19399 17781
rect 28257 17778 28323 17781
rect 31293 17778 31359 17781
rect 16113 17776 31359 17778
rect 16113 17720 16118 17776
rect 16174 17720 19338 17776
rect 19394 17720 28262 17776
rect 28318 17720 31298 17776
rect 31354 17720 31359 17776
rect 16113 17718 31359 17720
rect 16113 17715 16179 17718
rect 19333 17715 19399 17718
rect 28257 17715 28323 17718
rect 31293 17715 31359 17718
rect 33726 17716 33732 17780
rect 33796 17778 33802 17780
rect 36169 17778 36235 17781
rect 33796 17776 36235 17778
rect 33796 17720 36174 17776
rect 36230 17720 36235 17776
rect 33796 17718 36235 17720
rect 33796 17716 33802 17718
rect 36169 17715 36235 17718
rect 18229 17642 18295 17645
rect 18505 17642 18571 17645
rect 19057 17642 19123 17645
rect 29637 17642 29703 17645
rect 18229 17640 29703 17642
rect 18229 17584 18234 17640
rect 18290 17584 18510 17640
rect 18566 17584 19062 17640
rect 19118 17584 29642 17640
rect 29698 17584 29703 17640
rect 18229 17582 29703 17584
rect 18229 17579 18295 17582
rect 18505 17579 18571 17582
rect 19057 17579 19123 17582
rect 29637 17579 29703 17582
rect 17585 17506 17651 17509
rect 18873 17506 18939 17509
rect 17585 17504 18939 17506
rect 17585 17448 17590 17504
rect 17646 17448 18878 17504
rect 18934 17448 18939 17504
rect 17585 17446 18939 17448
rect 17585 17443 17651 17446
rect 18873 17443 18939 17446
rect 23013 17506 23079 17509
rect 23933 17506 23999 17509
rect 24342 17506 24348 17508
rect 23013 17504 24348 17506
rect 23013 17448 23018 17504
rect 23074 17448 23938 17504
rect 23994 17448 24348 17504
rect 23013 17446 24348 17448
rect 23013 17443 23079 17446
rect 23933 17443 23999 17446
rect 24342 17444 24348 17446
rect 24412 17444 24418 17508
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 21030 17308 21036 17372
rect 21100 17370 21106 17372
rect 26693 17370 26759 17373
rect 21100 17368 26759 17370
rect 21100 17312 26698 17368
rect 26754 17312 26759 17368
rect 21100 17310 26759 17312
rect 21100 17308 21106 17310
rect 26693 17307 26759 17310
rect 29862 17308 29868 17372
rect 29932 17370 29938 17372
rect 30005 17370 30071 17373
rect 35709 17370 35775 17373
rect 29932 17368 30071 17370
rect 29932 17312 30010 17368
rect 30066 17312 30071 17368
rect 29932 17310 30071 17312
rect 29932 17308 29938 17310
rect 30005 17307 30071 17310
rect 33366 17368 35775 17370
rect 33366 17312 35714 17368
rect 35770 17312 35775 17368
rect 33366 17310 35775 17312
rect 16430 17172 16436 17236
rect 16500 17234 16506 17236
rect 17217 17234 17283 17237
rect 16500 17232 17283 17234
rect 16500 17176 17222 17232
rect 17278 17176 17283 17232
rect 16500 17174 17283 17176
rect 16500 17172 16506 17174
rect 17217 17171 17283 17174
rect 22645 17234 22711 17237
rect 28625 17234 28691 17237
rect 22645 17232 28691 17234
rect 22645 17176 22650 17232
rect 22706 17176 28630 17232
rect 28686 17176 28691 17232
rect 22645 17174 28691 17176
rect 22645 17171 22711 17174
rect 28625 17171 28691 17174
rect 21909 17098 21975 17101
rect 26325 17098 26391 17101
rect 28073 17098 28139 17101
rect 21909 17096 28139 17098
rect 21909 17040 21914 17096
rect 21970 17040 26330 17096
rect 26386 17040 28078 17096
rect 28134 17040 28139 17096
rect 21909 17038 28139 17040
rect 21909 17035 21975 17038
rect 26325 17035 26391 17038
rect 28073 17035 28139 17038
rect 28574 17036 28580 17100
rect 28644 17098 28650 17100
rect 28901 17098 28967 17101
rect 28644 17096 28967 17098
rect 28644 17040 28906 17096
rect 28962 17040 28967 17096
rect 28644 17038 28967 17040
rect 33366 17098 33426 17310
rect 35709 17307 35775 17310
rect 33501 17234 33567 17237
rect 36537 17234 36603 17237
rect 33501 17232 36603 17234
rect 33501 17176 33506 17232
rect 33562 17176 36542 17232
rect 36598 17176 36603 17232
rect 33501 17174 36603 17176
rect 33501 17171 33567 17174
rect 36537 17171 36603 17174
rect 33501 17098 33567 17101
rect 38469 17098 38535 17101
rect 33366 17096 33567 17098
rect 33366 17040 33506 17096
rect 33562 17040 33567 17096
rect 33366 17038 33567 17040
rect 28644 17036 28650 17038
rect 28901 17035 28967 17038
rect 33501 17035 33567 17038
rect 34424 17096 38535 17098
rect 34424 17040 38474 17096
rect 38530 17040 38535 17096
rect 34424 17038 38535 17040
rect 20713 16962 20779 16965
rect 26049 16962 26115 16965
rect 20713 16960 26115 16962
rect 20713 16904 20718 16960
rect 20774 16904 26054 16960
rect 26110 16904 26115 16960
rect 20713 16902 26115 16904
rect 20713 16899 20779 16902
rect 26049 16899 26115 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 19885 16826 19951 16829
rect 23749 16826 23815 16829
rect 19885 16824 23815 16826
rect 19885 16768 19890 16824
rect 19946 16768 23754 16824
rect 23810 16768 23815 16824
rect 19885 16766 23815 16768
rect 19885 16763 19951 16766
rect 23749 16763 23815 16766
rect 32213 16826 32279 16829
rect 34424 16826 34484 17038
rect 38469 17035 38535 17038
rect 41749 17008 42549 17128
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 32213 16824 34484 16826
rect 32213 16768 32218 16824
rect 32274 16768 34484 16824
rect 32213 16766 34484 16768
rect 32213 16763 32279 16766
rect 23565 16692 23631 16693
rect 23565 16690 23612 16692
rect 23520 16688 23612 16690
rect 23520 16632 23570 16688
rect 23520 16630 23612 16632
rect 23565 16628 23612 16630
rect 23676 16628 23682 16692
rect 25865 16690 25931 16693
rect 26325 16690 26391 16693
rect 33409 16690 33475 16693
rect 25865 16688 26391 16690
rect 25865 16632 25870 16688
rect 25926 16632 26330 16688
rect 26386 16632 26391 16688
rect 25865 16630 26391 16632
rect 23565 16627 23631 16628
rect 25865 16627 25931 16630
rect 26325 16627 26391 16630
rect 30422 16688 33475 16690
rect 30422 16632 33414 16688
rect 33470 16632 33475 16688
rect 30422 16630 33475 16632
rect 10910 16492 10916 16556
rect 10980 16554 10986 16556
rect 11145 16554 11211 16557
rect 10980 16552 11211 16554
rect 10980 16496 11150 16552
rect 11206 16496 11211 16552
rect 10980 16494 11211 16496
rect 10980 16492 10986 16494
rect 11145 16491 11211 16494
rect 25998 16492 26004 16556
rect 26068 16554 26074 16556
rect 26141 16554 26207 16557
rect 26068 16552 26207 16554
rect 26068 16496 26146 16552
rect 26202 16496 26207 16552
rect 26068 16494 26207 16496
rect 26068 16492 26074 16494
rect 26141 16491 26207 16494
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 9029 16282 9095 16285
rect 9581 16282 9647 16285
rect 9029 16280 9647 16282
rect 9029 16224 9034 16280
rect 9090 16224 9586 16280
rect 9642 16224 9647 16280
rect 9029 16222 9647 16224
rect 9029 16219 9095 16222
rect 9581 16219 9647 16222
rect 19241 16146 19307 16149
rect 30422 16146 30482 16630
rect 33409 16627 33475 16630
rect 34053 16690 34119 16693
rect 34278 16690 34284 16692
rect 34053 16688 34284 16690
rect 34053 16632 34058 16688
rect 34114 16632 34284 16688
rect 34053 16630 34284 16632
rect 34053 16627 34119 16630
rect 34278 16628 34284 16630
rect 34348 16628 34354 16692
rect 36261 16690 36327 16693
rect 34470 16688 36327 16690
rect 34470 16632 36266 16688
rect 36322 16632 36327 16688
rect 34470 16630 36327 16632
rect 34470 16557 34530 16630
rect 36261 16627 36327 16630
rect 34421 16556 34530 16557
rect 34421 16554 34468 16556
rect 34380 16552 34468 16554
rect 34380 16496 34426 16552
rect 34380 16494 34468 16496
rect 34421 16492 34468 16494
rect 34532 16492 34538 16556
rect 34973 16554 35039 16557
rect 35750 16554 35756 16556
rect 34973 16552 35756 16554
rect 34973 16496 34978 16552
rect 35034 16496 35756 16552
rect 34973 16494 35756 16496
rect 34421 16491 34487 16492
rect 34973 16491 35039 16494
rect 35750 16492 35756 16494
rect 35820 16554 35826 16556
rect 36077 16554 36143 16557
rect 35820 16552 36143 16554
rect 35820 16496 36082 16552
rect 36138 16496 36143 16552
rect 35820 16494 36143 16496
rect 35820 16492 35826 16494
rect 36077 16491 36143 16494
rect 34513 16418 34579 16421
rect 35566 16418 35572 16420
rect 34513 16416 35572 16418
rect 34513 16360 34518 16416
rect 34574 16360 35572 16416
rect 34513 16358 35572 16360
rect 34513 16355 34579 16358
rect 35566 16356 35572 16358
rect 35636 16418 35642 16420
rect 36118 16418 36124 16420
rect 35636 16358 36124 16418
rect 35636 16356 35642 16358
rect 36118 16356 36124 16358
rect 36188 16356 36194 16420
rect 35433 16282 35499 16285
rect 36261 16282 36327 16285
rect 35433 16280 36327 16282
rect 35433 16224 35438 16280
rect 35494 16224 36266 16280
rect 36322 16224 36327 16280
rect 35433 16222 36327 16224
rect 35433 16219 35499 16222
rect 36261 16219 36327 16222
rect 19241 16144 30482 16146
rect 19241 16088 19246 16144
rect 19302 16088 30482 16144
rect 19241 16086 30482 16088
rect 31569 16146 31635 16149
rect 35433 16146 35499 16149
rect 37273 16148 37339 16149
rect 31569 16144 35499 16146
rect 31569 16088 31574 16144
rect 31630 16088 35438 16144
rect 35494 16088 35499 16144
rect 31569 16086 35499 16088
rect 19241 16083 19307 16086
rect 31569 16083 31635 16086
rect 35433 16083 35499 16086
rect 37222 16084 37228 16148
rect 37292 16146 37339 16148
rect 37292 16144 37384 16146
rect 37334 16088 37384 16144
rect 37292 16086 37384 16088
rect 37292 16084 37339 16086
rect 37273 16083 37339 16084
rect 21633 16010 21699 16013
rect 22870 16010 22876 16012
rect 21633 16008 22876 16010
rect 21633 15952 21638 16008
rect 21694 15952 22876 16008
rect 21633 15950 22876 15952
rect 21633 15947 21699 15950
rect 22870 15948 22876 15950
rect 22940 15948 22946 16012
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 22185 15740 22251 15741
rect 22134 15676 22140 15740
rect 22204 15738 22251 15740
rect 22204 15736 22296 15738
rect 22246 15680 22296 15736
rect 22204 15678 22296 15680
rect 22204 15676 22251 15678
rect 22185 15675 22251 15676
rect 15285 15466 15351 15469
rect 17125 15466 17191 15469
rect 19149 15466 19215 15469
rect 15285 15464 19215 15466
rect 15285 15408 15290 15464
rect 15346 15408 17130 15464
rect 17186 15408 19154 15464
rect 19210 15408 19215 15464
rect 15285 15406 19215 15408
rect 15285 15403 15351 15406
rect 17125 15403 17191 15406
rect 19149 15403 19215 15406
rect 26233 15330 26299 15333
rect 26877 15330 26943 15333
rect 26233 15328 26943 15330
rect 26233 15272 26238 15328
rect 26294 15272 26882 15328
rect 26938 15272 26943 15328
rect 26233 15270 26943 15272
rect 26233 15267 26299 15270
rect 26877 15267 26943 15270
rect 33910 15268 33916 15332
rect 33980 15330 33986 15332
rect 34789 15330 34855 15333
rect 33980 15328 34855 15330
rect 33980 15272 34794 15328
rect 34850 15272 34855 15328
rect 33980 15270 34855 15272
rect 33980 15268 33986 15270
rect 34789 15267 34855 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 1577 15194 1643 15197
rect 5349 15196 5415 15197
rect 5349 15194 5396 15196
rect 798 15192 1643 15194
rect 798 15136 1582 15192
rect 1638 15136 1643 15192
rect 798 15134 1643 15136
rect 5304 15192 5396 15194
rect 5304 15136 5354 15192
rect 5304 15134 5396 15136
rect 798 15088 858 15134
rect 1577 15131 1643 15134
rect 5349 15132 5396 15134
rect 5460 15132 5466 15196
rect 20161 15194 20227 15197
rect 20294 15194 20300 15196
rect 20161 15192 20300 15194
rect 20161 15136 20166 15192
rect 20222 15136 20300 15192
rect 20161 15134 20300 15136
rect 5349 15131 5415 15132
rect 20161 15131 20227 15134
rect 20294 15132 20300 15134
rect 20364 15132 20370 15196
rect 24577 15194 24643 15197
rect 25773 15196 25839 15197
rect 26877 15196 26943 15197
rect 24894 15194 24900 15196
rect 24577 15192 24900 15194
rect 24577 15136 24582 15192
rect 24638 15136 24900 15192
rect 24577 15134 24900 15136
rect 24577 15131 24643 15134
rect 24894 15132 24900 15134
rect 24964 15132 24970 15196
rect 25773 15194 25820 15196
rect 25728 15192 25820 15194
rect 25728 15136 25778 15192
rect 25728 15134 25820 15136
rect 25773 15132 25820 15134
rect 25884 15132 25890 15196
rect 26877 15194 26924 15196
rect 26832 15192 26924 15194
rect 26832 15136 26882 15192
rect 26832 15134 26924 15136
rect 26877 15132 26924 15134
rect 26988 15132 26994 15196
rect 27889 15194 27955 15197
rect 28206 15194 28212 15196
rect 27889 15192 28212 15194
rect 27889 15136 27894 15192
rect 27950 15136 28212 15192
rect 27889 15134 28212 15136
rect 25773 15131 25839 15132
rect 26877 15131 26943 15132
rect 27889 15131 27955 15134
rect 28206 15132 28212 15134
rect 28276 15132 28282 15196
rect 28441 15194 28507 15197
rect 28758 15194 28764 15196
rect 28441 15192 28764 15194
rect 28441 15136 28446 15192
rect 28502 15136 28764 15192
rect 28441 15134 28764 15136
rect 28441 15131 28507 15134
rect 28758 15132 28764 15134
rect 28828 15132 28834 15196
rect 29453 15194 29519 15197
rect 37549 15196 37615 15197
rect 30230 15194 30236 15196
rect 29453 15192 30236 15194
rect 29453 15136 29458 15192
rect 29514 15136 30236 15192
rect 29453 15134 30236 15136
rect 29453 15131 29519 15134
rect 30230 15132 30236 15134
rect 30300 15132 30306 15196
rect 37549 15192 37596 15196
rect 37660 15194 37666 15196
rect 37549 15136 37554 15192
rect 37549 15132 37596 15136
rect 37660 15134 37706 15194
rect 37660 15132 37666 15134
rect 37549 15131 37615 15132
rect 0 14998 858 15088
rect 0 14968 800 14998
rect 20110 14996 20116 15060
rect 20180 15058 20186 15060
rect 20897 15058 20963 15061
rect 20180 15056 20963 15058
rect 20180 15000 20902 15056
rect 20958 15000 20963 15056
rect 20180 14998 20963 15000
rect 20180 14996 20186 14998
rect 20897 14995 20963 14998
rect 21265 15058 21331 15061
rect 21909 15058 21975 15061
rect 21265 15056 21975 15058
rect 21265 15000 21270 15056
rect 21326 15000 21914 15056
rect 21970 15000 21975 15056
rect 21265 14998 21975 15000
rect 21265 14995 21331 14998
rect 21909 14995 21975 14998
rect 19425 14922 19491 14925
rect 21633 14922 21699 14925
rect 19425 14920 21699 14922
rect 19425 14864 19430 14920
rect 19486 14864 21638 14920
rect 21694 14864 21699 14920
rect 19425 14862 21699 14864
rect 19425 14859 19491 14862
rect 21633 14859 21699 14862
rect 22050 14862 35450 14922
rect 15653 14786 15719 14789
rect 21030 14786 21036 14788
rect 15653 14784 21036 14786
rect 15653 14728 15658 14784
rect 15714 14728 21036 14784
rect 15653 14726 21036 14728
rect 15653 14723 15719 14726
rect 21030 14724 21036 14726
rect 21100 14724 21106 14788
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 20345 14514 20411 14517
rect 22050 14514 22110 14862
rect 35390 14789 35450 14862
rect 30189 14786 30255 14789
rect 32765 14786 32831 14789
rect 35390 14788 35499 14789
rect 30189 14784 32831 14786
rect 30189 14728 30194 14784
rect 30250 14728 32770 14784
rect 32826 14728 32831 14784
rect 30189 14726 32831 14728
rect 30189 14723 30255 14726
rect 32765 14723 32831 14726
rect 35382 14724 35388 14788
rect 35452 14786 35499 14788
rect 35452 14784 35544 14786
rect 35494 14728 35544 14784
rect 35452 14726 35544 14728
rect 35452 14724 35499 14726
rect 35433 14723 35499 14724
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 22645 14650 22711 14653
rect 27429 14650 27495 14653
rect 22645 14648 27495 14650
rect 22645 14592 22650 14648
rect 22706 14592 27434 14648
rect 27490 14592 27495 14648
rect 22645 14590 27495 14592
rect 22645 14587 22711 14590
rect 27429 14587 27495 14590
rect 20345 14512 22110 14514
rect 20345 14456 20350 14512
rect 20406 14456 22110 14512
rect 20345 14454 22110 14456
rect 22737 14514 22803 14517
rect 28349 14514 28415 14517
rect 22737 14512 28415 14514
rect 22737 14456 22742 14512
rect 22798 14456 28354 14512
rect 28410 14456 28415 14512
rect 22737 14454 28415 14456
rect 20345 14451 20411 14454
rect 22737 14451 22803 14454
rect 28349 14451 28415 14454
rect 31937 14514 32003 14517
rect 39941 14514 40007 14517
rect 31937 14512 40007 14514
rect 31937 14456 31942 14512
rect 31998 14456 39946 14512
rect 40002 14456 40007 14512
rect 31937 14454 40007 14456
rect 31937 14451 32003 14454
rect 39941 14451 40007 14454
rect 19885 14378 19951 14381
rect 19382 14376 19951 14378
rect 19382 14320 19890 14376
rect 19946 14320 19951 14376
rect 19382 14318 19951 14320
rect 19382 13970 19442 14318
rect 19885 14315 19951 14318
rect 25497 14378 25563 14381
rect 27797 14378 27863 14381
rect 25497 14376 27863 14378
rect 25497 14320 25502 14376
rect 25558 14320 27802 14376
rect 27858 14320 27863 14376
rect 25497 14318 27863 14320
rect 25497 14315 25563 14318
rect 27797 14315 27863 14318
rect 29729 14378 29795 14381
rect 37774 14378 37780 14380
rect 29729 14376 37780 14378
rect 29729 14320 29734 14376
rect 29790 14320 37780 14376
rect 29729 14318 37780 14320
rect 29729 14315 29795 14318
rect 37774 14316 37780 14318
rect 37844 14378 37850 14380
rect 39757 14378 39823 14381
rect 37844 14376 39823 14378
rect 37844 14320 39762 14376
rect 39818 14320 39823 14376
rect 37844 14318 39823 14320
rect 37844 14316 37850 14318
rect 39757 14315 39823 14318
rect 26877 14242 26943 14245
rect 27797 14242 27863 14245
rect 37089 14244 37155 14245
rect 26877 14240 27863 14242
rect 26877 14184 26882 14240
rect 26938 14184 27802 14240
rect 27858 14184 27863 14240
rect 26877 14182 27863 14184
rect 26877 14179 26943 14182
rect 27797 14179 27863 14182
rect 37038 14180 37044 14244
rect 37108 14242 37155 14244
rect 37108 14240 37200 14242
rect 37150 14184 37200 14240
rect 37108 14182 37200 14184
rect 37108 14180 37155 14182
rect 37089 14179 37155 14180
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 25221 14106 25287 14109
rect 28349 14106 28415 14109
rect 25221 14104 28415 14106
rect 25221 14048 25226 14104
rect 25282 14048 28354 14104
rect 28410 14048 28415 14104
rect 25221 14046 28415 14048
rect 25221 14043 25287 14046
rect 28349 14043 28415 14046
rect 34646 14044 34652 14108
rect 34716 14106 34722 14108
rect 34789 14106 34855 14109
rect 34716 14104 34855 14106
rect 34716 14048 34794 14104
rect 34850 14048 34855 14104
rect 34716 14046 34855 14048
rect 34716 14044 34722 14046
rect 34789 14043 34855 14046
rect 19517 13970 19583 13973
rect 19382 13968 19583 13970
rect 19382 13912 19522 13968
rect 19578 13912 19583 13968
rect 19382 13910 19583 13912
rect 19517 13907 19583 13910
rect 19793 13970 19859 13973
rect 20846 13970 20852 13972
rect 19793 13968 20852 13970
rect 19793 13912 19798 13968
rect 19854 13912 20852 13968
rect 19793 13910 20852 13912
rect 19793 13907 19859 13910
rect 20846 13908 20852 13910
rect 20916 13908 20922 13972
rect 27061 13970 27127 13973
rect 28165 13970 28231 13973
rect 27061 13968 28231 13970
rect 27061 13912 27066 13968
rect 27122 13912 28170 13968
rect 28226 13912 28231 13968
rect 27061 13910 28231 13912
rect 27061 13907 27127 13910
rect 28165 13907 28231 13910
rect 16757 13834 16823 13837
rect 17534 13834 17540 13836
rect 16757 13832 17540 13834
rect 16757 13776 16762 13832
rect 16818 13776 17540 13832
rect 16757 13774 17540 13776
rect 16757 13771 16823 13774
rect 17534 13772 17540 13774
rect 17604 13772 17610 13836
rect 27245 13834 27311 13837
rect 27613 13834 27679 13837
rect 27245 13832 27679 13834
rect 27245 13776 27250 13832
rect 27306 13776 27618 13832
rect 27674 13776 27679 13832
rect 27245 13774 27679 13776
rect 27245 13771 27311 13774
rect 27613 13771 27679 13774
rect 32581 13834 32647 13837
rect 32990 13834 32996 13836
rect 32581 13832 32996 13834
rect 32581 13776 32586 13832
rect 32642 13776 32996 13832
rect 32581 13774 32996 13776
rect 32581 13771 32647 13774
rect 32990 13772 32996 13774
rect 33060 13772 33066 13836
rect 33777 13834 33843 13837
rect 34513 13834 34579 13837
rect 35065 13834 35131 13837
rect 33777 13832 35131 13834
rect 33777 13776 33782 13832
rect 33838 13776 34518 13832
rect 34574 13776 35070 13832
rect 35126 13776 35131 13832
rect 33777 13774 35131 13776
rect 33777 13771 33843 13774
rect 34513 13771 34579 13774
rect 35065 13771 35131 13774
rect 13537 13698 13603 13701
rect 17585 13698 17651 13701
rect 13537 13696 17651 13698
rect 13537 13640 13542 13696
rect 13598 13640 17590 13696
rect 17646 13640 17651 13696
rect 13537 13638 17651 13640
rect 13537 13635 13603 13638
rect 17585 13635 17651 13638
rect 24301 13698 24367 13701
rect 24710 13698 24716 13700
rect 24301 13696 24716 13698
rect 24301 13640 24306 13696
rect 24362 13640 24716 13696
rect 24301 13638 24716 13640
rect 24301 13635 24367 13638
rect 24710 13636 24716 13638
rect 24780 13636 24786 13700
rect 26550 13636 26556 13700
rect 26620 13698 26626 13700
rect 27245 13698 27311 13701
rect 26620 13696 27311 13698
rect 26620 13640 27250 13696
rect 27306 13640 27311 13696
rect 26620 13638 27311 13640
rect 26620 13636 26626 13638
rect 27245 13635 27311 13638
rect 37406 13636 37412 13700
rect 37476 13698 37482 13700
rect 37825 13698 37891 13701
rect 37476 13696 37891 13698
rect 37476 13640 37830 13696
rect 37886 13640 37891 13696
rect 37476 13638 37891 13640
rect 37476 13636 37482 13638
rect 37825 13635 37891 13638
rect 39021 13700 39087 13701
rect 39021 13696 39068 13700
rect 39132 13698 39138 13700
rect 41749 13698 42549 13728
rect 39021 13640 39026 13696
rect 39021 13636 39068 13640
rect 39132 13638 39178 13698
rect 39438 13638 42549 13698
rect 39132 13636 39138 13638
rect 39021 13635 39087 13636
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 12065 13562 12131 13565
rect 15745 13562 15811 13565
rect 16389 13562 16455 13565
rect 27429 13564 27495 13565
rect 27429 13562 27476 13564
rect 12065 13560 16455 13562
rect 12065 13504 12070 13560
rect 12126 13504 15750 13560
rect 15806 13504 16394 13560
rect 16450 13504 16455 13560
rect 12065 13502 16455 13504
rect 27384 13560 27476 13562
rect 27384 13504 27434 13560
rect 27384 13502 27476 13504
rect 12065 13499 12131 13502
rect 15745 13499 15811 13502
rect 16389 13499 16455 13502
rect 27429 13500 27476 13502
rect 27540 13500 27546 13564
rect 39113 13562 39179 13565
rect 39246 13562 39252 13564
rect 39113 13560 39252 13562
rect 39113 13504 39118 13560
rect 39174 13504 39252 13560
rect 39113 13502 39252 13504
rect 27429 13499 27495 13500
rect 39113 13499 39179 13502
rect 39246 13500 39252 13502
rect 39316 13500 39322 13564
rect 30833 13426 30899 13429
rect 37273 13426 37339 13429
rect 30833 13424 37339 13426
rect 30833 13368 30838 13424
rect 30894 13368 37278 13424
rect 37334 13368 37339 13424
rect 30833 13366 37339 13368
rect 30833 13363 30899 13366
rect 37273 13363 37339 13366
rect 38561 13426 38627 13429
rect 39438 13426 39498 13638
rect 41749 13608 42549 13638
rect 38561 13424 39498 13426
rect 38561 13368 38566 13424
rect 38622 13368 39498 13424
rect 38561 13366 39498 13368
rect 38561 13363 38627 13366
rect 10593 13290 10659 13293
rect 16665 13290 16731 13293
rect 10593 13288 16731 13290
rect 10593 13232 10598 13288
rect 10654 13232 16670 13288
rect 16726 13232 16731 13288
rect 10593 13230 16731 13232
rect 10593 13227 10659 13230
rect 16665 13227 16731 13230
rect 34513 13290 34579 13293
rect 36353 13290 36419 13293
rect 34513 13288 36419 13290
rect 34513 13232 34518 13288
rect 34574 13232 36358 13288
rect 36414 13232 36419 13288
rect 34513 13230 36419 13232
rect 34513 13227 34579 13230
rect 36353 13227 36419 13230
rect 16113 13154 16179 13157
rect 18413 13154 18479 13157
rect 16113 13152 18479 13154
rect 16113 13096 16118 13152
rect 16174 13096 18418 13152
rect 18474 13096 18479 13152
rect 16113 13094 18479 13096
rect 16113 13091 16179 13094
rect 18413 13091 18479 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 7373 13018 7439 13021
rect 7833 13018 7899 13021
rect 9213 13018 9279 13021
rect 11789 13018 11855 13021
rect 15469 13018 15535 13021
rect 17677 13018 17743 13021
rect 7373 13016 9279 13018
rect 7373 12960 7378 13016
rect 7434 12960 7838 13016
rect 7894 12960 9218 13016
rect 9274 12960 9279 13016
rect 7373 12958 9279 12960
rect 7373 12955 7439 12958
rect 7833 12955 7899 12958
rect 9213 12955 9279 12958
rect 9630 13016 17743 13018
rect 9630 12960 11794 13016
rect 11850 12960 15474 13016
rect 15530 12960 17682 13016
rect 17738 12960 17743 13016
rect 9630 12958 17743 12960
rect 8017 12882 8083 12885
rect 9121 12882 9187 12885
rect 8017 12880 9187 12882
rect 8017 12824 8022 12880
rect 8078 12824 9126 12880
rect 9182 12824 9187 12880
rect 8017 12822 9187 12824
rect 8017 12819 8083 12822
rect 9121 12819 9187 12822
rect 4889 12746 4955 12749
rect 5993 12746 6059 12749
rect 9630 12746 9690 12958
rect 11789 12955 11855 12958
rect 15469 12955 15535 12958
rect 17677 12955 17743 12958
rect 32581 13018 32647 13021
rect 37273 13018 37339 13021
rect 32581 13016 37339 13018
rect 32581 12960 32586 13016
rect 32642 12960 37278 13016
rect 37334 12960 37339 13016
rect 32581 12958 37339 12960
rect 32581 12955 32647 12958
rect 37273 12955 37339 12958
rect 10041 12882 10107 12885
rect 12617 12882 12683 12885
rect 10041 12880 12683 12882
rect 10041 12824 10046 12880
rect 10102 12824 12622 12880
rect 12678 12824 12683 12880
rect 10041 12822 12683 12824
rect 10041 12819 10107 12822
rect 12617 12819 12683 12822
rect 15561 12882 15627 12885
rect 23381 12882 23447 12885
rect 15561 12880 23447 12882
rect 15561 12824 15566 12880
rect 15622 12824 23386 12880
rect 23442 12824 23447 12880
rect 15561 12822 23447 12824
rect 15561 12819 15627 12822
rect 23381 12819 23447 12822
rect 30373 12882 30439 12885
rect 34053 12882 34119 12885
rect 30373 12880 34119 12882
rect 30373 12824 30378 12880
rect 30434 12824 34058 12880
rect 34114 12824 34119 12880
rect 30373 12822 34119 12824
rect 30373 12819 30439 12822
rect 34053 12819 34119 12822
rect 4889 12744 9690 12746
rect 4889 12688 4894 12744
rect 4950 12688 5998 12744
rect 6054 12688 9690 12744
rect 4889 12686 9690 12688
rect 11605 12746 11671 12749
rect 18781 12746 18847 12749
rect 11605 12744 18847 12746
rect 11605 12688 11610 12744
rect 11666 12688 18786 12744
rect 18842 12688 18847 12744
rect 11605 12686 18847 12688
rect 4889 12683 4955 12686
rect 5993 12683 6059 12686
rect 11605 12683 11671 12686
rect 18781 12683 18847 12686
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 24393 12474 24459 12477
rect 28625 12474 28691 12477
rect 24393 12472 28691 12474
rect 24393 12416 24398 12472
rect 24454 12416 28630 12472
rect 28686 12416 28691 12472
rect 24393 12414 28691 12416
rect 24393 12411 24459 12414
rect 28625 12411 28691 12414
rect 12525 12338 12591 12341
rect 14457 12338 14523 12341
rect 12525 12336 14523 12338
rect 12525 12280 12530 12336
rect 12586 12280 14462 12336
rect 14518 12280 14523 12336
rect 12525 12278 14523 12280
rect 12525 12275 12591 12278
rect 14457 12275 14523 12278
rect 23473 12338 23539 12341
rect 25589 12338 25655 12341
rect 23473 12336 25655 12338
rect 23473 12280 23478 12336
rect 23534 12280 25594 12336
rect 25650 12280 25655 12336
rect 23473 12278 25655 12280
rect 23473 12275 23539 12278
rect 25589 12275 25655 12278
rect 26509 12338 26575 12341
rect 27521 12338 27587 12341
rect 26509 12336 27587 12338
rect 26509 12280 26514 12336
rect 26570 12280 27526 12336
rect 27582 12280 27587 12336
rect 26509 12278 27587 12280
rect 26509 12275 26575 12278
rect 27521 12275 27587 12278
rect 32397 12338 32463 12341
rect 39389 12338 39455 12341
rect 40217 12338 40283 12341
rect 32397 12336 40283 12338
rect 32397 12280 32402 12336
rect 32458 12280 39394 12336
rect 39450 12280 40222 12336
rect 40278 12280 40283 12336
rect 32397 12278 40283 12280
rect 32397 12275 32463 12278
rect 39389 12275 39455 12278
rect 40217 12275 40283 12278
rect 13905 12202 13971 12205
rect 14641 12202 14707 12205
rect 30925 12202 30991 12205
rect 13905 12200 30991 12202
rect 13905 12144 13910 12200
rect 13966 12144 14646 12200
rect 14702 12144 30930 12200
rect 30986 12144 30991 12200
rect 13905 12142 30991 12144
rect 13905 12139 13971 12142
rect 14641 12139 14707 12142
rect 30925 12139 30991 12142
rect 11053 12068 11119 12069
rect 35985 12068 36051 12069
rect 11053 12064 11100 12068
rect 11164 12066 11170 12068
rect 35934 12066 35940 12068
rect 11053 12008 11058 12064
rect 11053 12004 11100 12008
rect 11164 12006 11210 12066
rect 35894 12006 35940 12066
rect 36004 12064 36051 12068
rect 36046 12008 36051 12064
rect 11164 12004 11170 12006
rect 35934 12004 35940 12006
rect 36004 12004 36051 12008
rect 11053 12003 11119 12004
rect 35985 12003 36051 12004
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 29269 11930 29335 11933
rect 38561 11930 38627 11933
rect 29269 11928 38627 11930
rect 29269 11872 29274 11928
rect 29330 11872 38566 11928
rect 38622 11872 38627 11928
rect 29269 11870 38627 11872
rect 29269 11867 29335 11870
rect 38561 11867 38627 11870
rect 15101 11794 15167 11797
rect 22737 11794 22803 11797
rect 15101 11792 22803 11794
rect 15101 11736 15106 11792
rect 15162 11736 22742 11792
rect 22798 11736 22803 11792
rect 15101 11734 22803 11736
rect 15101 11731 15167 11734
rect 22737 11731 22803 11734
rect 34421 11796 34487 11797
rect 34421 11792 34468 11796
rect 34532 11794 34538 11796
rect 35065 11794 35131 11797
rect 36813 11794 36879 11797
rect 34421 11736 34426 11792
rect 34421 11732 34468 11736
rect 34532 11734 34578 11794
rect 35065 11792 36879 11794
rect 35065 11736 35070 11792
rect 35126 11736 36818 11792
rect 36874 11736 36879 11792
rect 35065 11734 36879 11736
rect 34532 11732 34538 11734
rect 34421 11731 34487 11732
rect 35065 11731 35131 11734
rect 36813 11731 36879 11734
rect 0 11658 800 11688
rect 933 11658 999 11661
rect 0 11656 999 11658
rect 0 11600 938 11656
rect 994 11600 999 11656
rect 0 11598 999 11600
rect 0 11568 800 11598
rect 933 11595 999 11598
rect 39113 11658 39179 11661
rect 40033 11658 40099 11661
rect 39113 11656 40099 11658
rect 39113 11600 39118 11656
rect 39174 11600 40038 11656
rect 40094 11600 40099 11656
rect 39113 11598 40099 11600
rect 39113 11595 39179 11598
rect 40033 11595 40099 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 30281 11114 30347 11117
rect 33593 11114 33659 11117
rect 30281 11112 33659 11114
rect 30281 11056 30286 11112
rect 30342 11056 33598 11112
rect 33654 11056 33659 11112
rect 30281 11054 33659 11056
rect 30281 11051 30347 11054
rect 33593 11051 33659 11054
rect 11973 10980 12039 10981
rect 11973 10978 12020 10980
rect 11928 10976 12020 10978
rect 11928 10920 11978 10976
rect 11928 10918 12020 10920
rect 11973 10916 12020 10918
rect 12084 10916 12090 10980
rect 21398 10916 21404 10980
rect 21468 10978 21474 10980
rect 21633 10978 21699 10981
rect 21468 10976 21699 10978
rect 21468 10920 21638 10976
rect 21694 10920 21699 10976
rect 21468 10918 21699 10920
rect 21468 10916 21474 10918
rect 11973 10915 12039 10916
rect 21633 10915 21699 10918
rect 27429 10978 27495 10981
rect 29494 10978 29500 10980
rect 27429 10976 29500 10978
rect 27429 10920 27434 10976
rect 27490 10920 29500 10976
rect 27429 10918 29500 10920
rect 27429 10915 27495 10918
rect 29494 10916 29500 10918
rect 29564 10916 29570 10980
rect 32990 10916 32996 10980
rect 33060 10978 33066 10980
rect 38101 10978 38167 10981
rect 33060 10976 38167 10978
rect 33060 10920 38106 10976
rect 38162 10920 38167 10976
rect 33060 10918 38167 10920
rect 33060 10916 33066 10918
rect 38101 10915 38167 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 10358 10780 10364 10844
rect 10428 10842 10434 10844
rect 13445 10842 13511 10845
rect 10428 10840 13511 10842
rect 10428 10784 13450 10840
rect 13506 10784 13511 10840
rect 10428 10782 13511 10784
rect 10428 10780 10434 10782
rect 13445 10779 13511 10782
rect 16849 10842 16915 10845
rect 17718 10842 17724 10844
rect 16849 10840 17724 10842
rect 16849 10784 16854 10840
rect 16910 10784 17724 10840
rect 16849 10782 17724 10784
rect 16849 10779 16915 10782
rect 17718 10780 17724 10782
rect 17788 10780 17794 10844
rect 29637 10842 29703 10845
rect 33041 10842 33107 10845
rect 33174 10842 33180 10844
rect 29637 10840 33180 10842
rect 29637 10784 29642 10840
rect 29698 10784 33046 10840
rect 33102 10784 33180 10840
rect 29637 10782 33180 10784
rect 29637 10779 29703 10782
rect 33041 10779 33107 10782
rect 33174 10780 33180 10782
rect 33244 10780 33250 10844
rect 13077 10706 13143 10709
rect 19057 10706 19123 10709
rect 13077 10704 19123 10706
rect 13077 10648 13082 10704
rect 13138 10648 19062 10704
rect 19118 10648 19123 10704
rect 13077 10646 19123 10648
rect 13077 10643 13143 10646
rect 19057 10643 19123 10646
rect 24485 10436 24551 10437
rect 24485 10434 24532 10436
rect 24440 10432 24532 10434
rect 24440 10376 24490 10432
rect 24440 10374 24532 10376
rect 24485 10372 24532 10374
rect 24596 10372 24602 10436
rect 24485 10371 24551 10372
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 12934 10236 12940 10300
rect 13004 10298 13010 10300
rect 28993 10298 29059 10301
rect 13004 10296 29059 10298
rect 13004 10240 28998 10296
rect 29054 10240 29059 10296
rect 13004 10238 29059 10240
rect 13004 10236 13010 10238
rect 28993 10235 29059 10238
rect 27613 10162 27679 10165
rect 28533 10162 28599 10165
rect 27613 10160 28599 10162
rect 27613 10104 27618 10160
rect 27674 10104 28538 10160
rect 28594 10104 28599 10160
rect 27613 10102 28599 10104
rect 27613 10099 27679 10102
rect 28533 10099 28599 10102
rect 19425 10026 19491 10029
rect 22553 10026 22619 10029
rect 19425 10024 22619 10026
rect 19425 9968 19430 10024
rect 19486 9968 22558 10024
rect 22614 9968 22619 10024
rect 19425 9966 22619 9968
rect 19425 9963 19491 9966
rect 22553 9963 22619 9966
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 34278 9556 34284 9620
rect 34348 9618 34354 9620
rect 34605 9618 34671 9621
rect 34348 9616 34671 9618
rect 34348 9560 34610 9616
rect 34666 9560 34671 9616
rect 34348 9558 34671 9560
rect 34348 9556 34354 9558
rect 34605 9555 34671 9558
rect 37457 9618 37523 9621
rect 38878 9618 38884 9620
rect 37457 9616 38884 9618
rect 37457 9560 37462 9616
rect 37518 9560 38884 9616
rect 37457 9558 38884 9560
rect 37457 9555 37523 9558
rect 38878 9556 38884 9558
rect 38948 9556 38954 9620
rect 41597 9618 41663 9621
rect 41749 9618 42549 9648
rect 41597 9616 42549 9618
rect 41597 9560 41602 9616
rect 41658 9560 42549 9616
rect 41597 9558 42549 9560
rect 41597 9555 41663 9558
rect 41749 9528 42549 9558
rect 11605 9482 11671 9485
rect 12525 9482 12591 9485
rect 16941 9482 17007 9485
rect 11605 9480 17007 9482
rect 11605 9424 11610 9480
rect 11666 9424 12530 9480
rect 12586 9424 16946 9480
rect 17002 9424 17007 9480
rect 11605 9422 17007 9424
rect 11605 9419 11671 9422
rect 12525 9419 12591 9422
rect 16941 9419 17007 9422
rect 33961 9482 34027 9485
rect 35249 9482 35315 9485
rect 33961 9480 35315 9482
rect 33961 9424 33966 9480
rect 34022 9424 35254 9480
rect 35310 9424 35315 9480
rect 33961 9422 35315 9424
rect 33961 9419 34027 9422
rect 35249 9419 35315 9422
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 18086 9148 18092 9212
rect 18156 9210 18162 9212
rect 18413 9210 18479 9213
rect 18156 9208 18479 9210
rect 18156 9152 18418 9208
rect 18474 9152 18479 9208
rect 18156 9150 18479 9152
rect 18156 9148 18162 9150
rect 18413 9147 18479 9150
rect 30557 9210 30623 9213
rect 32765 9210 32831 9213
rect 30557 9208 32831 9210
rect 30557 9152 30562 9208
rect 30618 9152 32770 9208
rect 32826 9152 32831 9208
rect 30557 9150 32831 9152
rect 30557 9147 30623 9150
rect 32765 9147 32831 9150
rect 11237 9074 11303 9077
rect 11973 9074 12039 9077
rect 11237 9072 12039 9074
rect 11237 9016 11242 9072
rect 11298 9016 11978 9072
rect 12034 9016 12039 9072
rect 11237 9014 12039 9016
rect 11237 9011 11303 9014
rect 11973 9011 12039 9014
rect 11513 8802 11579 8805
rect 11973 8802 12039 8805
rect 11513 8800 12039 8802
rect 11513 8744 11518 8800
rect 11574 8744 11978 8800
rect 12034 8744 12039 8800
rect 11513 8742 12039 8744
rect 11513 8739 11579 8742
rect 11973 8739 12039 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 11513 8530 11579 8533
rect 14641 8530 14707 8533
rect 11513 8528 14707 8530
rect 11513 8472 11518 8528
rect 11574 8472 14646 8528
rect 14702 8472 14707 8528
rect 11513 8470 14707 8472
rect 11513 8467 11579 8470
rect 14641 8467 14707 8470
rect 18413 8530 18479 8533
rect 31293 8530 31359 8533
rect 31661 8530 31727 8533
rect 18413 8528 31727 8530
rect 18413 8472 18418 8528
rect 18474 8472 31298 8528
rect 31354 8472 31666 8528
rect 31722 8472 31727 8528
rect 18413 8470 31727 8472
rect 18413 8467 18479 8470
rect 31293 8467 31359 8470
rect 31661 8467 31727 8470
rect 32489 8394 32555 8397
rect 35893 8394 35959 8397
rect 32489 8392 35959 8394
rect 32489 8336 32494 8392
rect 32550 8336 35898 8392
rect 35954 8336 35959 8392
rect 32489 8334 35959 8336
rect 32489 8331 32555 8334
rect 35893 8331 35959 8334
rect 27429 8258 27495 8261
rect 28349 8258 28415 8261
rect 35617 8260 35683 8261
rect 27429 8256 28415 8258
rect 27429 8200 27434 8256
rect 27490 8200 28354 8256
rect 28410 8200 28415 8256
rect 27429 8198 28415 8200
rect 27429 8195 27495 8198
rect 28349 8195 28415 8198
rect 35566 8196 35572 8260
rect 35636 8258 35683 8260
rect 35636 8256 35728 8258
rect 35678 8200 35728 8256
rect 35636 8198 35728 8200
rect 35636 8196 35683 8198
rect 35617 8195 35683 8196
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 17534 8060 17540 8124
rect 17604 8122 17610 8124
rect 19057 8122 19123 8125
rect 17604 8120 19123 8122
rect 17604 8064 19062 8120
rect 19118 8064 19123 8120
rect 17604 8062 19123 8064
rect 17604 8060 17610 8062
rect 19057 8059 19123 8062
rect 30097 7986 30163 7989
rect 36077 7986 36143 7989
rect 30097 7984 36143 7986
rect 30097 7928 30102 7984
rect 30158 7928 36082 7984
rect 36138 7928 36143 7984
rect 30097 7926 36143 7928
rect 30097 7923 30163 7926
rect 36077 7923 36143 7926
rect 28165 7850 28231 7853
rect 31017 7850 31083 7853
rect 28165 7848 35450 7850
rect 28165 7792 28170 7848
rect 28226 7792 31022 7848
rect 31078 7792 35450 7848
rect 28165 7790 35450 7792
rect 28165 7787 28231 7790
rect 31017 7787 31083 7790
rect 19570 7648 19886 7649
rect 0 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 933 7578 999 7581
rect 0 7576 999 7578
rect 0 7520 938 7576
rect 994 7520 999 7576
rect 0 7518 999 7520
rect 0 7488 800 7518
rect 933 7515 999 7518
rect 30373 7578 30439 7581
rect 30373 7576 34898 7578
rect 30373 7520 30378 7576
rect 30434 7520 34898 7576
rect 30373 7518 34898 7520
rect 30373 7515 30439 7518
rect 28625 7442 28691 7445
rect 29729 7442 29795 7445
rect 33685 7442 33751 7445
rect 28625 7440 33751 7442
rect 28625 7384 28630 7440
rect 28686 7384 29734 7440
rect 29790 7384 33690 7440
rect 33746 7384 33751 7440
rect 28625 7382 33751 7384
rect 28625 7379 28691 7382
rect 29729 7379 29795 7382
rect 33685 7379 33751 7382
rect 12709 7306 12775 7309
rect 14457 7306 14523 7309
rect 15837 7306 15903 7309
rect 12709 7304 15903 7306
rect 12709 7248 12714 7304
rect 12770 7248 14462 7304
rect 14518 7248 15842 7304
rect 15898 7248 15903 7304
rect 12709 7246 15903 7248
rect 12709 7243 12775 7246
rect 14457 7243 14523 7246
rect 15837 7243 15903 7246
rect 20478 7244 20484 7308
rect 20548 7306 20554 7308
rect 20805 7306 20871 7309
rect 20548 7304 20871 7306
rect 20548 7248 20810 7304
rect 20866 7248 20871 7304
rect 20548 7246 20871 7248
rect 34838 7306 34898 7518
rect 35157 7442 35223 7445
rect 35390 7442 35450 7790
rect 35617 7442 35683 7445
rect 35157 7440 35683 7442
rect 35157 7384 35162 7440
rect 35218 7384 35622 7440
rect 35678 7384 35683 7440
rect 35157 7382 35683 7384
rect 35157 7379 35223 7382
rect 35617 7379 35683 7382
rect 35985 7306 36051 7309
rect 34838 7304 36051 7306
rect 34838 7248 35990 7304
rect 36046 7248 36051 7304
rect 34838 7246 36051 7248
rect 20548 7244 20554 7246
rect 20805 7243 20871 7246
rect 35985 7243 36051 7246
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 12617 6898 12683 6901
rect 15009 6898 15075 6901
rect 12617 6896 15075 6898
rect 12617 6840 12622 6896
rect 12678 6840 15014 6896
rect 15070 6840 15075 6896
rect 12617 6838 15075 6840
rect 12617 6835 12683 6838
rect 15009 6835 15075 6838
rect 33317 6898 33383 6901
rect 35801 6898 35867 6901
rect 33317 6896 35867 6898
rect 33317 6840 33322 6896
rect 33378 6840 35806 6896
rect 35862 6840 35867 6896
rect 33317 6838 35867 6840
rect 33317 6835 33383 6838
rect 35801 6835 35867 6838
rect 13629 6762 13695 6765
rect 15377 6762 15443 6765
rect 13629 6760 15443 6762
rect 13629 6704 13634 6760
rect 13690 6704 15382 6760
rect 15438 6704 15443 6760
rect 13629 6702 15443 6704
rect 13629 6699 13695 6702
rect 15377 6699 15443 6702
rect 33317 6762 33383 6765
rect 35433 6762 35499 6765
rect 33317 6760 35499 6762
rect 33317 6704 33322 6760
rect 33378 6704 35438 6760
rect 35494 6704 35499 6760
rect 33317 6702 35499 6704
rect 33317 6699 33383 6702
rect 35433 6699 35499 6702
rect 30373 6626 30439 6629
rect 33961 6626 34027 6629
rect 30373 6624 34027 6626
rect 30373 6568 30378 6624
rect 30434 6568 33966 6624
rect 34022 6568 34027 6624
rect 30373 6566 34027 6568
rect 30373 6563 30439 6566
rect 33961 6563 34027 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 12566 5612 12572 5676
rect 12636 5674 12642 5676
rect 17125 5674 17191 5677
rect 12636 5672 17191 5674
rect 12636 5616 17130 5672
rect 17186 5616 17191 5672
rect 12636 5614 17191 5616
rect 12636 5612 12642 5614
rect 17125 5611 17191 5614
rect 32581 5674 32647 5677
rect 35709 5674 35775 5677
rect 32581 5672 35775 5674
rect 32581 5616 32586 5672
rect 32642 5616 35714 5672
rect 35770 5616 35775 5672
rect 32581 5614 35775 5616
rect 32581 5611 32647 5614
rect 35709 5611 35775 5614
rect 16941 5540 17007 5541
rect 16941 5538 16988 5540
rect 16896 5536 16988 5538
rect 16896 5480 16946 5536
rect 16896 5478 16988 5480
rect 16941 5476 16988 5478
rect 17052 5476 17058 5540
rect 27470 5476 27476 5540
rect 27540 5538 27546 5540
rect 27705 5538 27771 5541
rect 27540 5536 27771 5538
rect 27540 5480 27710 5536
rect 27766 5480 27771 5536
rect 27540 5478 27771 5480
rect 27540 5476 27546 5478
rect 16941 5475 17007 5476
rect 27705 5475 27771 5478
rect 35985 5538 36051 5541
rect 36302 5538 36308 5540
rect 35985 5536 36308 5538
rect 35985 5480 35990 5536
rect 36046 5480 36308 5536
rect 35985 5478 36308 5480
rect 35985 5475 36051 5478
rect 36302 5476 36308 5478
rect 36372 5476 36378 5540
rect 41321 5538 41387 5541
rect 41749 5538 42549 5568
rect 41321 5536 42549 5538
rect 41321 5480 41326 5536
rect 41382 5480 42549 5536
rect 41321 5478 42549 5480
rect 41321 5475 41387 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 41749 5448 42549 5478
rect 19570 5407 19886 5408
rect 31661 5402 31727 5405
rect 34329 5402 34395 5405
rect 31661 5400 34395 5402
rect 31661 5344 31666 5400
rect 31722 5344 34334 5400
rect 34390 5344 34395 5400
rect 31661 5342 34395 5344
rect 31661 5339 31727 5342
rect 34329 5339 34395 5342
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 15009 4044 15075 4045
rect 14958 4042 14964 4044
rect 14918 3982 14964 4042
rect 15028 4040 15075 4044
rect 15070 3984 15075 4040
rect 14958 3980 14964 3982
rect 15028 3980 15075 3984
rect 15009 3979 15075 3980
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 14733 3634 14799 3637
rect 18638 3634 18644 3636
rect 14733 3632 18644 3634
rect 14733 3576 14738 3632
rect 14794 3576 18644 3632
rect 14733 3574 18644 3576
rect 14733 3571 14799 3574
rect 18638 3572 18644 3574
rect 18708 3572 18714 3636
rect 0 3498 800 3528
rect 933 3498 999 3501
rect 0 3496 999 3498
rect 0 3440 938 3496
rect 994 3440 999 3496
rect 0 3438 999 3440
rect 0 3408 800 3438
rect 933 3435 999 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 41749 1368 42549 1488
<< via3 >>
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 17724 42196 17788 42260
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 31340 41440 31404 41444
rect 31340 41384 31354 41440
rect 31354 41384 31404 41440
rect 31340 41380 31404 41384
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 17356 37300 17420 37364
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 31892 36076 31956 36140
rect 28764 35940 28828 36004
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 10916 35532 10980 35596
rect 29132 35532 29196 35596
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 22692 34988 22756 35052
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 20116 34716 20180 34780
rect 24532 34640 24596 34644
rect 24532 34584 24582 34640
rect 24582 34584 24596 34640
rect 24532 34580 24596 34584
rect 28948 34580 29012 34644
rect 29868 34640 29932 34644
rect 29868 34584 29918 34640
rect 29918 34584 29932 34640
rect 29868 34580 29932 34584
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 34652 34172 34716 34236
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 26740 33280 26804 33284
rect 26740 33224 26754 33280
rect 26754 33224 26804 33280
rect 26740 33220 26804 33224
rect 32444 33220 32508 33284
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 11836 32812 11900 32876
rect 20484 32812 20548 32876
rect 34468 32676 34532 32740
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 28028 32600 28092 32604
rect 28028 32544 28042 32600
rect 28042 32544 28092 32600
rect 28028 32540 28092 32544
rect 15884 32268 15948 32332
rect 30604 32192 30668 32196
rect 30604 32136 30654 32192
rect 30654 32136 30668 32192
rect 30604 32132 30668 32136
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 35940 31920 36004 31924
rect 35940 31864 35990 31920
rect 35990 31864 36004 31920
rect 35940 31860 36004 31864
rect 23244 31648 23308 31652
rect 23244 31592 23294 31648
rect 23294 31592 23308 31648
rect 23244 31588 23308 31592
rect 35388 31784 35452 31788
rect 35388 31728 35402 31784
rect 35402 31728 35452 31784
rect 35388 31724 35452 31728
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 22324 31240 22388 31244
rect 22324 31184 22338 31240
rect 22338 31184 22388 31240
rect 22324 31180 22388 31184
rect 32260 31044 32324 31108
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 16988 30908 17052 30972
rect 24900 30908 24964 30972
rect 17540 30636 17604 30700
rect 12020 30560 12084 30564
rect 12020 30504 12034 30560
rect 12034 30504 12084 30560
rect 12020 30500 12084 30504
rect 13676 30500 13740 30564
rect 26188 30500 26252 30564
rect 28580 30500 28644 30564
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 11100 30364 11164 30428
rect 12756 30424 12820 30428
rect 12756 30368 12770 30424
rect 12770 30368 12820 30424
rect 12756 30364 12820 30368
rect 25820 30424 25884 30428
rect 25820 30368 25870 30424
rect 25870 30368 25884 30424
rect 25820 30364 25884 30368
rect 33548 30364 33612 30428
rect 24348 30152 24412 30156
rect 24348 30096 24398 30152
rect 24398 30096 24412 30152
rect 24348 30092 24412 30096
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 18092 29684 18156 29748
rect 29868 29684 29932 29748
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 35388 29684 35452 29748
rect 9812 29412 9876 29476
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 31524 29276 31588 29340
rect 22140 29004 22204 29068
rect 25084 29004 25148 29068
rect 28396 29004 28460 29068
rect 30236 29004 30300 29068
rect 34100 29064 34164 29068
rect 34100 29008 34114 29064
rect 34114 29008 34164 29064
rect 34100 29004 34164 29008
rect 35388 29004 35452 29068
rect 37412 29064 37476 29068
rect 37412 29008 37426 29064
rect 37426 29008 37476 29064
rect 27292 28868 27356 28932
rect 37412 29004 37476 29008
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 22692 28732 22756 28796
rect 27844 28732 27908 28796
rect 23428 28596 23492 28660
rect 28212 28596 28276 28660
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 36860 28732 36924 28796
rect 20852 28460 20916 28524
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 34284 28460 34348 28524
rect 26740 28384 26804 28388
rect 26740 28328 26754 28384
rect 26754 28328 26804 28384
rect 26740 28324 26804 28328
rect 28948 28188 29012 28252
rect 31340 28188 31404 28252
rect 22324 27916 22388 27980
rect 24900 27916 24964 27980
rect 20852 27780 20916 27844
rect 24716 27780 24780 27844
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19380 27644 19444 27708
rect 20852 27704 20916 27708
rect 20852 27648 20866 27704
rect 20866 27648 20916 27704
rect 20852 27644 20916 27648
rect 26372 27644 26436 27708
rect 28028 27644 28092 27708
rect 29132 27644 29196 27708
rect 34468 27644 34532 27708
rect 39068 27644 39132 27708
rect 10916 27372 10980 27436
rect 24348 27508 24412 27572
rect 30972 27508 31036 27572
rect 21956 27296 22020 27300
rect 21956 27240 21970 27296
rect 21970 27240 22020 27296
rect 21956 27236 22020 27240
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 9812 27160 9876 27164
rect 9812 27104 9826 27160
rect 9826 27104 9876 27160
rect 9812 27100 9876 27104
rect 12572 27160 12636 27164
rect 12572 27104 12586 27160
rect 12586 27104 12636 27160
rect 12572 27100 12636 27104
rect 13676 27100 13740 27164
rect 16252 27160 16316 27164
rect 16252 27104 16302 27160
rect 16302 27104 16316 27160
rect 16252 27100 16316 27104
rect 35940 27100 36004 27164
rect 39252 27100 39316 27164
rect 9076 26752 9140 26756
rect 9076 26696 9126 26752
rect 9126 26696 9140 26752
rect 9076 26692 9140 26696
rect 15884 26692 15948 26756
rect 26188 26692 26252 26756
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19196 26556 19260 26620
rect 25268 26420 25332 26484
rect 10364 26344 10428 26348
rect 10364 26288 10378 26344
rect 10378 26288 10428 26344
rect 10364 26284 10428 26288
rect 11468 26344 11532 26348
rect 11468 26288 11482 26344
rect 11482 26288 11532 26344
rect 11468 26284 11532 26288
rect 16436 26284 16500 26348
rect 29500 26344 29564 26348
rect 29500 26288 29514 26344
rect 29514 26288 29564 26344
rect 29500 26284 29564 26288
rect 34468 26344 34532 26348
rect 34468 26288 34482 26344
rect 34482 26288 34532 26344
rect 34468 26284 34532 26288
rect 35756 26284 35820 26348
rect 28028 26208 28092 26212
rect 28028 26152 28042 26208
rect 28042 26152 28092 26208
rect 28028 26148 28092 26152
rect 31524 26148 31588 26212
rect 34652 26148 34716 26212
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 14780 25740 14844 25804
rect 20300 25604 20364 25668
rect 28212 25604 28276 25668
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 34284 25332 34348 25396
rect 37596 25332 37660 25396
rect 9812 25196 9876 25260
rect 18276 25196 18340 25260
rect 21220 25120 21284 25124
rect 21220 25064 21234 25120
rect 21234 25064 21284 25120
rect 21220 25060 21284 25064
rect 21956 25120 22020 25124
rect 21956 25064 22006 25120
rect 22006 25064 22020 25120
rect 21956 25060 22020 25064
rect 24532 25060 24596 25124
rect 29868 25060 29932 25124
rect 33364 25120 33428 25124
rect 33364 25064 33414 25120
rect 33414 25064 33428 25120
rect 33364 25060 33428 25064
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 9260 24984 9324 24988
rect 9260 24928 9274 24984
rect 9274 24928 9324 24984
rect 9260 24924 9324 24928
rect 13860 24924 13924 24988
rect 24900 24924 24964 24988
rect 37044 24984 37108 24988
rect 37044 24928 37094 24984
rect 37094 24928 37108 24984
rect 37044 24924 37108 24928
rect 12940 24576 13004 24580
rect 12940 24520 12990 24576
rect 12990 24520 13004 24576
rect 12940 24516 13004 24520
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 30052 24380 30116 24444
rect 30604 24440 30668 24444
rect 30604 24384 30618 24440
rect 30618 24384 30668 24440
rect 30604 24380 30668 24384
rect 20484 24244 20548 24308
rect 30604 24244 30668 24308
rect 27108 24108 27172 24172
rect 30236 24108 30300 24172
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 26556 23972 26620 24036
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 37596 23836 37660 23900
rect 25820 23700 25884 23764
rect 18644 23564 18708 23628
rect 23796 23564 23860 23628
rect 25084 23564 25148 23628
rect 26740 23564 26804 23628
rect 31524 23564 31588 23628
rect 11836 23428 11900 23492
rect 12572 23488 12636 23492
rect 12572 23432 12586 23488
rect 12586 23432 12636 23488
rect 12572 23428 12636 23432
rect 25636 23428 25700 23492
rect 26924 23428 26988 23492
rect 28580 23488 28644 23492
rect 28580 23432 28594 23488
rect 28594 23432 28644 23488
rect 28580 23428 28644 23432
rect 37228 23428 37292 23492
rect 37780 23488 37844 23492
rect 37780 23432 37794 23488
rect 37794 23432 37844 23488
rect 37780 23428 37844 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 23244 23156 23308 23220
rect 24716 23292 24780 23356
rect 5396 22884 5460 22948
rect 26372 22884 26436 22948
rect 29500 22884 29564 22948
rect 36124 22944 36188 22948
rect 36124 22888 36174 22944
rect 36174 22888 36188 22944
rect 36124 22884 36188 22888
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 23612 22748 23676 22812
rect 25820 22612 25884 22676
rect 35940 22612 36004 22676
rect 32260 22476 32324 22540
rect 34652 22476 34716 22540
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 20668 22068 20732 22132
rect 9076 21932 9140 21996
rect 12940 21992 13004 21996
rect 12940 21936 12954 21992
rect 12954 21936 13004 21992
rect 12940 21932 13004 21936
rect 13860 21932 13924 21996
rect 17540 21932 17604 21996
rect 22508 21992 22572 21996
rect 30052 22068 30116 22132
rect 30972 22068 31036 22132
rect 22508 21936 22522 21992
rect 22522 21936 22572 21992
rect 22508 21932 22572 21936
rect 24532 21932 24596 21996
rect 25636 21932 25700 21996
rect 26004 21992 26068 21996
rect 26004 21936 26018 21992
rect 26018 21936 26068 21992
rect 26004 21932 26068 21936
rect 21036 21796 21100 21860
rect 31708 21796 31772 21860
rect 36124 21796 36188 21860
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 34468 21660 34532 21724
rect 19380 21388 19444 21452
rect 21220 21252 21284 21316
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 9260 21116 9324 21180
rect 18276 21116 18340 21180
rect 27292 20980 27356 21044
rect 22876 20844 22940 20908
rect 16252 20768 16316 20772
rect 16252 20712 16266 20768
rect 16266 20712 16316 20768
rect 16252 20708 16316 20712
rect 33364 20708 33428 20772
rect 38884 20768 38948 20772
rect 38884 20712 38898 20768
rect 38898 20712 38948 20768
rect 38884 20708 38948 20712
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 23428 20572 23492 20636
rect 29500 20572 29564 20636
rect 32444 20436 32508 20500
rect 19196 20300 19260 20364
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 14780 20088 14844 20092
rect 14780 20032 14794 20088
rect 14794 20032 14844 20088
rect 14780 20028 14844 20032
rect 23612 19892 23676 19956
rect 28028 19620 28092 19684
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 29132 19544 29196 19548
rect 29132 19488 29182 19544
rect 29182 19488 29196 19544
rect 29132 19484 29196 19488
rect 30604 19544 30668 19548
rect 30604 19488 30654 19544
rect 30654 19488 30668 19544
rect 30604 19484 30668 19488
rect 17540 19408 17604 19412
rect 17540 19352 17554 19408
rect 17554 19352 17604 19408
rect 17540 19348 17604 19352
rect 24532 19408 24596 19412
rect 24532 19352 24582 19408
rect 24582 19352 24596 19408
rect 24532 19348 24596 19352
rect 33732 19348 33796 19412
rect 11468 19212 11532 19276
rect 20852 19212 20916 19276
rect 31524 19212 31588 19276
rect 14964 19076 15028 19140
rect 17908 19076 17972 19140
rect 21404 19076 21468 19140
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 33916 19076 33980 19140
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 25268 18940 25332 19004
rect 26740 18940 26804 19004
rect 35388 18668 35452 18732
rect 20852 18532 20916 18596
rect 22508 18532 22572 18596
rect 36860 18532 36924 18596
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 34100 18396 34164 18460
rect 36308 18396 36372 18460
rect 17356 18260 17420 18324
rect 15884 18124 15948 18188
rect 33548 18124 33612 18188
rect 35388 18124 35452 18188
rect 20668 18048 20732 18052
rect 20668 17992 20718 18048
rect 20718 17992 20732 18048
rect 20668 17988 20732 17992
rect 24900 17988 24964 18052
rect 33180 17988 33244 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 23796 17852 23860 17916
rect 27108 17852 27172 17916
rect 33732 17716 33796 17780
rect 24348 17444 24412 17508
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 21036 17308 21100 17372
rect 29868 17308 29932 17372
rect 16436 17172 16500 17236
rect 28580 17036 28644 17100
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 23612 16688 23676 16692
rect 23612 16632 23626 16688
rect 23626 16632 23676 16688
rect 23612 16628 23676 16632
rect 10916 16492 10980 16556
rect 26004 16492 26068 16556
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 34284 16628 34348 16692
rect 34468 16552 34532 16556
rect 34468 16496 34482 16552
rect 34482 16496 34532 16552
rect 34468 16492 34532 16496
rect 35756 16492 35820 16556
rect 35572 16356 35636 16420
rect 36124 16356 36188 16420
rect 37228 16144 37292 16148
rect 37228 16088 37278 16144
rect 37278 16088 37292 16144
rect 37228 16084 37292 16088
rect 22876 15948 22940 16012
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 22140 15736 22204 15740
rect 22140 15680 22190 15736
rect 22190 15680 22204 15736
rect 22140 15676 22204 15680
rect 33916 15268 33980 15332
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 5396 15192 5460 15196
rect 5396 15136 5410 15192
rect 5410 15136 5460 15192
rect 5396 15132 5460 15136
rect 20300 15132 20364 15196
rect 24900 15132 24964 15196
rect 25820 15192 25884 15196
rect 25820 15136 25834 15192
rect 25834 15136 25884 15192
rect 25820 15132 25884 15136
rect 26924 15192 26988 15196
rect 26924 15136 26938 15192
rect 26938 15136 26988 15192
rect 26924 15132 26988 15136
rect 28212 15132 28276 15196
rect 28764 15132 28828 15196
rect 30236 15132 30300 15196
rect 37596 15192 37660 15196
rect 37596 15136 37610 15192
rect 37610 15136 37660 15192
rect 37596 15132 37660 15136
rect 20116 14996 20180 15060
rect 21036 14724 21100 14788
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 35388 14784 35452 14788
rect 35388 14728 35438 14784
rect 35438 14728 35452 14784
rect 35388 14724 35452 14728
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 37780 14316 37844 14380
rect 37044 14240 37108 14244
rect 37044 14184 37094 14240
rect 37094 14184 37108 14240
rect 37044 14180 37108 14184
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 34652 14044 34716 14108
rect 20852 13908 20916 13972
rect 17540 13772 17604 13836
rect 32996 13772 33060 13836
rect 24716 13636 24780 13700
rect 26556 13636 26620 13700
rect 37412 13636 37476 13700
rect 39068 13696 39132 13700
rect 39068 13640 39082 13696
rect 39082 13640 39132 13696
rect 39068 13636 39132 13640
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 27476 13560 27540 13564
rect 27476 13504 27490 13560
rect 27490 13504 27540 13560
rect 27476 13500 27540 13504
rect 39252 13500 39316 13564
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 11100 12064 11164 12068
rect 11100 12008 11114 12064
rect 11114 12008 11164 12064
rect 11100 12004 11164 12008
rect 35940 12064 36004 12068
rect 35940 12008 35990 12064
rect 35990 12008 36004 12064
rect 35940 12004 36004 12008
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 34468 11792 34532 11796
rect 34468 11736 34482 11792
rect 34482 11736 34532 11792
rect 34468 11732 34532 11736
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 12020 10976 12084 10980
rect 12020 10920 12034 10976
rect 12034 10920 12084 10976
rect 12020 10916 12084 10920
rect 21404 10916 21468 10980
rect 29500 10916 29564 10980
rect 32996 10916 33060 10980
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 10364 10780 10428 10844
rect 17724 10780 17788 10844
rect 33180 10780 33244 10844
rect 24532 10432 24596 10436
rect 24532 10376 24546 10432
rect 24546 10376 24596 10432
rect 24532 10372 24596 10376
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 12940 10236 13004 10300
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 34284 9556 34348 9620
rect 38884 9556 38948 9620
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 18092 9148 18156 9212
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 35572 8256 35636 8260
rect 35572 8200 35622 8256
rect 35622 8200 35636 8256
rect 35572 8196 35636 8200
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 17540 8060 17604 8124
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 20484 7244 20548 7308
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 12572 5612 12636 5676
rect 16988 5536 17052 5540
rect 16988 5480 17002 5536
rect 17002 5480 17052 5536
rect 16988 5476 17052 5480
rect 27476 5476 27540 5540
rect 36308 5476 36372 5540
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 14964 4040 15028 4044
rect 14964 3984 15014 4040
rect 15014 3984 15028 4040
rect 14964 3980 15028 3984
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 18644 3572 18708 3636
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 41920 4528 42480
rect 19568 42464 19888 42480
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 17723 42260 17789 42261
rect 17723 42196 17724 42260
rect 17788 42196 17789 42260
rect 17723 42195 17789 42196
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 17355 37364 17421 37365
rect 17355 37300 17356 37364
rect 17420 37300 17421 37364
rect 17355 37299 17421 37300
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 10915 35596 10981 35597
rect 10915 35532 10916 35596
rect 10980 35532 10981 35596
rect 10915 35531 10981 35532
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 9811 29476 9877 29477
rect 9811 29412 9812 29476
rect 9876 29412 9877 29476
rect 9811 29411 9877 29412
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 9814 27165 9874 29411
rect 10918 27437 10978 35531
rect 11835 32876 11901 32877
rect 11835 32812 11836 32876
rect 11900 32812 11901 32876
rect 11835 32811 11901 32812
rect 11099 30428 11165 30429
rect 11099 30364 11100 30428
rect 11164 30364 11165 30428
rect 11099 30363 11165 30364
rect 10915 27436 10981 27437
rect 10915 27372 10916 27436
rect 10980 27372 10981 27436
rect 10915 27371 10981 27372
rect 9811 27164 9877 27165
rect 9811 27100 9812 27164
rect 9876 27100 9877 27164
rect 9811 27099 9877 27100
rect 9075 26756 9141 26757
rect 9075 26692 9076 26756
rect 9140 26692 9141 26756
rect 9075 26691 9141 26692
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 5395 22948 5461 22949
rect 5395 22884 5396 22948
rect 5460 22884 5461 22948
rect 5395 22883 5461 22884
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 5398 15197 5458 22883
rect 9078 21997 9138 26691
rect 9814 25261 9874 27099
rect 10363 26348 10429 26349
rect 10363 26284 10364 26348
rect 10428 26284 10429 26348
rect 10363 26283 10429 26284
rect 9811 25260 9877 25261
rect 9811 25196 9812 25260
rect 9876 25196 9877 25260
rect 9811 25195 9877 25196
rect 9259 24988 9325 24989
rect 9259 24924 9260 24988
rect 9324 24924 9325 24988
rect 9259 24923 9325 24924
rect 9075 21996 9141 21997
rect 9075 21932 9076 21996
rect 9140 21932 9141 21996
rect 9075 21931 9141 21932
rect 9262 21181 9322 24923
rect 9259 21180 9325 21181
rect 9259 21116 9260 21180
rect 9324 21116 9325 21180
rect 9259 21115 9325 21116
rect 5395 15196 5461 15197
rect 5395 15132 5396 15196
rect 5460 15132 5461 15196
rect 5395 15131 5461 15132
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 10366 10845 10426 26283
rect 10918 16557 10978 27371
rect 10915 16556 10981 16557
rect 10915 16492 10916 16556
rect 10980 16492 10981 16556
rect 10915 16491 10981 16492
rect 11102 12069 11162 30363
rect 11467 26348 11533 26349
rect 11467 26284 11468 26348
rect 11532 26284 11533 26348
rect 11467 26283 11533 26284
rect 11470 19277 11530 26283
rect 11838 23493 11898 32811
rect 15883 32332 15949 32333
rect 15883 32268 15884 32332
rect 15948 32268 15949 32332
rect 15883 32267 15949 32268
rect 12019 30564 12085 30565
rect 12019 30500 12020 30564
rect 12084 30500 12085 30564
rect 12019 30499 12085 30500
rect 13675 30564 13741 30565
rect 13675 30500 13676 30564
rect 13740 30500 13741 30564
rect 13675 30499 13741 30500
rect 11835 23492 11901 23493
rect 11835 23428 11836 23492
rect 11900 23428 11901 23492
rect 11835 23427 11901 23428
rect 11467 19276 11533 19277
rect 11467 19212 11468 19276
rect 11532 19212 11533 19276
rect 11467 19211 11533 19212
rect 11099 12068 11165 12069
rect 11099 12004 11100 12068
rect 11164 12004 11165 12068
rect 11099 12003 11165 12004
rect 12022 10981 12082 30499
rect 12755 30428 12821 30429
rect 12755 30364 12756 30428
rect 12820 30364 12821 30428
rect 12755 30363 12821 30364
rect 12571 27164 12637 27165
rect 12571 27100 12572 27164
rect 12636 27100 12637 27164
rect 12571 27099 12637 27100
rect 12574 23493 12634 27099
rect 12571 23492 12637 23493
rect 12571 23428 12572 23492
rect 12636 23428 12637 23492
rect 12571 23427 12637 23428
rect 12758 22110 12818 30363
rect 13678 27165 13738 30499
rect 13675 27164 13741 27165
rect 13675 27100 13676 27164
rect 13740 27100 13741 27164
rect 13675 27099 13741 27100
rect 15886 26757 15946 32267
rect 16987 30972 17053 30973
rect 16987 30908 16988 30972
rect 17052 30908 17053 30972
rect 16987 30907 17053 30908
rect 16251 27164 16317 27165
rect 16251 27100 16252 27164
rect 16316 27100 16317 27164
rect 16251 27099 16317 27100
rect 15883 26756 15949 26757
rect 15883 26692 15884 26756
rect 15948 26692 15949 26756
rect 15883 26691 15949 26692
rect 14779 25804 14845 25805
rect 14779 25740 14780 25804
rect 14844 25740 14845 25804
rect 14779 25739 14845 25740
rect 13859 24988 13925 24989
rect 13859 24924 13860 24988
rect 13924 24924 13925 24988
rect 13859 24923 13925 24924
rect 12939 24580 13005 24581
rect 12939 24516 12940 24580
rect 13004 24516 13005 24580
rect 12939 24515 13005 24516
rect 12574 22050 12818 22110
rect 12019 10980 12085 10981
rect 12019 10916 12020 10980
rect 12084 10916 12085 10980
rect 12019 10915 12085 10916
rect 10363 10844 10429 10845
rect 10363 10780 10364 10844
rect 10428 10780 10429 10844
rect 10363 10779 10429 10780
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 12574 5677 12634 22050
rect 12942 21997 13002 24515
rect 13862 21997 13922 24923
rect 12939 21996 13005 21997
rect 12939 21932 12940 21996
rect 13004 21932 13005 21996
rect 12939 21931 13005 21932
rect 13859 21996 13925 21997
rect 13859 21932 13860 21996
rect 13924 21932 13925 21996
rect 13859 21931 13925 21932
rect 12942 10301 13002 21931
rect 14782 20093 14842 25739
rect 14779 20092 14845 20093
rect 14779 20028 14780 20092
rect 14844 20028 14845 20092
rect 14779 20027 14845 20028
rect 14963 19140 15029 19141
rect 14963 19076 14964 19140
rect 15028 19076 15029 19140
rect 14963 19075 15029 19076
rect 12939 10300 13005 10301
rect 12939 10236 12940 10300
rect 13004 10236 13005 10300
rect 12939 10235 13005 10236
rect 12571 5676 12637 5677
rect 12571 5612 12572 5676
rect 12636 5612 12637 5676
rect 12571 5611 12637 5612
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 14966 4045 15026 19075
rect 15886 18189 15946 26691
rect 16254 20773 16314 27099
rect 16435 26348 16501 26349
rect 16435 26284 16436 26348
rect 16500 26284 16501 26348
rect 16435 26283 16501 26284
rect 16251 20772 16317 20773
rect 16251 20708 16252 20772
rect 16316 20708 16317 20772
rect 16251 20707 16317 20708
rect 15883 18188 15949 18189
rect 15883 18124 15884 18188
rect 15948 18124 15949 18188
rect 15883 18123 15949 18124
rect 16438 17237 16498 26283
rect 16435 17236 16501 17237
rect 16435 17172 16436 17236
rect 16500 17172 16501 17236
rect 16435 17171 16501 17172
rect 16990 5541 17050 30907
rect 17358 18325 17418 37299
rect 17726 31770 17786 42195
rect 19568 41376 19888 42400
rect 34928 41920 35248 42480
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 31339 41444 31405 41445
rect 31339 41380 31340 41444
rect 31404 41380 31405 41444
rect 31339 41379 31405 41380
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 28763 36004 28829 36005
rect 28763 35940 28764 36004
rect 28828 35940 28829 36004
rect 28763 35939 28829 35940
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 22691 35052 22757 35053
rect 22691 34988 22692 35052
rect 22756 34988 22757 35052
rect 22691 34987 22757 34988
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 20115 34780 20181 34781
rect 20115 34716 20116 34780
rect 20180 34716 20181 34780
rect 20115 34715 20181 34716
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 17726 31710 17970 31770
rect 17539 30700 17605 30701
rect 17539 30636 17540 30700
rect 17604 30636 17605 30700
rect 17539 30635 17605 30636
rect 17542 21997 17602 30635
rect 17539 21996 17605 21997
rect 17539 21932 17540 21996
rect 17604 21932 17605 21996
rect 17539 21931 17605 21932
rect 17542 20090 17602 21931
rect 17542 20030 17786 20090
rect 17539 19412 17605 19413
rect 17539 19348 17540 19412
rect 17604 19348 17605 19412
rect 17539 19347 17605 19348
rect 17355 18324 17421 18325
rect 17355 18260 17356 18324
rect 17420 18260 17421 18324
rect 17355 18259 17421 18260
rect 17542 13837 17602 19347
rect 17539 13836 17605 13837
rect 17539 13772 17540 13836
rect 17604 13772 17605 13836
rect 17539 13771 17605 13772
rect 17542 8125 17602 13771
rect 17726 10845 17786 20030
rect 17910 19141 17970 31710
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 18091 29748 18157 29749
rect 18091 29684 18092 29748
rect 18156 29684 18157 29748
rect 18091 29683 18157 29684
rect 17907 19140 17973 19141
rect 17907 19076 17908 19140
rect 17972 19076 17973 19140
rect 17907 19075 17973 19076
rect 17723 10844 17789 10845
rect 17723 10780 17724 10844
rect 17788 10780 17789 10844
rect 17723 10779 17789 10780
rect 18094 9213 18154 29683
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19379 27708 19445 27709
rect 19379 27644 19380 27708
rect 19444 27644 19445 27708
rect 19379 27643 19445 27644
rect 19195 26620 19261 26621
rect 19195 26556 19196 26620
rect 19260 26556 19261 26620
rect 19195 26555 19261 26556
rect 18275 25260 18341 25261
rect 18275 25196 18276 25260
rect 18340 25196 18341 25260
rect 18275 25195 18341 25196
rect 18278 21181 18338 25195
rect 18643 23628 18709 23629
rect 18643 23564 18644 23628
rect 18708 23564 18709 23628
rect 18643 23563 18709 23564
rect 18275 21180 18341 21181
rect 18275 21116 18276 21180
rect 18340 21116 18341 21180
rect 18275 21115 18341 21116
rect 18091 9212 18157 9213
rect 18091 9148 18092 9212
rect 18156 9148 18157 9212
rect 18091 9147 18157 9148
rect 17539 8124 17605 8125
rect 17539 8060 17540 8124
rect 17604 8060 17605 8124
rect 17539 8059 17605 8060
rect 16987 5540 17053 5541
rect 16987 5476 16988 5540
rect 17052 5476 17053 5540
rect 16987 5475 17053 5476
rect 14963 4044 15029 4045
rect 14963 3980 14964 4044
rect 15028 3980 15029 4044
rect 14963 3979 15029 3980
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 18646 3637 18706 23563
rect 19198 20365 19258 26555
rect 19382 21453 19442 27643
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19379 21452 19445 21453
rect 19379 21388 19380 21452
rect 19444 21388 19445 21452
rect 19379 21387 19445 21388
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19195 20364 19261 20365
rect 19195 20300 19196 20364
rect 19260 20300 19261 20364
rect 19195 20299 19261 20300
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 20118 15061 20178 34715
rect 20483 32876 20549 32877
rect 20483 32812 20484 32876
rect 20548 32812 20549 32876
rect 20483 32811 20549 32812
rect 20299 25668 20365 25669
rect 20299 25604 20300 25668
rect 20364 25604 20365 25668
rect 20299 25603 20365 25604
rect 20302 15197 20362 25603
rect 20486 24309 20546 32811
rect 22323 31244 22389 31245
rect 22323 31180 22324 31244
rect 22388 31180 22389 31244
rect 22323 31179 22389 31180
rect 22139 29068 22205 29069
rect 22139 29004 22140 29068
rect 22204 29004 22205 29068
rect 22139 29003 22205 29004
rect 20851 28524 20917 28525
rect 20851 28460 20852 28524
rect 20916 28460 20917 28524
rect 20851 28459 20917 28460
rect 20854 27845 20914 28459
rect 20851 27844 20917 27845
rect 20851 27780 20852 27844
rect 20916 27780 20917 27844
rect 20851 27779 20917 27780
rect 20851 27708 20917 27709
rect 20851 27644 20852 27708
rect 20916 27644 20917 27708
rect 20851 27643 20917 27644
rect 20483 24308 20549 24309
rect 20483 24244 20484 24308
rect 20548 24244 20549 24308
rect 20483 24243 20549 24244
rect 20299 15196 20365 15197
rect 20299 15132 20300 15196
rect 20364 15132 20365 15196
rect 20299 15131 20365 15132
rect 20115 15060 20181 15061
rect 20115 14996 20116 15060
rect 20180 14996 20181 15060
rect 20115 14995 20181 14996
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 20486 7309 20546 24243
rect 20667 22132 20733 22133
rect 20667 22068 20668 22132
rect 20732 22068 20733 22132
rect 20667 22067 20733 22068
rect 20670 18053 20730 22067
rect 20854 19277 20914 27643
rect 21955 27300 22021 27301
rect 21955 27236 21956 27300
rect 22020 27236 22021 27300
rect 21955 27235 22021 27236
rect 21958 25125 22018 27235
rect 21219 25124 21285 25125
rect 21219 25060 21220 25124
rect 21284 25060 21285 25124
rect 21219 25059 21285 25060
rect 21955 25124 22021 25125
rect 21955 25060 21956 25124
rect 22020 25060 22021 25124
rect 21955 25059 22021 25060
rect 21035 21860 21101 21861
rect 21035 21796 21036 21860
rect 21100 21796 21101 21860
rect 21035 21795 21101 21796
rect 20851 19276 20917 19277
rect 20851 19212 20852 19276
rect 20916 19212 20917 19276
rect 20851 19211 20917 19212
rect 20851 18596 20917 18597
rect 20851 18532 20852 18596
rect 20916 18532 20917 18596
rect 20851 18531 20917 18532
rect 20667 18052 20733 18053
rect 20667 17988 20668 18052
rect 20732 17988 20733 18052
rect 20667 17987 20733 17988
rect 20854 13973 20914 18531
rect 21038 17373 21098 21795
rect 21222 21317 21282 25059
rect 21219 21316 21285 21317
rect 21219 21252 21220 21316
rect 21284 21252 21285 21316
rect 21219 21251 21285 21252
rect 21403 19140 21469 19141
rect 21403 19076 21404 19140
rect 21468 19076 21469 19140
rect 21403 19075 21469 19076
rect 21035 17372 21101 17373
rect 21035 17308 21036 17372
rect 21100 17308 21101 17372
rect 21035 17307 21101 17308
rect 21038 14789 21098 17307
rect 21035 14788 21101 14789
rect 21035 14724 21036 14788
rect 21100 14724 21101 14788
rect 21035 14723 21101 14724
rect 20851 13972 20917 13973
rect 20851 13908 20852 13972
rect 20916 13908 20917 13972
rect 20851 13907 20917 13908
rect 21406 10981 21466 19075
rect 22142 15741 22202 29003
rect 22326 27981 22386 31179
rect 22694 28797 22754 34987
rect 24531 34644 24597 34645
rect 24531 34580 24532 34644
rect 24596 34580 24597 34644
rect 24531 34579 24597 34580
rect 23243 31652 23309 31653
rect 23243 31588 23244 31652
rect 23308 31588 23309 31652
rect 23243 31587 23309 31588
rect 22691 28796 22757 28797
rect 22691 28732 22692 28796
rect 22756 28732 22757 28796
rect 22691 28731 22757 28732
rect 22323 27980 22389 27981
rect 22323 27916 22324 27980
rect 22388 27916 22389 27980
rect 22323 27915 22389 27916
rect 23246 23221 23306 31587
rect 24347 30156 24413 30157
rect 24347 30092 24348 30156
rect 24412 30092 24413 30156
rect 24347 30091 24413 30092
rect 23427 28660 23493 28661
rect 23427 28596 23428 28660
rect 23492 28596 23493 28660
rect 23427 28595 23493 28596
rect 23243 23220 23309 23221
rect 23243 23156 23244 23220
rect 23308 23156 23309 23220
rect 23243 23155 23309 23156
rect 22507 21996 22573 21997
rect 22507 21932 22508 21996
rect 22572 21932 22573 21996
rect 22507 21931 22573 21932
rect 22510 18597 22570 21931
rect 22875 20908 22941 20909
rect 22875 20844 22876 20908
rect 22940 20844 22941 20908
rect 22875 20843 22941 20844
rect 22507 18596 22573 18597
rect 22507 18532 22508 18596
rect 22572 18532 22573 18596
rect 22507 18531 22573 18532
rect 22878 16013 22938 20843
rect 23430 20637 23490 28595
rect 24350 27573 24410 30091
rect 24347 27572 24413 27573
rect 24347 27508 24348 27572
rect 24412 27508 24413 27572
rect 24347 27507 24413 27508
rect 24534 25125 24594 34579
rect 26739 33284 26805 33285
rect 26739 33220 26740 33284
rect 26804 33220 26805 33284
rect 26739 33219 26805 33220
rect 24899 30972 24965 30973
rect 24899 30908 24900 30972
rect 24964 30908 24965 30972
rect 24899 30907 24965 30908
rect 24902 27981 24962 30907
rect 26187 30564 26253 30565
rect 26187 30500 26188 30564
rect 26252 30500 26253 30564
rect 26187 30499 26253 30500
rect 25819 30428 25885 30429
rect 25819 30364 25820 30428
rect 25884 30364 25885 30428
rect 25819 30363 25885 30364
rect 25083 29068 25149 29069
rect 25083 29004 25084 29068
rect 25148 29004 25149 29068
rect 25083 29003 25149 29004
rect 24899 27980 24965 27981
rect 24899 27916 24900 27980
rect 24964 27916 24965 27980
rect 24899 27915 24965 27916
rect 24715 27844 24781 27845
rect 24715 27780 24716 27844
rect 24780 27780 24781 27844
rect 24715 27779 24781 27780
rect 24531 25124 24597 25125
rect 24531 25060 24532 25124
rect 24596 25060 24597 25124
rect 24531 25059 24597 25060
rect 23795 23628 23861 23629
rect 23795 23564 23796 23628
rect 23860 23564 23861 23628
rect 23795 23563 23861 23564
rect 23611 22812 23677 22813
rect 23611 22748 23612 22812
rect 23676 22748 23677 22812
rect 23611 22747 23677 22748
rect 23427 20636 23493 20637
rect 23427 20572 23428 20636
rect 23492 20572 23493 20636
rect 23427 20571 23493 20572
rect 23614 19957 23674 22747
rect 23611 19956 23677 19957
rect 23611 19892 23612 19956
rect 23676 19892 23677 19956
rect 23611 19891 23677 19892
rect 23614 16693 23674 19891
rect 23798 17917 23858 23563
rect 24534 21997 24594 25059
rect 24718 23357 24778 27779
rect 24899 24988 24965 24989
rect 24899 24924 24900 24988
rect 24964 24924 24965 24988
rect 24899 24923 24965 24924
rect 24715 23356 24781 23357
rect 24715 23292 24716 23356
rect 24780 23292 24781 23356
rect 24715 23291 24781 23292
rect 24902 22110 24962 24923
rect 25086 23629 25146 29003
rect 25267 26484 25333 26485
rect 25267 26420 25268 26484
rect 25332 26420 25333 26484
rect 25267 26419 25333 26420
rect 25083 23628 25149 23629
rect 25083 23564 25084 23628
rect 25148 23564 25149 23628
rect 25083 23563 25149 23564
rect 24718 22050 24962 22110
rect 24531 21996 24597 21997
rect 24531 21994 24532 21996
rect 24350 21934 24532 21994
rect 23795 17916 23861 17917
rect 23795 17852 23796 17916
rect 23860 17852 23861 17916
rect 23795 17851 23861 17852
rect 24350 17509 24410 21934
rect 24531 21932 24532 21934
rect 24596 21932 24597 21996
rect 24531 21931 24597 21932
rect 24531 19412 24597 19413
rect 24531 19348 24532 19412
rect 24596 19348 24597 19412
rect 24531 19347 24597 19348
rect 24347 17508 24413 17509
rect 24347 17444 24348 17508
rect 24412 17444 24413 17508
rect 24347 17443 24413 17444
rect 23611 16692 23677 16693
rect 23611 16628 23612 16692
rect 23676 16628 23677 16692
rect 23611 16627 23677 16628
rect 22875 16012 22941 16013
rect 22875 15948 22876 16012
rect 22940 15948 22941 16012
rect 22875 15947 22941 15948
rect 22139 15740 22205 15741
rect 22139 15676 22140 15740
rect 22204 15676 22205 15740
rect 22139 15675 22205 15676
rect 21403 10980 21469 10981
rect 21403 10916 21404 10980
rect 21468 10916 21469 10980
rect 21403 10915 21469 10916
rect 24534 10437 24594 19347
rect 24718 13701 24778 22050
rect 25270 19005 25330 26419
rect 25822 23765 25882 30363
rect 26190 26757 26250 30499
rect 26742 28389 26802 33219
rect 28027 32604 28093 32605
rect 28027 32540 28028 32604
rect 28092 32540 28093 32604
rect 28027 32539 28093 32540
rect 27291 28932 27357 28933
rect 27291 28868 27292 28932
rect 27356 28868 27357 28932
rect 27291 28867 27357 28868
rect 26739 28388 26805 28389
rect 26739 28324 26740 28388
rect 26804 28324 26805 28388
rect 26739 28323 26805 28324
rect 26371 27708 26437 27709
rect 26371 27644 26372 27708
rect 26436 27644 26437 27708
rect 26371 27643 26437 27644
rect 26187 26756 26253 26757
rect 26187 26692 26188 26756
rect 26252 26692 26253 26756
rect 26187 26691 26253 26692
rect 25819 23764 25885 23765
rect 25819 23700 25820 23764
rect 25884 23700 25885 23764
rect 25819 23699 25885 23700
rect 25635 23492 25701 23493
rect 25635 23428 25636 23492
rect 25700 23428 25701 23492
rect 25635 23427 25701 23428
rect 25638 21997 25698 23427
rect 26374 22949 26434 27643
rect 27107 24172 27173 24173
rect 27107 24108 27108 24172
rect 27172 24108 27173 24172
rect 27107 24107 27173 24108
rect 26555 24036 26621 24037
rect 26555 23972 26556 24036
rect 26620 23972 26621 24036
rect 26555 23971 26621 23972
rect 26371 22948 26437 22949
rect 26371 22884 26372 22948
rect 26436 22884 26437 22948
rect 26371 22883 26437 22884
rect 25819 22676 25885 22677
rect 25819 22612 25820 22676
rect 25884 22612 25885 22676
rect 25819 22611 25885 22612
rect 25635 21996 25701 21997
rect 25635 21932 25636 21996
rect 25700 21932 25701 21996
rect 25635 21931 25701 21932
rect 25267 19004 25333 19005
rect 25267 18940 25268 19004
rect 25332 18940 25333 19004
rect 25267 18939 25333 18940
rect 24899 18052 24965 18053
rect 24899 17988 24900 18052
rect 24964 17988 24965 18052
rect 24899 17987 24965 17988
rect 24902 15197 24962 17987
rect 25822 15197 25882 22611
rect 26003 21996 26069 21997
rect 26003 21932 26004 21996
rect 26068 21932 26069 21996
rect 26003 21931 26069 21932
rect 26006 16557 26066 21931
rect 26003 16556 26069 16557
rect 26003 16492 26004 16556
rect 26068 16492 26069 16556
rect 26003 16491 26069 16492
rect 24899 15196 24965 15197
rect 24899 15132 24900 15196
rect 24964 15132 24965 15196
rect 24899 15131 24965 15132
rect 25819 15196 25885 15197
rect 25819 15132 25820 15196
rect 25884 15132 25885 15196
rect 25819 15131 25885 15132
rect 26558 13701 26618 23971
rect 26739 23628 26805 23629
rect 26739 23564 26740 23628
rect 26804 23564 26805 23628
rect 26739 23563 26805 23564
rect 26742 19005 26802 23563
rect 26923 23492 26989 23493
rect 26923 23428 26924 23492
rect 26988 23428 26989 23492
rect 26923 23427 26989 23428
rect 26739 19004 26805 19005
rect 26739 18940 26740 19004
rect 26804 18940 26805 19004
rect 26739 18939 26805 18940
rect 26926 15197 26986 23427
rect 27110 17917 27170 24107
rect 27294 21045 27354 28867
rect 27843 28796 27909 28797
rect 27843 28732 27844 28796
rect 27908 28732 27909 28796
rect 27843 28731 27909 28732
rect 27291 21044 27357 21045
rect 27291 20980 27292 21044
rect 27356 20980 27357 21044
rect 27291 20979 27357 20980
rect 27846 19350 27906 28731
rect 28030 27709 28090 32539
rect 28579 30564 28645 30565
rect 28579 30500 28580 30564
rect 28644 30500 28645 30564
rect 28579 30499 28645 30500
rect 28395 29068 28461 29069
rect 28395 29004 28396 29068
rect 28460 29004 28461 29068
rect 28395 29003 28461 29004
rect 28211 28660 28277 28661
rect 28211 28596 28212 28660
rect 28276 28596 28277 28660
rect 28211 28595 28277 28596
rect 28027 27708 28093 27709
rect 28027 27644 28028 27708
rect 28092 27644 28093 27708
rect 28027 27643 28093 27644
rect 28027 26212 28093 26213
rect 28027 26148 28028 26212
rect 28092 26148 28093 26212
rect 28027 26147 28093 26148
rect 28030 19685 28090 26147
rect 28214 25669 28274 28595
rect 28211 25668 28277 25669
rect 28211 25604 28212 25668
rect 28276 25604 28277 25668
rect 28211 25603 28277 25604
rect 28398 22110 28458 29003
rect 28582 23493 28642 30499
rect 28579 23492 28645 23493
rect 28579 23428 28580 23492
rect 28644 23428 28645 23492
rect 28579 23427 28645 23428
rect 28398 22050 28642 22110
rect 28027 19684 28093 19685
rect 28027 19620 28028 19684
rect 28092 19620 28093 19684
rect 28027 19619 28093 19620
rect 27846 19290 28274 19350
rect 27107 17916 27173 17917
rect 27107 17852 27108 17916
rect 27172 17852 27173 17916
rect 27107 17851 27173 17852
rect 28214 15197 28274 19290
rect 28582 17101 28642 22050
rect 28579 17100 28645 17101
rect 28579 17036 28580 17100
rect 28644 17036 28645 17100
rect 28579 17035 28645 17036
rect 28766 15197 28826 35939
rect 29131 35596 29197 35597
rect 29131 35532 29132 35596
rect 29196 35532 29197 35596
rect 29131 35531 29197 35532
rect 28947 34644 29013 34645
rect 28947 34580 28948 34644
rect 29012 34580 29013 34644
rect 28947 34579 29013 34580
rect 28950 28253 29010 34579
rect 28947 28252 29013 28253
rect 28947 28188 28948 28252
rect 29012 28188 29013 28252
rect 28947 28187 29013 28188
rect 29134 27709 29194 35531
rect 29867 34644 29933 34645
rect 29867 34580 29868 34644
rect 29932 34580 29933 34644
rect 29867 34579 29933 34580
rect 29870 29749 29930 34579
rect 30603 32196 30669 32197
rect 30603 32132 30604 32196
rect 30668 32132 30669 32196
rect 30603 32131 30669 32132
rect 29867 29748 29933 29749
rect 29867 29684 29868 29748
rect 29932 29684 29933 29748
rect 29867 29683 29933 29684
rect 30235 29068 30301 29069
rect 30235 29004 30236 29068
rect 30300 29004 30301 29068
rect 30235 29003 30301 29004
rect 29131 27708 29197 27709
rect 29131 27644 29132 27708
rect 29196 27644 29197 27708
rect 29131 27643 29197 27644
rect 29134 19549 29194 27643
rect 29499 26348 29565 26349
rect 29499 26284 29500 26348
rect 29564 26284 29565 26348
rect 29499 26283 29565 26284
rect 29502 22949 29562 26283
rect 29867 25124 29933 25125
rect 29867 25060 29868 25124
rect 29932 25060 29933 25124
rect 29867 25059 29933 25060
rect 29499 22948 29565 22949
rect 29499 22884 29500 22948
rect 29564 22884 29565 22948
rect 29499 22883 29565 22884
rect 29499 20636 29565 20637
rect 29499 20572 29500 20636
rect 29564 20572 29565 20636
rect 29499 20571 29565 20572
rect 29131 19548 29197 19549
rect 29131 19484 29132 19548
rect 29196 19484 29197 19548
rect 29131 19483 29197 19484
rect 26923 15196 26989 15197
rect 26923 15132 26924 15196
rect 26988 15132 26989 15196
rect 26923 15131 26989 15132
rect 28211 15196 28277 15197
rect 28211 15132 28212 15196
rect 28276 15132 28277 15196
rect 28211 15131 28277 15132
rect 28763 15196 28829 15197
rect 28763 15132 28764 15196
rect 28828 15132 28829 15196
rect 28763 15131 28829 15132
rect 24715 13700 24781 13701
rect 24715 13636 24716 13700
rect 24780 13636 24781 13700
rect 24715 13635 24781 13636
rect 26555 13700 26621 13701
rect 26555 13636 26556 13700
rect 26620 13636 26621 13700
rect 26555 13635 26621 13636
rect 27475 13564 27541 13565
rect 27475 13500 27476 13564
rect 27540 13500 27541 13564
rect 27475 13499 27541 13500
rect 24531 10436 24597 10437
rect 24531 10372 24532 10436
rect 24596 10372 24597 10436
rect 24531 10371 24597 10372
rect 20483 7308 20549 7309
rect 20483 7244 20484 7308
rect 20548 7244 20549 7308
rect 20483 7243 20549 7244
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 27478 5541 27538 13499
rect 29502 10981 29562 20571
rect 29870 17373 29930 25059
rect 30051 24444 30117 24445
rect 30051 24380 30052 24444
rect 30116 24380 30117 24444
rect 30051 24379 30117 24380
rect 30054 22133 30114 24379
rect 30238 24173 30298 29003
rect 30606 24445 30666 32131
rect 31342 28253 31402 41379
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 31891 36140 31957 36141
rect 31891 36076 31892 36140
rect 31956 36076 31957 36140
rect 31891 36075 31957 36076
rect 31523 29340 31589 29341
rect 31523 29276 31524 29340
rect 31588 29276 31589 29340
rect 31523 29275 31589 29276
rect 31339 28252 31405 28253
rect 31339 28188 31340 28252
rect 31404 28188 31405 28252
rect 31339 28187 31405 28188
rect 30971 27572 31037 27573
rect 30971 27508 30972 27572
rect 31036 27508 31037 27572
rect 30971 27507 31037 27508
rect 30603 24444 30669 24445
rect 30603 24380 30604 24444
rect 30668 24380 30669 24444
rect 30603 24379 30669 24380
rect 30603 24308 30669 24309
rect 30603 24244 30604 24308
rect 30668 24244 30669 24308
rect 30603 24243 30669 24244
rect 30235 24172 30301 24173
rect 30235 24108 30236 24172
rect 30300 24108 30301 24172
rect 30235 24107 30301 24108
rect 30051 22132 30117 22133
rect 30051 22068 30052 22132
rect 30116 22068 30117 22132
rect 30051 22067 30117 22068
rect 29867 17372 29933 17373
rect 29867 17308 29868 17372
rect 29932 17308 29933 17372
rect 29867 17307 29933 17308
rect 30238 15197 30298 24107
rect 30606 19549 30666 24243
rect 30974 22133 31034 27507
rect 31526 26213 31586 29275
rect 31523 26212 31589 26213
rect 31523 26148 31524 26212
rect 31588 26148 31589 26212
rect 31523 26147 31589 26148
rect 31523 23628 31589 23629
rect 31523 23564 31524 23628
rect 31588 23564 31589 23628
rect 31523 23563 31589 23564
rect 30971 22132 31037 22133
rect 30971 22068 30972 22132
rect 31036 22068 31037 22132
rect 30971 22067 31037 22068
rect 30603 19548 30669 19549
rect 30603 19484 30604 19548
rect 30668 19484 30669 19548
rect 30603 19483 30669 19484
rect 31526 19277 31586 23563
rect 31894 22266 31954 36075
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34651 34236 34717 34237
rect 34651 34172 34652 34236
rect 34716 34172 34717 34236
rect 34651 34171 34717 34172
rect 32443 33284 32509 33285
rect 32443 33220 32444 33284
rect 32508 33220 32509 33284
rect 32443 33219 32509 33220
rect 32259 31108 32325 31109
rect 32259 31044 32260 31108
rect 32324 31044 32325 31108
rect 32259 31043 32325 31044
rect 32262 22541 32322 31043
rect 32259 22540 32325 22541
rect 32259 22476 32260 22540
rect 32324 22476 32325 22540
rect 32259 22475 32325 22476
rect 31710 22206 31954 22266
rect 31710 21861 31770 22206
rect 31707 21860 31773 21861
rect 31707 21796 31708 21860
rect 31772 21796 31773 21860
rect 31707 21795 31773 21796
rect 32446 20501 32506 33219
rect 34467 32740 34533 32741
rect 34467 32676 34468 32740
rect 34532 32676 34533 32740
rect 34467 32675 34533 32676
rect 33547 30428 33613 30429
rect 33547 30364 33548 30428
rect 33612 30364 33613 30428
rect 33547 30363 33613 30364
rect 33363 25124 33429 25125
rect 33363 25060 33364 25124
rect 33428 25060 33429 25124
rect 33363 25059 33429 25060
rect 33366 20773 33426 25059
rect 33363 20772 33429 20773
rect 33363 20708 33364 20772
rect 33428 20708 33429 20772
rect 33363 20707 33429 20708
rect 32443 20500 32509 20501
rect 32443 20436 32444 20500
rect 32508 20436 32509 20500
rect 32443 20435 32509 20436
rect 31523 19276 31589 19277
rect 31523 19212 31524 19276
rect 31588 19212 31589 19276
rect 31523 19211 31589 19212
rect 33550 18189 33610 30363
rect 34099 29068 34165 29069
rect 34099 29004 34100 29068
rect 34164 29004 34165 29068
rect 34099 29003 34165 29004
rect 33731 19412 33797 19413
rect 33731 19348 33732 19412
rect 33796 19348 33797 19412
rect 33731 19347 33797 19348
rect 33547 18188 33613 18189
rect 33547 18124 33548 18188
rect 33612 18124 33613 18188
rect 33547 18123 33613 18124
rect 33179 18052 33245 18053
rect 33179 17988 33180 18052
rect 33244 17988 33245 18052
rect 33179 17987 33245 17988
rect 30235 15196 30301 15197
rect 30235 15132 30236 15196
rect 30300 15132 30301 15196
rect 30235 15131 30301 15132
rect 32995 13836 33061 13837
rect 32995 13772 32996 13836
rect 33060 13772 33061 13836
rect 32995 13771 33061 13772
rect 32998 10981 33058 13771
rect 29499 10980 29565 10981
rect 29499 10916 29500 10980
rect 29564 10916 29565 10980
rect 29499 10915 29565 10916
rect 32995 10980 33061 10981
rect 32995 10916 32996 10980
rect 33060 10916 33061 10980
rect 32995 10915 33061 10916
rect 33182 10845 33242 17987
rect 33734 17781 33794 19347
rect 33915 19140 33981 19141
rect 33915 19076 33916 19140
rect 33980 19076 33981 19140
rect 33915 19075 33981 19076
rect 33731 17780 33797 17781
rect 33731 17716 33732 17780
rect 33796 17716 33797 17780
rect 33731 17715 33797 17716
rect 33918 15333 33978 19075
rect 34102 18461 34162 29003
rect 34283 28524 34349 28525
rect 34283 28460 34284 28524
rect 34348 28460 34349 28524
rect 34283 28459 34349 28460
rect 34286 25397 34346 28459
rect 34470 27709 34530 32675
rect 34467 27708 34533 27709
rect 34467 27644 34468 27708
rect 34532 27644 34533 27708
rect 34467 27643 34533 27644
rect 34467 26348 34533 26349
rect 34467 26284 34468 26348
rect 34532 26284 34533 26348
rect 34467 26283 34533 26284
rect 34283 25396 34349 25397
rect 34283 25332 34284 25396
rect 34348 25332 34349 25396
rect 34283 25331 34349 25332
rect 34470 21725 34530 26283
rect 34654 26213 34714 34171
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 35939 31924 36005 31925
rect 35939 31860 35940 31924
rect 36004 31860 36005 31924
rect 35939 31859 36005 31860
rect 35387 31788 35453 31789
rect 35387 31724 35388 31788
rect 35452 31724 35453 31788
rect 35387 31723 35453 31724
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 35390 29749 35450 31723
rect 35387 29748 35453 29749
rect 35387 29684 35388 29748
rect 35452 29684 35453 29748
rect 35387 29683 35453 29684
rect 35387 29068 35453 29069
rect 35387 29004 35388 29068
rect 35452 29004 35453 29068
rect 35387 29003 35453 29004
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34651 26212 34717 26213
rect 34651 26148 34652 26212
rect 34716 26148 34717 26212
rect 34651 26147 34717 26148
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34651 22540 34717 22541
rect 34651 22476 34652 22540
rect 34716 22476 34717 22540
rect 34651 22475 34717 22476
rect 34467 21724 34533 21725
rect 34467 21660 34468 21724
rect 34532 21660 34533 21724
rect 34467 21659 34533 21660
rect 34099 18460 34165 18461
rect 34099 18396 34100 18460
rect 34164 18396 34165 18460
rect 34099 18395 34165 18396
rect 34283 16692 34349 16693
rect 34283 16628 34284 16692
rect 34348 16628 34349 16692
rect 34283 16627 34349 16628
rect 33915 15332 33981 15333
rect 33915 15268 33916 15332
rect 33980 15268 33981 15332
rect 33915 15267 33981 15268
rect 33179 10844 33245 10845
rect 33179 10780 33180 10844
rect 33244 10780 33245 10844
rect 33179 10779 33245 10780
rect 34286 9621 34346 16627
rect 34467 16556 34533 16557
rect 34467 16492 34468 16556
rect 34532 16492 34533 16556
rect 34467 16491 34533 16492
rect 34470 11797 34530 16491
rect 34654 14109 34714 22475
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 35390 18733 35450 29003
rect 35942 27165 36002 31859
rect 37411 29068 37477 29069
rect 37411 29004 37412 29068
rect 37476 29004 37477 29068
rect 37411 29003 37477 29004
rect 36859 28796 36925 28797
rect 36859 28732 36860 28796
rect 36924 28732 36925 28796
rect 36859 28731 36925 28732
rect 35939 27164 36005 27165
rect 35939 27100 35940 27164
rect 36004 27100 36005 27164
rect 35939 27099 36005 27100
rect 35755 26348 35821 26349
rect 35755 26284 35756 26348
rect 35820 26284 35821 26348
rect 35755 26283 35821 26284
rect 35387 18732 35453 18733
rect 35387 18668 35388 18732
rect 35452 18668 35453 18732
rect 35387 18667 35453 18668
rect 35387 18188 35453 18189
rect 35387 18124 35388 18188
rect 35452 18124 35453 18188
rect 35387 18123 35453 18124
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 35390 14789 35450 18123
rect 35758 16557 35818 26283
rect 36123 22948 36189 22949
rect 36123 22884 36124 22948
rect 36188 22884 36189 22948
rect 36123 22883 36189 22884
rect 35939 22676 36005 22677
rect 35939 22612 35940 22676
rect 36004 22612 36005 22676
rect 35939 22611 36005 22612
rect 35755 16556 35821 16557
rect 35755 16492 35756 16556
rect 35820 16492 35821 16556
rect 35755 16491 35821 16492
rect 35571 16420 35637 16421
rect 35571 16356 35572 16420
rect 35636 16356 35637 16420
rect 35571 16355 35637 16356
rect 35387 14788 35453 14789
rect 35387 14724 35388 14788
rect 35452 14724 35453 14788
rect 35387 14723 35453 14724
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34651 14108 34717 14109
rect 34651 14044 34652 14108
rect 34716 14044 34717 14108
rect 34651 14043 34717 14044
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34467 11796 34533 11797
rect 34467 11732 34468 11796
rect 34532 11732 34533 11796
rect 34467 11731 34533 11732
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34283 9620 34349 9621
rect 34283 9556 34284 9620
rect 34348 9556 34349 9620
rect 34283 9555 34349 9556
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 35574 8261 35634 16355
rect 35942 12069 36002 22611
rect 36126 21861 36186 22883
rect 36123 21860 36189 21861
rect 36123 21796 36124 21860
rect 36188 21796 36189 21860
rect 36123 21795 36189 21796
rect 36126 16421 36186 21795
rect 36862 18597 36922 28731
rect 37043 24988 37109 24989
rect 37043 24924 37044 24988
rect 37108 24924 37109 24988
rect 37043 24923 37109 24924
rect 36859 18596 36925 18597
rect 36859 18532 36860 18596
rect 36924 18532 36925 18596
rect 36859 18531 36925 18532
rect 36307 18460 36373 18461
rect 36307 18396 36308 18460
rect 36372 18396 36373 18460
rect 36307 18395 36373 18396
rect 36123 16420 36189 16421
rect 36123 16356 36124 16420
rect 36188 16356 36189 16420
rect 36123 16355 36189 16356
rect 35939 12068 36005 12069
rect 35939 12004 35940 12068
rect 36004 12004 36005 12068
rect 35939 12003 36005 12004
rect 35571 8260 35637 8261
rect 35571 8196 35572 8260
rect 35636 8196 35637 8260
rect 35571 8195 35637 8196
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 27475 5540 27541 5541
rect 27475 5476 27476 5540
rect 27540 5476 27541 5540
rect 27475 5475 27541 5476
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 18643 3636 18709 3637
rect 18643 3572 18644 3636
rect 18708 3572 18709 3636
rect 18643 3571 18709 3572
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 4928 35248 5952
rect 36310 5541 36370 18395
rect 37046 14245 37106 24923
rect 37227 23492 37293 23493
rect 37227 23428 37228 23492
rect 37292 23428 37293 23492
rect 37227 23427 37293 23428
rect 37230 16149 37290 23427
rect 37227 16148 37293 16149
rect 37227 16084 37228 16148
rect 37292 16084 37293 16148
rect 37227 16083 37293 16084
rect 37043 14244 37109 14245
rect 37043 14180 37044 14244
rect 37108 14180 37109 14244
rect 37043 14179 37109 14180
rect 37414 13701 37474 29003
rect 39067 27708 39133 27709
rect 39067 27644 39068 27708
rect 39132 27644 39133 27708
rect 39067 27643 39133 27644
rect 37595 25396 37661 25397
rect 37595 25332 37596 25396
rect 37660 25332 37661 25396
rect 37595 25331 37661 25332
rect 37598 23901 37658 25331
rect 37595 23900 37661 23901
rect 37595 23836 37596 23900
rect 37660 23836 37661 23900
rect 37595 23835 37661 23836
rect 37598 15197 37658 23835
rect 37779 23492 37845 23493
rect 37779 23428 37780 23492
rect 37844 23428 37845 23492
rect 37779 23427 37845 23428
rect 37595 15196 37661 15197
rect 37595 15132 37596 15196
rect 37660 15132 37661 15196
rect 37595 15131 37661 15132
rect 37782 14381 37842 23427
rect 38883 20772 38949 20773
rect 38883 20708 38884 20772
rect 38948 20708 38949 20772
rect 38883 20707 38949 20708
rect 37779 14380 37845 14381
rect 37779 14316 37780 14380
rect 37844 14316 37845 14380
rect 37779 14315 37845 14316
rect 37411 13700 37477 13701
rect 37411 13636 37412 13700
rect 37476 13636 37477 13700
rect 37411 13635 37477 13636
rect 38886 9621 38946 20707
rect 39070 13701 39130 27643
rect 39251 27164 39317 27165
rect 39251 27100 39252 27164
rect 39316 27100 39317 27164
rect 39251 27099 39317 27100
rect 39067 13700 39133 13701
rect 39067 13636 39068 13700
rect 39132 13636 39133 13700
rect 39067 13635 39133 13636
rect 39254 13565 39314 27099
rect 39251 13564 39317 13565
rect 39251 13500 39252 13564
rect 39316 13500 39317 13564
rect 39251 13499 39317 13500
rect 38883 9620 38949 9621
rect 38883 9556 38884 9620
rect 38948 9556 38949 9620
rect 38883 9555 38949 9556
rect 36307 5540 36373 5541
rect 36307 5476 36308 5540
rect 36372 5476 36373 5540
rect 36307 5475 36373 5476
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__clkbuf_4  _1509_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30268 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1510_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27232 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1511_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21344 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1512_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25208 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1513_
timestamp 1688980957
transform 1 0 29624 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1514_
timestamp 1688980957
transform 1 0 30452 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1515_
timestamp 1688980957
transform 1 0 38732 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1516_
timestamp 1688980957
transform 1 0 39284 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1517_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37996 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1518_
timestamp 1688980957
transform 1 0 37812 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1519_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 39284 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1520_
timestamp 1688980957
transform 1 0 38732 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1521_
timestamp 1688980957
transform 1 0 38088 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1522_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31372 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1523_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37628 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or4bb_1  _1524_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37720 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1525_
timestamp 1688980957
transform 1 0 37260 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1526_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32568 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1527_
timestamp 1688980957
transform 1 0 38640 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1528_
timestamp 1688980957
transform 1 0 38548 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _1529_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37720 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1530_
timestamp 1688980957
transform 1 0 38456 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1531_
timestamp 1688980957
transform 1 0 33672 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1532_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32752 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1533_
timestamp 1688980957
transform 1 0 37812 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1534_
timestamp 1688980957
transform 1 0 38456 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1535_
timestamp 1688980957
transform 1 0 34868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1536_
timestamp 1688980957
transform 1 0 38272 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1537_
timestamp 1688980957
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1538_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33948 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _1539_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33304 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_1  _1540_
timestamp 1688980957
transform 1 0 38364 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1541_
timestamp 1688980957
transform 1 0 38364 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1542_
timestamp 1688980957
transform 1 0 37260 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1543_
timestamp 1688980957
transform 1 0 31188 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1544_
timestamp 1688980957
transform 1 0 32660 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1545_
timestamp 1688980957
transform 1 0 36524 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1546_
timestamp 1688980957
transform 1 0 38640 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1547_
timestamp 1688980957
transform 1 0 35328 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1548_
timestamp 1688980957
transform 1 0 37812 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_2  _1549_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35328 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1550_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35328 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_2  _1551_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 36248 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_1  _1552_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35236 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_2  _1553_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 36156 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1554_
timestamp 1688980957
transform 1 0 29900 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _1555_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31096 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1556_
timestamp 1688980957
transform 1 0 37996 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1557_
timestamp 1688980957
transform 1 0 37536 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1558_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 38272 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand4b_4  _1559_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37260 0 -1 33728
box -38 -48 1786 592
use sky130_fd_sc_hd__or4bb_4  _1560_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 36616 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__a41o_1  _1561_
timestamp 1688980957
transform 1 0 37260 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1562_
timestamp 1688980957
transform 1 0 37536 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1563_
timestamp 1688980957
transform 1 0 36984 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1564_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24564 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _1565_
timestamp 1688980957
transform 1 0 37536 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _1566_
timestamp 1688980957
transform 1 0 39192 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1567_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37996 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _1568_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35972 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1569_
timestamp 1688980957
transform 1 0 36248 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1570_
timestamp 1688980957
transform 1 0 36340 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1571_
timestamp 1688980957
transform 1 0 36432 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1572_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31464 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1573_
timestamp 1688980957
transform 1 0 34132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1574_
timestamp 1688980957
transform 1 0 34684 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1575_
timestamp 1688980957
transform 1 0 31372 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _1576_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31280 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _1577_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _1578_
timestamp 1688980957
transform 1 0 36064 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1579_
timestamp 1688980957
transform 1 0 33764 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nand4b_4  _1580_
timestamp 1688980957
transform 1 0 32844 0 1 33728
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_2  _1581_
timestamp 1688980957
transform 1 0 33028 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1582_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27416 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1583_
timestamp 1688980957
transform 1 0 26128 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1584_
timestamp 1688980957
transform 1 0 35144 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1585_
timestamp 1688980957
transform 1 0 35604 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _1586_
timestamp 1688980957
transform 1 0 36064 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1587_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27140 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1588_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37076 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1589_
timestamp 1688980957
transform 1 0 37260 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1590_
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1591_
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _1592_
timestamp 1688980957
transform 1 0 33672 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _1593_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1594_
timestamp 1688980957
transform 1 0 26220 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1595_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26496 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _1596_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33856 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _1597_
timestamp 1688980957
transform 1 0 34684 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_2  _1598_
timestamp 1688980957
transform 1 0 33488 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _1599_
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1600_
timestamp 1688980957
transform 1 0 36064 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1601_
timestamp 1688980957
transform 1 0 34684 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1602_
timestamp 1688980957
transform 1 0 31188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1603_
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1604_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26312 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1605_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26312 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1606_
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1607_
timestamp 1688980957
transform 1 0 32936 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1608_
timestamp 1688980957
transform 1 0 33580 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1609_
timestamp 1688980957
transform 1 0 33304 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1610_
timestamp 1688980957
transform 1 0 30820 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1611_
timestamp 1688980957
transform 1 0 25852 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1612_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25300 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _1613_
timestamp 1688980957
transform 1 0 25760 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1614_
timestamp 1688980957
transform 1 0 37168 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _1615_
timestamp 1688980957
transform 1 0 37904 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _1616_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35052 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1617_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _1618_
timestamp 1688980957
transform 1 0 33580 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1619_
timestamp 1688980957
transform 1 0 34684 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _1620_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35696 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1621_
timestamp 1688980957
transform 1 0 34408 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1622_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _1623_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35604 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1624_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34040 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1625_
timestamp 1688980957
transform 1 0 32568 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1626_
timestamp 1688980957
transform 1 0 32660 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1627_
timestamp 1688980957
transform 1 0 33488 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1628_
timestamp 1688980957
transform 1 0 31648 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1629_
timestamp 1688980957
transform 1 0 35696 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1630_
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _1631_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33028 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1632_
timestamp 1688980957
transform 1 0 35512 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1633_
timestamp 1688980957
transform 1 0 32200 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1634_
timestamp 1688980957
transform 1 0 33764 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1635_
timestamp 1688980957
transform 1 0 31740 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_4  _1636_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33764 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__a21oi_1  _1637_
timestamp 1688980957
transform 1 0 31924 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1638_
timestamp 1688980957
transform 1 0 36156 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1639_
timestamp 1688980957
transform 1 0 33948 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1640_
timestamp 1688980957
transform 1 0 31096 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1641_
timestamp 1688980957
transform 1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1642_
timestamp 1688980957
transform 1 0 31372 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1643_
timestamp 1688980957
transform 1 0 31372 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _1644_
timestamp 1688980957
transform 1 0 32200 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _1645_
timestamp 1688980957
transform 1 0 33672 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1646_
timestamp 1688980957
transform 1 0 36708 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1647_
timestamp 1688980957
transform 1 0 33764 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1648_
timestamp 1688980957
transform 1 0 31004 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1649_
timestamp 1688980957
transform 1 0 31280 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1650_
timestamp 1688980957
transform 1 0 30912 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1651_
timestamp 1688980957
transform 1 0 31464 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1652_
timestamp 1688980957
transform 1 0 29624 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1653_
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1654_
timestamp 1688980957
transform 1 0 30912 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1655_
timestamp 1688980957
transform 1 0 29992 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1656_
timestamp 1688980957
transform 1 0 31924 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1657_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1658_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29624 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _1659_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30820 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1660_
timestamp 1688980957
transform 1 0 28428 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _1661_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30452 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1662_
timestamp 1688980957
transform 1 0 31464 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_2  _1663_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30912 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1664_
timestamp 1688980957
transform 1 0 22724 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1665_
timestamp 1688980957
transform 1 0 20792 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _1666_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33672 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _1667_
timestamp 1688980957
transform 1 0 27416 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_4  _1668_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20608 0 1 25024
box -38 -48 1326 592
use sky130_fd_sc_hd__o31ai_4  _1669_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25116 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__clkinv_4  _1670_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28704 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1671_
timestamp 1688980957
transform 1 0 20608 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1672_
timestamp 1688980957
transform 1 0 21160 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1673_
timestamp 1688980957
transform 1 0 19688 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1674_
timestamp 1688980957
transform 1 0 28060 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1675_
timestamp 1688980957
transform 1 0 30452 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1676_
timestamp 1688980957
transform 1 0 34776 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1677_
timestamp 1688980957
transform 1 0 28244 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1678_
timestamp 1688980957
transform 1 0 27324 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1679_
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1680_
timestamp 1688980957
transform 1 0 19964 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1681_
timestamp 1688980957
transform 1 0 19228 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1682_
timestamp 1688980957
transform 1 0 18676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1683_
timestamp 1688980957
transform 1 0 22356 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1684_
timestamp 1688980957
transform 1 0 25944 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1685_
timestamp 1688980957
transform 1 0 25668 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1686_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25944 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1687_
timestamp 1688980957
transform 1 0 26680 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1688_
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1689_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25944 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1690_
timestamp 1688980957
transform 1 0 28796 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1691_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1692_
timestamp 1688980957
transform 1 0 26312 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _1693_
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1694_
timestamp 1688980957
transform 1 0 27140 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1695_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1696_
timestamp 1688980957
transform 1 0 26864 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _1697_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27232 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1698_
timestamp 1688980957
transform 1 0 25484 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1699_
timestamp 1688980957
transform 1 0 27876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1700_
timestamp 1688980957
transform 1 0 21436 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1701_
timestamp 1688980957
transform 1 0 29256 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1702_
timestamp 1688980957
transform 1 0 29808 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1703_
timestamp 1688980957
transform 1 0 23276 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1704_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27232 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1705_
timestamp 1688980957
transform 1 0 28060 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1706_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1707_
timestamp 1688980957
transform 1 0 25024 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1708_
timestamp 1688980957
transform 1 0 21712 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1709_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27876 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1710_
timestamp 1688980957
transform 1 0 28520 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1711_
timestamp 1688980957
transform 1 0 25576 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1712_
timestamp 1688980957
transform 1 0 23092 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1713_
timestamp 1688980957
transform 1 0 27784 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1714_
timestamp 1688980957
transform 1 0 30728 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1715_
timestamp 1688980957
transform 1 0 27324 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1716_
timestamp 1688980957
transform 1 0 25576 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1717_
timestamp 1688980957
transform 1 0 27232 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1718_
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1719_
timestamp 1688980957
transform 1 0 25944 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1720_
timestamp 1688980957
transform 1 0 26496 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _1721_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22540 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_4  _1722_
timestamp 1688980957
transform 1 0 23368 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1723_
timestamp 1688980957
transform 1 0 32016 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1724_
timestamp 1688980957
transform 1 0 32200 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1725_
timestamp 1688980957
transform 1 0 18216 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1726_
timestamp 1688980957
transform 1 0 31280 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1727_
timestamp 1688980957
transform 1 0 31556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1728_
timestamp 1688980957
transform 1 0 30176 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1729_
timestamp 1688980957
transform 1 0 28704 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1730_
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1731_
timestamp 1688980957
transform 1 0 30176 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1732_
timestamp 1688980957
transform 1 0 30084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1733_
timestamp 1688980957
transform 1 0 26404 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1734_
timestamp 1688980957
transform 1 0 24840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1735_
timestamp 1688980957
transform 1 0 29992 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1736_
timestamp 1688980957
transform 1 0 30728 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1737_
timestamp 1688980957
transform 1 0 31372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1738_
timestamp 1688980957
transform 1 0 33580 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1739_
timestamp 1688980957
transform 1 0 38916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1740_
timestamp 1688980957
transform 1 0 35512 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1741_
timestamp 1688980957
transform 1 0 30636 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1742_
timestamp 1688980957
transform 1 0 34500 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1743_
timestamp 1688980957
transform 1 0 36432 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1744_
timestamp 1688980957
transform 1 0 32568 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1745_
timestamp 1688980957
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1746_
timestamp 1688980957
transform 1 0 29532 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1747_
timestamp 1688980957
transform 1 0 29624 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1748_
timestamp 1688980957
transform 1 0 29164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1749_
timestamp 1688980957
transform 1 0 28520 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1750_
timestamp 1688980957
transform 1 0 29440 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1751_
timestamp 1688980957
transform 1 0 28796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1752_
timestamp 1688980957
transform 1 0 28612 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1753_
timestamp 1688980957
transform 1 0 26312 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1754_
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _1755_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27968 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_2  _1756_
timestamp 1688980957
transform 1 0 31372 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1757_
timestamp 1688980957
transform 1 0 32108 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1758_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27692 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1759_
timestamp 1688980957
transform 1 0 29808 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1760_
timestamp 1688980957
transform 1 0 30084 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1761_
timestamp 1688980957
transform 1 0 35788 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1762_
timestamp 1688980957
transform 1 0 35144 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _1763_
timestamp 1688980957
transform 1 0 31280 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1764_
timestamp 1688980957
transform 1 0 32660 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1765_
timestamp 1688980957
transform 1 0 35512 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1766_
timestamp 1688980957
transform 1 0 35420 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1767_
timestamp 1688980957
transform 1 0 30820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1768_
timestamp 1688980957
transform 1 0 31556 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1769_
timestamp 1688980957
transform 1 0 34224 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1770_
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1771_
timestamp 1688980957
transform 1 0 29992 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1772_
timestamp 1688980957
transform 1 0 33764 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1773_
timestamp 1688980957
transform 1 0 33120 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1774_
timestamp 1688980957
transform 1 0 30544 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1775_
timestamp 1688980957
transform 1 0 31280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1776_
timestamp 1688980957
transform 1 0 31188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1777_
timestamp 1688980957
transform 1 0 30544 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1778_
timestamp 1688980957
transform 1 0 32844 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1779_
timestamp 1688980957
transform 1 0 32200 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1780_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32292 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1781_
timestamp 1688980957
transform 1 0 26036 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1782_
timestamp 1688980957
transform 1 0 26036 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1783_
timestamp 1688980957
transform 1 0 28428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1784_
timestamp 1688980957
transform 1 0 27048 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1785_
timestamp 1688980957
transform 1 0 34500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1786_
timestamp 1688980957
transform 1 0 35880 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1787_
timestamp 1688980957
transform 1 0 36340 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1788_
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1789_
timestamp 1688980957
transform 1 0 34868 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1790_
timestamp 1688980957
transform 1 0 33396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1791_
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1792_
timestamp 1688980957
transform 1 0 31556 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1793_
timestamp 1688980957
transform 1 0 30912 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1794_
timestamp 1688980957
transform 1 0 30544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1795_
timestamp 1688980957
transform 1 0 20516 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1796_
timestamp 1688980957
transform 1 0 19872 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1797_
timestamp 1688980957
transform 1 0 14076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_2  _1798_
timestamp 1688980957
transform 1 0 33028 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _1799_
timestamp 1688980957
transform 1 0 35420 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1800_
timestamp 1688980957
transform 1 0 33212 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1801_
timestamp 1688980957
transform 1 0 33948 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1802_
timestamp 1688980957
transform 1 0 31372 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _1803_
timestamp 1688980957
transform 1 0 30544 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1804_
timestamp 1688980957
transform 1 0 29348 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1805_
timestamp 1688980957
transform 1 0 36432 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1806_
timestamp 1688980957
transform 1 0 31280 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1807_
timestamp 1688980957
transform 1 0 37260 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1808_
timestamp 1688980957
transform 1 0 35696 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1809_
timestamp 1688980957
transform 1 0 33948 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1810_
timestamp 1688980957
transform 1 0 38088 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1811_
timestamp 1688980957
transform 1 0 33488 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1812_
timestamp 1688980957
transform 1 0 33580 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1813_
timestamp 1688980957
transform 1 0 35788 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _1814_
timestamp 1688980957
transform 1 0 31372 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1815_
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _1816_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33028 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _1817_
timestamp 1688980957
transform 1 0 34132 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1818_
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1819_
timestamp 1688980957
transform 1 0 33212 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_2  _1820_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and2_2  _1821_
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1822_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33764 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1823_
timestamp 1688980957
transform 1 0 35788 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1824_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35236 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_2  _1825_
timestamp 1688980957
transform 1 0 31096 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and3_2  _1826_
timestamp 1688980957
transform 1 0 32200 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1827_
timestamp 1688980957
transform 1 0 33488 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1828_
timestamp 1688980957
transform 1 0 32476 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _1829_
timestamp 1688980957
transform 1 0 31464 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1830_
timestamp 1688980957
transform 1 0 32476 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1831_
timestamp 1688980957
transform 1 0 32476 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1832_
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1833_
timestamp 1688980957
transform 1 0 33672 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1834_
timestamp 1688980957
transform 1 0 32936 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1835_
timestamp 1688980957
transform 1 0 32752 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1836_
timestamp 1688980957
transform 1 0 36432 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1837_
timestamp 1688980957
transform 1 0 38640 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1838_
timestamp 1688980957
transform 1 0 36892 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1839_
timestamp 1688980957
transform 1 0 31464 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1840_
timestamp 1688980957
transform 1 0 32016 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1841_
timestamp 1688980957
transform 1 0 38180 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1842_
timestamp 1688980957
transform 1 0 35052 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1843_
timestamp 1688980957
transform 1 0 37352 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1844_
timestamp 1688980957
transform 1 0 35420 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _1845_
timestamp 1688980957
transform 1 0 33120 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1846_
timestamp 1688980957
transform 1 0 32844 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1847_
timestamp 1688980957
transform 1 0 36708 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1848_
timestamp 1688980957
transform 1 0 35328 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1849_
timestamp 1688980957
transform 1 0 35420 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1850_
timestamp 1688980957
transform 1 0 35144 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1851_
timestamp 1688980957
transform 1 0 35512 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1852_
timestamp 1688980957
transform 1 0 38456 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1853_
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1854_
timestamp 1688980957
transform 1 0 32752 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1855_
timestamp 1688980957
transform 1 0 33120 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1856_
timestamp 1688980957
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1857_
timestamp 1688980957
transform 1 0 35604 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1858_
timestamp 1688980957
transform 1 0 35512 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _1859_
timestamp 1688980957
transform 1 0 33948 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1860_
timestamp 1688980957
transform 1 0 33948 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1861_
timestamp 1688980957
transform 1 0 38824 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1862_
timestamp 1688980957
transform 1 0 38732 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1863_
timestamp 1688980957
transform 1 0 39836 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1864_
timestamp 1688980957
transform 1 0 34960 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _1865_
timestamp 1688980957
transform 1 0 35052 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1866_
timestamp 1688980957
transform 1 0 34684 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1867_
timestamp 1688980957
transform 1 0 34776 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1868_
timestamp 1688980957
transform 1 0 35604 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1869_
timestamp 1688980957
transform 1 0 30728 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1870_
timestamp 1688980957
transform 1 0 30452 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1871_
timestamp 1688980957
transform 1 0 30912 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _1872_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29624 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1873_
timestamp 1688980957
transform 1 0 30360 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1874_
timestamp 1688980957
transform 1 0 35604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1875_
timestamp 1688980957
transform 1 0 36340 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1876_
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1877_
timestamp 1688980957
transform 1 0 30636 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1878_
timestamp 1688980957
transform 1 0 31280 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1879_
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1880_
timestamp 1688980957
transform 1 0 39836 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1881_
timestamp 1688980957
transform 1 0 40020 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1882_
timestamp 1688980957
transform 1 0 39836 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _1883_
timestamp 1688980957
transform 1 0 31556 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1884_
timestamp 1688980957
transform 1 0 34868 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1885_
timestamp 1688980957
transform 1 0 34868 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1886_
timestamp 1688980957
transform 1 0 33396 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1887_
timestamp 1688980957
transform 1 0 33672 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1888_
timestamp 1688980957
transform 1 0 34132 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1889_
timestamp 1688980957
transform 1 0 37260 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1890_
timestamp 1688980957
transform 1 0 39284 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1891_
timestamp 1688980957
transform 1 0 38272 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1892_
timestamp 1688980957
transform 1 0 38548 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1893_
timestamp 1688980957
transform 1 0 37352 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1894_
timestamp 1688980957
transform 1 0 31740 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_1  _1895_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1896_
timestamp 1688980957
transform 1 0 29532 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1897_
timestamp 1688980957
transform 1 0 33396 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1898_
timestamp 1688980957
transform 1 0 37720 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1899_
timestamp 1688980957
transform 1 0 36984 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1900_
timestamp 1688980957
transform 1 0 37444 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1901_
timestamp 1688980957
transform 1 0 38640 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1902_
timestamp 1688980957
transform 1 0 39836 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1903_
timestamp 1688980957
transform 1 0 30912 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1904_
timestamp 1688980957
transform 1 0 33120 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1905_
timestamp 1688980957
transform 1 0 31648 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1906_
timestamp 1688980957
transform 1 0 31004 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1907_
timestamp 1688980957
transform 1 0 31096 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1908_
timestamp 1688980957
transform 1 0 31188 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1909_
timestamp 1688980957
transform 1 0 40112 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1910_
timestamp 1688980957
transform 1 0 39560 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1911_
timestamp 1688980957
transform 1 0 40480 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1912_
timestamp 1688980957
transform 1 0 39836 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1913_
timestamp 1688980957
transform 1 0 35972 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1914_
timestamp 1688980957
transform 1 0 35696 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1915_
timestamp 1688980957
transform 1 0 37260 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1916_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1917_
timestamp 1688980957
transform 1 0 34224 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1918_
timestamp 1688980957
transform 1 0 37260 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1919_
timestamp 1688980957
transform 1 0 37444 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1920_
timestamp 1688980957
transform 1 0 38916 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1921_
timestamp 1688980957
transform 1 0 39192 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1922_
timestamp 1688980957
transform 1 0 34868 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1923_
timestamp 1688980957
transform 1 0 33856 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1924_
timestamp 1688980957
transform 1 0 39376 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1925_
timestamp 1688980957
transform 1 0 38456 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1926_
timestamp 1688980957
transform 1 0 39376 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1927_
timestamp 1688980957
transform 1 0 39836 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1928_
timestamp 1688980957
transform 1 0 39376 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1929_
timestamp 1688980957
transform 1 0 37444 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1930_
timestamp 1688980957
transform 1 0 37260 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1931_
timestamp 1688980957
transform 1 0 37260 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1932_
timestamp 1688980957
transform 1 0 36616 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1933_
timestamp 1688980957
transform 1 0 37260 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1934_
timestamp 1688980957
transform 1 0 37260 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1935_
timestamp 1688980957
transform 1 0 32108 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1936_
timestamp 1688980957
transform 1 0 31280 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1937_
timestamp 1688980957
transform 1 0 37720 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1938_
timestamp 1688980957
transform 1 0 37536 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1939_
timestamp 1688980957
transform 1 0 37260 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1940_
timestamp 1688980957
transform 1 0 37628 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1941_
timestamp 1688980957
transform 1 0 39468 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1942_
timestamp 1688980957
transform 1 0 39836 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1943_
timestamp 1688980957
transform 1 0 34224 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1944_
timestamp 1688980957
transform 1 0 37260 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1945_
timestamp 1688980957
transform 1 0 38548 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1946_
timestamp 1688980957
transform 1 0 39192 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1947_
timestamp 1688980957
transform 1 0 39836 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1948_
timestamp 1688980957
transform 1 0 35880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1949_
timestamp 1688980957
transform 1 0 38640 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1950_
timestamp 1688980957
transform 1 0 37260 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1951_
timestamp 1688980957
transform 1 0 33672 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1952_
timestamp 1688980957
transform 1 0 39376 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1953_
timestamp 1688980957
transform 1 0 39928 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1954_
timestamp 1688980957
transform 1 0 40112 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1955_
timestamp 1688980957
transform 1 0 39192 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _1956_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1957_
timestamp 1688980957
transform 1 0 36616 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1958_
timestamp 1688980957
transform 1 0 37904 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1959_
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1960_
timestamp 1688980957
transform 1 0 38088 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1961_
timestamp 1688980957
transform 1 0 39836 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1962_
timestamp 1688980957
transform 1 0 39836 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1963_
timestamp 1688980957
transform 1 0 40388 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1964_
timestamp 1688980957
transform 1 0 36156 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1965_
timestamp 1688980957
transform 1 0 38732 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1966_
timestamp 1688980957
transform 1 0 39928 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1967_
timestamp 1688980957
transform 1 0 39836 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1968_
timestamp 1688980957
transform 1 0 21160 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1969_
timestamp 1688980957
transform 1 0 21804 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1970_
timestamp 1688980957
transform 1 0 39836 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1971_
timestamp 1688980957
transform 1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1972_
timestamp 1688980957
transform 1 0 17572 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1973_
timestamp 1688980957
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1974_
timestamp 1688980957
transform 1 0 17664 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _1975_
timestamp 1688980957
transform 1 0 22264 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1976_
timestamp 1688980957
transform 1 0 28704 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1977_
timestamp 1688980957
transform 1 0 32292 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _1978_
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1979_
timestamp 1688980957
transform 1 0 20056 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1980_
timestamp 1688980957
transform 1 0 28612 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1981_
timestamp 1688980957
transform 1 0 30268 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1982_
timestamp 1688980957
transform 1 0 28336 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1983_
timestamp 1688980957
transform 1 0 28796 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1984_
timestamp 1688980957
transform 1 0 21712 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1985_
timestamp 1688980957
transform 1 0 28796 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1986_
timestamp 1688980957
transform 1 0 17296 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1987_
timestamp 1688980957
transform 1 0 19780 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _1988_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17480 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1989_
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1990_
timestamp 1688980957
transform 1 0 25852 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1991_
timestamp 1688980957
transform 1 0 24840 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _1992_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26404 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1993_
timestamp 1688980957
transform 1 0 25116 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_4  _1994_
timestamp 1688980957
transform 1 0 31740 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1995_
timestamp 1688980957
transform 1 0 26312 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1996_
timestamp 1688980957
transform 1 0 25576 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_4  _1997_
timestamp 1688980957
transform 1 0 32108 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_1  _1998_
timestamp 1688980957
transform 1 0 20976 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1999_
timestamp 1688980957
transform 1 0 23368 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _2000_
timestamp 1688980957
transform 1 0 25668 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _2001_
timestamp 1688980957
transform 1 0 25760 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _2002_
timestamp 1688980957
transform 1 0 26220 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2003_
timestamp 1688980957
transform 1 0 23276 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2004_
timestamp 1688980957
transform 1 0 23184 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2005_
timestamp 1688980957
transform 1 0 29624 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2006_
timestamp 1688980957
transform 1 0 28152 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2007_
timestamp 1688980957
transform 1 0 23736 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2008_
timestamp 1688980957
transform 1 0 31280 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2009_
timestamp 1688980957
transform 1 0 28520 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2010_
timestamp 1688980957
transform 1 0 22632 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _2011_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23368 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2012_
timestamp 1688980957
transform 1 0 20332 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2013_
timestamp 1688980957
transform 1 0 21160 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2014_
timestamp 1688980957
transform 1 0 21896 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2015_
timestamp 1688980957
transform 1 0 23184 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2016_
timestamp 1688980957
transform 1 0 20700 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2017_
timestamp 1688980957
transform 1 0 21160 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _2018_
timestamp 1688980957
transform 1 0 32936 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_1  _2019_
timestamp 1688980957
transform 1 0 28060 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2020_
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _2021_
timestamp 1688980957
transform 1 0 32752 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_4  _2022_
timestamp 1688980957
transform 1 0 33028 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_2  _2023_
timestamp 1688980957
transform 1 0 26312 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2024_
timestamp 1688980957
transform 1 0 20700 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _2025_
timestamp 1688980957
transform 1 0 20148 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2026_
timestamp 1688980957
transform 1 0 21068 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2027_
timestamp 1688980957
transform 1 0 21252 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _2028_
timestamp 1688980957
transform 1 0 25760 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2029_
timestamp 1688980957
transform 1 0 25576 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2030_
timestamp 1688980957
transform 1 0 25760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _2031_
timestamp 1688980957
transform 1 0 23276 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _2032_
timestamp 1688980957
transform 1 0 16008 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2033_
timestamp 1688980957
transform 1 0 27508 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2034_
timestamp 1688980957
transform 1 0 18124 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2035_
timestamp 1688980957
transform 1 0 29808 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2036_
timestamp 1688980957
transform 1 0 28244 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2037_
timestamp 1688980957
transform 1 0 28704 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _2038_
timestamp 1688980957
transform 1 0 27968 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _2039_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20424 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _2040_
timestamp 1688980957
transform 1 0 25668 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2041_
timestamp 1688980957
transform 1 0 26772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _2042_
timestamp 1688980957
transform 1 0 26220 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2043_
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2044_
timestamp 1688980957
transform 1 0 28888 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2045_
timestamp 1688980957
transform 1 0 29440 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _2046_
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _2047_
timestamp 1688980957
transform 1 0 28152 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_4  _2048_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__and2_1  _2049_
timestamp 1688980957
transform 1 0 28060 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _2050_
timestamp 1688980957
transform 1 0 28428 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2051_
timestamp 1688980957
transform 1 0 27416 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_2  _2052_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35880 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _2053_
timestamp 1688980957
transform 1 0 28060 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2054_
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2055_
timestamp 1688980957
transform 1 0 30084 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _2056_
timestamp 1688980957
transform 1 0 27876 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2057_
timestamp 1688980957
transform 1 0 28612 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _2058_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26036 0 1 21760
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_1  _2059_
timestamp 1688980957
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2060_
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2061_
timestamp 1688980957
transform 1 0 17756 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _2062_
timestamp 1688980957
transform 1 0 19872 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_2  _2063_
timestamp 1688980957
transform 1 0 20792 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _2064_
timestamp 1688980957
transform 1 0 25484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_2  _2065_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25760 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _2066_
timestamp 1688980957
transform 1 0 20700 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2067_
timestamp 1688980957
transform 1 0 20424 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _2068_
timestamp 1688980957
transform 1 0 17020 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _2069_
timestamp 1688980957
transform 1 0 16836 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _2070_
timestamp 1688980957
transform 1 0 14076 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__o41a_1  _2071_
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2072_
timestamp 1688980957
transform 1 0 27968 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _2073_
timestamp 1688980957
transform 1 0 31096 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _2074_
timestamp 1688980957
transform 1 0 30268 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2075_
timestamp 1688980957
transform 1 0 28520 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _2076_
timestamp 1688980957
transform 1 0 28888 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2077_
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2078_
timestamp 1688980957
transform 1 0 29072 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _2079_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _2080_
timestamp 1688980957
transform 1 0 28428 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _2081_
timestamp 1688980957
transform 1 0 27324 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2082_
timestamp 1688980957
transform 1 0 26036 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _2083_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25300 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _2084_
timestamp 1688980957
transform 1 0 28244 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _2085_
timestamp 1688980957
transform 1 0 28520 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2086_
timestamp 1688980957
transform 1 0 28244 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2087_
timestamp 1688980957
transform 1 0 27600 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_2  _2088_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20056 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_1  _2089_
timestamp 1688980957
transform 1 0 29808 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _2090_
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2091_
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _2092_
timestamp 1688980957
transform 1 0 27324 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2093_
timestamp 1688980957
transform 1 0 26680 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2094_
timestamp 1688980957
transform 1 0 26680 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _2095_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _2096_
timestamp 1688980957
transform 1 0 30544 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _2097_
timestamp 1688980957
transform 1 0 26128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2098_
timestamp 1688980957
transform 1 0 27784 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2099_
timestamp 1688980957
transform 1 0 26956 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _2100_
timestamp 1688980957
transform 1 0 18952 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2101_
timestamp 1688980957
transform 1 0 26956 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2102_
timestamp 1688980957
transform 1 0 30544 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2103_
timestamp 1688980957
transform 1 0 28612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _2104_
timestamp 1688980957
transform 1 0 25300 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o41ai_4  _2105_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25576 0 1 22848
box -38 -48 2062 592
use sky130_fd_sc_hd__and4bb_1  _2106_
timestamp 1688980957
transform 1 0 15824 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _2107_
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _2108_
timestamp 1688980957
transform 1 0 16744 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2109_
timestamp 1688980957
transform 1 0 14996 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2110_
timestamp 1688980957
transform 1 0 16100 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _2111_
timestamp 1688980957
transform 1 0 14996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _2112_
timestamp 1688980957
transform 1 0 14904 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _2113_
timestamp 1688980957
transform 1 0 14352 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2114_
timestamp 1688980957
transform 1 0 14996 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _2115_
timestamp 1688980957
transform 1 0 15088 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _2116_
timestamp 1688980957
transform 1 0 15456 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _2117_
timestamp 1688980957
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _2118_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15272 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2119_
timestamp 1688980957
transform 1 0 5060 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2120_
timestamp 1688980957
transform 1 0 4232 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2121_
timestamp 1688980957
transform 1 0 5612 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a2111oi_1  _2122_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15548 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _2123_
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2124_
timestamp 1688980957
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _2125_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _2126_
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _2127_
timestamp 1688980957
transform 1 0 28888 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a311oi_1  _2128_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32936 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2129_
timestamp 1688980957
transform 1 0 29440 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2130_
timestamp 1688980957
transform 1 0 33304 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _2131_
timestamp 1688980957
transform 1 0 33764 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _2132_
timestamp 1688980957
transform 1 0 33120 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _2133_
timestamp 1688980957
transform 1 0 29900 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _2134_
timestamp 1688980957
transform 1 0 30728 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _2135_
timestamp 1688980957
transform 1 0 23644 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2136_
timestamp 1688980957
transform 1 0 24932 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2137_
timestamp 1688980957
transform 1 0 28980 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _2138_
timestamp 1688980957
transform 1 0 32292 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2139_
timestamp 1688980957
transform 1 0 26772 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _2140_
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _2141_
timestamp 1688980957
transform 1 0 26036 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2142_
timestamp 1688980957
transform 1 0 27140 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2143_
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2144_
timestamp 1688980957
transform 1 0 26588 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _2145_
timestamp 1688980957
transform 1 0 24472 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2146_
timestamp 1688980957
transform 1 0 22540 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2147_
timestamp 1688980957
transform 1 0 25116 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2148_
timestamp 1688980957
transform 1 0 24288 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _2149_
timestamp 1688980957
transform 1 0 24196 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2150_
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2151_
timestamp 1688980957
transform 1 0 23276 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _2152_
timestamp 1688980957
transform 1 0 21528 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2153_
timestamp 1688980957
transform 1 0 23920 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2154_
timestamp 1688980957
transform 1 0 22264 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2155_
timestamp 1688980957
transform 1 0 25392 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2156_
timestamp 1688980957
transform 1 0 23644 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2157_
timestamp 1688980957
transform 1 0 25024 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2158_
timestamp 1688980957
transform 1 0 23736 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _2159_
timestamp 1688980957
transform 1 0 21988 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2160_
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2161_
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2162_
timestamp 1688980957
transform 1 0 18584 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_1  _2163_
timestamp 1688980957
transform 1 0 20700 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2164_
timestamp 1688980957
transform 1 0 20884 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2165_
timestamp 1688980957
transform 1 0 20240 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_2  _2166_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17664 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__nor4_1  _2167_
timestamp 1688980957
transform 1 0 15548 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2168_
timestamp 1688980957
transform 1 0 7912 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2169_
timestamp 1688980957
transform 1 0 5520 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2170_
timestamp 1688980957
transform 1 0 26128 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2171_
timestamp 1688980957
transform 1 0 26772 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2172_
timestamp 1688980957
transform 1 0 25392 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2173_
timestamp 1688980957
transform 1 0 23184 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2174_
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2175_
timestamp 1688980957
transform 1 0 24564 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2176_
timestamp 1688980957
transform 1 0 24380 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2177_
timestamp 1688980957
transform 1 0 23920 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2178_
timestamp 1688980957
transform 1 0 23920 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2179_
timestamp 1688980957
transform 1 0 29532 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2180_
timestamp 1688980957
transform 1 0 27876 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2181_
timestamp 1688980957
transform 1 0 27324 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2182_
timestamp 1688980957
transform 1 0 27324 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _2183_
timestamp 1688980957
transform 1 0 27416 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _2184_
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_2  _2185_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24840 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2186_
timestamp 1688980957
transform 1 0 21252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2187_
timestamp 1688980957
transform 1 0 20608 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2188_
timestamp 1688980957
transform 1 0 26864 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2189_
timestamp 1688980957
transform 1 0 26220 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2190_
timestamp 1688980957
transform 1 0 26496 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2191_
timestamp 1688980957
transform 1 0 26036 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _2192_
timestamp 1688980957
transform 1 0 25760 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _2193_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2194_
timestamp 1688980957
transform 1 0 18032 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _2195_
timestamp 1688980957
transform 1 0 17480 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _2196_
timestamp 1688980957
transform 1 0 17296 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2197_
timestamp 1688980957
transform 1 0 21988 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _2198_
timestamp 1688980957
transform 1 0 20884 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2199_
timestamp 1688980957
transform 1 0 19136 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2200_
timestamp 1688980957
transform 1 0 18676 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _2201_
timestamp 1688980957
transform 1 0 17848 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _2202_
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_4  _2203_
timestamp 1688980957
transform 1 0 17572 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__nor4_1  _2204_
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _2205_
timestamp 1688980957
transform 1 0 18584 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2206_
timestamp 1688980957
transform 1 0 7820 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2207_
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2208_
timestamp 1688980957
transform 1 0 8188 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _2209_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5428 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2210_
timestamp 1688980957
transform 1 0 8464 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2211_
timestamp 1688980957
transform 1 0 18308 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__a2111oi_2  _2212_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_1  _2213_
timestamp 1688980957
transform 1 0 22816 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _2214_
timestamp 1688980957
transform 1 0 22080 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _2215_
timestamp 1688980957
transform 1 0 22448 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a221oi_2  _2216_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22448 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _2217_
timestamp 1688980957
transform 1 0 23644 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2218_
timestamp 1688980957
transform 1 0 23460 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _2219_
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _2220_
timestamp 1688980957
transform 1 0 13616 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _2221_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _2222_
timestamp 1688980957
transform 1 0 10580 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _2223_
timestamp 1688980957
transform 1 0 21804 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2224_
timestamp 1688980957
transform 1 0 19872 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2225_
timestamp 1688980957
transform 1 0 26680 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2226_
timestamp 1688980957
transform 1 0 25484 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2227_
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2228_
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2229_
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2230_
timestamp 1688980957
transform 1 0 21436 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2231_
timestamp 1688980957
transform 1 0 25208 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2232_
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2233_
timestamp 1688980957
transform 1 0 19504 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2234_
timestamp 1688980957
transform 1 0 23184 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2235_
timestamp 1688980957
transform 1 0 22724 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_2  _2236_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nor3_1  _2237_
timestamp 1688980957
transform 1 0 17940 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2238_
timestamp 1688980957
transform 1 0 24932 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _2239_
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2240_
timestamp 1688980957
transform 1 0 18860 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2241_
timestamp 1688980957
transform 1 0 17572 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _2242_
timestamp 1688980957
transform 1 0 18032 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _2243_
timestamp 1688980957
transform 1 0 18124 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _2244_
timestamp 1688980957
transform 1 0 17480 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _2245_
timestamp 1688980957
transform 1 0 13616 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2246_
timestamp 1688980957
transform 1 0 17296 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2247_
timestamp 1688980957
transform 1 0 17480 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2248_
timestamp 1688980957
transform 1 0 17296 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2249_
timestamp 1688980957
transform 1 0 17020 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2250_
timestamp 1688980957
transform 1 0 17848 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2251_
timestamp 1688980957
transform 1 0 9016 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_2  _2252_
timestamp 1688980957
transform 1 0 9936 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _2253_
timestamp 1688980957
transform 1 0 11040 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2254_
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2255_
timestamp 1688980957
transform 1 0 20700 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2256_
timestamp 1688980957
transform 1 0 16836 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2257_
timestamp 1688980957
transform 1 0 17388 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2258_
timestamp 1688980957
transform 1 0 10304 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _2259_
timestamp 1688980957
transform 1 0 8004 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2260_
timestamp 1688980957
transform 1 0 5244 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2261_
timestamp 1688980957
transform 1 0 4968 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2262_
timestamp 1688980957
transform 1 0 4324 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _2263_
timestamp 1688980957
transform 1 0 5336 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2264_
timestamp 1688980957
transform 1 0 8004 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2265_
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2266_
timestamp 1688980957
transform 1 0 7820 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2267_
timestamp 1688980957
transform 1 0 8648 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _2268_
timestamp 1688980957
transform 1 0 7544 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _2269_
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2270_
timestamp 1688980957
transform 1 0 8096 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _2271_
timestamp 1688980957
transform 1 0 5704 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2272_
timestamp 1688980957
transform 1 0 10396 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _2273_
timestamp 1688980957
transform 1 0 10488 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2274_
timestamp 1688980957
transform 1 0 8832 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_2  _2275_
timestamp 1688980957
transform 1 0 9752 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _2276_
timestamp 1688980957
transform 1 0 10580 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2277_
timestamp 1688980957
transform 1 0 12144 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2278_
timestamp 1688980957
transform 1 0 10856 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _2279_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9476 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2280_
timestamp 1688980957
transform 1 0 5428 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2281_
timestamp 1688980957
transform 1 0 7176 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2282_
timestamp 1688980957
transform 1 0 8188 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2283_
timestamp 1688980957
transform 1 0 15456 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2284_
timestamp 1688980957
transform 1 0 7176 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2285_
timestamp 1688980957
transform 1 0 8004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2286_
timestamp 1688980957
transform 1 0 7268 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _2287_
timestamp 1688980957
transform 1 0 19872 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _2288_
timestamp 1688980957
transform 1 0 19780 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2289_
timestamp 1688980957
transform 1 0 16100 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2290_
timestamp 1688980957
transform 1 0 7912 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2291_
timestamp 1688980957
transform 1 0 7268 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _2292_
timestamp 1688980957
transform 1 0 7176 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2293_
timestamp 1688980957
transform 1 0 7820 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _2294_
timestamp 1688980957
transform 1 0 7268 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2295_
timestamp 1688980957
transform 1 0 11224 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _2296_
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _2297_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9936 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_4  _2298_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2299_
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _2300_
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2301_
timestamp 1688980957
transform 1 0 12972 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2302_
timestamp 1688980957
transform 1 0 12880 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _2303_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14260 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2304_
timestamp 1688980957
transform 1 0 13432 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2305_
timestamp 1688980957
transform 1 0 11868 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2306_
timestamp 1688980957
transform 1 0 12052 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _2307_
timestamp 1688980957
transform 1 0 13064 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2308_
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2309_
timestamp 1688980957
transform 1 0 12788 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2310_
timestamp 1688980957
transform 1 0 12880 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _2311_
timestamp 1688980957
transform 1 0 12972 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2312_
timestamp 1688980957
transform 1 0 12236 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2313_
timestamp 1688980957
transform 1 0 12052 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _2314_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13616 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2315_
timestamp 1688980957
transform 1 0 12512 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _2316_
timestamp 1688980957
transform 1 0 11960 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2317_
timestamp 1688980957
transform 1 0 12696 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _2318_
timestamp 1688980957
transform 1 0 13432 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2319_
timestamp 1688980957
transform 1 0 13432 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2320_
timestamp 1688980957
transform 1 0 11684 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2321_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10948 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2322_
timestamp 1688980957
transform 1 0 12236 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2323_
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2324_
timestamp 1688980957
transform 1 0 9200 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _2325_
timestamp 1688980957
transform 1 0 10120 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2326_
timestamp 1688980957
transform 1 0 10488 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2327_
timestamp 1688980957
transform 1 0 7636 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2328_
timestamp 1688980957
transform 1 0 7728 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2329_
timestamp 1688980957
transform 1 0 8280 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _2330_
timestamp 1688980957
transform 1 0 9292 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2331_
timestamp 1688980957
transform 1 0 9476 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2332_
timestamp 1688980957
transform 1 0 9844 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _2333_
timestamp 1688980957
transform 1 0 10212 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _2334_
timestamp 1688980957
transform 1 0 12880 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _2335_
timestamp 1688980957
transform 1 0 10948 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2336_
timestamp 1688980957
transform 1 0 14904 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o2111ai_2  _2337_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18032 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _2338_
timestamp 1688980957
transform 1 0 9936 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2339_
timestamp 1688980957
transform 1 0 10856 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_2  _2340_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17204 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _2341_
timestamp 1688980957
transform 1 0 14076 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_4  _2342_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13248 0 -1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _2343_
timestamp 1688980957
transform 1 0 11868 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2344_
timestamp 1688980957
transform 1 0 9016 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_4  _2345_
timestamp 1688980957
transform 1 0 9660 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _2346_
timestamp 1688980957
transform 1 0 12328 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a311oi_1  _2347_
timestamp 1688980957
transform 1 0 10764 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2348_
timestamp 1688980957
transform 1 0 16192 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _2349_
timestamp 1688980957
transform 1 0 16008 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2350_
timestamp 1688980957
transform 1 0 11500 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2351_
timestamp 1688980957
transform 1 0 11960 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2352_
timestamp 1688980957
transform 1 0 10396 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2353_
timestamp 1688980957
transform 1 0 11224 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2354_
timestamp 1688980957
transform 1 0 12420 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_2  _2355_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11960 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_2  _2356_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11684 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2357_
timestamp 1688980957
transform 1 0 11776 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _2358_
timestamp 1688980957
transform 1 0 18124 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2359_
timestamp 1688980957
transform 1 0 12512 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2360_
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _2361_
timestamp 1688980957
transform 1 0 14536 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _2362_
timestamp 1688980957
transform 1 0 14536 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_4  _2363_
timestamp 1688980957
transform 1 0 11500 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__o21ai_1  _2364_
timestamp 1688980957
transform 1 0 12512 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2365_
timestamp 1688980957
transform 1 0 12880 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2366_
timestamp 1688980957
transform 1 0 13156 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _2367_
timestamp 1688980957
transform 1 0 15088 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2368_
timestamp 1688980957
transform 1 0 18124 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _2369_
timestamp 1688980957
transform 1 0 29624 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2370_
timestamp 1688980957
transform 1 0 28060 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2371_
timestamp 1688980957
transform 1 0 27048 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2372_
timestamp 1688980957
transform 1 0 27600 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2373_
timestamp 1688980957
transform 1 0 27508 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _2374_
timestamp 1688980957
transform 1 0 25484 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2375_
timestamp 1688980957
transform 1 0 25024 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _2376_
timestamp 1688980957
transform 1 0 24012 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2377_
timestamp 1688980957
transform 1 0 14168 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _2378_
timestamp 1688980957
transform 1 0 14812 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2379_
timestamp 1688980957
transform 1 0 14444 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2380_
timestamp 1688980957
transform 1 0 15088 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_2  _2381_
timestamp 1688980957
transform 1 0 15640 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _2382_
timestamp 1688980957
transform 1 0 15088 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a32oi_4  _2383_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14536 0 -1 19584
box -38 -48 2062 592
use sky130_fd_sc_hd__a22oi_2  _2384_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15180 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _2385_
timestamp 1688980957
transform 1 0 14352 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a41oi_4  _2386_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 -1 23936
box -38 -48 2062 592
use sky130_fd_sc_hd__a221o_1  _2387_
timestamp 1688980957
transform 1 0 15272 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2388_
timestamp 1688980957
transform 1 0 14904 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _2389_
timestamp 1688980957
transform 1 0 14352 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _2390_
timestamp 1688980957
transform 1 0 15456 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2391_
timestamp 1688980957
transform 1 0 14812 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _2392_
timestamp 1688980957
transform 1 0 15824 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2393_
timestamp 1688980957
transform 1 0 17020 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _2394_
timestamp 1688980957
transform 1 0 18400 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2395_
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2396_
timestamp 1688980957
transform 1 0 16836 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_2  _2397_
timestamp 1688980957
transform 1 0 17296 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _2398_
timestamp 1688980957
transform 1 0 15732 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_4  _2399_
timestamp 1688980957
transform 1 0 14720 0 1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _2400_
timestamp 1688980957
transform 1 0 16192 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2401_
timestamp 1688980957
transform 1 0 15272 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _2402_
timestamp 1688980957
transform 1 0 14812 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _2403_
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _2404_
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _2405_
timestamp 1688980957
transform 1 0 11960 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _2406_
timestamp 1688980957
transform 1 0 10672 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _2407_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_2  _2408_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15272 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _2409_
timestamp 1688980957
transform 1 0 13156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_2  _2410_
timestamp 1688980957
transform 1 0 11684 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _2411_
timestamp 1688980957
transform 1 0 9200 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2412_
timestamp 1688980957
transform 1 0 9108 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2413_
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2414_
timestamp 1688980957
transform 1 0 8188 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2415_
timestamp 1688980957
transform 1 0 9660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2416_
timestamp 1688980957
transform 1 0 9752 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _2417_
timestamp 1688980957
transform 1 0 7912 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2418_
timestamp 1688980957
transform 1 0 6808 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2419_
timestamp 1688980957
transform 1 0 8464 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2420_
timestamp 1688980957
transform 1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2421_
timestamp 1688980957
transform 1 0 8832 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2422_
timestamp 1688980957
transform 1 0 6440 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2423_
timestamp 1688980957
transform 1 0 5244 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2424_
timestamp 1688980957
transform 1 0 4876 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2425_
timestamp 1688980957
transform 1 0 5244 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2426_
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _2427_
timestamp 1688980957
transform 1 0 9292 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2428_
timestamp 1688980957
transform 1 0 4692 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2429_
timestamp 1688980957
transform 1 0 9200 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2430_
timestamp 1688980957
transform 1 0 9936 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2431_
timestamp 1688980957
transform 1 0 9476 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _2432_
timestamp 1688980957
transform 1 0 5336 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2433_
timestamp 1688980957
transform 1 0 8188 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _2434_
timestamp 1688980957
transform 1 0 4784 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2435_
timestamp 1688980957
transform 1 0 10764 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _2436_
timestamp 1688980957
transform 1 0 9016 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2437_
timestamp 1688980957
transform 1 0 10120 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_4  _2438_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _2439_
timestamp 1688980957
transform 1 0 9752 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2440_
timestamp 1688980957
transform 1 0 9660 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _2441_
timestamp 1688980957
transform 1 0 9200 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2442_
timestamp 1688980957
transform 1 0 7728 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2443_
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2444_
timestamp 1688980957
transform 1 0 6900 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _2445_
timestamp 1688980957
transform 1 0 6992 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _2446_
timestamp 1688980957
transform 1 0 6440 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _2447_
timestamp 1688980957
transform 1 0 6440 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _2448_
timestamp 1688980957
transform 1 0 5520 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2449_
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2450_
timestamp 1688980957
transform 1 0 7084 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2451_
timestamp 1688980957
transform 1 0 6532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2452_
timestamp 1688980957
transform 1 0 7360 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2453_
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2454_
timestamp 1688980957
transform 1 0 7360 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2455_
timestamp 1688980957
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2456_
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2457_
timestamp 1688980957
transform 1 0 12972 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2458_
timestamp 1688980957
transform 1 0 17572 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2459_
timestamp 1688980957
transform 1 0 16744 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2460_
timestamp 1688980957
transform 1 0 21252 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a2111oi_1  _2461_
timestamp 1688980957
transform 1 0 22540 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2462_
timestamp 1688980957
transform 1 0 23644 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2463_
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2464_
timestamp 1688980957
transform 1 0 24012 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2465_
timestamp 1688980957
transform 1 0 23644 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2466_
timestamp 1688980957
transform 1 0 24012 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_1  _2467_
timestamp 1688980957
transform 1 0 23276 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _2468_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20792 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2469_
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _2470_
timestamp 1688980957
transform 1 0 12052 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2471_
timestamp 1688980957
transform 1 0 29348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2472_
timestamp 1688980957
transform 1 0 18584 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2473_
timestamp 1688980957
transform 1 0 16468 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2474_
timestamp 1688980957
transform 1 0 11776 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_2  _2475_
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _2476_
timestamp 1688980957
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2477_
timestamp 1688980957
transform 1 0 26312 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2478_
timestamp 1688980957
transform 1 0 18308 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _2479_
timestamp 1688980957
transform 1 0 18492 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _2480_
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _2481_
timestamp 1688980957
transform 1 0 20056 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _2482_
timestamp 1688980957
transform 1 0 20332 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _2483_
timestamp 1688980957
transform 1 0 21528 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2484_
timestamp 1688980957
transform 1 0 18952 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _2485_
timestamp 1688980957
transform 1 0 17572 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2486_
timestamp 1688980957
transform 1 0 18124 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2487_
timestamp 1688980957
transform 1 0 18032 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2488_
timestamp 1688980957
transform 1 0 29256 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2489_
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2490_
timestamp 1688980957
transform 1 0 30176 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2491_
timestamp 1688980957
transform 1 0 28980 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _2492_
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2493_
timestamp 1688980957
transform 1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _2494_
timestamp 1688980957
transform 1 0 15732 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2495_
timestamp 1688980957
transform 1 0 15824 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2496_
timestamp 1688980957
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2497_
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _2498_
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2499_
timestamp 1688980957
transform 1 0 20516 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2500_
timestamp 1688980957
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2501_
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2502_
timestamp 1688980957
transform 1 0 18308 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2503_
timestamp 1688980957
transform 1 0 17388 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2504_
timestamp 1688980957
transform 1 0 33396 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2505_
timestamp 1688980957
transform 1 0 17940 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _2506_
timestamp 1688980957
transform 1 0 17940 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2507_
timestamp 1688980957
transform 1 0 16836 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2508_
timestamp 1688980957
transform 1 0 18216 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2509_
timestamp 1688980957
transform 1 0 20424 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _2510_
timestamp 1688980957
transform 1 0 19872 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _2511_
timestamp 1688980957
transform 1 0 21804 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2512_
timestamp 1688980957
transform 1 0 19320 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _2513_
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2514_
timestamp 1688980957
transform 1 0 12696 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _2515_
timestamp 1688980957
transform 1 0 12236 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _2516_
timestamp 1688980957
transform 1 0 18492 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2517_
timestamp 1688980957
transform 1 0 18584 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _2518_
timestamp 1688980957
transform 1 0 19872 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _2519_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1840 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _2520_
timestamp 1688980957
transform 1 0 14628 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2521_
timestamp 1688980957
transform 1 0 18676 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _2522_
timestamp 1688980957
transform 1 0 18308 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2523_
timestamp 1688980957
transform 1 0 19964 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2524_
timestamp 1688980957
transform 1 0 23552 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _2525_
timestamp 1688980957
transform 1 0 21528 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2526_
timestamp 1688980957
transform 1 0 20884 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2527_
timestamp 1688980957
transform 1 0 20700 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2528_
timestamp 1688980957
transform 1 0 22264 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2529_
timestamp 1688980957
transform 1 0 21988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2530_
timestamp 1688980957
transform 1 0 20792 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2531_
timestamp 1688980957
transform 1 0 19136 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2532_
timestamp 1688980957
transform 1 0 19228 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _2533_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2534_
timestamp 1688980957
transform 1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _2535_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19688 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2536_
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _2537_
timestamp 1688980957
transform 1 0 18308 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2538_
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _2539_
timestamp 1688980957
transform -1 0 20792 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _2540_
timestamp 1688980957
transform 1 0 19320 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2541_
timestamp 1688980957
transform 1 0 26404 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2542_
timestamp 1688980957
transform 1 0 22356 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2543_
timestamp 1688980957
transform 1 0 22540 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2544_
timestamp 1688980957
transform 1 0 23644 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _2545_
timestamp 1688980957
transform 1 0 23092 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2546_
timestamp 1688980957
transform 1 0 22172 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2547_
timestamp 1688980957
transform 1 0 22448 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2548_
timestamp 1688980957
transform 1 0 20148 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2549_
timestamp 1688980957
transform 1 0 20976 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2550_
timestamp 1688980957
transform 1 0 2852 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2551_
timestamp 1688980957
transform 1 0 2208 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2552_
timestamp 1688980957
transform 1 0 19504 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2553_
timestamp 1688980957
transform 1 0 19320 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2554_
timestamp 1688980957
transform 1 0 18308 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2555_
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2556_
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2557_
timestamp 1688980957
transform 1 0 5520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2558_
timestamp 1688980957
transform 1 0 23000 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2559_
timestamp 1688980957
transform 1 0 22908 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2560_
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2561_
timestamp 1688980957
transform 1 0 3404 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2562_
timestamp 1688980957
transform 1 0 25668 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o221ai_1  _2563_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22816 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _2564_
timestamp 1688980957
transform 1 0 22264 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _2565_
timestamp 1688980957
transform 1 0 21528 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _2566_
timestamp 1688980957
transform 1 0 17940 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2oi_4  _2567_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21436 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__a31o_1  _2568_
timestamp 1688980957
transform 1 0 21160 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2569_
timestamp 1688980957
transform 1 0 31648 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2570_
timestamp 1688980957
transform 1 0 24380 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _2571_
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _2572_
timestamp 1688980957
transform 1 0 25668 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2573_
timestamp 1688980957
transform 1 0 24748 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2574_
timestamp 1688980957
transform 1 0 28152 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2575_
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _2576_
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2577_
timestamp 1688980957
transform 1 0 22632 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2578_
timestamp 1688980957
transform 1 0 23736 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2579_
timestamp 1688980957
transform 1 0 24196 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2580_
timestamp 1688980957
transform 1 0 23460 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2581_
timestamp 1688980957
transform 1 0 23828 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _2582_
timestamp 1688980957
transform 1 0 23460 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _2583_
timestamp 1688980957
transform 1 0 22540 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2b_2  _2584_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _2585_
timestamp 1688980957
transform 1 0 16928 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2586_
timestamp 1688980957
transform 1 0 7912 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2587_
timestamp 1688980957
transform 1 0 12236 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _2588_
timestamp 1688980957
transform 1 0 16928 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2b_2  _2589_
timestamp 1688980957
transform 1 0 10488 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2590_
timestamp 1688980957
transform 1 0 11868 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _2591_
timestamp 1688980957
transform 1 0 10672 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _2592_
timestamp 1688980957
transform 1 0 10764 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2593_
timestamp 1688980957
transform 1 0 12512 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _2594_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11960 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2595_
timestamp 1688980957
transform 1 0 20240 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2596_
timestamp 1688980957
transform 1 0 19780 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2597_
timestamp 1688980957
transform 1 0 15916 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2598_
timestamp 1688980957
transform 1 0 10764 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2599_
timestamp 1688980957
transform 1 0 7728 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2600_
timestamp 1688980957
transform 1 0 14996 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2601_
timestamp 1688980957
transform 1 0 15824 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2602_
timestamp 1688980957
transform 1 0 15272 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _2603_
timestamp 1688980957
transform 1 0 12420 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _2604_
timestamp 1688980957
transform 1 0 12144 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2605_
timestamp 1688980957
transform 1 0 11224 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2606_
timestamp 1688980957
transform 1 0 10856 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2607_
timestamp 1688980957
transform 1 0 16284 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2608_
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2609_
timestamp 1688980957
transform 1 0 15180 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2610_
timestamp 1688980957
transform 1 0 14352 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2611_
timestamp 1688980957
transform 1 0 14076 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2612_
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2613_
timestamp 1688980957
transform 1 0 16928 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2614_
timestamp 1688980957
transform 1 0 10856 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2615_
timestamp 1688980957
transform 1 0 10580 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2616_
timestamp 1688980957
transform 1 0 9752 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2617_
timestamp 1688980957
transform 1 0 17480 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2618_
timestamp 1688980957
transform 1 0 7912 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2619_
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2620_
timestamp 1688980957
transform 1 0 11224 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2621_
timestamp 1688980957
transform 1 0 11132 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2622_
timestamp 1688980957
transform 1 0 15824 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2623_
timestamp 1688980957
transform 1 0 14720 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2624_
timestamp 1688980957
transform 1 0 14260 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2625_
timestamp 1688980957
transform 1 0 14536 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2626_
timestamp 1688980957
transform 1 0 15548 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2627_
timestamp 1688980957
transform 1 0 14720 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2628_
timestamp 1688980957
transform 1 0 15824 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2629_
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2630_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18952 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2631_
timestamp 1688980957
transform 1 0 20424 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2632_
timestamp 1688980957
transform 1 0 19872 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2633_
timestamp 1688980957
transform 1 0 19688 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2634_
timestamp 1688980957
transform 1 0 18124 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2635_
timestamp 1688980957
transform 1 0 19412 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _2636_
timestamp 1688980957
transform 1 0 18400 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2637_
timestamp 1688980957
transform 1 0 17204 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2638_
timestamp 1688980957
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_4  _2639_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14996 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_1  _2640_
timestamp 1688980957
transform 1 0 16652 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _2641_
timestamp 1688980957
transform 1 0 15088 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2642_
timestamp 1688980957
transform 1 0 10580 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2643_
timestamp 1688980957
transform 1 0 9844 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _2644_
timestamp 1688980957
transform 1 0 16744 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _2645_
timestamp 1688980957
transform 1 0 10120 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2646_
timestamp 1688980957
transform 1 0 10396 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2647_
timestamp 1688980957
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2648_
timestamp 1688980957
transform 1 0 10856 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2649_
timestamp 1688980957
transform 1 0 11316 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2650_
timestamp 1688980957
transform 1 0 11776 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2651_
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2652_
timestamp 1688980957
transform 1 0 13800 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _2653_
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2654_
timestamp 1688980957
transform 1 0 10488 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2655_
timestamp 1688980957
transform 1 0 9568 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2656_
timestamp 1688980957
transform 1 0 9844 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2657_
timestamp 1688980957
transform 1 0 10212 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2658_
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2659_
timestamp 1688980957
transform 1 0 11960 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2660_
timestamp 1688980957
transform 1 0 9384 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _2661_
timestamp 1688980957
transform 1 0 9660 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _2662_
timestamp 1688980957
transform 1 0 9844 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2663_
timestamp 1688980957
transform 1 0 9476 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2664_
timestamp 1688980957
transform 1 0 9660 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2665_
timestamp 1688980957
transform 1 0 9568 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2666_
timestamp 1688980957
transform 1 0 8096 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2667_
timestamp 1688980957
transform 1 0 7360 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2668_
timestamp 1688980957
transform 1 0 10856 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _2669_
timestamp 1688980957
transform 1 0 11040 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2670_
timestamp 1688980957
transform 1 0 7360 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2671_
timestamp 1688980957
transform 1 0 8464 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _2672_
timestamp 1688980957
transform 1 0 7820 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2673_
timestamp 1688980957
transform 1 0 8372 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2674_
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2675_
timestamp 1688980957
transform 1 0 7268 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2676_
timestamp 1688980957
transform 1 0 6808 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _2677_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7544 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _2678_
timestamp 1688980957
transform 1 0 6256 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2679_
timestamp 1688980957
transform 1 0 13524 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _2680_
timestamp 1688980957
transform 1 0 13156 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2681_
timestamp 1688980957
transform 1 0 13432 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2682_
timestamp 1688980957
transform 1 0 11776 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2683_
timestamp 1688980957
transform 1 0 16100 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _2684_
timestamp 1688980957
transform 1 0 11500 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _2685_
timestamp 1688980957
transform 1 0 9936 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_1  _2686_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2687_
timestamp 1688980957
transform 1 0 9568 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2688_
timestamp 1688980957
transform 1 0 8740 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2689_
timestamp 1688980957
transform 1 0 9384 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2690_
timestamp 1688980957
transform 1 0 6900 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2691_
timestamp 1688980957
transform 1 0 5244 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2692_
timestamp 1688980957
transform 1 0 4692 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2693_
timestamp 1688980957
transform 1 0 6348 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2694_
timestamp 1688980957
transform 1 0 6716 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2695_
timestamp 1688980957
transform 1 0 7636 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2696_
timestamp 1688980957
transform 1 0 6716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _2697_
timestamp 1688980957
transform 1 0 8648 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _2698_
timestamp 1688980957
transform 1 0 7176 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2699_
timestamp 1688980957
transform 1 0 8740 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2700_
timestamp 1688980957
transform 1 0 6716 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2701_
timestamp 1688980957
transform 1 0 7544 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2702_
timestamp 1688980957
transform 1 0 6992 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2703_
timestamp 1688980957
transform 1 0 6808 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2704_
timestamp 1688980957
transform 1 0 7268 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2705_
timestamp 1688980957
transform 1 0 6440 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2706_
timestamp 1688980957
transform 1 0 6624 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2707_
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2708_
timestamp 1688980957
transform 1 0 7268 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2709_
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2710_
timestamp 1688980957
transform 1 0 4508 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2711_
timestamp 1688980957
transform 1 0 4140 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2712_
timestamp 1688980957
transform 1 0 5336 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2713_
timestamp 1688980957
transform 1 0 5888 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2714_
timestamp 1688980957
transform 1 0 4784 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _2715_
timestamp 1688980957
transform 1 0 5152 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2716_
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2717_
timestamp 1688980957
transform 1 0 4232 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2718_
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2719_
timestamp 1688980957
transform 1 0 6532 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2720_
timestamp 1688980957
transform 1 0 6348 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2721_
timestamp 1688980957
transform 1 0 5060 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2722_
timestamp 1688980957
transform 1 0 4232 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2723_
timestamp 1688980957
transform 1 0 4508 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _2724_
timestamp 1688980957
transform 1 0 4968 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _2725_
timestamp 1688980957
transform 1 0 5336 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _2726_
timestamp 1688980957
transform 1 0 4600 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2727_
timestamp 1688980957
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2728_
timestamp 1688980957
transform 1 0 6992 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _2729_
timestamp 1688980957
transform 1 0 7176 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _2730_
timestamp 1688980957
transform 1 0 7912 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _2731_
timestamp 1688980957
transform 1 0 8740 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2732_
timestamp 1688980957
transform 1 0 9752 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2733_
timestamp 1688980957
transform 1 0 5244 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2734_
timestamp 1688980957
transform 1 0 4784 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2735_
timestamp 1688980957
transform 1 0 6072 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2736_
timestamp 1688980957
transform 1 0 4784 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _2737_
timestamp 1688980957
transform 1 0 4876 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2738_
timestamp 1688980957
transform 1 0 5888 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _2739_
timestamp 1688980957
transform 1 0 9016 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2740_
timestamp 1688980957
transform 1 0 27784 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_2  _2741_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28060 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _2742_
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2743_
timestamp 1688980957
transform 1 0 8372 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2744_
timestamp 1688980957
transform 1 0 7176 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2745_
timestamp 1688980957
transform 1 0 15088 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2746_
timestamp 1688980957
transform 1 0 14996 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2747_
timestamp 1688980957
transform 1 0 6716 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2748_
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2749_
timestamp 1688980957
transform 1 0 11224 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2750_
timestamp 1688980957
transform 1 0 10580 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2751_
timestamp 1688980957
transform 1 0 4784 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2752_
timestamp 1688980957
transform 1 0 4508 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2753_
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2754_
timestamp 1688980957
transform 1 0 2392 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2755_
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2756_
timestamp 1688980957
transform 1 0 1840 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2757_
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2758_
timestamp 1688980957
transform 1 0 1840 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2759_
timestamp 1688980957
transform 1 0 31004 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2760_
timestamp 1688980957
transform 1 0 30360 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2761_
timestamp 1688980957
transform 1 0 16928 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2762_
timestamp 1688980957
transform 1 0 16376 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2763_
timestamp 1688980957
transform 1 0 8740 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2764_
timestamp 1688980957
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2765_
timestamp 1688980957
transform 1 0 14076 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2766_
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2767_
timestamp 1688980957
transform 1 0 6900 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2768_
timestamp 1688980957
transform 1 0 7084 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2769_
timestamp 1688980957
transform 1 0 11776 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2770_
timestamp 1688980957
transform 1 0 10488 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2771_
timestamp 1688980957
transform 1 0 4968 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2772_
timestamp 1688980957
transform 1 0 4692 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2773_
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2774_
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2775_
timestamp 1688980957
transform 1 0 2208 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2776_
timestamp 1688980957
transform 1 0 1840 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2777_
timestamp 1688980957
transform 1 0 2484 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2778_
timestamp 1688980957
transform 1 0 1840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2779_
timestamp 1688980957
transform 1 0 21528 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2780_
timestamp 1688980957
transform 1 0 24564 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2781_
timestamp 1688980957
transform 1 0 25392 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2782_
timestamp 1688980957
transform 1 0 24932 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2783_
timestamp 1688980957
transform 1 0 23000 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2784_
timestamp 1688980957
transform 1 0 31464 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _2785_
timestamp 1688980957
transform 1 0 24472 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2786_
timestamp 1688980957
transform 1 0 25208 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2787_
timestamp 1688980957
transform 1 0 25116 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2788_
timestamp 1688980957
transform 1 0 23828 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2789_
timestamp 1688980957
transform 1 0 27508 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _2790_
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _2791_
timestamp 1688980957
transform 1 0 27232 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2792_
timestamp 1688980957
transform 1 0 27692 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2793_
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_4  _2794_
timestamp 1688980957
transform 1 0 24196 0 -1 29376
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _2795_
timestamp 1688980957
transform 1 0 2116 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2796_
timestamp 1688980957
transform 1 0 1840 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2797_
timestamp 1688980957
transform 1 0 2484 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2798_
timestamp 1688980957
transform 1 0 2024 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2799_
timestamp 1688980957
transform 1 0 2944 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2800_
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2801_
timestamp 1688980957
transform 1 0 19412 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2802_
timestamp 1688980957
transform 1 0 19504 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2803_
timestamp 1688980957
transform 1 0 2760 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2804_
timestamp 1688980957
transform 1 0 2300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2805_
timestamp 1688980957
transform 1 0 2392 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2806_
timestamp 1688980957
transform 1 0 1840 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2807_
timestamp 1688980957
transform 1 0 4600 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2808_
timestamp 1688980957
transform 1 0 4232 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2809_
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2810_
timestamp 1688980957
transform 1 0 2760 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2811_
timestamp 1688980957
transform 1 0 17848 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2812_
timestamp 1688980957
transform 1 0 18308 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2813_
timestamp 1688980957
transform 1 0 18676 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2814_
timestamp 1688980957
transform 1 0 15732 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2815_
timestamp 1688980957
transform 1 0 15824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2816_
timestamp 1688980957
transform 1 0 15916 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2817_
timestamp 1688980957
transform 1 0 19136 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2818_
timestamp 1688980957
transform 1 0 17572 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2819_
timestamp 1688980957
transform 1 0 17664 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2820_
timestamp 1688980957
transform 1 0 16928 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2821_
timestamp 1688980957
transform 1 0 16376 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2822_
timestamp 1688980957
transform 1 0 17940 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2823_
timestamp 1688980957
transform 1 0 18768 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2824_
timestamp 1688980957
transform 1 0 18400 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2825_
timestamp 1688980957
transform 1 0 15456 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2826_
timestamp 1688980957
transform 1 0 16284 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _2827_
timestamp 1688980957
transform 1 0 17020 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2828_
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2829_
timestamp 1688980957
transform 1 0 18860 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2830_
timestamp 1688980957
transform 1 0 17756 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _2831_
timestamp 1688980957
transform 1 0 18124 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _2832_
timestamp 1688980957
transform 1 0 14444 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _2833_
timestamp 1688980957
transform 1 0 14168 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2834_
timestamp 1688980957
transform 1 0 17480 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2835_
timestamp 1688980957
transform 1 0 17204 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2836_
timestamp 1688980957
transform 1 0 17848 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2837_
timestamp 1688980957
transform 1 0 13800 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2838_
timestamp 1688980957
transform 1 0 12880 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2839_
timestamp 1688980957
transform 1 0 14536 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2840_
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _2841_
timestamp 1688980957
transform 1 0 13432 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2842_
timestamp 1688980957
transform 1 0 16192 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2843_
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2844_
timestamp 1688980957
transform 1 0 14168 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2845_
timestamp 1688980957
transform 1 0 12880 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2846_
timestamp 1688980957
transform 1 0 12420 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2847_
timestamp 1688980957
transform 1 0 15180 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2848_
timestamp 1688980957
transform 1 0 14260 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2849_
timestamp 1688980957
transform 1 0 14536 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2850_
timestamp 1688980957
transform 1 0 14352 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2851_
timestamp 1688980957
transform 1 0 13156 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2852_
timestamp 1688980957
transform 1 0 12420 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2853_
timestamp 1688980957
transform 1 0 11776 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2854_
timestamp 1688980957
transform 1 0 11684 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2855_
timestamp 1688980957
transform 1 0 11960 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2856_
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2857_
timestamp 1688980957
transform 1 0 11776 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2858_
timestamp 1688980957
transform 1 0 13064 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2859_
timestamp 1688980957
transform 1 0 15272 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2860_
timestamp 1688980957
transform 1 0 15364 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _2861_
timestamp 1688980957
transform 1 0 15824 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2862_
timestamp 1688980957
transform 1 0 12788 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2863_
timestamp 1688980957
transform 1 0 14812 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2864_
timestamp 1688980957
transform 1 0 15732 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2865_
timestamp 1688980957
transform 1 0 16284 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2866_
timestamp 1688980957
transform 1 0 12512 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2867_
timestamp 1688980957
transform 1 0 16284 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2868_
timestamp 1688980957
transform 1 0 17020 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2869_
timestamp 1688980957
transform 1 0 16836 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2870_
timestamp 1688980957
transform 1 0 17296 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _2871_
timestamp 1688980957
transform 1 0 30268 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2872_
timestamp 1688980957
transform 1 0 30176 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_4  _2873_
timestamp 1688980957
transform 1 0 29256 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _2874_
timestamp 1688980957
transform 1 0 8832 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2875_
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2876_
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2877_
timestamp 1688980957
transform 1 0 13524 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2878_
timestamp 1688980957
transform 1 0 6624 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2879_
timestamp 1688980957
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2880_
timestamp 1688980957
transform 1 0 12144 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2881_
timestamp 1688980957
transform 1 0 12512 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2882_
timestamp 1688980957
transform 1 0 4140 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2883_
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2884_
timestamp 1688980957
transform 1 0 2852 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2885_
timestamp 1688980957
transform 1 0 2116 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2886_
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2887_
timestamp 1688980957
transform 1 0 1840 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2888_
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2889_
timestamp 1688980957
transform 1 0 2760 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2890_
timestamp 1688980957
transform 1 0 23460 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2891_
timestamp 1688980957
transform 1 0 23368 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _2892_
timestamp 1688980957
transform 1 0 22540 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _2893_
timestamp 1688980957
transform 1 0 22908 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2894_
timestamp 1688980957
transform 1 0 24472 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2895_
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _2896_
timestamp 1688980957
transform 1 0 23460 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o41a_1  _2897_
timestamp 1688980957
transform 1 0 23276 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _2898_
timestamp 1688980957
transform 1 0 22448 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _2899_
timestamp 1688980957
transform 1 0 21160 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _2900_
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2901_
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2902_
timestamp 1688980957
transform 1 0 12512 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2903_
timestamp 1688980957
transform 1 0 12788 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2904_
timestamp 1688980957
transform 1 0 22632 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2905_
timestamp 1688980957
transform 1 0 22356 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2906_
timestamp 1688980957
transform 1 0 12604 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2907_
timestamp 1688980957
transform 1 0 12236 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2908_
timestamp 1688980957
transform 1 0 14812 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2909_
timestamp 1688980957
transform 1 0 14076 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2910_
timestamp 1688980957
transform 1 0 22264 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2911_
timestamp 1688980957
transform 1 0 21528 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2912_
timestamp 1688980957
transform 1 0 21068 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _2913_
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _2914_
timestamp 1688980957
transform 1 0 21712 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_4  _2915_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21436 0 1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__or2b_1  _2916_
timestamp 1688980957
transform 1 0 14720 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _2917_
timestamp 1688980957
transform 1 0 14076 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2918_
timestamp 1688980957
transform 1 0 14260 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2919_
timestamp 1688980957
transform 1 0 16008 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _2920_
timestamp 1688980957
transform 1 0 19136 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2921_
timestamp 1688980957
transform 1 0 15272 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _2922_
timestamp 1688980957
transform 1 0 15456 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _2923_
timestamp 1688980957
transform 1 0 14536 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2924_
timestamp 1688980957
transform 1 0 13984 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2925_
timestamp 1688980957
transform 1 0 11408 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2926_
timestamp 1688980957
transform 1 0 16100 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2927_
timestamp 1688980957
transform 1 0 15088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2928_
timestamp 1688980957
transform 1 0 16744 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _2929_
timestamp 1688980957
transform 1 0 15548 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _2930_
timestamp 1688980957
transform 1 0 16468 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _2931_
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _2932_
timestamp 1688980957
transform 1 0 15732 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2933_
timestamp 1688980957
transform 1 0 16100 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _2934_
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2935_
timestamp 1688980957
transform 1 0 15456 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2936_
timestamp 1688980957
transform 1 0 13524 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2937_
timestamp 1688980957
transform 1 0 12788 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2938_
timestamp 1688980957
transform 1 0 12420 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _2939_
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2940_
timestamp 1688980957
transform 1 0 13984 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _2941_
timestamp 1688980957
transform 1 0 17296 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2942_
timestamp 1688980957
transform 1 0 13248 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2943_
timestamp 1688980957
transform 1 0 13524 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2944_
timestamp 1688980957
transform 1 0 14904 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _2945_
timestamp 1688980957
transform 1 0 13892 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2946_
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2947_
timestamp 1688980957
transform 1 0 10396 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2948_
timestamp 1688980957
transform 1 0 9568 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2949_
timestamp 1688980957
transform 1 0 12788 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2950_
timestamp 1688980957
transform 1 0 12052 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _2951_
timestamp 1688980957
transform 1 0 12052 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2952_
timestamp 1688980957
transform 1 0 11040 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2953_
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2954_
timestamp 1688980957
transform 1 0 10948 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2955_
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _2956_
timestamp 1688980957
transform 1 0 11592 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2957_
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2958_
timestamp 1688980957
transform 1 0 11316 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2959_
timestamp 1688980957
transform 1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2960_
timestamp 1688980957
transform 1 0 8740 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2961_
timestamp 1688980957
transform 1 0 9568 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2962_
timestamp 1688980957
transform 1 0 8832 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2963_
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2964_
timestamp 1688980957
transform 1 0 7084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _2965_
timestamp 1688980957
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _2966_
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2967_
timestamp 1688980957
transform 1 0 8004 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2968_
timestamp 1688980957
transform 1 0 7820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _2969_
timestamp 1688980957
transform 1 0 7912 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2970_
timestamp 1688980957
transform 1 0 8924 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _2971_
timestamp 1688980957
transform 1 0 8372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2972_
timestamp 1688980957
transform 1 0 7912 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _2973_
timestamp 1688980957
transform 1 0 7176 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _2974_
timestamp 1688980957
transform 1 0 6716 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2975_
timestamp 1688980957
transform 1 0 5152 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2976_
timestamp 1688980957
transform 1 0 4692 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2977_
timestamp 1688980957
transform 1 0 5796 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2978_
timestamp 1688980957
transform 1 0 5612 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2979_
timestamp 1688980957
transform 1 0 8372 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2980_
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2981_
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2982_
timestamp 1688980957
transform 1 0 8004 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2983_
timestamp 1688980957
transform 1 0 7544 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2984_
timestamp 1688980957
transform 1 0 7360 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2985_
timestamp 1688980957
transform 1 0 6256 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2986_
timestamp 1688980957
transform 1 0 2852 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2987_
timestamp 1688980957
transform 1 0 3496 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2988_
timestamp 1688980957
transform 1 0 5704 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _2989_
timestamp 1688980957
transform 1 0 5244 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a311oi_1  _2990_
timestamp 1688980957
transform 1 0 3956 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2991_
timestamp 1688980957
transform 1 0 4692 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _2992_
timestamp 1688980957
transform 1 0 4324 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2993_
timestamp 1688980957
transform 1 0 4600 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2994_
timestamp 1688980957
transform 1 0 5428 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2995_
timestamp 1688980957
transform 1 0 10304 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2996_
timestamp 1688980957
transform 1 0 10396 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2997_
timestamp 1688980957
transform 1 0 10856 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _2998_
timestamp 1688980957
transform 1 0 12328 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2999_
timestamp 1688980957
transform 1 0 10580 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _3000_
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _3001_
timestamp 1688980957
transform 1 0 9844 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _3002_
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _3003_
timestamp 1688980957
transform 1 0 30176 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _3004_
timestamp 1688980957
transform 1 0 29624 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _3005_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _3006_
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _3007_
timestamp 1688980957
transform 1 0 8464 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _3008_
timestamp 1688980957
transform 1 0 14076 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _3009_
timestamp 1688980957
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _3010_
timestamp 1688980957
transform 1 0 7084 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _3011_
timestamp 1688980957
transform 1 0 6716 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _3012_
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _3013_
timestamp 1688980957
transform 1 0 10948 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _3014_
timestamp 1688980957
transform 1 0 5428 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _3015_
timestamp 1688980957
transform 1 0 5888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _3016_
timestamp 1688980957
transform 1 0 4324 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _3017_
timestamp 1688980957
transform 1 0 3956 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _3018_
timestamp 1688980957
transform 1 0 2668 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _3019_
timestamp 1688980957
transform 1 0 2024 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _3020_
timestamp 1688980957
transform 1 0 2760 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _3021_
timestamp 1688980957
transform 1 0 2208 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _3022_
timestamp 1688980957
transform 1 0 17940 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _3023_
timestamp 1688980957
transform 1 0 17572 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _3024_
timestamp 1688980957
transform 1 0 33856 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _3025_
timestamp 1688980957
transform 1 0 27600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _3026_
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _3027_
timestamp 1688980957
transform 1 0 20792 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _3028_
timestamp 1688980957
transform 1 0 19412 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _3029_
timestamp 1688980957
transform 1 0 16928 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _3030_
timestamp 1688980957
transform 1 0 17204 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _3031_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31832 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _3032_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _3033_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33304 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3034_
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3035_
timestamp 1688980957
transform 1 0 24472 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _3036_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28336 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3037_
timestamp 1688980957
transform 1 0 27416 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _3038_
timestamp 1688980957
transform 1 0 24196 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3039_
timestamp 1688980957
transform 1 0 35144 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3040_
timestamp 1688980957
transform 1 0 29992 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3041_
timestamp 1688980957
transform 1 0 26036 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3042_
timestamp 1688980957
transform 1 0 26036 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _3043_
timestamp 1688980957
transform 1 0 23460 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _3044_
timestamp 1688980957
transform 1 0 29808 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _3045_
timestamp 1688980957
transform 1 0 23736 0 -1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _3046_
timestamp 1688980957
transform 1 0 27600 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3047_
timestamp 1688980957
transform 1 0 25852 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _3048_
timestamp 1688980957
transform 1 0 27876 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _3049_
timestamp 1688980957
transform 1 0 24656 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _3050_
timestamp 1688980957
transform 1 0 26956 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _3051_
timestamp 1688980957
transform 1 0 18768 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _3052_
timestamp 1688980957
transform 1 0 39008 0 -1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _3053_
timestamp 1688980957
transform 1 0 39284 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3054_
timestamp 1688980957
transform 1 0 39008 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3055_
timestamp 1688980957
transform 1 0 39284 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3056_
timestamp 1688980957
transform 1 0 39284 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3057_
timestamp 1688980957
transform 1 0 39284 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _3058_
timestamp 1688980957
transform 1 0 17572 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3059_
timestamp 1688980957
transform 1 0 15364 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _3060_
timestamp 1688980957
transform 1 0 17388 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _3061_
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _3062_
timestamp 1688980957
transform 1 0 18400 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _3063_
timestamp 1688980957
transform 1 0 19596 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _3064_
timestamp 1688980957
transform 1 0 22264 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _3065_
timestamp 1688980957
transform 1 0 17296 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3066_
timestamp 1688980957
transform 1 0 20792 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _3067_
timestamp 1688980957
transform 1 0 19964 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _3068_
timestamp 1688980957
transform 1 0 18124 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3069_
timestamp 1688980957
transform 1 0 19596 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _3070_
timestamp 1688980957
transform 1 0 38824 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _3071_
timestamp 1688980957
transform 1 0 39192 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _3072_
timestamp 1688980957
transform 1 0 1840 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3073_
timestamp 1688980957
transform 1 0 16008 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3074_
timestamp 1688980957
transform 1 0 21988 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3075_
timestamp 1688980957
transform 1 0 19320 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3076_
timestamp 1688980957
transform 1 0 1472 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3077_
timestamp 1688980957
transform 1 0 19596 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3078_
timestamp 1688980957
transform 1 0 18124 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3079_
timestamp 1688980957
transform 1 0 5152 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3080_
timestamp 1688980957
transform 1 0 23184 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3081_
timestamp 1688980957
transform 1 0 2300 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _3082_
timestamp 1688980957
transform 1 0 9844 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _3083_
timestamp 1688980957
transform 1 0 12604 0 -1 39168
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3084_
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3085_
timestamp 1688980957
transform 1 0 4140 0 -1 39168
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _3086_
timestamp 1688980957
transform 1 0 4324 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _3087_
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _3088_
timestamp 1688980957
transform 1 0 6624 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _3089_
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _3090_
timestamp 1688980957
transform 1 0 6532 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3091_
timestamp 1688980957
transform 1 0 14720 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3092_
timestamp 1688980957
transform 1 0 5888 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3093_
timestamp 1688980957
transform 1 0 10212 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3094_
timestamp 1688980957
transform 1 0 4140 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3095_
timestamp 1688980957
transform 1 0 2668 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3096_
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3097_
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3098_
timestamp 1688980957
transform 1 0 8004 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3099_
timestamp 1688980957
transform 1 0 13156 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3100_
timestamp 1688980957
transform 1 0 6072 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3101_
timestamp 1688980957
transform 1 0 9936 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3102_
timestamp 1688980957
transform 1 0 4232 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3103_
timestamp 1688980957
transform 1 0 3036 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3104_
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3105_
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _3106_
timestamp 1688980957
transform 1 0 21712 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3107_
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3108_
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3109_
timestamp 1688980957
transform 1 0 1564 0 1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3110_
timestamp 1688980957
transform 1 0 19320 0 1 41344
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3111_
timestamp 1688980957
transform 1 0 1748 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3112_
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3113_
timestamp 1688980957
transform 1 0 3772 0 -1 41344
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3114_
timestamp 1688980957
transform 1 0 2208 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3115_
timestamp 1688980957
transform 1 0 19412 0 1 40256
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3116_
timestamp 1688980957
transform 1 0 16928 0 1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3117_
timestamp 1688980957
transform 1 0 19596 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3118_
timestamp 1688980957
transform 1 0 18032 0 -1 39168
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _3119_
timestamp 1688980957
transform 1 0 14168 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _3120_
timestamp 1688980957
transform 1 0 12052 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3121_
timestamp 1688980957
transform 1 0 12880 0 -1 40256
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3122_
timestamp 1688980957
transform 1 0 16836 0 1 41344
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _3123_
timestamp 1688980957
transform 1 0 8096 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _3124_
timestamp 1688980957
transform 1 0 13064 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3125_
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3126_
timestamp 1688980957
transform 1 0 11592 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3127_
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3128_
timestamp 1688980957
transform 1 0 1472 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3129_
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3130_
timestamp 1688980957
transform 1 0 2392 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _3131_
timestamp 1688980957
transform 1 0 21804 0 -1 41344
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3132_
timestamp 1688980957
transform 1 0 21160 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3133_
timestamp 1688980957
transform 1 0 16100 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3134_
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3135_
timestamp 1688980957
transform 1 0 22172 0 1 41344
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3136_
timestamp 1688980957
transform 1 0 11776 0 1 41344
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3137_
timestamp 1688980957
transform 1 0 14076 0 1 41344
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _3138_
timestamp 1688980957
transform 1 0 21804 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _3139_
timestamp 1688980957
transform 1 0 12144 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _3140_
timestamp 1688980957
transform 1 0 15640 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _3141_
timestamp 1688980957
transform 1 0 9108 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3142_
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _3143_
timestamp 1688980957
transform 1 0 8280 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _3144_
timestamp 1688980957
transform 1 0 4140 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _3145_
timestamp 1688980957
transform 1 0 3404 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _3146_
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3147_
timestamp 1688980957
transform 1 0 20240 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3148_
timestamp 1688980957
transform 1 0 21160 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3149_
timestamp 1688980957
transform 1 0 8004 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3150_
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3151_
timestamp 1688980957
transform 1 0 6256 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3152_
timestamp 1688980957
transform 1 0 10396 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3153_
timestamp 1688980957
transform 1 0 4600 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3154_
timestamp 1688980957
transform 1 0 3496 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3155_
timestamp 1688980957
transform 1 0 1564 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3156_
timestamp 1688980957
transform 1 0 1748 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _3157_
timestamp 1688980957
transform 1 0 16928 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _3158_
timestamp 1688980957
transform 1 0 26128 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _3159_
timestamp 1688980957
transform 1 0 16928 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__buf_2  _3160_
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23092 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 34868 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform -1 0 35144 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1688980957
transform -1 0 19872 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1688980957
transform 1 0 35604 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21252 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2668 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1688980957
transform 1 0 2944 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1688980957
transform 1 0 5888 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1688980957
transform 1 0 10028 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1688980957
transform 1 0 7820 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1688980957
transform 1 0 7452 0 -1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1688980957
transform 1 0 17848 0 1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1688980957
transform 1 0 19964 0 -1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1688980957
transform 1 0 19136 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1688980957
transform 1 0 21896 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1688980957
transform 1 0 24288 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1688980957
transform 1 0 25852 0 -1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1688980957
transform 1 0 35696 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1688980957
transform 1 0 34868 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout34
timestamp 1688980957
transform 1 0 5612 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout35
timestamp 1688980957
transform 1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout36
timestamp 1688980957
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout38
timestamp 1688980957
transform 1 0 20056 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout39
timestamp 1688980957
transform 1 0 19780 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout40
timestamp 1688980957
transform 1 0 7452 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout41
timestamp 1688980957
transform 1 0 6716 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout42
timestamp 1688980957
transform 1 0 20792 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout43
timestamp 1688980957
transform 1 0 16560 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout44
timestamp 1688980957
transform 1 0 18124 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout45
timestamp 1688980957
transform 1 0 25392 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout46
timestamp 1688980957
transform 1 0 28612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout47
timestamp 1688980957
transform 1 0 35972 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout48
timestamp 1688980957
transform 1 0 31740 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 1688980957
transform 1 0 40572 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout50
timestamp 1688980957
transform 1 0 40572 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_72
timestamp 1688980957
transform 1 0 7728 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_225 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_233
timestamp 1688980957
transform 1 0 22540 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_245 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1688980957
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1688980957
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1688980957
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_315
timestamp 1688980957
transform 1 0 30084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_327
timestamp 1688980957
transform 1 0 31188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_335
timestamp 1688980957
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_345
timestamp 1688980957
transform 1 0 32844 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_352
timestamp 1688980957
transform 1 0 33488 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 1688980957
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_393
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_405
timestamp 1688980957
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_417
timestamp 1688980957
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_144
timestamp 1688980957
transform 1 0 14352 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_156
timestamp 1688980957
transform 1 0 15456 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_429
timestamp 1688980957
transform 1 0 40572 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_152
timestamp 1688980957
transform 1 0 15088 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_164
timestamp 1688980957
transform 1 0 16192 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_176
timestamp 1688980957
transform 1 0 17296 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_188
timestamp 1688980957
transform 1 0 18400 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_7
timestamp 1688980957
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_11
timestamp 1688980957
transform 1 0 2116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_23
timestamp 1688980957
transform 1 0 3220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_35
timestamp 1688980957
transform 1 0 4324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_47
timestamp 1688980957
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_109
timestamp 1688980957
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_323
timestamp 1688980957
transform 1 0 30820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_429
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_7
timestamp 1688980957
transform 1 0 1748 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_161
timestamp 1688980957
transform 1 0 15916 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_182
timestamp 1688980957
transform 1 0 17848 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_194
timestamp 1688980957
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_271
timestamp 1688980957
transform 1 0 26036 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_293
timestamp 1688980957
transform 1 0 28060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_305
timestamp 1688980957
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_313
timestamp 1688980957
transform 1 0 29900 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_355
timestamp 1688980957
transform 1 0 33764 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_383
timestamp 1688980957
transform 1 0 36340 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_395
timestamp 1688980957
transform 1 0 37444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_407
timestamp 1688980957
transform 1 0 38548 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_89
timestamp 1688980957
transform 1 0 9292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_95
timestamp 1688980957
transform 1 0 9844 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_104
timestamp 1688980957
transform 1 0 10672 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_133
timestamp 1688980957
transform 1 0 13340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_145
timestamp 1688980957
transform 1 0 14444 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_157
timestamp 1688980957
transform 1 0 15548 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_165
timestamp 1688980957
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_175
timestamp 1688980957
transform 1 0 17204 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_183
timestamp 1688980957
transform 1 0 17940 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_233
timestamp 1688980957
transform 1 0 22540 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_245
timestamp 1688980957
transform 1 0 23644 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_257
timestamp 1688980957
transform 1 0 24748 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_269
timestamp 1688980957
transform 1 0 25852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_277
timestamp 1688980957
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_292
timestamp 1688980957
transform 1 0 27968 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_319
timestamp 1688980957
transform 1 0 30452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_323
timestamp 1688980957
transform 1 0 30820 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_333
timestamp 1688980957
transform 1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_347
timestamp 1688980957
transform 1 0 33028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_390
timestamp 1688980957
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_107
timestamp 1688980957
transform 1 0 10948 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_119
timestamp 1688980957
transform 1 0 12052 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_131
timestamp 1688980957
transform 1 0 13156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_161
timestamp 1688980957
transform 1 0 15916 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_186
timestamp 1688980957
transform 1 0 18216 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_194
timestamp 1688980957
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_241
timestamp 1688980957
transform 1 0 23276 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_249
timestamp 1688980957
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_285
timestamp 1688980957
transform 1 0 27324 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_303
timestamp 1688980957
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_327
timestamp 1688980957
transform 1 0 31188 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_339
timestamp 1688980957
transform 1 0 32292 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_347
timestamp 1688980957
transform 1 0 33028 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_362
timestamp 1688980957
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_369
timestamp 1688980957
transform 1 0 35052 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_376
timestamp 1688980957
transform 1 0 35696 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_380
timestamp 1688980957
transform 1 0 36064 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_429
timestamp 1688980957
transform 1 0 40572 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_47
timestamp 1688980957
transform 1 0 5428 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_66
timestamp 1688980957
transform 1 0 7176 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_72
timestamp 1688980957
transform 1 0 7728 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_76
timestamp 1688980957
transform 1 0 8096 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1688980957
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_124
timestamp 1688980957
transform 1 0 12512 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_130
timestamp 1688980957
transform 1 0 13064 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_134
timestamp 1688980957
transform 1 0 13432 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_138
timestamp 1688980957
transform 1 0 13800 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_146
timestamp 1688980957
transform 1 0 14536 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_158
timestamp 1688980957
transform 1 0 15640 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 1688980957
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_219
timestamp 1688980957
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_229
timestamp 1688980957
transform 1 0 22172 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_233
timestamp 1688980957
transform 1 0 22540 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_245
timestamp 1688980957
transform 1 0 23644 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_253
timestamp 1688980957
transform 1 0 24380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_311
timestamp 1688980957
transform 1 0 29716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_323
timestamp 1688980957
transform 1 0 30820 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_330
timestamp 1688980957
transform 1 0 31464 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_353
timestamp 1688980957
transform 1 0 33580 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_359
timestamp 1688980957
transform 1 0 34132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_365
timestamp 1688980957
transform 1 0 34684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_380
timestamp 1688980957
transform 1 0 36064 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1688980957
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_429
timestamp 1688980957
transform 1 0 40572 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_72
timestamp 1688980957
transform 1 0 7728 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_155
timestamp 1688980957
transform 1 0 15364 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_179
timestamp 1688980957
transform 1 0 17572 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_185
timestamp 1688980957
transform 1 0 18124 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_192
timestamp 1688980957
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_200
timestamp 1688980957
transform 1 0 19504 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_204
timestamp 1688980957
transform 1 0 19872 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_213
timestamp 1688980957
transform 1 0 20700 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_248
timestamp 1688980957
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_261
timestamp 1688980957
transform 1 0 25116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_291
timestamp 1688980957
transform 1 0 27876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_304
timestamp 1688980957
transform 1 0 29072 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_320
timestamp 1688980957
transform 1 0 30544 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_328
timestamp 1688980957
transform 1 0 31280 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_344
timestamp 1688980957
transform 1 0 32752 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_372
timestamp 1688980957
transform 1 0 35328 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_383
timestamp 1688980957
transform 1 0 36340 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_395
timestamp 1688980957
transform 1 0 37444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_407
timestamp 1688980957
transform 1 0 38548 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1688980957
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_89
timestamp 1688980957
transform 1 0 9292 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_101
timestamp 1688980957
transform 1 0 10396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_128
timestamp 1688980957
transform 1 0 12880 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_148
timestamp 1688980957
transform 1 0 14720 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_208
timestamp 1688980957
transform 1 0 20240 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_229
timestamp 1688980957
transform 1 0 22172 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_241
timestamp 1688980957
transform 1 0 23276 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_266
timestamp 1688980957
transform 1 0 25576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_270
timestamp 1688980957
transform 1 0 25944 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_278
timestamp 1688980957
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_296
timestamp 1688980957
transform 1 0 28336 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_326
timestamp 1688980957
transform 1 0 31096 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_354
timestamp 1688980957
transform 1 0 33672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_362
timestamp 1688980957
transform 1 0 34408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_389
timestamp 1688980957
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1688980957
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_429
timestamp 1688980957
transform 1 0 40572 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_9
timestamp 1688980957
transform 1 0 1932 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_21
timestamp 1688980957
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_73
timestamp 1688980957
transform 1 0 7820 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1688980957
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_105
timestamp 1688980957
transform 1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_119
timestamp 1688980957
transform 1 0 12052 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_134
timestamp 1688980957
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_185
timestamp 1688980957
transform 1 0 18124 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_194
timestamp 1688980957
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_237
timestamp 1688980957
transform 1 0 22908 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_241
timestamp 1688980957
transform 1 0 23276 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_248
timestamp 1688980957
transform 1 0 23920 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_273
timestamp 1688980957
transform 1 0 26220 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_285
timestamp 1688980957
transform 1 0 27324 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_297
timestamp 1688980957
transform 1 0 28428 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_305
timestamp 1688980957
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_313
timestamp 1688980957
transform 1 0 29900 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_325
timestamp 1688980957
transform 1 0 31004 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_337
timestamp 1688980957
transform 1 0 32108 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_349
timestamp 1688980957
transform 1 0 33212 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_361
timestamp 1688980957
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_379
timestamp 1688980957
transform 1 0 35972 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_385
timestamp 1688980957
transform 1 0 36524 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_393
timestamp 1688980957
transform 1 0 37260 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_405
timestamp 1688980957
transform 1 0 38364 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_417
timestamp 1688980957
transform 1 0 39468 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_433
timestamp 1688980957
transform 1 0 40940 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_90
timestamp 1688980957
transform 1 0 9384 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_102
timestamp 1688980957
transform 1 0 10488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp 1688980957
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_124
timestamp 1688980957
transform 1 0 12512 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_147
timestamp 1688980957
transform 1 0 14628 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_153
timestamp 1688980957
transform 1 0 15180 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_177
timestamp 1688980957
transform 1 0 17388 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_189
timestamp 1688980957
transform 1 0 18492 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_204
timestamp 1688980957
transform 1 0 19872 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_216
timestamp 1688980957
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1688980957
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_304
timestamp 1688980957
transform 1 0 29072 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_334
timestamp 1688980957
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_343
timestamp 1688980957
transform 1 0 32660 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_356
timestamp 1688980957
transform 1 0 33856 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_363
timestamp 1688980957
transform 1 0 34500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_375
timestamp 1688980957
transform 1 0 35604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_387
timestamp 1688980957
transform 1 0 36708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_406
timestamp 1688980957
transform 1 0 38456 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_418
timestamp 1688980957
transform 1 0 39560 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_430
timestamp 1688980957
transform 1 0 40664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_434
timestamp 1688980957
transform 1 0 41032 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_54
timestamp 1688980957
transform 1 0 6072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_78
timestamp 1688980957
transform 1 0 8280 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_105
timestamp 1688980957
transform 1 0 10764 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_162
timestamp 1688980957
transform 1 0 16008 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_166
timestamp 1688980957
transform 1 0 16376 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_174
timestamp 1688980957
transform 1 0 17112 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_207
timestamp 1688980957
transform 1 0 20148 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_213
timestamp 1688980957
transform 1 0 20700 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_219
timestamp 1688980957
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_223
timestamp 1688980957
transform 1 0 21620 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_247
timestamp 1688980957
transform 1 0 23828 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_257
timestamp 1688980957
transform 1 0 24748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_261
timestamp 1688980957
transform 1 0 25116 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_269
timestamp 1688980957
transform 1 0 25852 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_291
timestamp 1688980957
transform 1 0 27876 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_302
timestamp 1688980957
transform 1 0 28888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_324
timestamp 1688980957
transform 1 0 30912 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_340
timestamp 1688980957
transform 1 0 32384 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_373
timestamp 1688980957
transform 1 0 35420 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_380
timestamp 1688980957
transform 1 0 36064 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_392
timestamp 1688980957
transform 1 0 37168 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_402
timestamp 1688980957
transform 1 0 38088 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_414
timestamp 1688980957
transform 1 0 39192 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1688980957
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_433
timestamp 1688980957
transform 1 0 40940 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_63
timestamp 1688980957
transform 1 0 6900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_74
timestamp 1688980957
transform 1 0 7912 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_82
timestamp 1688980957
transform 1 0 8648 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_98
timestamp 1688980957
transform 1 0 10120 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_106
timestamp 1688980957
transform 1 0 10856 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_122
timestamp 1688980957
transform 1 0 12328 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_157
timestamp 1688980957
transform 1 0 15548 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_177
timestamp 1688980957
transform 1 0 17388 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_189
timestamp 1688980957
transform 1 0 18492 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_195
timestamp 1688980957
transform 1 0 19044 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_278
timestamp 1688980957
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_297
timestamp 1688980957
transform 1 0 28428 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_309
timestamp 1688980957
transform 1 0 29532 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_321
timestamp 1688980957
transform 1 0 30636 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_327
timestamp 1688980957
transform 1 0 31188 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_331
timestamp 1688980957
transform 1 0 31556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1688980957
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_342
timestamp 1688980957
transform 1 0 32568 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_350
timestamp 1688980957
transform 1 0 33304 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_365
timestamp 1688980957
transform 1 0 34684 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_377
timestamp 1688980957
transform 1 0 35788 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_389
timestamp 1688980957
transform 1 0 36892 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_405
timestamp 1688980957
transform 1 0 38364 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_417
timestamp 1688980957
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_429
timestamp 1688980957
transform 1 0 40572 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_37
timestamp 1688980957
transform 1 0 4508 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_48
timestamp 1688980957
transform 1 0 5520 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_56
timestamp 1688980957
transform 1 0 6256 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_68
timestamp 1688980957
transform 1 0 7360 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_78
timestamp 1688980957
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_96
timestamp 1688980957
transform 1 0 9936 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_108
timestamp 1688980957
transform 1 0 11040 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_116
timestamp 1688980957
transform 1 0 11776 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_122
timestamp 1688980957
transform 1 0 12328 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_134
timestamp 1688980957
transform 1 0 13432 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_146
timestamp 1688980957
transform 1 0 14536 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_175
timestamp 1688980957
transform 1 0 17204 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_187
timestamp 1688980957
transform 1 0 18308 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1688980957
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_201
timestamp 1688980957
transform 1 0 19596 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_204
timestamp 1688980957
transform 1 0 19872 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_229
timestamp 1688980957
transform 1 0 22172 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_246
timestamp 1688980957
transform 1 0 23736 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_274
timestamp 1688980957
transform 1 0 26312 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_284
timestamp 1688980957
transform 1 0 27232 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_292
timestamp 1688980957
transform 1 0 27968 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_296
timestamp 1688980957
transform 1 0 28336 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_303
timestamp 1688980957
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1688980957
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_319
timestamp 1688980957
transform 1 0 30452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_334
timestamp 1688980957
transform 1 0 31832 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_342
timestamp 1688980957
transform 1 0 32568 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_347
timestamp 1688980957
transform 1 0 33028 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_355
timestamp 1688980957
transform 1 0 33764 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 1688980957
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_365
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_377
timestamp 1688980957
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_389
timestamp 1688980957
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_401
timestamp 1688980957
transform 1 0 37996 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_408
timestamp 1688980957
transform 1 0 38640 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_421
timestamp 1688980957
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_433
timestamp 1688980957
transform 1 0 40940 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1688980957
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_68
timestamp 1688980957
transform 1 0 7360 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_100
timestamp 1688980957
transform 1 0 10304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_108
timestamp 1688980957
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_122
timestamp 1688980957
transform 1 0 12328 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_126
timestamp 1688980957
transform 1 0 12696 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_130
timestamp 1688980957
transform 1 0 13064 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_142
timestamp 1688980957
transform 1 0 14168 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_154
timestamp 1688980957
transform 1 0 15272 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_158
timestamp 1688980957
transform 1 0 15640 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_212
timestamp 1688980957
transform 1 0 20608 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_237
timestamp 1688980957
transform 1 0 22908 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_248
timestamp 1688980957
transform 1 0 23920 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_260
timestamp 1688980957
transform 1 0 25024 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_276
timestamp 1688980957
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_285
timestamp 1688980957
transform 1 0 27324 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_322
timestamp 1688980957
transform 1 0 30728 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_337
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_341
timestamp 1688980957
transform 1 0 32476 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_360
timestamp 1688980957
transform 1 0 34224 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_372
timestamp 1688980957
transform 1 0 35328 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_384
timestamp 1688980957
transform 1 0 36432 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_400
timestamp 1688980957
transform 1 0 37904 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_412
timestamp 1688980957
transform 1 0 39008 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_424
timestamp 1688980957
transform 1 0 40112 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_432
timestamp 1688980957
transform 1 0 40848 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_47
timestamp 1688980957
transform 1 0 5428 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_59
timestamp 1688980957
transform 1 0 6532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_67
timestamp 1688980957
transform 1 0 7268 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_100
timestamp 1688980957
transform 1 0 10304 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_119
timestamp 1688980957
transform 1 0 12052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_126
timestamp 1688980957
transform 1 0 12696 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1688980957
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_153
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_162
timestamp 1688980957
transform 1 0 16008 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_170
timestamp 1688980957
transform 1 0 16744 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_182
timestamp 1688980957
transform 1 0 17848 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_194
timestamp 1688980957
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_242
timestamp 1688980957
transform 1 0 23368 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_250
timestamp 1688980957
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_265
timestamp 1688980957
transform 1 0 25484 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_273
timestamp 1688980957
transform 1 0 26220 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_282
timestamp 1688980957
transform 1 0 27048 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_294
timestamp 1688980957
transform 1 0 28152 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_302
timestamp 1688980957
transform 1 0 28888 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_317
timestamp 1688980957
transform 1 0 30268 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_327
timestamp 1688980957
transform 1 0 31188 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_339
timestamp 1688980957
transform 1 0 32292 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_345
timestamp 1688980957
transform 1 0 32844 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_357
timestamp 1688980957
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 1688980957
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_365
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_390
timestamp 1688980957
transform 1 0 36984 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_394
timestamp 1688980957
transform 1 0 37352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_416
timestamp 1688980957
transform 1 0 39376 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_421
timestamp 1688980957
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_433
timestamp 1688980957
transform 1 0 40940 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_9
timestamp 1688980957
transform 1 0 1932 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_17
timestamp 1688980957
transform 1 0 2668 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_33
timestamp 1688980957
transform 1 0 4140 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_42
timestamp 1688980957
transform 1 0 4968 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 1688980957
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_63
timestamp 1688980957
transform 1 0 6900 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_78
timestamp 1688980957
transform 1 0 8280 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_90
timestamp 1688980957
transform 1 0 9384 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_102
timestamp 1688980957
transform 1 0 10488 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_125
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_131
timestamp 1688980957
transform 1 0 13156 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_147
timestamp 1688980957
transform 1 0 14628 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_159
timestamp 1688980957
transform 1 0 15732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1688980957
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_181
timestamp 1688980957
transform 1 0 17756 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_187
timestamp 1688980957
transform 1 0 18308 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_211
timestamp 1688980957
transform 1 0 20516 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_216
timestamp 1688980957
transform 1 0 20976 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_237
timestamp 1688980957
transform 1 0 22908 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_252
timestamp 1688980957
transform 1 0 24288 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_264
timestamp 1688980957
transform 1 0 25392 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1688980957
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_287
timestamp 1688980957
transform 1 0 27508 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_299
timestamp 1688980957
transform 1 0 28612 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_312
timestamp 1688980957
transform 1 0 29808 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 1688980957
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 1688980957
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_349
timestamp 1688980957
transform 1 0 33212 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_363
timestamp 1688980957
transform 1 0 34500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_373
timestamp 1688980957
transform 1 0 35420 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_383
timestamp 1688980957
transform 1 0 36340 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_391
timestamp 1688980957
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_393
timestamp 1688980957
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_405
timestamp 1688980957
transform 1 0 38364 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_413
timestamp 1688980957
transform 1 0 39100 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_427
timestamp 1688980957
transform 1 0 40388 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_68
timestamp 1688980957
transform 1 0 7360 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_80
timestamp 1688980957
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_90
timestamp 1688980957
transform 1 0 9384 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_98
timestamp 1688980957
transform 1 0 10120 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_105
timestamp 1688980957
transform 1 0 10764 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_117
timestamp 1688980957
transform 1 0 11868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_155
timestamp 1688980957
transform 1 0 15364 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_167
timestamp 1688980957
transform 1 0 16468 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_175
timestamp 1688980957
transform 1 0 17204 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_181
timestamp 1688980957
transform 1 0 17756 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_189
timestamp 1688980957
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_207
timestamp 1688980957
transform 1 0 20148 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_230
timestamp 1688980957
transform 1 0 22264 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_238
timestamp 1688980957
transform 1 0 23000 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_250
timestamp 1688980957
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_260
timestamp 1688980957
transform 1 0 25024 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_292
timestamp 1688980957
transform 1 0 27968 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_304
timestamp 1688980957
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_340
timestamp 1688980957
transform 1 0 32384 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_354
timestamp 1688980957
transform 1 0 33672 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_361
timestamp 1688980957
transform 1 0 34316 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 1688980957
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 1688980957
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_401
timestamp 1688980957
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_413
timestamp 1688980957
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_419
timestamp 1688980957
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_421
timestamp 1688980957
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_433
timestamp 1688980957
transform 1 0 40940 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1688980957
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_74
timestamp 1688980957
transform 1 0 7912 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_78
timestamp 1688980957
transform 1 0 8280 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_87
timestamp 1688980957
transform 1 0 9108 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_130
timestamp 1688980957
transform 1 0 13064 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_138
timestamp 1688980957
transform 1 0 13800 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_148
timestamp 1688980957
transform 1 0 14720 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_164
timestamp 1688980957
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_174
timestamp 1688980957
transform 1 0 17112 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_183
timestamp 1688980957
transform 1 0 17940 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_194
timestamp 1688980957
transform 1 0 18952 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_206
timestamp 1688980957
transform 1 0 20056 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_218
timestamp 1688980957
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_232
timestamp 1688980957
transform 1 0 22448 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_244
timestamp 1688980957
transform 1 0 23552 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_260
timestamp 1688980957
transform 1 0 25024 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_268
timestamp 1688980957
transform 1 0 25760 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_277
timestamp 1688980957
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_293
timestamp 1688980957
transform 1 0 28060 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_307
timestamp 1688980957
transform 1 0 29348 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_318
timestamp 1688980957
transform 1 0 30360 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_330
timestamp 1688980957
transform 1 0 31464 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_337
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_351
timestamp 1688980957
transform 1 0 33396 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_368
timestamp 1688980957
transform 1 0 34960 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_380
timestamp 1688980957
transform 1 0 36064 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_388
timestamp 1688980957
transform 1 0 36800 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_393
timestamp 1688980957
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_405
timestamp 1688980957
transform 1 0 38364 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_409
timestamp 1688980957
transform 1 0 38732 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_417
timestamp 1688980957
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_429
timestamp 1688980957
transform 1 0 40572 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_11
timestamp 1688980957
transform 1 0 2116 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_37
timestamp 1688980957
transform 1 0 4508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_46
timestamp 1688980957
transform 1 0 5336 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_50
timestamp 1688980957
transform 1 0 5704 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_58
timestamp 1688980957
transform 1 0 6440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_62
timestamp 1688980957
transform 1 0 6808 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_72
timestamp 1688980957
transform 1 0 7728 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_94
timestamp 1688980957
transform 1 0 9752 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_112
timestamp 1688980957
transform 1 0 11408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_132
timestamp 1688980957
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_147
timestamp 1688980957
transform 1 0 14628 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_176
timestamp 1688980957
transform 1 0 17296 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_187
timestamp 1688980957
transform 1 0 18308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_209
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_213
timestamp 1688980957
transform 1 0 20700 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_238
timestamp 1688980957
transform 1 0 23000 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_250
timestamp 1688980957
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1688980957
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_277
timestamp 1688980957
transform 1 0 26588 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_286
timestamp 1688980957
transform 1 0 27416 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_298
timestamp 1688980957
transform 1 0 28520 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_306
timestamp 1688980957
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_315
timestamp 1688980957
transform 1 0 30084 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 1688980957
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_333
timestamp 1688980957
transform 1 0 31740 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_337
timestamp 1688980957
transform 1 0 32108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_344
timestamp 1688980957
transform 1 0 32752 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_356
timestamp 1688980957
transform 1 0 33856 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_390
timestamp 1688980957
transform 1 0 36984 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_400
timestamp 1688980957
transform 1 0 37904 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_408
timestamp 1688980957
transform 1 0 38640 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_416
timestamp 1688980957
transform 1 0 39376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_426
timestamp 1688980957
transform 1 0 40296 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_434
timestamp 1688980957
transform 1 0 41032 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_24
timestamp 1688980957
transform 1 0 3312 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp 1688980957
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_64
timestamp 1688980957
transform 1 0 6992 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_85
timestamp 1688980957
transform 1 0 8924 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_98
timestamp 1688980957
transform 1 0 10120 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1688980957
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_130
timestamp 1688980957
transform 1 0 13064 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_142
timestamp 1688980957
transform 1 0 14168 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_154
timestamp 1688980957
transform 1 0 15272 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_166
timestamp 1688980957
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_205
timestamp 1688980957
transform 1 0 19964 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_218
timestamp 1688980957
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1688980957
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1688980957
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_261
timestamp 1688980957
transform 1 0 25116 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_270
timestamp 1688980957
transform 1 0 25944 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_297
timestamp 1688980957
transform 1 0 28428 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_305
timestamp 1688980957
transform 1 0 29164 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_318
timestamp 1688980957
transform 1 0 30360 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_324
timestamp 1688980957
transform 1 0 30912 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_332
timestamp 1688980957
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_343
timestamp 1688980957
transform 1 0 32660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_355
timestamp 1688980957
transform 1 0 33764 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_359
timestamp 1688980957
transform 1 0 34132 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_366
timestamp 1688980957
transform 1 0 34776 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_374
timestamp 1688980957
transform 1 0 35512 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_383
timestamp 1688980957
transform 1 0 36340 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 1688980957
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_400
timestamp 1688980957
transform 1 0 37904 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_412
timestamp 1688980957
transform 1 0 39008 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_424
timestamp 1688980957
transform 1 0 40112 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_432
timestamp 1688980957
transform 1 0 40848 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_37
timestamp 1688980957
transform 1 0 4508 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_49
timestamp 1688980957
transform 1 0 5612 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_61
timestamp 1688980957
transform 1 0 6716 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_72
timestamp 1688980957
transform 1 0 7728 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_109
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_115
timestamp 1688980957
transform 1 0 11684 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_119
timestamp 1688980957
transform 1 0 12052 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_131
timestamp 1688980957
transform 1 0 13156 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1688980957
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_156
timestamp 1688980957
transform 1 0 15456 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_168
timestamp 1688980957
transform 1 0 16560 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_184
timestamp 1688980957
transform 1 0 18032 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_212
timestamp 1688980957
transform 1 0 20608 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_228
timestamp 1688980957
transform 1 0 22080 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_236
timestamp 1688980957
transform 1 0 22816 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_241
timestamp 1688980957
transform 1 0 23276 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_249
timestamp 1688980957
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_257
timestamp 1688980957
transform 1 0 24748 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_290
timestamp 1688980957
transform 1 0 27784 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_298
timestamp 1688980957
transform 1 0 28520 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_306
timestamp 1688980957
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_336
timestamp 1688980957
transform 1 0 32016 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_348
timestamp 1688980957
transform 1 0 33120 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_359
timestamp 1688980957
transform 1 0 34132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 1688980957
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_373
timestamp 1688980957
transform 1 0 35420 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_385
timestamp 1688980957
transform 1 0 36524 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_393
timestamp 1688980957
transform 1 0 37260 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_405
timestamp 1688980957
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_413
timestamp 1688980957
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_419
timestamp 1688980957
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_427
timestamp 1688980957
transform 1 0 40388 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_25
timestamp 1688980957
transform 1 0 3404 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_37
timestamp 1688980957
transform 1 0 4508 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_49
timestamp 1688980957
transform 1 0 5612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_83
timestamp 1688980957
transform 1 0 8740 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_91
timestamp 1688980957
transform 1 0 9476 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_133
timestamp 1688980957
transform 1 0 13340 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_159
timestamp 1688980957
transform 1 0 15732 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_190
timestamp 1688980957
transform 1 0 18584 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_206
timestamp 1688980957
transform 1 0 20056 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_214
timestamp 1688980957
transform 1 0 20792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_220
timestamp 1688980957
transform 1 0 21344 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_237
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_257
timestamp 1688980957
transform 1 0 24748 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_269
timestamp 1688980957
transform 1 0 25852 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_277
timestamp 1688980957
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_289
timestamp 1688980957
transform 1 0 27692 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_298
timestamp 1688980957
transform 1 0 28520 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_313
timestamp 1688980957
transform 1 0 29900 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_325
timestamp 1688980957
transform 1 0 31004 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_333
timestamp 1688980957
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_345
timestamp 1688980957
transform 1 0 32844 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_366
timestamp 1688980957
transform 1 0 34776 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_378
timestamp 1688980957
transform 1 0 35880 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_390
timestamp 1688980957
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_393
timestamp 1688980957
transform 1 0 37260 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_401
timestamp 1688980957
transform 1 0 37996 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_411
timestamp 1688980957
transform 1 0 38916 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_423
timestamp 1688980957
transform 1 0 40020 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_9
timestamp 1688980957
transform 1 0 1932 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_13
timestamp 1688980957
transform 1 0 2300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_26
timestamp 1688980957
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_34
timestamp 1688980957
transform 1 0 4232 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_58
timestamp 1688980957
transform 1 0 6440 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_70
timestamp 1688980957
transform 1 0 7544 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_79
timestamp 1688980957
transform 1 0 8372 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_114
timestamp 1688980957
transform 1 0 11592 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_126
timestamp 1688980957
transform 1 0 12696 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_130
timestamp 1688980957
transform 1 0 13064 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 1688980957
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1688980957
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_165
timestamp 1688980957
transform 1 0 16284 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_191
timestamp 1688980957
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1688980957
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_209
timestamp 1688980957
transform 1 0 20332 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_217
timestamp 1688980957
transform 1 0 21068 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_230
timestamp 1688980957
transform 1 0 22264 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_242
timestamp 1688980957
transform 1 0 23368 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_282
timestamp 1688980957
transform 1 0 27048 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_294
timestamp 1688980957
transform 1 0 28152 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_306
timestamp 1688980957
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_309
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 1688980957
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_333
timestamp 1688980957
transform 1 0 31740 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_346
timestamp 1688980957
transform 1 0 32936 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_358
timestamp 1688980957
transform 1 0 34040 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_365
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_381
timestamp 1688980957
transform 1 0 36156 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_401
timestamp 1688980957
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_413
timestamp 1688980957
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_419
timestamp 1688980957
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_427
timestamp 1688980957
transform 1 0 40388 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_15
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_23
timestamp 1688980957
transform 1 0 3220 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_46
timestamp 1688980957
transform 1 0 5336 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_65
timestamp 1688980957
transform 1 0 7084 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_73
timestamp 1688980957
transform 1 0 7820 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_103
timestamp 1688980957
transform 1 0 10580 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1688980957
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_121
timestamp 1688980957
transform 1 0 12236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_136
timestamp 1688980957
transform 1 0 13616 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_140
timestamp 1688980957
transform 1 0 13984 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_150
timestamp 1688980957
transform 1 0 14904 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_166
timestamp 1688980957
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_176
timestamp 1688980957
transform 1 0 17296 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_182
timestamp 1688980957
transform 1 0 17848 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_200
timestamp 1688980957
transform 1 0 19504 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_212
timestamp 1688980957
transform 1 0 20608 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_237
timestamp 1688980957
transform 1 0 22908 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_243
timestamp 1688980957
transform 1 0 23460 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_252
timestamp 1688980957
transform 1 0 24288 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_264
timestamp 1688980957
transform 1 0 25392 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 1688980957
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1688980957
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1688980957
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1688980957
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_317
timestamp 1688980957
transform 1 0 30268 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_325
timestamp 1688980957
transform 1 0 31004 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_332
timestamp 1688980957
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 1688980957
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_361
timestamp 1688980957
transform 1 0 34316 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_369
timestamp 1688980957
transform 1 0 35052 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_378
timestamp 1688980957
transform 1 0 35880 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_390
timestamp 1688980957
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_399
timestamp 1688980957
transform 1 0 37812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_411
timestamp 1688980957
transform 1 0 38916 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_420
timestamp 1688980957
transform 1 0 39744 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_432
timestamp 1688980957
transform 1 0 40848 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_55
timestamp 1688980957
transform 1 0 6164 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_76
timestamp 1688980957
transform 1 0 8096 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_94
timestamp 1688980957
transform 1 0 9752 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_100
timestamp 1688980957
transform 1 0 10304 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1688980957
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_133
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_161
timestamp 1688980957
transform 1 0 15916 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_173
timestamp 1688980957
transform 1 0 17020 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_185
timestamp 1688980957
transform 1 0 18124 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_193
timestamp 1688980957
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_208
timestamp 1688980957
transform 1 0 20240 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_216
timestamp 1688980957
transform 1 0 20976 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_230
timestamp 1688980957
transform 1 0 22264 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_238
timestamp 1688980957
transform 1 0 23000 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_246
timestamp 1688980957
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_259
timestamp 1688980957
transform 1 0 24932 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_276
timestamp 1688980957
transform 1 0 26496 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_288
timestamp 1688980957
transform 1 0 27600 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_302
timestamp 1688980957
transform 1 0 28888 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_322
timestamp 1688980957
transform 1 0 30728 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_334
timestamp 1688980957
transform 1 0 31832 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_344
timestamp 1688980957
transform 1 0 32752 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_350
timestamp 1688980957
transform 1 0 33304 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_357
timestamp 1688980957
transform 1 0 33948 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_365
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_375
timestamp 1688980957
transform 1 0 35604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_387
timestamp 1688980957
transform 1 0 36708 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_398
timestamp 1688980957
transform 1 0 37720 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_410
timestamp 1688980957
transform 1 0 38824 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_418
timestamp 1688980957
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_427
timestamp 1688980957
transform 1 0 40388 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_7
timestamp 1688980957
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_11
timestamp 1688980957
transform 1 0 2116 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_35
timestamp 1688980957
transform 1 0 4324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_47
timestamp 1688980957
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_64
timestamp 1688980957
transform 1 0 6992 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_74
timestamp 1688980957
transform 1 0 7912 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_95
timestamp 1688980957
transform 1 0 9844 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_101
timestamp 1688980957
transform 1 0 10396 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_105
timestamp 1688980957
transform 1 0 10764 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_110
timestamp 1688980957
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_130
timestamp 1688980957
transform 1 0 13064 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_151
timestamp 1688980957
transform 1 0 14996 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_159
timestamp 1688980957
transform 1 0 15732 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 1688980957
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_178
timestamp 1688980957
transform 1 0 17480 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_202
timestamp 1688980957
transform 1 0 19688 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_217
timestamp 1688980957
transform 1 0 21068 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_231
timestamp 1688980957
transform 1 0 22356 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_257
timestamp 1688980957
transform 1 0 24748 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_269
timestamp 1688980957
transform 1 0 25852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_273
timestamp 1688980957
transform 1 0 26220 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_318
timestamp 1688980957
transform 1 0 30360 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_330
timestamp 1688980957
transform 1 0 31464 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_364
timestamp 1688980957
transform 1 0 34592 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_376
timestamp 1688980957
transform 1 0 35696 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_388
timestamp 1688980957
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_393
timestamp 1688980957
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_405
timestamp 1688980957
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_417
timestamp 1688980957
transform 1 0 39468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_429
timestamp 1688980957
transform 1 0 40572 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_23
timestamp 1688980957
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_33
timestamp 1688980957
transform 1 0 4140 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_54
timestamp 1688980957
transform 1 0 6072 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_66
timestamp 1688980957
transform 1 0 7176 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_72
timestamp 1688980957
transform 1 0 7728 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_93
timestamp 1688980957
transform 1 0 9660 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_144
timestamp 1688980957
transform 1 0 14352 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_152
timestamp 1688980957
transform 1 0 15088 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_178
timestamp 1688980957
transform 1 0 17480 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_192
timestamp 1688980957
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_209
timestamp 1688980957
transform 1 0 20332 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_222
timestamp 1688980957
transform 1 0 21528 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_234
timestamp 1688980957
transform 1 0 22632 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_246
timestamp 1688980957
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_261
timestamp 1688980957
transform 1 0 25116 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_273
timestamp 1688980957
transform 1 0 26220 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_285
timestamp 1688980957
transform 1 0 27324 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_305
timestamp 1688980957
transform 1 0 29164 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_321
timestamp 1688980957
transform 1 0 30636 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_333
timestamp 1688980957
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_345
timestamp 1688980957
transform 1 0 32844 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_353
timestamp 1688980957
transform 1 0 33580 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_362
timestamp 1688980957
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_365
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_379
timestamp 1688980957
transform 1 0 35972 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_391
timestamp 1688980957
transform 1 0 37076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_401
timestamp 1688980957
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_407
timestamp 1688980957
transform 1 0 38548 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_414
timestamp 1688980957
transform 1 0 39192 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_421
timestamp 1688980957
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_433
timestamp 1688980957
transform 1 0 40940 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_32
timestamp 1688980957
transform 1 0 4048 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_38
timestamp 1688980957
transform 1 0 4600 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1688980957
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1688980957
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_68
timestamp 1688980957
transform 1 0 7360 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_80
timestamp 1688980957
transform 1 0 8464 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_92
timestamp 1688980957
transform 1 0 9568 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_104
timestamp 1688980957
transform 1 0 10672 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1688980957
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_137
timestamp 1688980957
transform 1 0 13708 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_150
timestamp 1688980957
transform 1 0 14904 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_158
timestamp 1688980957
transform 1 0 15640 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_176
timestamp 1688980957
transform 1 0 17296 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_192
timestamp 1688980957
transform 1 0 18768 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_203
timestamp 1688980957
transform 1 0 19780 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_215
timestamp 1688980957
transform 1 0 20884 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1688980957
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1688980957
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1688980957
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1688980957
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 1688980957
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1688980957
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1688980957
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_305
timestamp 1688980957
transform 1 0 29164 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_309
timestamp 1688980957
transform 1 0 29532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_322
timestamp 1688980957
transform 1 0 30728 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_328
timestamp 1688980957
transform 1 0 31280 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_332
timestamp 1688980957
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_349
timestamp 1688980957
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_361
timestamp 1688980957
transform 1 0 34316 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_375
timestamp 1688980957
transform 1 0 35604 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_383
timestamp 1688980957
transform 1 0 36340 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_390
timestamp 1688980957
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_393
timestamp 1688980957
transform 1 0 37260 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_403
timestamp 1688980957
transform 1 0 38180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_415
timestamp 1688980957
transform 1 0 39284 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_433
timestamp 1688980957
transform 1 0 40940 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_46
timestamp 1688980957
transform 1 0 5336 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_82
timestamp 1688980957
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_127
timestamp 1688980957
transform 1 0 12788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1688980957
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_165
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1688980957
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_193
timestamp 1688980957
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_209
timestamp 1688980957
transform 1 0 20332 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_228
timestamp 1688980957
transform 1 0 22080 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_240
timestamp 1688980957
transform 1 0 23184 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_249
timestamp 1688980957
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_279
timestamp 1688980957
transform 1 0 26772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_291
timestamp 1688980957
transform 1 0 27876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_303
timestamp 1688980957
transform 1 0 28980 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1688980957
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_321
timestamp 1688980957
transform 1 0 30636 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_327
timestamp 1688980957
transform 1 0 31188 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_336
timestamp 1688980957
transform 1 0 32016 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_344
timestamp 1688980957
transform 1 0 32752 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_359
timestamp 1688980957
transform 1 0 34132 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 1688980957
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_365
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_380
timestamp 1688980957
transform 1 0 36064 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_392
timestamp 1688980957
transform 1 0 37168 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_404
timestamp 1688980957
transform 1 0 38272 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_412
timestamp 1688980957
transform 1 0 39008 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_426
timestamp 1688980957
transform 1 0 40296 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_434
timestamp 1688980957
transform 1 0 41032 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_7
timestamp 1688980957
transform 1 0 1748 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_11
timestamp 1688980957
transform 1 0 2116 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_49
timestamp 1688980957
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_72
timestamp 1688980957
transform 1 0 7728 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_108
timestamp 1688980957
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_119
timestamp 1688980957
transform 1 0 12052 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_129
timestamp 1688980957
transform 1 0 12972 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_141
timestamp 1688980957
transform 1 0 14076 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_145
timestamp 1688980957
transform 1 0 14444 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_181
timestamp 1688980957
transform 1 0 17756 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_191
timestamp 1688980957
transform 1 0 18676 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_197
timestamp 1688980957
transform 1 0 19228 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_209
timestamp 1688980957
transform 1 0 20332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_221
timestamp 1688980957
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_237
timestamp 1688980957
transform 1 0 22908 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_247
timestamp 1688980957
transform 1 0 23828 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_270
timestamp 1688980957
transform 1 0 25944 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_290
timestamp 1688980957
transform 1 0 27784 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_297
timestamp 1688980957
transform 1 0 28428 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_303
timestamp 1688980957
transform 1 0 28980 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_315
timestamp 1688980957
transform 1 0 30084 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_330
timestamp 1688980957
transform 1 0 31464 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_349
timestamp 1688980957
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_361
timestamp 1688980957
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_373
timestamp 1688980957
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_385
timestamp 1688980957
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_391
timestamp 1688980957
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_393
timestamp 1688980957
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_405
timestamp 1688980957
transform 1 0 38364 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_413
timestamp 1688980957
transform 1 0 39100 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_422
timestamp 1688980957
transform 1 0 39928 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_434
timestamp 1688980957
transform 1 0 41032 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_23
timestamp 1688980957
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_32
timestamp 1688980957
transform 1 0 4048 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_50
timestamp 1688980957
transform 1 0 5704 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_62
timestamp 1688980957
transform 1 0 6808 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_70
timestamp 1688980957
transform 1 0 7544 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_134
timestamp 1688980957
transform 1 0 13432 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_138
timestamp 1688980957
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_150
timestamp 1688980957
transform 1 0 14904 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_158
timestamp 1688980957
transform 1 0 15640 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_170
timestamp 1688980957
transform 1 0 16744 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_214
timestamp 1688980957
transform 1 0 20792 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_226
timestamp 1688980957
transform 1 0 21896 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_238
timestamp 1688980957
transform 1 0 23000 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_248
timestamp 1688980957
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_267
timestamp 1688980957
transform 1 0 25668 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_279
timestamp 1688980957
transform 1 0 26772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_285
timestamp 1688980957
transform 1 0 27324 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_291
timestamp 1688980957
transform 1 0 27876 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_318
timestamp 1688980957
transform 1 0 30360 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_326
timestamp 1688980957
transform 1 0 31096 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_336
timestamp 1688980957
transform 1 0 32016 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 1688980957
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_372
timestamp 1688980957
transform 1 0 35328 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_384
timestamp 1688980957
transform 1 0 36432 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_396
timestamp 1688980957
transform 1 0 37536 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_408
timestamp 1688980957
transform 1 0 38640 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_421
timestamp 1688980957
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_433
timestamp 1688980957
transform 1 0 40940 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_36
timestamp 1688980957
transform 1 0 4416 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_44
timestamp 1688980957
transform 1 0 5152 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_52
timestamp 1688980957
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_78
timestamp 1688980957
transform 1 0 8280 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_97
timestamp 1688980957
transform 1 0 10028 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_127
timestamp 1688980957
transform 1 0 12788 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_150
timestamp 1688980957
transform 1 0 14904 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_178
timestamp 1688980957
transform 1 0 17480 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_190
timestamp 1688980957
transform 1 0 18584 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_202
timestamp 1688980957
transform 1 0 19688 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_208
timestamp 1688980957
transform 1 0 20240 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_219
timestamp 1688980957
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1688980957
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_233
timestamp 1688980957
transform 1 0 22540 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_242
timestamp 1688980957
transform 1 0 23368 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_254
timestamp 1688980957
transform 1 0 24472 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_262
timestamp 1688980957
transform 1 0 25208 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_271
timestamp 1688980957
transform 1 0 26036 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1688980957
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_285
timestamp 1688980957
transform 1 0 27324 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_291
timestamp 1688980957
transform 1 0 27876 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_299
timestamp 1688980957
transform 1 0 28612 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_311
timestamp 1688980957
transform 1 0 29716 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_323
timestamp 1688980957
transform 1 0 30820 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_334
timestamp 1688980957
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 1688980957
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_361
timestamp 1688980957
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_373
timestamp 1688980957
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_385
timestamp 1688980957
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 1688980957
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_399
timestamp 1688980957
transform 1 0 37812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_411
timestamp 1688980957
transform 1 0 38916 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_415
timestamp 1688980957
transform 1 0 39284 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_421
timestamp 1688980957
transform 1 0 39836 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_427
timestamp 1688980957
transform 1 0 40388 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_23
timestamp 1688980957
transform 1 0 3220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_38
timestamp 1688980957
transform 1 0 4600 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_44
timestamp 1688980957
transform 1 0 5152 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_72
timestamp 1688980957
transform 1 0 7728 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 1688980957
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_109
timestamp 1688980957
transform 1 0 11132 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_119
timestamp 1688980957
transform 1 0 12052 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_131
timestamp 1688980957
transform 1 0 13156 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 1688980957
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_189
timestamp 1688980957
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1688980957
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_203
timestamp 1688980957
transform 1 0 19780 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_215
timestamp 1688980957
transform 1 0 20884 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_224
timestamp 1688980957
transform 1 0 21712 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_244
timestamp 1688980957
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 1688980957
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_277
timestamp 1688980957
transform 1 0 26588 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_285
timestamp 1688980957
transform 1 0 27324 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_297
timestamp 1688980957
transform 1 0 28428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_305
timestamp 1688980957
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_317
timestamp 1688980957
transform 1 0 30268 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_334
timestamp 1688980957
transform 1 0 31832 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_340
timestamp 1688980957
transform 1 0 32384 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_348
timestamp 1688980957
transform 1 0 33120 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_360
timestamp 1688980957
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_365
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_382
timestamp 1688980957
transform 1 0 36248 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_402
timestamp 1688980957
transform 1 0 38088 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_408
timestamp 1688980957
transform 1 0 38640 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_415
timestamp 1688980957
transform 1 0 39284 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_419
timestamp 1688980957
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_432
timestamp 1688980957
transform 1 0 40848 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_7
timestamp 1688980957
transform 1 0 1748 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_11
timestamp 1688980957
transform 1 0 2116 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_37
timestamp 1688980957
transform 1 0 4508 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_49
timestamp 1688980957
transform 1 0 5612 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_60
timestamp 1688980957
transform 1 0 6624 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_70
timestamp 1688980957
transform 1 0 7544 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_82
timestamp 1688980957
transform 1 0 8648 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_92
timestamp 1688980957
transform 1 0 9568 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_106
timestamp 1688980957
transform 1 0 10856 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_125
timestamp 1688980957
transform 1 0 12604 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_133
timestamp 1688980957
transform 1 0 13340 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_138
timestamp 1688980957
transform 1 0 13800 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_150
timestamp 1688980957
transform 1 0 14904 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_164
timestamp 1688980957
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_183
timestamp 1688980957
transform 1 0 17940 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_187
timestamp 1688980957
transform 1 0 18308 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_200
timestamp 1688980957
transform 1 0 19504 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_206
timestamp 1688980957
transform 1 0 20056 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_220
timestamp 1688980957
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_233
timestamp 1688980957
transform 1 0 22540 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_245
timestamp 1688980957
transform 1 0 23644 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_254
timestamp 1688980957
transform 1 0 24472 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_266
timestamp 1688980957
transform 1 0 25576 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_274
timestamp 1688980957
transform 1 0 26312 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_306
timestamp 1688980957
transform 1 0 29256 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_318
timestamp 1688980957
transform 1 0 30360 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_330
timestamp 1688980957
transform 1 0 31464 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_349
timestamp 1688980957
transform 1 0 33212 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_359
timestamp 1688980957
transform 1 0 34132 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_367
timestamp 1688980957
transform 1 0 34868 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_377
timestamp 1688980957
transform 1 0 35788 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_389
timestamp 1688980957
transform 1 0 36892 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_399
timestamp 1688980957
transform 1 0 37812 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_416
timestamp 1688980957
transform 1 0 39376 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_428
timestamp 1688980957
transform 1 0 40480 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_24
timestamp 1688980957
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_55
timestamp 1688980957
transform 1 0 6164 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_63
timestamp 1688980957
transform 1 0 6900 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_69
timestamp 1688980957
transform 1 0 7452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_81
timestamp 1688980957
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_114
timestamp 1688980957
transform 1 0 11592 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_149
timestamp 1688980957
transform 1 0 14812 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_161
timestamp 1688980957
transform 1 0 15916 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_173
timestamp 1688980957
transform 1 0 17020 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_211
timestamp 1688980957
transform 1 0 20516 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_225
timestamp 1688980957
transform 1 0 21804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_241
timestamp 1688980957
transform 1 0 23276 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_245
timestamp 1688980957
transform 1 0 23644 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1688980957
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_260
timestamp 1688980957
transform 1 0 25024 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_302
timestamp 1688980957
transform 1 0 28888 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_318
timestamp 1688980957
transform 1 0 30360 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_326
timestamp 1688980957
transform 1 0 31096 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_335
timestamp 1688980957
transform 1 0 31924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_347
timestamp 1688980957
transform 1 0 33028 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_353
timestamp 1688980957
transform 1 0 33580 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_362
timestamp 1688980957
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_365
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_377
timestamp 1688980957
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_389
timestamp 1688980957
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_401
timestamp 1688980957
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_413
timestamp 1688980957
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_419
timestamp 1688980957
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_421
timestamp 1688980957
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_433
timestamp 1688980957
transform 1 0 40940 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_7
timestamp 1688980957
transform 1 0 1748 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_11
timestamp 1688980957
transform 1 0 2116 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_24
timestamp 1688980957
transform 1 0 3312 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_32
timestamp 1688980957
transform 1 0 4048 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_53
timestamp 1688980957
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_88
timestamp 1688980957
transform 1 0 9200 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_103
timestamp 1688980957
transform 1 0 10580 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_131
timestamp 1688980957
transform 1 0 13156 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_135
timestamp 1688980957
transform 1 0 13524 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_142
timestamp 1688980957
transform 1 0 14168 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_151
timestamp 1688980957
transform 1 0 14996 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_179
timestamp 1688980957
transform 1 0 17572 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 1688980957
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 1688980957
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 1688980957
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_235
timestamp 1688980957
transform 1 0 22724 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_243
timestamp 1688980957
transform 1 0 23460 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_263
timestamp 1688980957
transform 1 0 25300 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_275
timestamp 1688980957
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1688980957
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_298
timestamp 1688980957
transform 1 0 28520 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_306
timestamp 1688980957
transform 1 0 29256 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_332
timestamp 1688980957
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_337
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_344
timestamp 1688980957
transform 1 0 32752 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_356
timestamp 1688980957
transform 1 0 33856 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_364
timestamp 1688980957
transform 1 0 34592 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_368
timestamp 1688980957
transform 1 0 34960 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_384
timestamp 1688980957
transform 1 0 36432 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_393
timestamp 1688980957
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_405
timestamp 1688980957
transform 1 0 38364 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_414
timestamp 1688980957
transform 1 0 39192 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_422
timestamp 1688980957
transform 1 0 39928 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_434
timestamp 1688980957
transform 1 0 41032 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_23
timestamp 1688980957
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_50
timestamp 1688980957
transform 1 0 5704 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_62
timestamp 1688980957
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_73
timestamp 1688980957
transform 1 0 7820 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_81
timestamp 1688980957
transform 1 0 8556 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_93
timestamp 1688980957
transform 1 0 9660 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_120
timestamp 1688980957
transform 1 0 12144 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_132
timestamp 1688980957
transform 1 0 13248 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_150
timestamp 1688980957
transform 1 0 14904 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_165
timestamp 1688980957
transform 1 0 16284 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_173
timestamp 1688980957
transform 1 0 17020 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_188
timestamp 1688980957
transform 1 0 18400 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_209
timestamp 1688980957
transform 1 0 20332 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_239
timestamp 1688980957
transform 1 0 23092 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_245
timestamp 1688980957
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1688980957
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_265
timestamp 1688980957
transform 1 0 25484 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_288
timestamp 1688980957
transform 1 0 27600 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_298
timestamp 1688980957
transform 1 0 28520 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_306
timestamp 1688980957
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_321
timestamp 1688980957
transform 1 0 30636 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_329
timestamp 1688980957
transform 1 0 31372 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_336
timestamp 1688980957
transform 1 0 32016 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_347
timestamp 1688980957
transform 1 0 33028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_359
timestamp 1688980957
transform 1 0 34132 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 1688980957
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_365
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_377
timestamp 1688980957
transform 1 0 35788 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_387
timestamp 1688980957
transform 1 0 36708 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_399
timestamp 1688980957
transform 1 0 37812 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_407
timestamp 1688980957
transform 1 0 38548 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_415
timestamp 1688980957
transform 1 0 39284 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_419
timestamp 1688980957
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_421
timestamp 1688980957
transform 1 0 39836 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_427
timestamp 1688980957
transform 1 0 40388 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_11
timestamp 1688980957
transform 1 0 2116 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_34
timestamp 1688980957
transform 1 0 4232 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_46
timestamp 1688980957
transform 1 0 5336 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_54
timestamp 1688980957
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_65
timestamp 1688980957
transform 1 0 7084 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_73
timestamp 1688980957
transform 1 0 7820 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_85
timestamp 1688980957
transform 1 0 8924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_94
timestamp 1688980957
transform 1 0 9752 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_108
timestamp 1688980957
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_131
timestamp 1688980957
transform 1 0 13156 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_139
timestamp 1688980957
transform 1 0 13892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_164
timestamp 1688980957
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_176
timestamp 1688980957
transform 1 0 17296 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_184
timestamp 1688980957
transform 1 0 18032 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_191
timestamp 1688980957
transform 1 0 18676 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_203
timestamp 1688980957
transform 1 0 19780 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_222
timestamp 1688980957
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_233
timestamp 1688980957
transform 1 0 22540 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_245
timestamp 1688980957
transform 1 0 23644 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_253
timestamp 1688980957
transform 1 0 24380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_263
timestamp 1688980957
transform 1 0 25300 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_278
timestamp 1688980957
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_293
timestamp 1688980957
transform 1 0 28060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_297
timestamp 1688980957
transform 1 0 28428 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_305
timestamp 1688980957
transform 1 0 29164 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_315
timestamp 1688980957
transform 1 0 30084 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_323
timestamp 1688980957
transform 1 0 30820 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_331
timestamp 1688980957
transform 1 0 31556 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 1688980957
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_337
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_345
timestamp 1688980957
transform 1 0 32844 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_359
timestamp 1688980957
transform 1 0 34132 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_367
timestamp 1688980957
transform 1 0 34868 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_373
timestamp 1688980957
transform 1 0 35420 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_387
timestamp 1688980957
transform 1 0 36708 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_401
timestamp 1688980957
transform 1 0 37996 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_421
timestamp 1688980957
transform 1 0 39836 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_433
timestamp 1688980957
transform 1 0 40940 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_21
timestamp 1688980957
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_38
timestamp 1688980957
transform 1 0 4600 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_76
timestamp 1688980957
transform 1 0 8096 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_82
timestamp 1688980957
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_92
timestamp 1688980957
transform 1 0 9568 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_104
timestamp 1688980957
transform 1 0 10672 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_112
timestamp 1688980957
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_138
timestamp 1688980957
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_148
timestamp 1688980957
transform 1 0 14720 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_162
timestamp 1688980957
transform 1 0 16008 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_170
timestamp 1688980957
transform 1 0 16744 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1688980957
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_203
timestamp 1688980957
transform 1 0 19780 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_210
timestamp 1688980957
transform 1 0 20424 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_222
timestamp 1688980957
transform 1 0 21528 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_230
timestamp 1688980957
transform 1 0 22264 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_238
timestamp 1688980957
transform 1 0 23000 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_250
timestamp 1688980957
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_270
timestamp 1688980957
transform 1 0 25944 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_278
timestamp 1688980957
transform 1 0 26680 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_298
timestamp 1688980957
transform 1 0 28520 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_306
timestamp 1688980957
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_318
timestamp 1688980957
transform 1 0 30360 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_326
timestamp 1688980957
transform 1 0 31096 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_334
timestamp 1688980957
transform 1 0 31832 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_346
timestamp 1688980957
transform 1 0 32936 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_361
timestamp 1688980957
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_370
timestamp 1688980957
transform 1 0 35144 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_382
timestamp 1688980957
transform 1 0 36248 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_402
timestamp 1688980957
transform 1 0 38088 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_407
timestamp 1688980957
transform 1 0 38548 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_419
timestamp 1688980957
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_421
timestamp 1688980957
transform 1 0 39836 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_427
timestamp 1688980957
transform 1 0 40388 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_7
timestamp 1688980957
transform 1 0 1748 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_11
timestamp 1688980957
transform 1 0 2116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_24
timestamp 1688980957
transform 1 0 3312 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_32
timestamp 1688980957
transform 1 0 4048 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_85
timestamp 1688980957
transform 1 0 8924 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_96
timestamp 1688980957
transform 1 0 9936 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_104
timestamp 1688980957
transform 1 0 10672 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_123
timestamp 1688980957
transform 1 0 12420 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_141
timestamp 1688980957
transform 1 0 14076 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 1688980957
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1688980957
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_175
timestamp 1688980957
transform 1 0 17204 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_191
timestamp 1688980957
transform 1 0 18676 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_205
timestamp 1688980957
transform 1 0 19964 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_209
timestamp 1688980957
transform 1 0 20332 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1688980957
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_232
timestamp 1688980957
transform 1 0 22448 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_241
timestamp 1688980957
transform 1 0 23276 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_253
timestamp 1688980957
transform 1 0 24380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_265
timestamp 1688980957
transform 1 0 25484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_277
timestamp 1688980957
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_285
timestamp 1688980957
transform 1 0 27324 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_291
timestamp 1688980957
transform 1 0 27876 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_299
timestamp 1688980957
transform 1 0 28612 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_311
timestamp 1688980957
transform 1 0 29716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_323
timestamp 1688980957
transform 1 0 30820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 1688980957
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_340
timestamp 1688980957
transform 1 0 32384 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_352
timestamp 1688980957
transform 1 0 33488 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_356
timestamp 1688980957
transform 1 0 33856 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_363
timestamp 1688980957
transform 1 0 34500 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_371
timestamp 1688980957
transform 1 0 35236 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_375
timestamp 1688980957
transform 1 0 35604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_387
timestamp 1688980957
transform 1 0 36708 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_391
timestamp 1688980957
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_393
timestamp 1688980957
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_405
timestamp 1688980957
transform 1 0 38364 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_413
timestamp 1688980957
transform 1 0 39100 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_23
timestamp 1688980957
transform 1 0 3220 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_32
timestamp 1688980957
transform 1 0 4048 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_44
timestamp 1688980957
transform 1 0 5152 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_56
timestamp 1688980957
transform 1 0 6256 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_75
timestamp 1688980957
transform 1 0 8004 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_95
timestamp 1688980957
transform 1 0 9844 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_114
timestamp 1688980957
transform 1 0 11592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_124
timestamp 1688980957
transform 1 0 12512 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_132
timestamp 1688980957
transform 1 0 13248 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_147
timestamp 1688980957
transform 1 0 14628 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_174
timestamp 1688980957
transform 1 0 17112 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_182
timestamp 1688980957
transform 1 0 17848 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_187
timestamp 1688980957
transform 1 0 18308 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_226
timestamp 1688980957
transform 1 0 21896 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_238
timestamp 1688980957
transform 1 0 23000 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_250
timestamp 1688980957
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_257
timestamp 1688980957
transform 1 0 24748 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_266
timestamp 1688980957
transform 1 0 25576 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_278
timestamp 1688980957
transform 1 0 26680 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_284
timestamp 1688980957
transform 1 0 27232 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_292
timestamp 1688980957
transform 1 0 27968 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_304
timestamp 1688980957
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_316
timestamp 1688980957
transform 1 0 30176 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_324
timestamp 1688980957
transform 1 0 30912 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_331
timestamp 1688980957
transform 1 0 31556 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_339
timestamp 1688980957
transform 1 0 32292 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_343
timestamp 1688980957
transform 1 0 32660 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_352
timestamp 1688980957
transform 1 0 33488 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_362
timestamp 1688980957
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_365
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_370
timestamp 1688980957
transform 1 0 35144 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_381
timestamp 1688980957
transform 1 0 36156 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_389
timestamp 1688980957
transform 1 0 36892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_403
timestamp 1688980957
transform 1 0 38180 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_407
timestamp 1688980957
transform 1 0 38548 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_414
timestamp 1688980957
transform 1 0 39192 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_424
timestamp 1688980957
transform 1 0 40112 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_428
timestamp 1688980957
transform 1 0 40480 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_19
timestamp 1688980957
transform 1 0 2852 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_31
timestamp 1688980957
transform 1 0 3956 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_42
timestamp 1688980957
transform 1 0 4968 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_54
timestamp 1688980957
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_80
timestamp 1688980957
transform 1 0 8464 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_92
timestamp 1688980957
transform 1 0 9568 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_100
timestamp 1688980957
transform 1 0 10304 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_108
timestamp 1688980957
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_154
timestamp 1688980957
transform 1 0 15272 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_166
timestamp 1688980957
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_178
timestamp 1688980957
transform 1 0 17480 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_190
timestamp 1688980957
transform 1 0 18584 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_200
timestamp 1688980957
transform 1 0 19504 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_221
timestamp 1688980957
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_249
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_257
timestamp 1688980957
transform 1 0 24748 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_268
timestamp 1688980957
transform 1 0 25760 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_275
timestamp 1688980957
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1688980957
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_300
timestamp 1688980957
transform 1 0 28704 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_323
timestamp 1688980957
transform 1 0 30820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_335
timestamp 1688980957
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_337
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 1688980957
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_361
timestamp 1688980957
transform 1 0 34316 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_369
timestamp 1688980957
transform 1 0 35052 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_375
timestamp 1688980957
transform 1 0 35604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_387
timestamp 1688980957
transform 1 0 36708 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 1688980957
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_412
timestamp 1688980957
transform 1 0 39008 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_14
timestamp 1688980957
transform 1 0 2392 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_18
timestamp 1688980957
transform 1 0 2760 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_49
timestamp 1688980957
transform 1 0 5612 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_59
timestamp 1688980957
transform 1 0 6532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_71
timestamp 1688980957
transform 1 0 7636 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_81
timestamp 1688980957
transform 1 0 8556 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_93
timestamp 1688980957
transform 1 0 9660 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_101
timestamp 1688980957
transform 1 0 10396 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_105
timestamp 1688980957
transform 1 0 10764 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_127
timestamp 1688980957
transform 1 0 12788 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_137
timestamp 1688980957
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_161
timestamp 1688980957
transform 1 0 15916 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_170
timestamp 1688980957
transform 1 0 16744 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_178
timestamp 1688980957
transform 1 0 17480 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_204
timestamp 1688980957
transform 1 0 19872 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_212
timestamp 1688980957
transform 1 0 20608 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_216
timestamp 1688980957
transform 1 0 20976 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_230
timestamp 1688980957
transform 1 0 22264 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_236
timestamp 1688980957
transform 1 0 22816 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_240
timestamp 1688980957
transform 1 0 23184 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_245
timestamp 1688980957
transform 1 0 23644 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1688980957
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_266
timestamp 1688980957
transform 1 0 25576 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_282
timestamp 1688980957
transform 1 0 27048 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_292
timestamp 1688980957
transform 1 0 27968 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_300
timestamp 1688980957
transform 1 0 28704 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_323
timestamp 1688980957
transform 1 0 30820 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_331
timestamp 1688980957
transform 1 0 31556 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 1688980957
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_365
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_377
timestamp 1688980957
transform 1 0 35788 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_386
timestamp 1688980957
transform 1 0 36616 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_398
timestamp 1688980957
transform 1 0 37720 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_406
timestamp 1688980957
transform 1 0 38456 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_421
timestamp 1688980957
transform 1 0 39836 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_24
timestamp 1688980957
transform 1 0 3312 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_36
timestamp 1688980957
transform 1 0 4416 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_44
timestamp 1688980957
transform 1 0 5152 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_66
timestamp 1688980957
transform 1 0 7176 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_104
timestamp 1688980957
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_127
timestamp 1688980957
transform 1 0 12788 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1688980957
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_173
timestamp 1688980957
transform 1 0 17020 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_190
timestamp 1688980957
transform 1 0 18584 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_208
timestamp 1688980957
transform 1 0 20240 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_220
timestamp 1688980957
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_244
timestamp 1688980957
transform 1 0 23552 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_250
timestamp 1688980957
transform 1 0 24104 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_256
timestamp 1688980957
transform 1 0 24656 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_270
timestamp 1688980957
transform 1 0 25944 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_278
timestamp 1688980957
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_287
timestamp 1688980957
transform 1 0 27508 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_299
timestamp 1688980957
transform 1 0 28612 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_305
timestamp 1688980957
transform 1 0 29164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_312
timestamp 1688980957
transform 1 0 29808 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_324
timestamp 1688980957
transform 1 0 30912 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_334
timestamp 1688980957
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_349
timestamp 1688980957
transform 1 0 33212 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_370
timestamp 1688980957
transform 1 0 35144 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_382
timestamp 1688980957
transform 1 0 36248 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_390
timestamp 1688980957
transform 1 0 36984 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_393
timestamp 1688980957
transform 1 0 37260 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_399
timestamp 1688980957
transform 1 0 37812 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_404
timestamp 1688980957
transform 1 0 38272 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_432
timestamp 1688980957
transform 1 0 40848 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_37
timestamp 1688980957
transform 1 0 4508 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_61
timestamp 1688980957
transform 1 0 6716 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_69
timestamp 1688980957
transform 1 0 7452 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_104
timestamp 1688980957
transform 1 0 10672 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_116
timestamp 1688980957
transform 1 0 11776 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_128
timestamp 1688980957
transform 1 0 12880 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_137
timestamp 1688980957
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_149
timestamp 1688980957
transform 1 0 14812 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_155
timestamp 1688980957
transform 1 0 15364 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_171
timestamp 1688980957
transform 1 0 16836 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_177
timestamp 1688980957
transform 1 0 17388 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_183
timestamp 1688980957
transform 1 0 17940 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_189
timestamp 1688980957
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1688980957
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_202
timestamp 1688980957
transform 1 0 19688 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_214
timestamp 1688980957
transform 1 0 20792 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_226
timestamp 1688980957
transform 1 0 21896 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_231
timestamp 1688980957
transform 1 0 22356 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_237
timestamp 1688980957
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_249
timestamp 1688980957
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_278
timestamp 1688980957
transform 1 0 26680 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_286
timestamp 1688980957
transform 1 0 27416 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_298
timestamp 1688980957
transform 1 0 28520 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_306
timestamp 1688980957
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_340
timestamp 1688980957
transform 1 0 32384 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_346
timestamp 1688980957
transform 1 0 32936 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_368
timestamp 1688980957
transform 1 0 34960 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_372
timestamp 1688980957
transform 1 0 35328 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_376
timestamp 1688980957
transform 1 0 35696 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_388
timestamp 1688980957
transform 1 0 36800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_408
timestamp 1688980957
transform 1 0 38640 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_419
timestamp 1688980957
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_424
timestamp 1688980957
transform 1 0 40112 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_432
timestamp 1688980957
transform 1 0 40848 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_26
timestamp 1688980957
transform 1 0 3496 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_38
timestamp 1688980957
transform 1 0 4600 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 1688980957
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 1688980957
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_109
timestamp 1688980957
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_117
timestamp 1688980957
transform 1 0 11868 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_127
timestamp 1688980957
transform 1 0 12788 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_139
timestamp 1688980957
transform 1 0 13892 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_151
timestamp 1688980957
transform 1 0 14996 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_163
timestamp 1688980957
transform 1 0 16100 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1688980957
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 1688980957
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_205
timestamp 1688980957
transform 1 0 19964 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_211
timestamp 1688980957
transform 1 0 20516 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_219
timestamp 1688980957
transform 1 0 21252 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1688980957
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 1688980957
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 1688980957
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 1688980957
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_276
timestamp 1688980957
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_287
timestamp 1688980957
transform 1 0 27508 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 1688980957
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 1688980957
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_329
timestamp 1688980957
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 1688980957
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_349
timestamp 1688980957
transform 1 0 33212 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_361
timestamp 1688980957
transform 1 0 34316 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_388
timestamp 1688980957
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_410
timestamp 1688980957
transform 1 0 38824 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_55
timestamp 1688980957
transform 1 0 6164 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_63
timestamp 1688980957
transform 1 0 6900 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_75
timestamp 1688980957
transform 1 0 8004 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1688980957
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_93
timestamp 1688980957
transform 1 0 9660 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_102
timestamp 1688980957
transform 1 0 10488 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_111
timestamp 1688980957
transform 1 0 11316 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_120
timestamp 1688980957
transform 1 0 12144 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_135
timestamp 1688980957
transform 1 0 13524 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_155
timestamp 1688980957
transform 1 0 15364 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_162
timestamp 1688980957
transform 1 0 16008 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_167
timestamp 1688980957
transform 1 0 16468 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_171
timestamp 1688980957
transform 1 0 16836 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_188
timestamp 1688980957
transform 1 0 18400 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_202
timestamp 1688980957
transform 1 0 19688 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_231
timestamp 1688980957
transform 1 0 22356 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_235
timestamp 1688980957
transform 1 0 22724 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_250
timestamp 1688980957
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_260
timestamp 1688980957
transform 1 0 25024 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_286
timestamp 1688980957
transform 1 0 27416 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1688980957
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_321
timestamp 1688980957
transform 1 0 30636 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_335
timestamp 1688980957
transform 1 0 31924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_343
timestamp 1688980957
transform 1 0 32660 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_351
timestamp 1688980957
transform 1 0 33396 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_357
timestamp 1688980957
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 1688980957
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_373
timestamp 1688980957
transform 1 0 35420 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_381
timestamp 1688980957
transform 1 0 36156 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_392
timestamp 1688980957
transform 1 0 37168 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_404
timestamp 1688980957
transform 1 0 38272 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_416
timestamp 1688980957
transform 1 0 39376 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_421
timestamp 1688980957
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_433
timestamp 1688980957
transform 1 0 40940 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_7
timestamp 1688980957
transform 1 0 1748 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_29
timestamp 1688980957
transform 1 0 3772 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_64
timestamp 1688980957
transform 1 0 6992 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_88
timestamp 1688980957
transform 1 0 9200 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_109
timestamp 1688980957
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_117
timestamp 1688980957
transform 1 0 11868 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_203
timestamp 1688980957
transform 1 0 19780 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_209
timestamp 1688980957
transform 1 0 20332 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_221
timestamp 1688980957
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_234
timestamp 1688980957
transform 1 0 22632 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_238
timestamp 1688980957
transform 1 0 23000 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_241
timestamp 1688980957
transform 1 0 23276 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_265
timestamp 1688980957
transform 1 0 25484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_277
timestamp 1688980957
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1688980957
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_305
timestamp 1688980957
transform 1 0 29164 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_316
timestamp 1688980957
transform 1 0 30176 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_322
timestamp 1688980957
transform 1 0 30728 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 1688980957
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_337
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_372
timestamp 1688980957
transform 1 0 35328 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_384
timestamp 1688980957
transform 1 0 36432 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_398
timestamp 1688980957
transform 1 0 37720 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_404
timestamp 1688980957
transform 1 0 38272 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_409
timestamp 1688980957
transform 1 0 38732 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_421
timestamp 1688980957
transform 1 0 39836 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_433
timestamp 1688980957
transform 1 0 40940 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_18
timestamp 1688980957
transform 1 0 2760 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_26
timestamp 1688980957
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_37
timestamp 1688980957
transform 1 0 4508 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_62
timestamp 1688980957
transform 1 0 6808 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1688980957
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_99
timestamp 1688980957
transform 1 0 10212 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_111
timestamp 1688980957
transform 1 0 11316 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_119
timestamp 1688980957
transform 1 0 12052 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_126
timestamp 1688980957
transform 1 0 12696 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_130
timestamp 1688980957
transform 1 0 13064 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_161
timestamp 1688980957
transform 1 0 15916 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_169
timestamp 1688980957
transform 1 0 16652 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_177
timestamp 1688980957
transform 1 0 17388 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_186
timestamp 1688980957
transform 1 0 18216 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_194
timestamp 1688980957
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_221
timestamp 1688980957
transform 1 0 21436 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_229
timestamp 1688980957
transform 1 0 22172 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_236
timestamp 1688980957
transform 1 0 22816 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_247
timestamp 1688980957
transform 1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 1688980957
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_265
timestamp 1688980957
transform 1 0 25484 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_281
timestamp 1688980957
transform 1 0 26956 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_293
timestamp 1688980957
transform 1 0 28060 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_317
timestamp 1688980957
transform 1 0 30268 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_328
timestamp 1688980957
transform 1 0 31280 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_333
timestamp 1688980957
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_345
timestamp 1688980957
transform 1 0 32844 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_353
timestamp 1688980957
transform 1 0 33580 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_371
timestamp 1688980957
transform 1 0 35236 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_386
timestamp 1688980957
transform 1 0 36616 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_392
timestamp 1688980957
transform 1 0 37168 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_419
timestamp 1688980957
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_424
timestamp 1688980957
transform 1 0 40112 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_432
timestamp 1688980957
transform 1 0 40848 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_11
timestamp 1688980957
transform 1 0 2116 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_23
timestamp 1688980957
transform 1 0 3220 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_35
timestamp 1688980957
transform 1 0 4324 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_47
timestamp 1688980957
transform 1 0 5428 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_69
timestamp 1688980957
transform 1 0 7452 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_83
timestamp 1688980957
transform 1 0 8740 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_97
timestamp 1688980957
transform 1 0 10028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_109
timestamp 1688980957
transform 1 0 11132 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 1688980957
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1688980957
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 1688980957
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_181
timestamp 1688980957
transform 1 0 17756 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_190
timestamp 1688980957
transform 1 0 18584 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_194
timestamp 1688980957
transform 1 0 18952 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_202
timestamp 1688980957
transform 1 0 19688 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 1688980957
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 1688980957
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 1688980957
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1688980957
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_281
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 1688980957
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_305
timestamp 1688980957
transform 1 0 29164 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_316
timestamp 1688980957
transform 1 0 30176 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_328
timestamp 1688980957
transform 1 0 31280 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_337
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_341
timestamp 1688980957
transform 1 0 32476 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 1688980957
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_361
timestamp 1688980957
transform 1 0 34316 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_369
timestamp 1688980957
transform 1 0 35052 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_385
timestamp 1688980957
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_391
timestamp 1688980957
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_414
timestamp 1688980957
transform 1 0 39192 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_26
timestamp 1688980957
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_38
timestamp 1688980957
transform 1 0 4600 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_50
timestamp 1688980957
transform 1 0 5704 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_62
timestamp 1688980957
transform 1 0 6808 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_74
timestamp 1688980957
transform 1 0 7912 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_82
timestamp 1688980957
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_97
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_130
timestamp 1688980957
transform 1 0 13064 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_138
timestamp 1688980957
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 1688980957
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_165
timestamp 1688980957
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_177
timestamp 1688980957
transform 1 0 17388 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 1688980957
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_212
timestamp 1688980957
transform 1 0 20608 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_221
timestamp 1688980957
transform 1 0 21436 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_230
timestamp 1688980957
transform 1 0 22264 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_242
timestamp 1688980957
transform 1 0 23368 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_250
timestamp 1688980957
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_267
timestamp 1688980957
transform 1 0 25668 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_281
timestamp 1688980957
transform 1 0 26956 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_293
timestamp 1688980957
transform 1 0 28060 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_303
timestamp 1688980957
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1688980957
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_321
timestamp 1688980957
transform 1 0 30636 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_332
timestamp 1688980957
transform 1 0 31648 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_341
timestamp 1688980957
transform 1 0 32476 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_353
timestamp 1688980957
transform 1 0 33580 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_358
timestamp 1688980957
transform 1 0 34040 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_365
timestamp 1688980957
transform 1 0 34684 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_373
timestamp 1688980957
transform 1 0 35420 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_381
timestamp 1688980957
transform 1 0 36156 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_385
timestamp 1688980957
transform 1 0 36524 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_419
timestamp 1688980957
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_424
timestamp 1688980957
transform 1 0 40112 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_432
timestamp 1688980957
transform 1 0 40848 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_7
timestamp 1688980957
transform 1 0 1748 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_11
timestamp 1688980957
transform 1 0 2116 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_35
timestamp 1688980957
transform 1 0 4324 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_46
timestamp 1688980957
transform 1 0 5336 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_54
timestamp 1688980957
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_81
timestamp 1688980957
transform 1 0 8556 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_90
timestamp 1688980957
transform 1 0 9384 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_102
timestamp 1688980957
transform 1 0 10488 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_110
timestamp 1688980957
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_136
timestamp 1688980957
transform 1 0 13616 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_149
timestamp 1688980957
transform 1 0 14812 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_153
timestamp 1688980957
transform 1 0 15180 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_159
timestamp 1688980957
transform 1 0 15732 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1688980957
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_234
timestamp 1688980957
transform 1 0 22632 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_241
timestamp 1688980957
transform 1 0 23276 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_258
timestamp 1688980957
transform 1 0 24840 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_290
timestamp 1688980957
transform 1 0 27784 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_302
timestamp 1688980957
transform 1 0 28888 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_319
timestamp 1688980957
transform 1 0 30452 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_327
timestamp 1688980957
transform 1 0 31188 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1688980957
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_345
timestamp 1688980957
transform 1 0 32844 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_356
timestamp 1688980957
transform 1 0 33856 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_371
timestamp 1688980957
transform 1 0 35236 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_383
timestamp 1688980957
transform 1 0 36340 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_391
timestamp 1688980957
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_393
timestamp 1688980957
transform 1 0 37260 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_413
timestamp 1688980957
transform 1 0 39100 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_21
timestamp 1688980957
transform 1 0 3036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_37
timestamp 1688980957
transform 1 0 4508 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_56
timestamp 1688980957
transform 1 0 6256 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_72
timestamp 1688980957
transform 1 0 7728 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_106
timestamp 1688980957
transform 1 0 10856 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_118
timestamp 1688980957
transform 1 0 11960 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_122
timestamp 1688980957
transform 1 0 12328 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_127
timestamp 1688980957
transform 1 0 12788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_163
timestamp 1688980957
transform 1 0 16100 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_172
timestamp 1688980957
transform 1 0 16928 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_180
timestamp 1688980957
transform 1 0 17664 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_193
timestamp 1688980957
transform 1 0 18860 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 1688980957
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_229
timestamp 1688980957
transform 1 0 22172 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_250
timestamp 1688980957
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_264
timestamp 1688980957
transform 1 0 25392 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_272
timestamp 1688980957
transform 1 0 26128 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_294
timestamp 1688980957
transform 1 0 28152 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_314
timestamp 1688980957
transform 1 0 29992 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_340
timestamp 1688980957
transform 1 0 32384 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_348
timestamp 1688980957
transform 1 0 33120 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 1688980957
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_370
timestamp 1688980957
transform 1 0 35144 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_374
timestamp 1688980957
transform 1 0 35512 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_390
timestamp 1688980957
transform 1 0 36984 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_412
timestamp 1688980957
transform 1 0 39008 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_421
timestamp 1688980957
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_433
timestamp 1688980957
transform 1 0 40940 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_44
timestamp 1688980957
transform 1 0 5152 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_52
timestamp 1688980957
transform 1 0 5888 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_64
timestamp 1688980957
transform 1 0 6992 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_73
timestamp 1688980957
transform 1 0 7820 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_82
timestamp 1688980957
transform 1 0 8648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_101
timestamp 1688980957
transform 1 0 10396 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_109
timestamp 1688980957
transform 1 0 11132 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_119
timestamp 1688980957
transform 1 0 12052 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_131
timestamp 1688980957
transform 1 0 13156 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_137
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_149
timestamp 1688980957
transform 1 0 14812 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_157
timestamp 1688980957
transform 1 0 15548 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_163
timestamp 1688980957
transform 1 0 16100 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1688980957
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_181
timestamp 1688980957
transform 1 0 17756 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_189
timestamp 1688980957
transform 1 0 18492 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_201
timestamp 1688980957
transform 1 0 19596 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_213
timestamp 1688980957
transform 1 0 20700 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_221
timestamp 1688980957
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 1688980957
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_249
timestamp 1688980957
transform 1 0 24012 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_257
timestamp 1688980957
transform 1 0 24748 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_269
timestamp 1688980957
transform 1 0 25852 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_273
timestamp 1688980957
transform 1 0 26220 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_290
timestamp 1688980957
transform 1 0 27784 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_301
timestamp 1688980957
transform 1 0 28796 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_331
timestamp 1688980957
transform 1 0 31556 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1688980957
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_347
timestamp 1688980957
transform 1 0 33028 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_359
timestamp 1688980957
transform 1 0 34132 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_371
timestamp 1688980957
transform 1 0 35236 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_379
timestamp 1688980957
transform 1 0 35972 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_389
timestamp 1688980957
transform 1 0 36892 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_393
timestamp 1688980957
transform 1 0 37260 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_405
timestamp 1688980957
transform 1 0 38364 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_409
timestamp 1688980957
transform 1 0 38732 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_430
timestamp 1688980957
transform 1 0 40664 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1688980957
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_72
timestamp 1688980957
transform 1 0 7728 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_109
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_122
timestamp 1688980957
transform 1 0 12328 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_134
timestamp 1688980957
transform 1 0 13432 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_153
timestamp 1688980957
transform 1 0 15180 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_168
timestamp 1688980957
transform 1 0 16560 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_176
timestamp 1688980957
transform 1 0 17296 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_181
timestamp 1688980957
transform 1 0 17756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_193
timestamp 1688980957
transform 1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_209
timestamp 1688980957
transform 1 0 20332 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_213
timestamp 1688980957
transform 1 0 20700 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_220
timestamp 1688980957
transform 1 0 21344 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_232
timestamp 1688980957
transform 1 0 22448 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_237
timestamp 1688980957
transform 1 0 22908 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_249
timestamp 1688980957
transform 1 0 24012 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_259
timestamp 1688980957
transform 1 0 24932 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_267
timestamp 1688980957
transform 1 0 25668 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_275
timestamp 1688980957
transform 1 0 26404 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_287
timestamp 1688980957
transform 1 0 27508 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_299
timestamp 1688980957
transform 1 0 28612 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1688980957
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_317
timestamp 1688980957
transform 1 0 30268 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_325
timestamp 1688980957
transform 1 0 31004 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_337
timestamp 1688980957
transform 1 0 32108 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_349
timestamp 1688980957
transform 1 0 33212 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_361
timestamp 1688980957
transform 1 0 34316 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_371
timestamp 1688980957
transform 1 0 35236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_424
timestamp 1688980957
transform 1 0 40112 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_33
timestamp 1688980957
transform 1 0 4140 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_48
timestamp 1688980957
transform 1 0 5520 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_61
timestamp 1688980957
transform 1 0 6716 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_84
timestamp 1688980957
transform 1 0 8832 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_90
timestamp 1688980957
transform 1 0 9384 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_102
timestamp 1688980957
transform 1 0 10488 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_110
timestamp 1688980957
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_117
timestamp 1688980957
transform 1 0 11868 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_126
timestamp 1688980957
transform 1 0 12696 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_133
timestamp 1688980957
transform 1 0 13340 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_150
timestamp 1688980957
transform 1 0 14904 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_158
timestamp 1688980957
transform 1 0 15640 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_182
timestamp 1688980957
transform 1 0 17848 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_194
timestamp 1688980957
transform 1 0 18952 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_221
timestamp 1688980957
transform 1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_231
timestamp 1688980957
transform 1 0 22356 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_243
timestamp 1688980957
transform 1 0 23460 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_247
timestamp 1688980957
transform 1 0 23828 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_254
timestamp 1688980957
transform 1 0 24472 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_262
timestamp 1688980957
transform 1 0 25208 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_270
timestamp 1688980957
transform 1 0 25944 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_278
timestamp 1688980957
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_281
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_288
timestamp 1688980957
transform 1 0 27600 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_300
timestamp 1688980957
transform 1 0 28704 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_312
timestamp 1688980957
transform 1 0 29808 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_324
timestamp 1688980957
transform 1 0 30912 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_343
timestamp 1688980957
transform 1 0 32660 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_362
timestamp 1688980957
transform 1 0 34408 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_370
timestamp 1688980957
transform 1 0 35144 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_389
timestamp 1688980957
transform 1 0 36892 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_412
timestamp 1688980957
transform 1 0 39008 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_36
timestamp 1688980957
transform 1 0 4416 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_57
timestamp 1688980957
transform 1 0 6348 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_80
timestamp 1688980957
transform 1 0 8464 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_96
timestamp 1688980957
transform 1 0 9936 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_108
timestamp 1688980957
transform 1 0 11040 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_115
timestamp 1688980957
transform 1 0 11684 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_120
timestamp 1688980957
transform 1 0 12144 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_147
timestamp 1688980957
transform 1 0 14628 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_159
timestamp 1688980957
transform 1 0 15732 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_165
timestamp 1688980957
transform 1 0 16284 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1688980957
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_215
timestamp 1688980957
transform 1 0 20884 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_225
timestamp 1688980957
transform 1 0 21804 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_229
timestamp 1688980957
transform 1 0 22172 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_238
timestamp 1688980957
transform 1 0 23000 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_260
timestamp 1688980957
transform 1 0 25024 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_272
timestamp 1688980957
transform 1 0 26128 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_296
timestamp 1688980957
transform 1 0 28336 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_306
timestamp 1688980957
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_324
timestamp 1688980957
transform 1 0 30912 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_340
timestamp 1688980957
transform 1 0 32384 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_344
timestamp 1688980957
transform 1 0 32752 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_371
timestamp 1688980957
transform 1 0 35236 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_391
timestamp 1688980957
transform 1 0 37076 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_403
timestamp 1688980957
transform 1 0 38180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_415
timestamp 1688980957
transform 1 0 39284 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_419
timestamp 1688980957
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_421
timestamp 1688980957
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_433
timestamp 1688980957
transform 1 0 40940 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_7
timestamp 1688980957
transform 1 0 1748 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_11
timestamp 1688980957
transform 1 0 2116 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_23
timestamp 1688980957
transform 1 0 3220 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_35
timestamp 1688980957
transform 1 0 4324 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_47
timestamp 1688980957
transform 1 0 5428 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_61
timestamp 1688980957
transform 1 0 6716 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_70
timestamp 1688980957
transform 1 0 7544 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_82
timestamp 1688980957
transform 1 0 8648 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_95
timestamp 1688980957
transform 1 0 9844 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_103
timestamp 1688980957
transform 1 0 10580 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_109
timestamp 1688980957
transform 1 0 11132 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_133
timestamp 1688980957
transform 1 0 13340 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_141
timestamp 1688980957
transform 1 0 14076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_150
timestamp 1688980957
transform 1 0 14904 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_162
timestamp 1688980957
transform 1 0 16008 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_185
timestamp 1688980957
transform 1 0 18124 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_193
timestamp 1688980957
transform 1 0 18860 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_213
timestamp 1688980957
transform 1 0 20700 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_221
timestamp 1688980957
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_225
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_249
timestamp 1688980957
transform 1 0 24012 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_262
timestamp 1688980957
transform 1 0 25208 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_270
timestamp 1688980957
transform 1 0 25944 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_289
timestamp 1688980957
transform 1 0 27692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_301
timestamp 1688980957
transform 1 0 28796 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_315
timestamp 1688980957
transform 1 0 30084 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_323
timestamp 1688980957
transform 1 0 30820 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_330
timestamp 1688980957
transform 1 0 31464 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_354
timestamp 1688980957
transform 1 0 33672 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_366
timestamp 1688980957
transform 1 0 34776 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_377
timestamp 1688980957
transform 1 0 35788 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_381
timestamp 1688980957
transform 1 0 36156 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_388
timestamp 1688980957
transform 1 0 36800 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_393
timestamp 1688980957
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_405
timestamp 1688980957
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_417
timestamp 1688980957
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_429
timestamp 1688980957
transform 1 0 40572 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1688980957
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_68
timestamp 1688980957
transform 1 0 7360 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_91
timestamp 1688980957
transform 1 0 9476 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_102
timestamp 1688980957
transform 1 0 10488 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_112
timestamp 1688980957
transform 1 0 11408 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_118
timestamp 1688980957
transform 1 0 11960 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_130
timestamp 1688980957
transform 1 0 13064 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_138
timestamp 1688980957
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_163
timestamp 1688980957
transform 1 0 16100 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_172
timestamp 1688980957
transform 1 0 16928 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_184
timestamp 1688980957
transform 1 0 18032 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_203
timestamp 1688980957
transform 1 0 19780 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_210
timestamp 1688980957
transform 1 0 20424 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_234
timestamp 1688980957
transform 1 0 22632 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_249
timestamp 1688980957
transform 1 0 24012 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_269
timestamp 1688980957
transform 1 0 25852 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 1688980957
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_301
timestamp 1688980957
transform 1 0 28796 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1688980957
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_321
timestamp 1688980957
transform 1 0 30636 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_328
timestamp 1688980957
transform 1 0 31280 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_340
timestamp 1688980957
transform 1 0 32384 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_348
timestamp 1688980957
transform 1 0 33120 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 1688980957
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_377
timestamp 1688980957
transform 1 0 35788 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_385
timestamp 1688980957
transform 1 0 36524 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_397
timestamp 1688980957
transform 1 0 37628 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_409
timestamp 1688980957
transform 1 0 38732 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_417
timestamp 1688980957
transform 1 0 39468 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_421
timestamp 1688980957
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_433
timestamp 1688980957
transform 1 0 40940 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_33
timestamp 1688980957
transform 1 0 4140 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_37
timestamp 1688980957
transform 1 0 4508 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_48
timestamp 1688980957
transform 1 0 5520 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_66
timestamp 1688980957
transform 1 0 7176 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_78
timestamp 1688980957
transform 1 0 8280 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_90
timestamp 1688980957
transform 1 0 9384 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_94
timestamp 1688980957
transform 1 0 9752 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_107
timestamp 1688980957
transform 1 0 10948 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 1688980957
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_137
timestamp 1688980957
transform 1 0 13708 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_153
timestamp 1688980957
transform 1 0 15180 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_160
timestamp 1688980957
transform 1 0 15824 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1688980957
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_193
timestamp 1688980957
transform 1 0 18860 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_201
timestamp 1688980957
transform 1 0 19596 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_207
timestamp 1688980957
transform 1 0 20148 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_219
timestamp 1688980957
transform 1 0 21252 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_272
timestamp 1688980957
transform 1 0 26128 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1688980957
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_305
timestamp 1688980957
transform 1 0 29164 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_309
timestamp 1688980957
transform 1 0 29532 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_318
timestamp 1688980957
transform 1 0 30360 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_349
timestamp 1688980957
transform 1 0 33212 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_371
timestamp 1688980957
transform 1 0 35236 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_383
timestamp 1688980957
transform 1 0 36340 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 1688980957
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 1688980957
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_405
timestamp 1688980957
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_417
timestamp 1688980957
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_429
timestamp 1688980957
transform 1 0 40572 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_11
timestamp 1688980957
transform 1 0 2116 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_16
timestamp 1688980957
transform 1 0 2576 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_50
timestamp 1688980957
transform 1 0 5704 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_56
timestamp 1688980957
transform 1 0 6256 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_64
timestamp 1688980957
transform 1 0 6992 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 1688980957
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1688980957
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_91
timestamp 1688980957
transform 1 0 9476 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_107
timestamp 1688980957
transform 1 0 10948 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_119
timestamp 1688980957
transform 1 0 12052 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_130
timestamp 1688980957
transform 1 0 13064 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_157
timestamp 1688980957
transform 1 0 15548 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_163
timestamp 1688980957
transform 1 0 16100 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_169
timestamp 1688980957
transform 1 0 16652 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_181
timestamp 1688980957
transform 1 0 17756 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_190
timestamp 1688980957
transform 1 0 18584 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_195
timestamp 1688980957
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_200
timestamp 1688980957
transform 1 0 19504 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_212
timestamp 1688980957
transform 1 0 20608 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_224
timestamp 1688980957
transform 1 0 21712 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_236
timestamp 1688980957
transform 1 0 22816 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_248
timestamp 1688980957
transform 1 0 23920 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_265
timestamp 1688980957
transform 1 0 25484 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_272
timestamp 1688980957
transform 1 0 26128 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_302
timestamp 1688980957
transform 1 0 28888 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_323
timestamp 1688980957
transform 1 0 30820 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_331
timestamp 1688980957
transform 1 0 31556 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_338
timestamp 1688980957
transform 1 0 32200 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_350
timestamp 1688980957
transform 1 0 33304 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_358
timestamp 1688980957
transform 1 0 34040 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1688980957
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1688980957
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 1688980957
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_401
timestamp 1688980957
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_413
timestamp 1688980957
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_419
timestamp 1688980957
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_421
timestamp 1688980957
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_433
timestamp 1688980957
transform 1 0 40940 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_30
timestamp 1688980957
transform 1 0 3864 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_34
timestamp 1688980957
transform 1 0 4232 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_76
timestamp 1688980957
transform 1 0 8096 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_88
timestamp 1688980957
transform 1 0 9200 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_101
timestamp 1688980957
transform 1 0 10396 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_109
timestamp 1688980957
transform 1 0 11132 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_142
timestamp 1688980957
transform 1 0 14168 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_157
timestamp 1688980957
transform 1 0 15548 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 1688980957
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_178
timestamp 1688980957
transform 1 0 17480 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_182
timestamp 1688980957
transform 1 0 17848 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_238
timestamp 1688980957
transform 1 0 23000 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_250
timestamp 1688980957
transform 1 0 24104 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_262
timestamp 1688980957
transform 1 0 25208 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_274
timestamp 1688980957
transform 1 0 26312 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_281
timestamp 1688980957
transform 1 0 26956 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_319
timestamp 1688980957
transform 1 0 30452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_331
timestamp 1688980957
transform 1 0 31556 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 1688980957
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 1688980957
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 1688980957
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_361
timestamp 1688980957
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_373
timestamp 1688980957
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_385
timestamp 1688980957
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 1688980957
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_393
timestamp 1688980957
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_405
timestamp 1688980957
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_417
timestamp 1688980957
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_429
timestamp 1688980957
transform 1 0 40572 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1688980957
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 1688980957
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_77
timestamp 1688980957
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 1688980957
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_97
timestamp 1688980957
transform 1 0 10028 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_106
timestamp 1688980957
transform 1 0 10856 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_112
timestamp 1688980957
transform 1 0 11408 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_120
timestamp 1688980957
transform 1 0 12144 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_132
timestamp 1688980957
transform 1 0 13248 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_136
timestamp 1688980957
transform 1 0 13616 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_175
timestamp 1688980957
transform 1 0 17204 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_187
timestamp 1688980957
transform 1 0 18308 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_202
timestamp 1688980957
transform 1 0 19688 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_214
timestamp 1688980957
transform 1 0 20792 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_226
timestamp 1688980957
transform 1 0 21896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_247
timestamp 1688980957
transform 1 0 23828 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_251
timestamp 1688980957
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_266
timestamp 1688980957
transform 1 0 25576 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_277
timestamp 1688980957
transform 1 0 26588 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_292
timestamp 1688980957
transform 1 0 27968 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_304
timestamp 1688980957
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_339
timestamp 1688980957
transform 1 0 32292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_351
timestamp 1688980957
transform 1 0 33396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 1688980957
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1688980957
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1688980957
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_389
timestamp 1688980957
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_401
timestamp 1688980957
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_413
timestamp 1688980957
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_419
timestamp 1688980957
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_421
timestamp 1688980957
transform 1 0 39836 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_429
timestamp 1688980957
transform 1 0 40572 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1688980957
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 1688980957
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 1688980957
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 1688980957
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 1688980957
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_60
timestamp 1688980957
transform 1 0 6624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_78
timestamp 1688980957
transform 1 0 8280 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_82
timestamp 1688980957
transform 1 0 8648 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_93
timestamp 1688980957
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_109
timestamp 1688980957
transform 1 0 11132 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_116
timestamp 1688980957
transform 1 0 11776 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_128
timestamp 1688980957
transform 1 0 12880 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_140
timestamp 1688980957
transform 1 0 13984 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_149
timestamp 1688980957
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_165
timestamp 1688980957
transform 1 0 16284 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_169
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_192
timestamp 1688980957
transform 1 0 18768 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_204
timestamp 1688980957
transform 1 0 19872 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_212
timestamp 1688980957
transform 1 0 20608 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_217
timestamp 1688980957
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_223
timestamp 1688980957
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_230
timestamp 1688980957
transform 1 0 22264 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_235
timestamp 1688980957
transform 1 0 22724 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_275
timestamp 1688980957
transform 1 0 26404 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_279
timestamp 1688980957
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_302
timestamp 1688980957
transform 1 0 28888 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_314
timestamp 1688980957
transform 1 0 29992 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_326
timestamp 1688980957
transform 1 0 31096 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_334
timestamp 1688980957
transform 1 0 31832 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_337
timestamp 1688980957
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_349
timestamp 1688980957
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_361
timestamp 1688980957
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_373
timestamp 1688980957
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_385
timestamp 1688980957
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_391
timestamp 1688980957
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_393
timestamp 1688980957
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_405
timestamp 1688980957
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_417
timestamp 1688980957
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_429
timestamp 1688980957
transform 1 0 40572 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_15
timestamp 1688980957
transform 1 0 2484 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_23
timestamp 1688980957
transform 1 0 3220 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_38
timestamp 1688980957
transform 1 0 4600 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_42
timestamp 1688980957
transform 1 0 4968 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_54
timestamp 1688980957
transform 1 0 6072 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_76
timestamp 1688980957
transform 1 0 8096 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_97
timestamp 1688980957
transform 1 0 10028 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_105
timestamp 1688980957
transform 1 0 10764 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_114
timestamp 1688980957
transform 1 0 11592 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_126
timestamp 1688980957
transform 1 0 12696 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_138
timestamp 1688980957
transform 1 0 13800 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 1688980957
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_165
timestamp 1688980957
transform 1 0 16284 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_171
timestamp 1688980957
transform 1 0 16836 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_185
timestamp 1688980957
transform 1 0 18124 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_193
timestamp 1688980957
transform 1 0 18860 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_197
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_205
timestamp 1688980957
transform 1 0 19964 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_228
timestamp 1688980957
transform 1 0 22080 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_240
timestamp 1688980957
transform 1 0 23184 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_253
timestamp 1688980957
transform 1 0 24380 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_277
timestamp 1688980957
transform 1 0 26588 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_285
timestamp 1688980957
transform 1 0 27324 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_309
timestamp 1688980957
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_321
timestamp 1688980957
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_333
timestamp 1688980957
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_345
timestamp 1688980957
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_357
timestamp 1688980957
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_363
timestamp 1688980957
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_365
timestamp 1688980957
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_377
timestamp 1688980957
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_389
timestamp 1688980957
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_401
timestamp 1688980957
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_413
timestamp 1688980957
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_419
timestamp 1688980957
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_421
timestamp 1688980957
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_433
timestamp 1688980957
transform 1 0 40940 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_3
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_11
timestamp 1688980957
transform 1 0 2116 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_61
timestamp 1688980957
transform 1 0 6716 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_75
timestamp 1688980957
transform 1 0 8004 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_87
timestamp 1688980957
transform 1 0 9108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_99
timestamp 1688980957
transform 1 0 10212 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_105
timestamp 1688980957
transform 1 0 10764 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 1688980957
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_120
timestamp 1688980957
transform 1 0 12144 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_124
timestamp 1688980957
transform 1 0 12512 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_156
timestamp 1688980957
transform 1 0 15456 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_169
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_207
timestamp 1688980957
transform 1 0 20148 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_215
timestamp 1688980957
transform 1 0 20884 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_225
timestamp 1688980957
transform 1 0 21804 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_240
timestamp 1688980957
transform 1 0 23184 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_252
timestamp 1688980957
transform 1 0 24288 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_264
timestamp 1688980957
transform 1 0 25392 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_273
timestamp 1688980957
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_279
timestamp 1688980957
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_289
timestamp 1688980957
transform 1 0 27692 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_301
timestamp 1688980957
transform 1 0 28796 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_313
timestamp 1688980957
transform 1 0 29900 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_325
timestamp 1688980957
transform 1 0 31004 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_333
timestamp 1688980957
transform 1 0 31740 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_337
timestamp 1688980957
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_349
timestamp 1688980957
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_361
timestamp 1688980957
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_373
timestamp 1688980957
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_385
timestamp 1688980957
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_391
timestamp 1688980957
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_393
timestamp 1688980957
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_405
timestamp 1688980957
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_417
timestamp 1688980957
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_429
timestamp 1688980957
transform 1 0 40572 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_3
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_15
timestamp 1688980957
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 1688980957
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_37
timestamp 1688980957
transform 1 0 4508 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_49
timestamp 1688980957
transform 1 0 5612 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_61
timestamp 1688980957
transform 1 0 6716 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_67
timestamp 1688980957
transform 1 0 7268 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_80
timestamp 1688980957
transform 1 0 8464 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_120
timestamp 1688980957
transform 1 0 12144 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_126
timestamp 1688980957
transform 1 0 12696 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_135
timestamp 1688980957
transform 1 0 13524 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_139
timestamp 1688980957
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_147
timestamp 1688980957
transform 1 0 14628 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_153
timestamp 1688980957
transform 1 0 15180 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_165
timestamp 1688980957
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_177
timestamp 1688980957
transform 1 0 17388 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_181
timestamp 1688980957
transform 1 0 17756 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_185
timestamp 1688980957
transform 1 0 18124 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_193
timestamp 1688980957
transform 1 0 18860 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_197
timestamp 1688980957
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_209
timestamp 1688980957
transform 1 0 20332 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_217
timestamp 1688980957
transform 1 0 21068 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_247
timestamp 1688980957
transform 1 0 23828 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_251
timestamp 1688980957
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_253
timestamp 1688980957
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_265
timestamp 1688980957
transform 1 0 25484 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_289
timestamp 1688980957
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_301
timestamp 1688980957
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_307
timestamp 1688980957
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_309
timestamp 1688980957
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_321
timestamp 1688980957
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_333
timestamp 1688980957
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_345
timestamp 1688980957
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_357
timestamp 1688980957
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_363
timestamp 1688980957
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_365
timestamp 1688980957
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_377
timestamp 1688980957
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_389
timestamp 1688980957
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_401
timestamp 1688980957
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_413
timestamp 1688980957
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_419
timestamp 1688980957
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_421
timestamp 1688980957
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_433
timestamp 1688980957
transform 1 0 40940 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_3
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_15
timestamp 1688980957
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_27
timestamp 1688980957
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_39
timestamp 1688980957
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_51
timestamp 1688980957
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_55
timestamp 1688980957
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_85
timestamp 1688980957
transform 1 0 8924 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_93
timestamp 1688980957
transform 1 0 9660 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_108
timestamp 1688980957
transform 1 0 11040 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_118
timestamp 1688980957
transform 1 0 11960 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_126
timestamp 1688980957
transform 1 0 12696 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_151
timestamp 1688980957
transform 1 0 14996 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_167
timestamp 1688980957
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_174
timestamp 1688980957
transform 1 0 17112 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_186
timestamp 1688980957
transform 1 0 18216 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_190
timestamp 1688980957
transform 1 0 18584 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_198
timestamp 1688980957
transform 1 0 19320 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_204
timestamp 1688980957
transform 1 0 19872 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_216
timestamp 1688980957
transform 1 0 20976 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_228
timestamp 1688980957
transform 1 0 22080 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_236
timestamp 1688980957
transform 1 0 22816 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_260
timestamp 1688980957
transform 1 0 25024 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_272
timestamp 1688980957
transform 1 0 26128 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_281
timestamp 1688980957
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_293
timestamp 1688980957
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_305
timestamp 1688980957
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_317
timestamp 1688980957
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_329
timestamp 1688980957
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_335
timestamp 1688980957
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_337
timestamp 1688980957
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_349
timestamp 1688980957
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_361
timestamp 1688980957
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_373
timestamp 1688980957
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_385
timestamp 1688980957
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_391
timestamp 1688980957
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_393
timestamp 1688980957
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_405
timestamp 1688980957
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_417
timestamp 1688980957
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_429
timestamp 1688980957
transform 1 0 40572 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_3
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_9
timestamp 1688980957
transform 1 0 1932 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_13
timestamp 1688980957
transform 1 0 2300 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_24
timestamp 1688980957
transform 1 0 3312 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_29
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_33
timestamp 1688980957
transform 1 0 4140 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_37
timestamp 1688980957
transform 1 0 4508 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_47
timestamp 1688980957
transform 1 0 5428 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_59
timestamp 1688980957
transform 1 0 6532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_71
timestamp 1688980957
transform 1 0 7636 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_80
timestamp 1688980957
transform 1 0 8464 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_85
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_97
timestamp 1688980957
transform 1 0 10028 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_109
timestamp 1688980957
transform 1 0 11132 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_113
timestamp 1688980957
transform 1 0 11500 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_125
timestamp 1688980957
transform 1 0 12604 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_137
timestamp 1688980957
transform 1 0 13708 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_141
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_152
timestamp 1688980957
transform 1 0 15088 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_172
timestamp 1688980957
transform 1 0 16928 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_185
timestamp 1688980957
transform 1 0 18124 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_197
timestamp 1688980957
transform 1 0 19228 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_222
timestamp 1688980957
transform 1 0 21528 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_230
timestamp 1688980957
transform 1 0 22264 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_237
timestamp 1688980957
transform 1 0 22908 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_249
timestamp 1688980957
transform 1 0 24012 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_253
timestamp 1688980957
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_265
timestamp 1688980957
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_277
timestamp 1688980957
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_289
timestamp 1688980957
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_301
timestamp 1688980957
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_307
timestamp 1688980957
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_309
timestamp 1688980957
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_321
timestamp 1688980957
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_333
timestamp 1688980957
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_345
timestamp 1688980957
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_357
timestamp 1688980957
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_363
timestamp 1688980957
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_365
timestamp 1688980957
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_377
timestamp 1688980957
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_389
timestamp 1688980957
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_401
timestamp 1688980957
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_413
timestamp 1688980957
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_419
timestamp 1688980957
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_421
timestamp 1688980957
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_433
timestamp 1688980957
transform 1 0 40940 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_26
timestamp 1688980957
transform 1 0 3496 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_52
timestamp 1688980957
transform 1 0 5888 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_69
timestamp 1688980957
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_81
timestamp 1688980957
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_93
timestamp 1688980957
transform 1 0 9660 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_109
timestamp 1688980957
transform 1 0 11132 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_113
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_124
timestamp 1688980957
transform 1 0 12512 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_128
timestamp 1688980957
transform 1 0 12880 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_140
timestamp 1688980957
transform 1 0 13984 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_144
timestamp 1688980957
transform 1 0 14352 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_148
timestamp 1688980957
transform 1 0 14720 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_152
timestamp 1688980957
transform 1 0 15088 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_164
timestamp 1688980957
transform 1 0 16192 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_169
timestamp 1688980957
transform 1 0 16652 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_180
timestamp 1688980957
transform 1 0 17664 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_192
timestamp 1688980957
transform 1 0 18768 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_198
timestamp 1688980957
transform 1 0 19320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_208
timestamp 1688980957
transform 1 0 20240 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_216
timestamp 1688980957
transform 1 0 20976 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_248
timestamp 1688980957
transform 1 0 23920 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_260
timestamp 1688980957
transform 1 0 25024 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_272
timestamp 1688980957
transform 1 0 26128 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_281
timestamp 1688980957
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_293
timestamp 1688980957
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_305
timestamp 1688980957
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_317
timestamp 1688980957
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_329
timestamp 1688980957
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_335
timestamp 1688980957
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_337
timestamp 1688980957
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_349
timestamp 1688980957
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_361
timestamp 1688980957
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_373
timestamp 1688980957
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_385
timestamp 1688980957
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_391
timestamp 1688980957
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_393
timestamp 1688980957
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_405
timestamp 1688980957
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_417
timestamp 1688980957
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_429
timestamp 1688980957
transform 1 0 40572 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_3
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_15
timestamp 1688980957
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 1688980957
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 1688980957
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 1688980957
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_65
timestamp 1688980957
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_77
timestamp 1688980957
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_83
timestamp 1688980957
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_93
timestamp 1688980957
transform 1 0 9660 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_139
timestamp 1688980957
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_164
timestamp 1688980957
transform 1 0 16192 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_170
timestamp 1688980957
transform 1 0 16744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_194
timestamp 1688980957
transform 1 0 18952 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_197
timestamp 1688980957
transform 1 0 19228 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_221
timestamp 1688980957
transform 1 0 21436 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_253
timestamp 1688980957
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_265
timestamp 1688980957
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_277
timestamp 1688980957
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_289
timestamp 1688980957
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_301
timestamp 1688980957
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_307
timestamp 1688980957
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_309
timestamp 1688980957
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_321
timestamp 1688980957
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_333
timestamp 1688980957
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_345
timestamp 1688980957
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_357
timestamp 1688980957
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_363
timestamp 1688980957
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_365
timestamp 1688980957
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_377
timestamp 1688980957
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_389
timestamp 1688980957
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_401
timestamp 1688980957
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_413
timestamp 1688980957
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_419
timestamp 1688980957
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_421
timestamp 1688980957
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_433
timestamp 1688980957
transform 1 0 40940 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_9
timestamp 1688980957
transform 1 0 1932 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_21
timestamp 1688980957
transform 1 0 3036 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_27
timestamp 1688980957
transform 1 0 3588 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_29
timestamp 1688980957
transform 1 0 3772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_41
timestamp 1688980957
transform 1 0 4876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_53
timestamp 1688980957
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_57
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_69
timestamp 1688980957
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_81
timestamp 1688980957
transform 1 0 8556 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_85
timestamp 1688980957
transform 1 0 8924 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_93
timestamp 1688980957
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_105
timestamp 1688980957
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_111
timestamp 1688980957
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 1688980957
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_137
timestamp 1688980957
transform 1 0 13708 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_141
timestamp 1688980957
transform 1 0 14076 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_153
timestamp 1688980957
transform 1 0 15180 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_165
timestamp 1688980957
transform 1 0 16284 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_169
timestamp 1688980957
transform 1 0 16652 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_175
timestamp 1688980957
transform 1 0 17204 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_179
timestamp 1688980957
transform 1 0 17572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_191
timestamp 1688980957
transform 1 0 18676 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_195
timestamp 1688980957
transform 1 0 19044 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_197
timestamp 1688980957
transform 1 0 19228 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_203
timestamp 1688980957
transform 1 0 19780 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_215
timestamp 1688980957
transform 1 0 20884 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_223
timestamp 1688980957
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_225
timestamp 1688980957
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_237
timestamp 1688980957
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_249
timestamp 1688980957
transform 1 0 24012 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_253
timestamp 1688980957
transform 1 0 24380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_265
timestamp 1688980957
transform 1 0 25484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_277
timestamp 1688980957
transform 1 0 26588 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_281
timestamp 1688980957
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_293
timestamp 1688980957
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_305
timestamp 1688980957
transform 1 0 29164 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_309
timestamp 1688980957
transform 1 0 29532 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_321
timestamp 1688980957
transform 1 0 30636 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_331
timestamp 1688980957
transform 1 0 31556 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_335
timestamp 1688980957
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_337
timestamp 1688980957
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_349
timestamp 1688980957
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_361
timestamp 1688980957
transform 1 0 34316 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_365
timestamp 1688980957
transform 1 0 34684 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_373
timestamp 1688980957
transform 1 0 35420 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_377
timestamp 1688980957
transform 1 0 35788 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_389
timestamp 1688980957
transform 1 0 36892 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_393
timestamp 1688980957
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_405
timestamp 1688980957
transform 1 0 38364 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_415
timestamp 1688980957
transform 1 0 39284 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_419
timestamp 1688980957
transform 1 0 39652 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_421
timestamp 1688980957
transform 1 0 39836 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_433
timestamp 1688980957
transform 1 0 40940 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 40388 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 9936 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 19412 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 36156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 23184 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 20608 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 33120 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 25300 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 27692 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform 1 0 20792 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 5336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 21988 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 3680 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform 1 0 20332 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform 1 0 7912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 4876 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform 1 0 12328 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform 1 0 4600 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform 1 0 12604 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform 1 0 26956 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 13248 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform 1 0 10396 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform 1 0 7084 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform 1 0 27600 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 6992 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform 1 0 9844 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform 1 0 3312 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform 1 0 22540 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform 1 0 7820 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform 1 0 19964 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform 1 0 6992 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform 1 0 14444 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform 1 0 3588 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform 1 0 14720 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform 1 0 34776 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform 1 0 5152 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input2
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input3
timestamp 1688980957
transform 1 0 38732 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1688980957
transform 1 0 40572 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input5
timestamp 1688980957
transform 1 0 31004 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1688980957
transform 1 0 9108 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input7
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1688980957
transform 1 0 40756 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 40848 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap1
timestamp 1688980957
transform 1 0 14628 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap2
timestamp 1688980957
transform 1 0 16560 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap19
timestamp 1688980957
transform 1 0 15548 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap20
timestamp 1688980957
transform 1 0 12052 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap21
timestamp 1688980957
transform 1 0 14352 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  max_cap22
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  max_cap24
timestamp 1688980957
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  max_cap26
timestamp 1688980957
transform 1 0 34040 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap27
timestamp 1688980957
transform 1 0 22080 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap30
timestamp 1688980957
transform 1 0 22632 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap32
timestamp 1688980957
transform 1 0 22724 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1688980957
transform 1 0 40756 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 1688980957
transform 1 0 21988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1688980957
transform 1 0 40756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 1688980957
transform 1 0 32936 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 1688980957
transform 1 0 7176 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1688980957
transform 1 0 40756 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1688980957
transform 1 0 34868 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 41400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 41400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 41400 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 41400 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 41400 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 41400 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 41400 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 41400 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 41400 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 41400 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 41400 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 41400 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 41400 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 41400 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 41400 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 41400 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 41400 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 41400 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 41400 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 41400 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 41400 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 41400 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 41400 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 41400 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 41400 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 41400 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 41400 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 41400 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 41400 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 41400 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 41400 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 41400 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 41400 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 41400 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 41400 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 41400 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 41400 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 41400 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 41400 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 41400 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 41400 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 41400 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 41400 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 41400 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 41400 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 41400 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 41400 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 41400 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 41400 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 41400 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 41400 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 41400 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 41400 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 41400 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 41400 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 41400 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 41400 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 41400 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 41400 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 41400 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 41400 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 41400 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 41400 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 41400 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 41400 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 41400 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 41400 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 41400 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 41400 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 41400 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 41400 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 41400 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 41400 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1688980957
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1688980957
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1688980957
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1688980957
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1688980957
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1688980957
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1688980957
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1688980957
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1688980957
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1688980957
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1688980957
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1688980957
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1688980957
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1688980957
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1688980957
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1688980957
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1688980957
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1688980957
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1688980957
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1688980957
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1688980957
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1688980957
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1688980957
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1688980957
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1688980957
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1688980957
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1688980957
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1688980957
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1688980957
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1688980957
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1688980957
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1688980957
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1688980957
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1688980957
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1688980957
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1688980957
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1688980957
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1688980957
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1688980957
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1688980957
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1688980957
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1688980957
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1688980957
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1688980957
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1688980957
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1688980957
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1688980957
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1688980957
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1688980957
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1688980957
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1688980957
transform 1 0 3680 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1688980957
transform 1 0 8832 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1688980957
transform 1 0 13984 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1688980957
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1688980957
transform 1 0 19136 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1688980957
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1688980957
transform 1 0 24288 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1688980957
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1688980957
transform 1 0 29440 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1688980957
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1688980957
transform 1 0 34592 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1688980957
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1688980957
transform 1 0 39744 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire23
timestamp 1688980957
transform 1 0 23000 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  wire25
timestamp 1688980957
transform 1 0 14996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  wire28
timestamp 1688980957
transform 1 0 23184 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  wire29
timestamp 1688980957
transform 1 0 28612 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  wire31
timestamp 1688980957
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  wire33
timestamp 1688980957
transform 1 0 28704 0 1 5440
box -38 -48 314 592
<< labels >>
flabel metal4 s 19568 2128 19888 42480 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 42480 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 34928 2128 35248 42480 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 41749 9528 42549 9648 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 41749 1368 42549 1488 0 FreeSans 480 0 0 0 cs
port 3 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 dataBusIn[0]
port 4 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 dataBusIn[1]
port 5 nsew signal input
flabel metal2 s 38658 43893 38714 44693 0 FreeSans 224 90 0 0 dataBusIn[2]
port 6 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 dataBusIn[3]
port 7 nsew signal input
flabel metal2 s 30930 43893 30986 44693 0 FreeSans 224 90 0 0 dataBusIn[4]
port 8 nsew signal input
flabel metal2 s 9034 43893 9090 44693 0 FreeSans 224 90 0 0 dataBusIn[5]
port 9 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 dataBusIn[6]
port 10 nsew signal input
flabel metal3 s 41749 5448 42549 5568 0 FreeSans 480 0 0 0 dataBusIn[7]
port 11 nsew signal input
flabel metal3 s 41749 36728 42549 36848 0 FreeSans 480 0 0 0 dataBusOut[0]
port 12 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 dataBusOut[1]
port 13 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 dataBusOut[2]
port 14 nsew signal tristate
flabel metal3 s 41749 32648 42549 32768 0 FreeSans 480 0 0 0 dataBusOut[3]
port 15 nsew signal tristate
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 dataBusOut[4]
port 16 nsew signal tristate
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 dataBusOut[5]
port 17 nsew signal tristate
flabel metal3 s 41749 40808 42549 40928 0 FreeSans 480 0 0 0 dataBusOut[6]
port 18 nsew signal tristate
flabel metal2 s 1306 43893 1362 44693 0 FreeSans 224 90 0 0 dataBusOut[7]
port 19 nsew signal tristate
flabel metal2 s 34794 43893 34850 44693 0 FreeSans 224 90 0 0 dataBusSelect
port 20 nsew signal tristate
flabel metal2 s 23846 43893 23902 44693 0 FreeSans 224 90 0 0 gpio[0]
port 21 nsew signal bidirectional
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 gpio[10]
port 22 nsew signal bidirectional
flabel metal2 s 19982 43893 20038 44693 0 FreeSans 224 90 0 0 gpio[11]
port 23 nsew signal bidirectional
flabel metal3 s 0 38768 800 38888 0 FreeSans 480 0 0 0 gpio[12]
port 24 nsew signal bidirectional
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 gpio[13]
port 25 nsew signal bidirectional
flabel metal2 s 5170 43893 5226 44693 0 FreeSans 224 90 0 0 gpio[14]
port 26 nsew signal bidirectional
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 gpio[15]
port 27 nsew signal bidirectional
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 gpio[16]
port 28 nsew signal bidirectional
flabel metal3 s 41749 29248 42549 29368 0 FreeSans 480 0 0 0 gpio[17]
port 29 nsew signal bidirectional
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 gpio[18]
port 30 nsew signal bidirectional
flabel metal3 s 41749 25168 42549 25288 0 FreeSans 480 0 0 0 gpio[19]
port 31 nsew signal bidirectional
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 gpio[1]
port 32 nsew signal bidirectional
flabel metal2 s 27710 43893 27766 44693 0 FreeSans 224 90 0 0 gpio[20]
port 33 nsew signal bidirectional
flabel metal3 s 41749 13608 42549 13728 0 FreeSans 480 0 0 0 gpio[21]
port 34 nsew signal bidirectional
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 gpio[22]
port 35 nsew signal bidirectional
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 gpio[23]
port 36 nsew signal bidirectional
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 gpio[24]
port 37 nsew signal bidirectional
flabel metal3 s 41749 17008 42549 17128 0 FreeSans 480 0 0 0 gpio[25]
port 38 nsew signal bidirectional
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 gpio[2]
port 39 nsew signal bidirectional
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 gpio[3]
port 40 nsew signal bidirectional
flabel metal2 s 41878 43893 41934 44693 0 FreeSans 224 90 0 0 gpio[4]
port 41 nsew signal bidirectional
flabel metal2 s 12898 43893 12954 44693 0 FreeSans 224 90 0 0 gpio[5]
port 42 nsew signal bidirectional
flabel metal2 s 16118 43893 16174 44693 0 FreeSans 224 90 0 0 gpio[6]
port 43 nsew signal bidirectional
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 gpio[7]
port 44 nsew signal bidirectional
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 gpio[8]
port 45 nsew signal bidirectional
flabel metal3 s 0 42848 800 42968 0 FreeSans 480 0 0 0 gpio[9]
port 46 nsew signal bidirectional
flabel metal3 s 41749 21088 42549 21208 0 FreeSans 480 0 0 0 nrst
port 47 nsew signal input
rlabel metal1 21252 42432 21252 42432 0 VGND
rlabel metal1 21252 41888 21252 41888 0 VPWR
rlabel metal1 32614 4658 32614 4658 0 _0000_
rlabel metal1 26949 6970 26949 6970 0 _0001_
rlabel metal1 27002 9010 27002 9010 0 _0002_
rlabel metal1 24472 7310 24472 7310 0 _0003_
rlabel metal1 26404 9418 26404 9418 0 _0004_
rlabel metal1 33580 5270 33580 5270 0 _0005_
rlabel metal1 26220 7922 26220 7922 0 _0006_
rlabel metal1 25576 6222 25576 6222 0 _0007_
rlabel metal1 29302 5134 29302 5134 0 _0008_
rlabel metal1 27738 10744 27738 10744 0 _0009_
rlabel metal1 24702 9146 24702 9146 0 _0010_
rlabel metal1 35420 5270 35420 5270 0 _0011_
rlabel metal2 30590 4386 30590 4386 0 _0012_
rlabel metal1 30084 37230 30084 37230 0 _0013_
rlabel metal1 23874 37774 23874 37774 0 _0014_
rlabel metal2 27922 37842 27922 37842 0 _0015_
rlabel metal1 26128 39066 26128 39066 0 _0016_
rlabel metal2 28198 36788 28198 36788 0 _0017_
rlabel metal2 25024 37366 25024 37366 0 _0018_
rlabel metal1 26910 37434 26910 37434 0 _0019_
rlabel metal1 39606 27642 39606 27642 0 _0020_
rlabel metal1 39744 30906 39744 30906 0 _0021_
rlabel metal1 39330 27064 39330 27064 0 _0022_
rlabel metal1 39744 29818 39744 29818 0 _0023_
rlabel metal1 39882 24378 39882 24378 0 _0024_
rlabel metal1 39744 25466 39744 25466 0 _0025_
rlabel metal1 19826 30906 19826 30906 0 _0026_
rlabel metal1 20102 11186 20102 11186 0 _0027_
rlabel metal1 22540 9554 22540 9554 0 _0028_
rlabel metal1 18722 8330 18722 8330 0 _0029_
rlabel metal1 21482 35122 21482 35122 0 _0030_
rlabel metal1 20700 7514 20700 7514 0 _0031_
rlabel metal1 18584 7446 18584 7446 0 _0032_
rlabel metal1 19964 9622 19964 9622 0 _0033_
rlabel metal1 22356 37298 22356 37298 0 _0034_
rlabel metal1 20332 5746 20332 5746 0 _0035_
rlabel metal1 2024 13498 2024 13498 0 _0036_
rlabel metal1 19632 33286 19632 33286 0 _0037_
rlabel metal1 18584 5270 18584 5270 0 _0038_
rlabel metal2 5566 6562 5566 6562 0 _0039_
rlabel metal1 23506 40120 23506 40120 0 _0040_
rlabel metal1 3266 38522 3266 38522 0 _0041_
rlabel metal1 10672 41650 10672 41650 0 _0042_
rlabel metal1 12788 38522 12788 38522 0 _0043_
rlabel metal1 9154 39066 9154 39066 0 _0044_
rlabel metal2 4738 38760 4738 38760 0 _0045_
rlabel metal1 5842 36686 5842 36686 0 _0046_
rlabel metal1 4232 35802 4232 35802 0 _0047_
rlabel metal2 7682 31450 7682 31450 0 _0048_
rlabel metal1 9476 31858 9476 31858 0 _0049_
rlabel metal2 7222 22372 7222 22372 0 _0050_
rlabel metal2 15042 25500 15042 25500 0 _0051_
rlabel metal1 6256 20978 6256 20978 0 _0052_
rlabel metal1 10580 18802 10580 18802 0 _0053_
rlabel metal1 4600 22202 4600 22202 0 _0054_
rlabel metal1 2806 21420 2806 21420 0 _0055_
rlabel metal1 1794 22746 1794 22746 0 _0056_
rlabel metal1 1787 21114 1787 21114 0 _0057_
rlabel metal1 8464 17238 8464 17238 0 _0058_
rlabel metal1 13478 17272 13478 17272 0 _0059_
rlabel metal2 7130 18496 7130 18496 0 _0060_
rlabel metal1 10396 17306 10396 17306 0 _0061_
rlabel metal1 4554 17544 4554 17544 0 _0062_
rlabel metal1 3496 19414 3496 19414 0 _0063_
rlabel metal1 1794 19482 1794 19482 0 _0064_
rlabel metal1 1794 17306 1794 17306 0 _0065_
rlabel metal2 22126 9588 22126 9588 0 _0066_
rlabel metal1 1794 28118 1794 28118 0 _0067_
rlabel metal1 1886 40698 1886 40698 0 _0068_
rlabel metal1 2208 28594 2208 28594 0 _0069_
rlabel metal2 19642 41820 19642 41820 0 _0070_
rlabel metal1 2208 36346 2208 36346 0 _0071_
rlabel metal1 1748 30770 1748 30770 0 _0072_
rlabel metal1 4186 40698 4186 40698 0 _0073_
rlabel metal2 2806 31518 2806 31518 0 _0074_
rlabel metal1 19366 40154 19366 40154 0 _0075_
rlabel metal1 16836 33898 16836 33898 0 _0076_
rlabel metal1 19642 36346 19642 36346 0 _0077_
rlabel metal1 18308 38998 18308 38998 0 _0078_
rlabel metal1 14812 34442 14812 34442 0 _0079_
rlabel metal1 12282 36686 12282 36686 0 _0080_
rlabel metal1 13340 39610 13340 39610 0 _0081_
rlabel metal1 17243 41786 17243 41786 0 _0082_
rlabel metal1 8510 19414 8510 19414 0 _0083_
rlabel metal1 13478 20026 13478 20026 0 _0084_
rlabel metal1 6348 24718 6348 24718 0 _0085_
rlabel metal2 12558 20060 12558 20060 0 _0086_
rlabel metal1 3910 25466 3910 25466 0 _0087_
rlabel metal1 1978 26554 1978 26554 0 _0088_
rlabel metal1 1794 24922 1794 24922 0 _0089_
rlabel metal1 2714 23800 2714 23800 0 _0090_
rlabel metal1 22034 41038 22034 41038 0 _0091_
rlabel metal1 21482 5576 21482 5576 0 _0092_
rlabel metal2 16698 5440 16698 5440 0 _0093_
rlabel metal2 11822 31076 11822 31076 0 _0094_
rlabel metal2 22494 41106 22494 41106 0 _0095_
rlabel metal1 12236 41242 12236 41242 0 _0096_
rlabel metal1 14352 41242 14352 41242 0 _0097_
rlabel metal1 21896 6698 21896 6698 0 _0098_
rlabel metal1 13662 11866 13662 11866 0 _0099_
rlabel metal1 15722 6970 15722 6970 0 _0100_
rlabel metal1 9522 5338 9522 5338 0 _0101_
rlabel metal1 11822 5304 11822 5304 0 _0102_
rlabel metal1 8510 6222 8510 6222 0 _0103_
rlabel metal1 5329 9146 5329 9146 0 _0104_
rlabel metal1 4232 13498 4232 13498 0 _0105_
rlabel metal1 6854 14042 6854 14042 0 _0106_
rlabel metal1 8418 15674 8418 15674 0 _0107_
rlabel metal1 14398 16456 14398 16456 0 _0108_
rlabel metal1 6624 16626 6624 16626 0 _0109_
rlabel metal1 10764 16626 10764 16626 0 _0110_
rlabel metal1 5191 15674 5191 15674 0 _0111_
rlabel metal1 3910 15674 3910 15674 0 _0112_
rlabel metal1 1886 15096 1886 15096 0 _0113_
rlabel metal1 2116 16626 2116 16626 0 _0114_
rlabel metal1 17434 30906 17434 30906 0 _0115_
rlabel metal1 26772 4658 26772 4658 0 _0116_
rlabel via1 17243 20026 17243 20026 0 _0117_
rlabel metal1 18768 24922 18768 24922 0 _0118_
rlabel metal1 17986 24174 17986 24174 0 _0119_
rlabel metal2 24978 24752 24978 24752 0 _0120_
rlabel metal1 20148 24718 20148 24718 0 _0121_
rlabel metal1 18492 24650 18492 24650 0 _0122_
rlabel metal1 18032 24242 18032 24242 0 _0123_
rlabel metal1 18446 23766 18446 23766 0 _0124_
rlabel metal1 9246 21590 9246 21590 0 _0125_
rlabel metal2 18078 22039 18078 22039 0 _0126_
rlabel metal1 13156 24922 13156 24922 0 _0127_
rlabel metal1 17204 24242 17204 24242 0 _0128_
rlabel metal2 17434 23137 17434 23137 0 _0129_
rlabel via1 17411 22610 17411 22610 0 _0130_
rlabel metal1 18032 23018 18032 23018 0 _0131_
rlabel metal1 18078 22610 18078 22610 0 _0132_
rlabel metal1 9844 23630 9844 23630 0 _0133_
rlabel metal1 11270 33966 11270 33966 0 _0134_
rlabel metal1 10856 14246 10856 14246 0 _0135_
rlabel metal1 21206 21556 21206 21556 0 _0136_
rlabel metal1 17020 16082 17020 16082 0 _0137_
rlabel metal1 17480 15402 17480 15402 0 _0138_
rlabel metal1 14950 15062 14950 15062 0 _0139_
rlabel metal1 8878 13906 8878 13906 0 _0140_
rlabel metal2 9062 12512 9062 12512 0 _0141_
rlabel metal1 5014 19856 5014 19856 0 _0142_
rlabel metal1 5244 19958 5244 19958 0 _0143_
rlabel metal1 4784 24582 4784 24582 0 _0144_
rlabel metal1 5980 26282 5980 26282 0 _0145_
rlabel metal2 6578 29614 6578 29614 0 _0146_
rlabel metal1 6808 27030 6808 27030 0 _0147_
rlabel metal1 8694 26554 8694 26554 0 _0148_
rlabel metal1 8510 27098 8510 27098 0 _0149_
rlabel metal1 6992 27098 6992 27098 0 _0150_
rlabel metal1 4830 16592 4830 16592 0 _0151_
rlabel metal1 9154 15334 9154 15334 0 _0152_
rlabel metal1 13294 17068 13294 17068 0 _0153_
rlabel metal1 10626 10506 10626 10506 0 _0154_
rlabel metal1 10212 10642 10212 10642 0 _0155_
rlabel metal1 9660 21658 9660 21658 0 _0156_
rlabel metal1 10028 22066 10028 22066 0 _0157_
rlabel metal1 12190 30736 12190 30736 0 _0158_
rlabel metal1 12604 36142 12604 36142 0 _0159_
rlabel metal1 10258 10506 10258 10506 0 _0160_
rlabel metal1 9798 10030 9798 10030 0 _0161_
rlabel metal1 6716 18938 6716 18938 0 _0162_
rlabel metal1 7636 23290 7636 23290 0 _0163_
rlabel metal1 7590 23766 7590 23766 0 _0164_
rlabel metal1 9338 23800 9338 23800 0 _0165_
rlabel metal1 7452 24106 7452 24106 0 _0166_
rlabel metal1 7498 29172 7498 29172 0 _0167_
rlabel metal1 7820 28594 7820 28594 0 _0168_
rlabel metal1 20010 21930 20010 21930 0 _0169_
rlabel metal1 19596 22066 19596 22066 0 _0170_
rlabel metal2 16698 26707 16698 26707 0 _0171_
rlabel metal1 7866 26928 7866 26928 0 _0172_
rlabel metal1 7590 26758 7590 26758 0 _0173_
rlabel metal1 5980 16014 5980 16014 0 _0174_
rlabel metal2 8832 13226 8832 13226 0 _0175_
rlabel metal1 18400 6358 18400 6358 0 _0176_
rlabel metal1 11592 10778 11592 10778 0 _0177_
rlabel metal1 9798 23086 9798 23086 0 _0178_
rlabel metal2 11776 28356 11776 28356 0 _0179_
rlabel metal2 22494 39440 22494 39440 0 _0180_
rlabel metal1 9430 10064 9430 10064 0 _0181_
rlabel metal1 9246 8908 9246 8908 0 _0182_
rlabel metal1 13570 24616 13570 24616 0 _0183_
rlabel metal1 14260 26894 14260 26894 0 _0184_
rlabel metal1 13478 27404 13478 27404 0 _0185_
rlabel metal1 13892 26962 13892 26962 0 _0186_
rlabel via1 12742 18819 12742 18819 0 _0187_
rlabel metal1 12788 18938 12788 18938 0 _0188_
rlabel metal2 13018 23868 13018 23868 0 _0189_
rlabel metal2 14122 26384 14122 26384 0 _0190_
rlabel metal1 13432 29274 13432 29274 0 _0191_
rlabel metal2 13294 27370 13294 27370 0 _0192_
rlabel metal2 12558 15827 12558 15827 0 _0193_
rlabel metal1 12834 10608 12834 10608 0 _0194_
rlabel metal2 12190 9418 12190 9418 0 _0195_
rlabel metal3 17963 32300 17963 32300 0 _0196_
rlabel metal1 12328 15130 12328 15130 0 _0197_
rlabel metal1 12742 21930 12742 21930 0 _0198_
rlabel metal1 13432 21998 13432 21998 0 _0199_
rlabel metal1 13478 21556 13478 21556 0 _0200_
rlabel metal1 12926 15062 12926 15062 0 _0201_
rlabel via2 11270 9027 11270 9027 0 _0202_
rlabel metal1 11592 8942 11592 8942 0 _0203_
rlabel metal1 12466 7446 12466 7446 0 _0204_
rlabel metal2 9522 25602 9522 25602 0 _0205_
rlabel metal2 9890 27268 9890 27268 0 _0206_
rlabel metal1 10488 27642 10488 27642 0 _0207_
rlabel via1 10810 25347 10810 25347 0 _0208_
rlabel metal1 7774 19856 7774 19856 0 _0209_
rlabel metal1 8372 20026 8372 20026 0 _0210_
rlabel metal1 8832 24378 8832 24378 0 _0211_
rlabel metal1 11454 25228 11454 25228 0 _0212_
rlabel metal1 10120 29478 10120 29478 0 _0213_
rlabel metal2 10534 26826 10534 26826 0 _0214_
rlabel metal1 7498 19346 7498 19346 0 _0215_
rlabel metal2 13846 9350 13846 9350 0 _0216_
rlabel metal2 15594 14722 15594 14722 0 _0217_
rlabel metal1 14950 14892 14950 14892 0 _0218_
rlabel metal2 17986 21760 17986 21760 0 _0219_
rlabel metal2 10856 21998 10856 21998 0 _0220_
rlabel metal1 16238 21522 16238 21522 0 _0221_
rlabel metal1 14858 14994 14858 14994 0 _0222_
rlabel metal1 14306 9554 14306 9554 0 _0223_
rlabel metal1 13800 8466 13800 8466 0 _0224_
rlabel metal1 12006 24242 12006 24242 0 _0225_
rlabel metal1 9706 19754 9706 19754 0 _0226_
rlabel metal1 10120 19958 10120 19958 0 _0227_
rlabel metal1 11592 24582 11592 24582 0 _0228_
rlabel metal1 11684 24922 11684 24922 0 _0229_
rlabel metal1 16284 28730 16284 28730 0 _0230_
rlabel metal1 12466 28084 12466 28084 0 _0231_
rlabel metal1 12190 28730 12190 28730 0 _0232_
rlabel metal2 12190 26554 12190 26554 0 _0233_
rlabel metal1 11132 26010 11132 26010 0 _0234_
rlabel metal2 11914 26724 11914 26724 0 _0235_
rlabel metal1 12466 26452 12466 26452 0 _0236_
rlabel metal2 13570 16864 13570 16864 0 _0237_
rlabel metal1 10810 14416 10810 14416 0 _0238_
rlabel metal1 15410 14416 15410 14416 0 _0239_
rlabel metal1 14674 22576 14674 22576 0 _0240_
rlabel metal2 14030 21998 14030 21998 0 _0241_
rlabel metal2 14766 22406 14766 22406 0 _0242_
rlabel metal1 14904 14586 14904 14586 0 _0243_
rlabel metal1 14720 14246 14720 14246 0 _0244_
rlabel metal1 13064 24310 13064 24310 0 _0245_
rlabel metal1 13064 15470 13064 15470 0 _0246_
rlabel metal1 13662 15504 13662 15504 0 _0247_
rlabel metal1 14398 14382 14398 14382 0 _0248_
rlabel metal1 15686 12852 15686 12852 0 _0249_
rlabel metal2 28566 16932 28566 16932 0 _0250_
rlabel metal1 29072 17850 29072 17850 0 _0251_
rlabel metal1 27968 17850 27968 17850 0 _0252_
rlabel metal2 27738 18428 27738 18428 0 _0253_
rlabel metal1 27784 17306 27784 17306 0 _0254_
rlabel metal1 24426 17204 24426 17204 0 _0255_
rlabel metal1 25392 16218 25392 16218 0 _0256_
rlabel metal1 25116 16762 25116 16762 0 _0257_
rlabel metal1 15502 12818 15502 12818 0 _0258_
rlabel metal1 14766 13498 14766 13498 0 _0259_
rlabel metal1 15134 12614 15134 12614 0 _0260_
rlabel metal1 15088 24582 15088 24582 0 _0261_
rlabel metal2 15778 27268 15778 27268 0 _0262_
rlabel metal2 15134 28764 15134 28764 0 _0263_
rlabel metal1 15088 28594 15088 28594 0 _0264_
rlabel metal1 15042 19210 15042 19210 0 _0265_
rlabel metal1 15548 22678 15548 22678 0 _0266_
rlabel metal1 14490 23188 14490 23188 0 _0267_
rlabel metal1 14720 26962 14720 26962 0 _0268_
rlabel metal1 14812 29546 14812 29546 0 _0269_
rlabel metal1 14674 28492 14674 28492 0 _0270_
rlabel metal1 14490 18326 14490 18326 0 _0271_
rlabel via1 15975 12818 15975 12818 0 _0272_
rlabel viali 16426 26962 16426 26962 0 _0273_
rlabel metal2 17250 17153 17250 17153 0 _0274_
rlabel metal1 16606 10642 16606 10642 0 _0275_
rlabel metal1 18354 21658 18354 21658 0 _0276_
rlabel metal1 16790 22610 16790 22610 0 _0277_
rlabel metal1 17480 22406 17480 22406 0 _0278_
rlabel metal4 17664 20060 17664 20060 0 _0279_
rlabel metal1 16146 9996 16146 9996 0 _0280_
rlabel metal1 15962 9010 15962 9010 0 _0281_
rlabel metal1 16790 10064 16790 10064 0 _0282_
rlabel metal1 16606 8942 16606 8942 0 _0283_
rlabel metal2 13570 8772 13570 8772 0 _0284_
rlabel metal1 14214 8942 14214 8942 0 _0285_
rlabel metal1 12926 7854 12926 7854 0 _0286_
rlabel metal1 12006 7820 12006 7820 0 _0287_
rlabel metal1 9246 7412 9246 7412 0 _0288_
rlabel metal1 14122 6256 14122 6256 0 _0289_
rlabel metal2 16330 7786 16330 7786 0 _0290_
rlabel metal1 12926 6970 12926 6970 0 _0291_
rlabel metal1 8602 7378 8602 7378 0 _0292_
rlabel metal1 9062 9588 9062 9588 0 _0293_
rlabel metal1 8878 8432 8878 8432 0 _0294_
rlabel metal1 9200 8262 9200 8262 0 _0295_
rlabel metal1 7222 8942 7222 8942 0 _0296_
rlabel metal1 9154 10234 9154 10234 0 _0297_
rlabel metal1 9154 10574 9154 10574 0 _0298_
rlabel metal1 8602 10574 8602 10574 0 _0299_
rlabel metal1 6854 9554 6854 9554 0 _0300_
rlabel metal1 9154 13328 9154 13328 0 _0301_
rlabel viali 8878 12817 8878 12817 0 _0302_
rlabel metal1 8652 12818 8652 12818 0 _0303_
rlabel metal1 6670 12852 6670 12852 0 _0304_
rlabel metal1 4922 19380 4922 19380 0 _0305_
rlabel metal1 5428 23766 5428 23766 0 _0306_
rlabel metal1 5244 24174 5244 24174 0 _0307_
rlabel metal1 5060 27370 5060 27370 0 _0308_
rlabel metal2 6486 29818 6486 29818 0 _0309_
rlabel metal2 5750 28560 5750 28560 0 _0310_
rlabel metal1 9890 25466 9890 25466 0 _0311_
rlabel metal1 10350 27098 10350 27098 0 _0312_
rlabel metal1 7130 28118 7130 28118 0 _0313_
rlabel metal1 3634 17238 3634 17238 0 _0314_
rlabel metal1 9246 13906 9246 13906 0 _0315_
rlabel metal1 16284 17170 16284 17170 0 _0316_
rlabel metal1 10488 15130 10488 15130 0 _0317_
rlabel metal2 9706 21692 9706 21692 0 _0318_
rlabel metal1 11132 21658 11132 21658 0 _0319_
rlabel via2 16514 35037 16514 35037 0 _0320_
rlabel metal2 9430 14348 9430 14348 0 _0321_
rlabel metal1 7958 13974 7958 13974 0 _0322_
rlabel metal1 7820 13906 7820 13906 0 _0323_
rlabel metal1 10672 12818 10672 12818 0 _0324_
rlabel metal1 6578 12614 6578 12614 0 _0325_
rlabel metal1 7038 11730 7038 11730 0 _0326_
rlabel metal1 6302 11084 6302 11084 0 _0327_
rlabel metal2 6578 9350 6578 9350 0 _0328_
rlabel metal1 5244 9962 5244 9962 0 _0329_
rlabel metal1 5612 11322 5612 11322 0 _0330_
rlabel metal1 4278 12070 4278 12070 0 _0331_
rlabel metal1 7084 12818 7084 12818 0 _0332_
rlabel metal2 6762 12988 6762 12988 0 _0333_
rlabel metal1 8234 12682 8234 12682 0 _0334_
rlabel metal1 8007 7854 8007 7854 0 _0335_
rlabel metal1 7774 11084 7774 11084 0 _0336_
rlabel viali 8050 11729 8050 11729 0 _0337_
rlabel metal1 11270 13294 11270 13294 0 _0338_
rlabel metal1 12926 13838 12926 13838 0 _0339_
rlabel metal1 16790 12852 16790 12852 0 _0340_
rlabel metal2 14214 9452 14214 9452 0 _0341_
rlabel metal2 21206 14246 21206 14246 0 _0342_
rlabel metal1 21712 14994 21712 14994 0 _0343_
rlabel metal2 24242 21862 24242 21862 0 _0344_
rlabel metal1 24242 21522 24242 21522 0 _0345_
rlabel metal2 24150 15793 24150 15793 0 _0346_
rlabel metal1 24058 15028 24058 15028 0 _0347_
rlabel metal1 23966 14858 23966 14858 0 _0348_
rlabel metal1 23276 14382 23276 14382 0 _0349_
rlabel metal2 20838 12823 20838 12823 0 _0350_
rlabel metal2 8142 7956 8142 7956 0 _0351_
rlabel metal1 12236 12818 12236 12818 0 _0352_
rlabel metal1 22402 14314 22402 14314 0 _0353_
rlabel metal2 16146 12971 16146 12971 0 _0354_
rlabel metal1 15732 11050 15732 11050 0 _0355_
rlabel metal2 12098 12801 12098 12801 0 _0356_
rlabel metal2 18998 21828 18998 21828 0 _0357_
rlabel metal2 17986 18122 17986 18122 0 _0358_
rlabel metal1 20562 18734 20562 18734 0 _0359_
rlabel metal1 18676 18394 18676 18394 0 _0360_
rlabel metal1 17618 15470 17618 15470 0 _0361_
rlabel metal1 19504 17850 19504 17850 0 _0362_
rlabel metal1 18262 15368 18262 15368 0 _0363_
rlabel metal1 18492 16218 18492 16218 0 _0364_
rlabel metal1 20608 18190 20608 18190 0 _0365_
rlabel metal2 17802 17765 17802 17765 0 _0366_
rlabel metal1 18768 17646 18768 17646 0 _0367_
rlabel metal1 18400 18054 18400 18054 0 _0368_
rlabel metal1 29578 26350 29578 26350 0 _0369_
rlabel metal1 29624 25466 29624 25466 0 _0370_
rlabel metal1 29118 26350 29118 26350 0 _0371_
rlabel metal1 29486 26282 29486 26282 0 _0372_
rlabel metal2 19734 20145 19734 20145 0 _0373_
rlabel metal1 16882 18156 16882 18156 0 _0374_
rlabel metal1 16514 18224 16514 18224 0 _0375_
rlabel metal2 16330 17782 16330 17782 0 _0376_
rlabel metal1 16836 17306 16836 17306 0 _0377_
rlabel metal1 16928 16966 16928 16966 0 _0378_
rlabel metal1 20424 20230 20424 20230 0 _0379_
rlabel metal1 18768 12682 18768 12682 0 _0380_
rlabel metal1 19228 12750 19228 12750 0 _0381_
rlabel metal1 17618 12784 17618 12784 0 _0382_
rlabel metal1 18538 16082 18538 16082 0 _0383_
rlabel metal1 18367 15470 18367 15470 0 _0384_
rlabel metal1 17066 15436 17066 15436 0 _0385_
rlabel metal1 19633 14960 19633 14960 0 _0386_
rlabel metal2 20562 14586 20562 14586 0 _0387_
rlabel metal1 19872 14518 19872 14518 0 _0388_
rlabel metal1 20125 15062 20125 15062 0 _0389_
rlabel metal1 18906 13940 18906 13940 0 _0390_
rlabel metal1 18906 13736 18906 13736 0 _0391_
rlabel metal1 12926 13430 12926 13430 0 _0392_
rlabel metal1 18538 13974 18538 13974 0 _0393_
rlabel metal2 18998 13124 18998 13124 0 _0394_
rlabel via2 1886 34595 1886 34595 0 _0395_
rlabel metal1 20378 30634 20378 30634 0 _0396_
rlabel metal1 19596 30634 19596 30634 0 _0397_
rlabel metal1 22034 15504 22034 15504 0 _0398_
rlabel metal2 21574 13804 21574 13804 0 _0399_
rlabel metal1 20930 11798 20930 11798 0 _0400_
rlabel metal2 22402 10676 22402 10676 0 _0401_
rlabel metal1 20194 9078 20194 9078 0 _0402_
rlabel metal1 19458 8534 19458 8534 0 _0403_
rlabel metal1 21712 7174 21712 7174 0 _0404_
rlabel metal1 19918 10642 19918 10642 0 _0405_
rlabel metal1 19090 7718 19090 7718 0 _0406_
rlabel metal1 19734 10234 19734 10234 0 _0407_
rlabel metal1 25898 23834 25898 23834 0 _0408_
rlabel metal1 22494 24378 22494 24378 0 _0409_
rlabel via1 23882 24038 23882 24038 0 _0410_
rlabel metal1 23598 24174 23598 24174 0 _0411_
rlabel metal2 19642 36448 19642 36448 0 _0412_
rlabel metal1 22448 36890 22448 36890 0 _0413_
rlabel metal1 21068 6290 21068 6290 0 _0414_
rlabel metal2 2806 13770 2806 13770 0 _0415_
rlabel metal2 19550 33286 19550 33286 0 _0416_
rlabel metal1 18906 6426 18906 6426 0 _0417_
rlabel metal1 6072 6290 6072 6290 0 _0418_
rlabel metal1 23092 39610 23092 39610 0 _0419_
rlabel metal1 3726 38318 3726 38318 0 _0420_
rlabel metal1 23966 29614 23966 29614 0 _0421_
rlabel metal2 22034 30498 22034 30498 0 _0422_
rlabel metal1 21850 30736 21850 30736 0 _0423_
rlabel metal1 17802 32878 17802 32878 0 _0424_
rlabel metal1 17802 35462 17802 35462 0 _0425_
rlabel metal1 19228 16422 19228 16422 0 _0426_
rlabel metal1 15594 33626 15594 33626 0 _0427_
rlabel metal2 32062 26639 32062 26639 0 _0428_
rlabel metal1 24012 31994 24012 31994 0 _0429_
rlabel metal2 24426 31620 24426 31620 0 _0430_
rlabel metal1 25484 35734 25484 35734 0 _0431_
rlabel metal1 24472 34510 24472 34510 0 _0432_
rlabel metal1 26956 31314 26956 31314 0 _0433_
rlabel metal1 24564 34170 24564 34170 0 _0434_
rlabel metal1 24196 34034 24196 34034 0 _0435_
rlabel metal1 23506 33898 23506 33898 0 _0436_
rlabel metal2 24242 33150 24242 33150 0 _0437_
rlabel metal1 23736 32538 23736 32538 0 _0438_
rlabel metal2 23690 29002 23690 29002 0 _0439_
rlabel metal2 23506 28832 23506 28832 0 _0440_
rlabel metal2 23598 31892 23598 31892 0 _0441_
rlabel metal2 20470 33626 20470 33626 0 _0442_
rlabel metal2 17342 33184 17342 33184 0 _0443_
rlabel metal1 17572 38862 17572 38862 0 _0444_
rlabel via1 13296 39406 13296 39406 0 _0445_
rlabel metal2 12374 29342 12374 29342 0 _0446_
rlabel metal1 6877 29614 6877 29614 0 _0447_
rlabel metal1 6716 29546 6716 29546 0 _0448_
rlabel metal2 12374 27370 12374 27370 0 _0449_
rlabel metal1 11086 28118 11086 28118 0 _0450_
rlabel metal1 4508 29546 4508 29546 0 _0451_
rlabel metal1 12604 28186 12604 28186 0 _0452_
rlabel metal2 4554 29495 4554 29495 0 _0453_
rlabel metal2 20654 35190 20654 35190 0 _0454_
rlabel metal1 19366 36686 19366 36686 0 _0455_
rlabel metal1 14260 40494 14260 40494 0 _0456_
rlabel metal1 11040 37978 11040 37978 0 _0457_
rlabel metal1 6394 37876 6394 37876 0 _0458_
rlabel metal1 8418 32300 8418 32300 0 _0459_
rlabel metal1 16054 32334 16054 32334 0 _0460_
rlabel metal1 13340 32198 13340 32198 0 _0461_
rlabel metal1 12788 33490 12788 33490 0 _0462_
rlabel metal1 12558 34578 12558 34578 0 _0463_
rlabel metal1 11684 34170 11684 34170 0 _0464_
rlabel metal1 10856 35666 10856 35666 0 _0465_
rlabel metal1 16928 5202 16928 5202 0 _0466_
rlabel metal1 16100 31790 16100 31790 0 _0467_
rlabel metal1 14904 32402 14904 32402 0 _0468_
rlabel metal2 14858 33014 14858 33014 0 _0469_
rlabel metal1 11960 33490 11960 33490 0 _0470_
rlabel metal1 11592 34714 11592 34714 0 _0471_
rlabel metal1 16422 37264 16422 37264 0 _0472_
rlabel metal1 10258 34986 10258 34986 0 _0473_
rlabel metal2 10810 36516 10810 36516 0 _0474_
rlabel metal1 10534 36890 10534 36890 0 _0475_
rlabel metal1 8050 34000 8050 34000 0 _0476_
rlabel metal1 7590 36176 7590 36176 0 _0477_
rlabel metal1 11776 39950 11776 39950 0 _0478_
rlabel metal1 11178 40052 11178 40052 0 _0479_
rlabel via2 10810 40035 10810 40035 0 _0480_
rlabel metal2 15502 39712 15502 39712 0 _0481_
rlabel metal2 14904 40494 14904 40494 0 _0482_
rlabel metal1 14582 40528 14582 40528 0 _0483_
rlabel metal1 15272 40494 15272 40494 0 _0484_
rlabel metal1 16146 36754 16146 36754 0 _0485_
rlabel metal1 15502 37264 15502 37264 0 _0486_
rlabel metal1 17158 36652 17158 36652 0 _0487_
rlabel metal2 19274 37570 19274 37570 0 _0488_
rlabel metal1 18400 37162 18400 37162 0 _0489_
rlabel metal1 20194 34476 20194 34476 0 _0490_
rlabel metal1 19550 34578 19550 34578 0 _0491_
rlabel metal1 18814 36108 18814 36108 0 _0492_
rlabel metal1 18998 37264 18998 37264 0 _0493_
rlabel metal1 19366 37910 19366 37910 0 _0494_
rlabel metal1 17250 36788 17250 36788 0 _0495_
rlabel metal1 16790 36210 16790 36210 0 _0496_
rlabel metal1 15042 37196 15042 37196 0 _0497_
rlabel metal1 15364 39338 15364 39338 0 _0498_
rlabel metal1 15778 40052 15778 40052 0 _0499_
rlabel metal1 12420 39406 12420 39406 0 _0500_
rlabel via1 10179 40086 10179 40086 0 _0501_
rlabel metal1 10166 39814 10166 39814 0 _0502_
rlabel metal1 16192 36142 16192 36142 0 _0503_
rlabel via1 10534 40171 10534 40171 0 _0504_
rlabel metal1 11362 37434 11362 37434 0 _0505_
rlabel metal1 11454 38454 11454 38454 0 _0506_
rlabel metal1 11546 38522 11546 38522 0 _0507_
rlabel metal1 11822 38964 11822 38964 0 _0508_
rlabel metal2 12282 38522 12282 38522 0 _0509_
rlabel metal1 14030 29274 14030 29274 0 _0510_
rlabel metal1 9522 33388 9522 33388 0 _0511_
rlabel metal1 10534 35462 10534 35462 0 _0512_
rlabel metal1 10350 36176 10350 36176 0 _0513_
rlabel metal1 10120 36346 10120 36346 0 _0514_
rlabel metal1 10902 37434 10902 37434 0 _0515_
rlabel metal1 11822 37978 11822 37978 0 _0516_
rlabel metal1 9706 29172 9706 29172 0 _0517_
rlabel metal2 10074 34357 10074 34357 0 _0518_
rlabel metal1 9844 35258 9844 35258 0 _0519_
rlabel metal1 9798 33626 9798 33626 0 _0520_
rlabel metal2 9798 34544 9798 34544 0 _0521_
rlabel metal1 9982 35156 9982 35156 0 _0522_
rlabel metal1 8740 35258 8740 35258 0 _0523_
rlabel metal1 7360 39474 7360 39474 0 _0524_
rlabel metal2 11270 39236 11270 39236 0 _0525_
rlabel metal2 8510 39746 8510 39746 0 _0526_
rlabel metal1 7406 39270 7406 39270 0 _0527_
rlabel metal1 8188 39338 8188 39338 0 _0528_
rlabel metal1 8418 38998 8418 38998 0 _0529_
rlabel metal1 6854 38318 6854 38318 0 _0530_
rlabel metal1 6670 37230 6670 37230 0 _0531_
rlabel metal1 6808 38726 6808 38726 0 _0532_
rlabel metal1 7544 38386 7544 38386 0 _0533_
rlabel metal1 6992 38386 6992 38386 0 _0534_
rlabel metal2 13202 29665 13202 29665 0 _0535_
rlabel metal1 17986 40902 17986 40902 0 _0536_
rlabel metal1 12995 32538 12995 32538 0 _0537_
rlabel metal1 12052 32538 12052 32538 0 _0538_
rlabel metal1 14720 31858 14720 31858 0 _0539_
rlabel metal1 11730 33014 11730 33014 0 _0540_
rlabel metal1 10120 34578 10120 34578 0 _0541_
rlabel metal1 9614 34612 9614 34612 0 _0542_
rlabel metal2 9706 36244 9706 36244 0 _0543_
rlabel metal1 9338 37842 9338 37842 0 _0544_
rlabel metal1 9476 37978 9476 37978 0 _0545_
rlabel metal1 6302 38250 6302 38250 0 _0546_
rlabel metal1 5106 38318 5106 38318 0 _0547_
rlabel metal2 6946 36448 6946 36448 0 _0548_
rlabel metal1 6808 37434 6808 37434 0 _0549_
rlabel via1 7314 36754 7314 36754 0 _0550_
rlabel metal2 7222 36890 7222 36890 0 _0551_
rlabel metal1 9108 29070 9108 29070 0 _0552_
rlabel metal1 7130 35054 7130 35054 0 _0553_
rlabel metal1 7314 35122 7314 35122 0 _0554_
rlabel metal1 7498 35258 7498 35258 0 _0555_
rlabel metal1 7866 36346 7866 36346 0 _0556_
rlabel metal1 6900 33966 6900 33966 0 _0557_
rlabel metal1 7498 34034 7498 34034 0 _0558_
rlabel metal1 6670 35666 6670 35666 0 _0559_
rlabel metal2 7038 34221 7038 34221 0 _0560_
rlabel metal1 6118 33354 6118 33354 0 _0561_
rlabel metal1 5566 33966 5566 33966 0 _0562_
rlabel metal1 4554 33898 4554 33898 0 _0563_
rlabel metal1 4830 33830 4830 33830 0 _0564_
rlabel metal1 5014 29274 5014 29274 0 _0565_
rlabel metal1 4462 29818 4462 29818 0 _0566_
rlabel metal1 6072 33966 6072 33966 0 _0567_
rlabel metal2 5750 34017 5750 34017 0 _0568_
rlabel metal1 5152 34170 5152 34170 0 _0569_
rlabel metal1 4600 35666 4600 35666 0 _0570_
rlabel metal1 7130 32538 7130 32538 0 _0571_
rlabel metal2 7222 33354 7222 33354 0 _0572_
rlabel metal1 7130 31654 7130 31654 0 _0573_
rlabel metal1 4738 33388 4738 33388 0 _0574_
rlabel metal1 4462 33558 4462 33558 0 _0575_
rlabel metal1 4922 32402 4922 32402 0 _0576_
rlabel metal1 5428 28730 5428 28730 0 _0577_
rlabel metal1 4876 31858 4876 31858 0 _0578_
rlabel metal1 5612 31994 5612 31994 0 _0579_
rlabel metal1 7038 31824 7038 31824 0 _0580_
rlabel metal1 7820 32538 7820 32538 0 _0581_
rlabel metal1 8740 31246 8740 31246 0 _0582_
rlabel metal1 9614 31246 9614 31246 0 _0583_
rlabel metal1 9844 32470 9844 32470 0 _0584_
rlabel metal1 5382 31926 5382 31926 0 _0585_
rlabel metal1 6118 29648 6118 29648 0 _0586_
rlabel metal1 5934 31110 5934 31110 0 _0587_
rlabel metal1 6118 31892 6118 31892 0 _0588_
rlabel metal1 5750 31178 5750 31178 0 _0589_
rlabel metal1 8280 32402 8280 32402 0 _0590_
rlabel metal2 28382 28288 28382 28288 0 _0591_
rlabel metal2 16974 26979 16974 26979 0 _0592_
rlabel metal1 14674 21046 14674 21046 0 _0593_
rlabel metal1 7912 21998 7912 21998 0 _0594_
rlabel metal1 15180 24922 15180 24922 0 _0595_
rlabel metal1 6670 21522 6670 21522 0 _0596_
rlabel metal1 10810 20468 10810 20468 0 _0597_
rlabel metal1 4784 21862 4784 21862 0 _0598_
rlabel metal1 2622 21556 2622 21556 0 _0599_
rlabel metal1 2300 22610 2300 22610 0 _0600_
rlabel metal1 2300 21522 2300 21522 0 _0601_
rlabel metal1 30590 19448 30590 19448 0 _0602_
rlabel metal1 17158 18768 17158 18768 0 _0603_
rlabel metal1 16928 18666 16928 18666 0 _0604_
rlabel metal1 7498 19210 7498 19210 0 _0605_
rlabel metal2 8786 17850 8786 17850 0 _0606_
rlabel metal1 14214 17646 14214 17646 0 _0607_
rlabel metal1 7130 18258 7130 18258 0 _0608_
rlabel metal1 10718 17136 10718 17136 0 _0609_
rlabel metal1 4968 18258 4968 18258 0 _0610_
rlabel metal1 3910 18938 3910 18938 0 _0611_
rlabel metal1 2162 19346 2162 19346 0 _0612_
rlabel metal1 2070 17204 2070 17204 0 _0613_
rlabel metal1 25530 23494 25530 23494 0 _0614_
rlabel metal1 25300 19482 25300 19482 0 _0615_
rlabel metal1 25162 20026 25162 20026 0 _0616_
rlabel metal1 24012 32266 24012 32266 0 _0617_
rlabel metal1 24978 35700 24978 35700 0 _0618_
rlabel metal1 24334 35632 24334 35632 0 _0619_
rlabel via1 25328 35054 25328 35054 0 _0620_
rlabel metal1 25484 35258 25484 35258 0 _0621_
rlabel metal2 24518 33660 24518 33660 0 _0622_
rlabel metal1 27416 30362 27416 30362 0 _0623_
rlabel metal1 27140 31450 27140 31450 0 _0624_
rlabel metal1 27692 31790 27692 31790 0 _0625_
rlabel metal1 24518 31790 24518 31790 0 _0626_
rlabel metal2 24886 30396 24886 30396 0 _0627_
rlabel metal1 20608 41038 20608 41038 0 _0628_
rlabel metal1 2116 29138 2116 29138 0 _0629_
rlabel metal1 2392 40494 2392 40494 0 _0630_
rlabel metal2 2714 29444 2714 29444 0 _0631_
rlabel metal1 19596 42194 19596 42194 0 _0632_
rlabel metal1 2806 36074 2806 36074 0 _0633_
rlabel metal1 2254 30362 2254 30362 0 _0634_
rlabel metal1 4554 40494 4554 40494 0 _0635_
rlabel metal1 3404 30906 3404 30906 0 _0636_
rlabel metal1 18814 40630 18814 40630 0 _0637_
rlabel metal1 18584 39950 18584 39950 0 _0638_
rlabel metal1 16054 33082 16054 33082 0 _0639_
rlabel metal2 16054 32980 16054 32980 0 _0640_
rlabel metal1 16698 33626 16698 33626 0 _0641_
rlabel metal1 17710 34544 17710 34544 0 _0642_
rlabel metal2 17710 34170 17710 34170 0 _0643_
rlabel metal1 17158 34510 17158 34510 0 _0644_
rlabel metal1 16698 33966 16698 33966 0 _0645_
rlabel metal1 18170 37706 18170 37706 0 _0646_
rlabel metal1 18630 36346 18630 36346 0 _0647_
rlabel metal1 19458 36176 19458 36176 0 _0648_
rlabel metal1 16238 31926 16238 31926 0 _0649_
rlabel metal1 17158 31926 17158 31926 0 _0650_
rlabel metal1 18170 35530 18170 35530 0 _0651_
rlabel metal1 18538 37672 18538 37672 0 _0652_
rlabel metal1 17940 37978 17940 37978 0 _0653_
rlabel metal2 18170 38148 18170 38148 0 _0654_
rlabel metal2 14490 31450 14490 31450 0 _0655_
rlabel metal1 15502 31110 15502 31110 0 _0656_
rlabel metal1 18032 38522 18032 38522 0 _0657_
rlabel metal2 17250 39236 17250 39236 0 _0658_
rlabel metal1 13892 32538 13892 32538 0 _0659_
rlabel metal1 13110 33932 13110 33932 0 _0660_
rlabel metal1 14585 33626 14585 33626 0 _0661_
rlabel metal1 13800 34034 13800 34034 0 _0662_
rlabel metal1 14122 34170 14122 34170 0 _0663_
rlabel metal1 16744 36346 16744 36346 0 _0664_
rlabel metal1 14214 34646 14214 34646 0 _0665_
rlabel metal1 12834 34170 12834 34170 0 _0666_
rlabel metal1 13294 36074 13294 36074 0 _0667_
rlabel metal1 15226 36346 15226 36346 0 _0668_
rlabel metal1 14628 37434 14628 37434 0 _0669_
rlabel metal2 14674 37162 14674 37162 0 _0670_
rlabel metal1 13662 36244 13662 36244 0 _0671_
rlabel metal1 13018 36346 13018 36346 0 _0672_
rlabel metal2 12466 36958 12466 36958 0 _0673_
rlabel metal1 12052 34578 12052 34578 0 _0674_
rlabel metal1 12834 34680 12834 34680 0 _0675_
rlabel metal1 11779 33626 11779 33626 0 _0676_
rlabel metal2 12834 34272 12834 34272 0 _0677_
rlabel metal1 13156 34714 13156 34714 0 _0678_
rlabel metal1 15272 40630 15272 40630 0 _0679_
rlabel metal1 16008 39610 16008 39610 0 _0680_
rlabel metal1 12834 39440 12834 39440 0 _0681_
rlabel metal1 16146 40494 16146 40494 0 _0682_
rlabel metal1 16330 40562 16330 40562 0 _0683_
rlabel metal1 17158 40358 17158 40358 0 _0684_
rlabel metal1 13340 34442 13340 34442 0 _0685_
rlabel metal1 17158 35258 17158 35258 0 _0686_
rlabel metal1 17158 40698 17158 40698 0 _0687_
rlabel metal1 17204 41242 17204 41242 0 _0688_
rlabel metal1 30130 25466 30130 25466 0 _0689_
rlabel metal2 30222 29036 30222 29036 0 _0690_
rlabel metal2 14766 19975 14766 19975 0 _0691_
rlabel metal1 8832 20434 8832 20434 0 _0692_
rlabel metal1 13938 19822 13938 19822 0 _0693_
rlabel metal1 6210 24820 6210 24820 0 _0694_
rlabel metal2 12742 19958 12742 19958 0 _0695_
rlabel metal1 4048 25262 4048 25262 0 _0696_
rlabel metal1 2553 26350 2553 26350 0 _0697_
rlabel metal1 2300 24786 2300 24786 0 _0698_
rlabel metal1 3404 24174 3404 24174 0 _0699_
rlabel metal1 23368 35258 23368 35258 0 _0700_
rlabel metal1 23276 34714 23276 34714 0 _0701_
rlabel metal1 22770 34714 22770 34714 0 _0702_
rlabel metal2 23690 33456 23690 33456 0 _0703_
rlabel metal2 16330 17068 16330 17068 0 _0704_
rlabel metal1 24702 29206 24702 29206 0 _0705_
rlabel metal1 23828 29274 23828 29274 0 _0706_
rlabel metal1 22770 31824 22770 31824 0 _0707_
rlabel metal2 17158 5423 17158 5423 0 _0708_
rlabel metal1 12834 30736 12834 30736 0 _0709_
rlabel metal1 22402 40460 22402 40460 0 _0710_
rlabel metal1 12282 41140 12282 41140 0 _0711_
rlabel metal1 14122 41140 14122 41140 0 _0712_
rlabel metal1 21574 6693 21574 6693 0 _0713_
rlabel via1 22034 15011 22034 15011 0 _0714_
rlabel metal1 21758 14416 21758 14416 0 _0715_
rlabel metal1 21390 13294 21390 13294 0 _0716_
rlabel metal1 14766 11730 14766 11730 0 _0717_
rlabel metal1 14766 13158 14766 13158 0 _0718_
rlabel metal1 14536 12614 14536 12614 0 _0719_
rlabel metal1 14490 11798 14490 11798 0 _0720_
rlabel metal1 8648 13294 8648 13294 0 _0721_
rlabel metal2 19734 13566 19734 13566 0 _0722_
rlabel metal1 15226 12342 15226 12342 0 _0723_
rlabel metal1 15318 12682 15318 12682 0 _0724_
rlabel metal1 14076 11730 14076 11730 0 _0725_
rlabel metal1 11822 6970 11822 6970 0 _0726_
rlabel metal1 15824 7378 15824 7378 0 _0727_
rlabel metal1 15686 7412 15686 7412 0 _0728_
rlabel metal2 16974 9724 16974 9724 0 _0729_
rlabel metal1 15318 13498 15318 13498 0 _0730_
rlabel metal1 16652 13430 16652 13430 0 _0731_
rlabel viali 16422 9555 16422 9555 0 _0732_
rlabel metal1 16652 8398 16652 8398 0 _0733_
rlabel metal1 16606 8466 16606 8466 0 _0734_
rlabel metal1 15962 7344 15962 7344 0 _0735_
rlabel metal1 13018 9588 13018 9588 0 _0736_
rlabel metal1 12466 9588 12466 9588 0 _0737_
rlabel metal1 14582 8976 14582 8976 0 _0738_
rlabel metal1 14168 7378 14168 7378 0 _0739_
rlabel metal1 14260 6766 14260 6766 0 _0740_
rlabel metal2 13754 7565 13754 7565 0 _0741_
rlabel metal1 13616 6834 13616 6834 0 _0742_
rlabel metal1 14950 6732 14950 6732 0 _0743_
rlabel metal1 14766 6222 14766 6222 0 _0744_
rlabel metal1 14536 6426 14536 6426 0 _0745_
rlabel metal1 13294 6120 13294 6120 0 _0746_
rlabel metal1 10120 5202 10120 5202 0 _0747_
rlabel metal1 12834 6834 12834 6834 0 _0748_
rlabel metal2 12098 6562 12098 6562 0 _0749_
rlabel metal1 11638 6800 11638 6800 0 _0750_
rlabel metal1 11408 6290 11408 6290 0 _0751_
rlabel metal2 11546 6596 11546 6596 0 _0752_
rlabel metal1 11730 9588 11730 9588 0 _0753_
rlabel metal1 12098 9010 12098 9010 0 _0754_
rlabel metal2 11960 8466 11960 8466 0 _0755_
rlabel metal2 11362 7548 11362 7548 0 _0756_
rlabel metal1 8970 7412 8970 7412 0 _0757_
rlabel metal1 8050 7242 8050 7242 0 _0758_
rlabel metal1 9154 8976 9154 8976 0 _0759_
rlabel metal1 8970 9010 8970 9010 0 _0760_
rlabel metal1 7406 7412 7406 7412 0 _0761_
rlabel metal1 7820 6698 7820 6698 0 _0762_
rlabel metal1 7636 7378 7636 7378 0 _0763_
rlabel metal1 7774 6766 7774 6766 0 _0764_
rlabel metal1 8050 6324 8050 6324 0 _0765_
rlabel metal1 7406 9520 7406 9520 0 _0766_
rlabel metal1 8602 10676 8602 10676 0 _0767_
rlabel metal1 7958 10064 7958 10064 0 _0768_
rlabel metal2 7774 9860 7774 9860 0 _0769_
rlabel metal1 5842 9520 5842 9520 0 _0770_
rlabel metal1 5934 12682 5934 12682 0 _0771_
rlabel metal1 5520 10234 5520 10234 0 _0772_
rlabel metal1 5842 10064 5842 10064 0 _0773_
rlabel metal1 5704 9554 5704 9554 0 _0774_
rlabel metal1 8602 12954 8602 12954 0 _0775_
rlabel viali 8234 13293 8234 13293 0 _0776_
rlabel metal1 7866 13226 7866 13226 0 _0777_
rlabel metal1 8096 11186 8096 11186 0 _0778_
rlabel metal1 7636 11322 7636 11322 0 _0779_
rlabel metal1 5198 13260 5198 13260 0 _0780_
rlabel metal1 5750 12172 5750 12172 0 _0781_
rlabel metal1 3450 11628 3450 11628 0 _0782_
rlabel metal1 4002 12138 4002 12138 0 _0783_
rlabel metal1 5566 12138 5566 12138 0 _0784_
rlabel metal1 4830 12410 4830 12410 0 _0785_
rlabel metal1 4462 12104 4462 12104 0 _0786_
rlabel metal1 4876 11866 4876 11866 0 _0787_
rlabel metal1 5060 12070 5060 12070 0 _0788_
rlabel metal1 6072 13498 6072 13498 0 _0789_
rlabel metal2 10442 13192 10442 13192 0 _0790_
rlabel metal1 10764 12410 10764 12410 0 _0791_
rlabel metal1 10166 12614 10166 12614 0 _0792_
rlabel metal1 11730 12954 11730 12954 0 _0793_
rlabel metal1 10580 12954 10580 12954 0 _0794_
rlabel metal1 9798 12818 9798 12818 0 _0795_
rlabel metal1 7314 12682 7314 12682 0 _0796_
rlabel metal1 30544 17646 30544 17646 0 _0797_
rlabel metal2 30406 17884 30406 17884 0 _0798_
rlabel metal2 14766 16388 14766 16388 0 _0799_
rlabel metal1 8832 15470 8832 15470 0 _0800_
rlabel metal1 14030 16218 14030 16218 0 _0801_
rlabel metal1 7038 17170 7038 17170 0 _0802_
rlabel metal1 11362 17170 11362 17170 0 _0803_
rlabel metal1 5796 16218 5796 16218 0 _0804_
rlabel metal2 4186 15521 4186 15521 0 _0805_
rlabel metal1 2484 15470 2484 15470 0 _0806_
rlabel metal1 2806 17102 2806 17102 0 _0807_
rlabel metal1 18308 30362 18308 30362 0 _0808_
rlabel metal1 27646 5273 27646 5273 0 _0809_
rlabel metal1 27186 5168 27186 5168 0 _0810_
rlabel metal2 21482 19482 21482 19482 0 _0811_
rlabel metal1 17618 19244 17618 19244 0 _0812_
rlabel metal1 17204 19482 17204 19482 0 _0813_
rlabel metal1 27094 17170 27094 17170 0 _0814_
rlabel metal1 27140 33286 27140 33286 0 _0815_
rlabel metal2 24978 30957 24978 30957 0 _0816_
rlabel metal1 25346 27506 25346 27506 0 _0817_
rlabel metal1 27370 19822 27370 19822 0 _0818_
rlabel metal1 31326 26962 31326 26962 0 _0819_
rlabel metal1 38962 31212 38962 31212 0 _0820_
rlabel metal1 36248 33082 36248 33082 0 _0821_
rlabel metal1 37950 30158 37950 30158 0 _0822_
rlabel metal2 34454 23290 34454 23290 0 _0823_
rlabel metal1 39284 26350 39284 26350 0 _0824_
rlabel metal1 34132 27438 34132 27438 0 _0825_
rlabel metal1 38088 25330 38088 25330 0 _0826_
rlabel metal2 19642 17884 19642 17884 0 _0827_
rlabel metal1 38364 30702 38364 30702 0 _0828_
rlabel metal1 37950 30294 37950 30294 0 _0829_
rlabel metal1 35374 30260 35374 30260 0 _0830_
rlabel metal1 32936 24582 32936 24582 0 _0831_
rlabel via1 20838 19907 20838 19907 0 _0832_
rlabel metal1 37766 29648 37766 29648 0 _0833_
rlabel metal1 32430 27438 32430 27438 0 _0834_
rlabel metal1 33718 25330 33718 25330 0 _0835_
rlabel metal1 33442 25194 33442 25194 0 _0836_
rlabel metal1 32844 26350 32844 26350 0 _0837_
rlabel metal1 38594 31858 38594 31858 0 _0838_
rlabel metal1 37352 32402 37352 32402 0 _0839_
rlabel metal2 36294 14246 36294 14246 0 _0840_
rlabel metal1 39146 29546 39146 29546 0 _0841_
rlabel metal1 38548 27438 38548 27438 0 _0842_
rlabel metal1 34086 24106 34086 24106 0 _0843_
rlabel metal1 32706 26418 32706 26418 0 _0844_
rlabel metal1 38778 29138 38778 29138 0 _0845_
rlabel metal1 33580 29478 33580 29478 0 _0846_
rlabel metal1 36708 25398 36708 25398 0 _0847_
rlabel metal1 31970 35700 31970 35700 0 _0848_
rlabel metal1 35006 17578 35006 17578 0 _0849_
rlabel metal1 36156 33422 36156 33422 0 _0850_
rlabel metal1 37950 33456 37950 33456 0 _0851_
rlabel metal1 31694 34068 31694 34068 0 _0852_
rlabel metal1 37697 33966 37697 33966 0 _0853_
rlabel metal1 35512 33830 35512 33830 0 _0854_
rlabel metal1 35834 24582 35834 24582 0 _0855_
rlabel metal2 35374 21835 35374 21835 0 _0856_
rlabel via1 36107 25262 36107 25262 0 _0857_
rlabel metal1 32154 26350 32154 26350 0 _0858_
rlabel metal1 27784 26010 27784 26010 0 _0859_
rlabel metal2 31142 27234 31142 27234 0 _0860_
rlabel metal1 38456 26758 38456 26758 0 _0861_
rlabel metal2 37766 21495 37766 21495 0 _0862_
rlabel metal1 37950 27540 37950 27540 0 _0863_
rlabel metal2 32890 33796 32890 33796 0 _0864_
rlabel metal1 36984 28050 36984 28050 0 _0865_
rlabel metal1 37444 27438 37444 27438 0 _0866_
rlabel metal1 37674 27370 37674 27370 0 _0867_
rlabel metal1 18906 30158 18906 30158 0 _0868_
rlabel metal1 24886 27370 24886 27370 0 _0869_
rlabel metal1 38502 32538 38502 32538 0 _0870_
rlabel metal1 38502 28016 38502 28016 0 _0871_
rlabel via3 39077 13668 39077 13668 0 _0872_
rlabel metal1 36340 34578 36340 34578 0 _0873_
rlabel metal1 34868 28526 34868 28526 0 _0874_
rlabel metal1 36800 31790 36800 31790 0 _0875_
rlabel metal2 36662 31867 36662 31867 0 _0876_
rlabel metal1 29210 29580 29210 29580 0 _0877_
rlabel metal1 34684 35666 34684 35666 0 _0878_
rlabel metal1 34822 35598 34822 35598 0 _0879_
rlabel metal1 30360 29750 30360 29750 0 _0880_
rlabel metal2 29762 23052 29762 23052 0 _0881_
rlabel metal1 26266 29682 26266 29682 0 _0882_
rlabel metal1 32982 24786 32982 24786 0 _0883_
rlabel metal2 34086 29257 34086 29257 0 _0884_
rlabel metal1 34178 26452 34178 26452 0 _0885_
rlabel metal1 34132 18802 34132 18802 0 _0886_
rlabel metal2 21114 28101 21114 28101 0 _0887_
rlabel metal1 26128 29818 26128 29818 0 _0888_
rlabel metal1 35052 30090 35052 30090 0 _0889_
rlabel metal2 36248 27302 36248 27302 0 _0890_
rlabel metal3 39215 13532 39215 13532 0 _0891_
rlabel metal1 27002 34000 27002 34000 0 _0892_
rlabel metal1 37582 33082 37582 33082 0 _0893_
rlabel metal1 34776 31246 34776 31246 0 _0894_
rlabel metal1 32200 35734 32200 35734 0 _0895_
rlabel metal1 21666 28526 21666 28526 0 _0896_
rlabel metal1 34638 33626 34638 33626 0 _0897_
rlabel via1 35282 18275 35282 18275 0 _0898_
rlabel metal2 26818 34986 26818 34986 0 _0899_
rlabel metal1 26312 33082 26312 33082 0 _0900_
rlabel metal1 25622 28730 25622 28730 0 _0901_
rlabel metal1 30130 15606 30130 15606 0 _0902_
rlabel metal2 22126 32895 22126 32895 0 _0903_
rlabel via1 39974 17323 39974 17323 0 _0904_
rlabel metal1 35236 31858 35236 31858 0 _0905_
rlabel metal1 27738 32368 27738 32368 0 _0906_
rlabel metal2 31786 31586 31786 31586 0 _0907_
rlabel metal1 28842 13940 28842 13940 0 _0908_
rlabel metal1 25990 32402 25990 32402 0 _0909_
rlabel metal1 26772 32266 26772 32266 0 _0910_
rlabel metal1 35190 29614 35190 29614 0 _0911_
rlabel metal1 21712 28730 21712 28730 0 _0912_
rlabel metal1 33718 35054 33718 35054 0 _0913_
rlabel metal2 33534 35411 33534 35411 0 _0914_
rlabel metal1 30452 25874 30452 25874 0 _0915_
rlabel metal1 20976 20434 20976 20434 0 _0916_
rlabel metal1 25576 32878 25576 32878 0 _0917_
rlabel metal1 25944 27438 25944 27438 0 _0918_
rlabel metal1 37904 31790 37904 31790 0 _0919_
rlabel metal2 37030 24378 37030 24378 0 _0920_
rlabel metal1 35558 17680 35558 17680 0 _0921_
rlabel metal1 34086 28084 34086 28084 0 _0922_
rlabel metal1 33534 15062 33534 15062 0 _0923_
rlabel metal2 20378 14433 20378 14433 0 _0924_
rlabel metal1 35926 26384 35926 26384 0 _0925_
rlabel metal2 21482 21097 21482 21097 0 _0926_
rlabel metal1 31510 27438 31510 27438 0 _0927_
rlabel metal1 33534 28492 33534 28492 0 _0928_
rlabel metal1 32568 31314 32568 31314 0 _0929_
rlabel metal1 32246 30770 32246 30770 0 _0930_
rlabel metal1 32430 32436 32430 32436 0 _0931_
rlabel metal1 32913 14450 32913 14450 0 _0932_
rlabel metal1 31740 32334 31740 32334 0 _0933_
rlabel metal1 30590 20978 30590 20978 0 _0934_
rlabel metal1 32430 30906 32430 30906 0 _0935_
rlabel metal1 32982 31790 32982 31790 0 _0936_
rlabel metal1 36294 29478 36294 29478 0 _0937_
rlabel metal2 32246 27166 32246 27166 0 _0938_
rlabel metal3 33511 18156 33511 18156 0 _0939_
rlabel metal1 32108 27574 32108 27574 0 _0940_
rlabel metal2 28842 25007 28842 25007 0 _0941_
rlabel metal1 31855 25398 31855 25398 0 _0942_
rlabel metal1 36524 18326 36524 18326 0 _0943_
rlabel metal2 32982 18666 32982 18666 0 _0944_
rlabel metal2 31510 26486 31510 26486 0 _0945_
rlabel metal3 36892 20740 36892 20740 0 _0946_
rlabel metal2 31924 18292 31924 18292 0 _0947_
rlabel metal1 31602 20774 31602 20774 0 _0948_
rlabel metal2 22494 23001 22494 23001 0 _0949_
rlabel metal1 20838 18734 20838 18734 0 _0950_
rlabel metal1 37904 29478 37904 29478 0 _0951_
rlabel metal1 33166 15130 33166 15130 0 _0952_
rlabel metal1 31418 23834 31418 23834 0 _0953_
rlabel metal1 31832 24378 31832 24378 0 _0954_
rlabel metal1 30912 22610 30912 22610 0 _0955_
rlabel metal1 26220 27438 26220 27438 0 _0956_
rlabel metal1 33396 27302 33396 27302 0 _0957_
rlabel metal1 29670 30838 29670 30838 0 _0958_
rlabel metal1 30958 35122 30958 35122 0 _0959_
rlabel metal1 31602 35054 31602 35054 0 _0960_
rlabel metal1 31326 34952 31326 34952 0 _0961_
rlabel metal1 30038 35700 30038 35700 0 _0962_
rlabel metal1 31188 35054 31188 35054 0 _0963_
rlabel metal2 31188 30702 31188 30702 0 _0964_
rlabel metal1 24472 22066 24472 22066 0 _0965_
rlabel metal2 30498 30124 30498 30124 0 _0966_
rlabel metal2 31510 30906 31510 30906 0 _0967_
rlabel metal1 29256 30566 29256 30566 0 _0968_
rlabel metal1 19320 21522 19320 21522 0 _0969_
rlabel metal1 28750 6120 28750 6120 0 _0970_
rlabel metal1 27922 5678 27922 5678 0 _0971_
rlabel metal2 17342 22916 17342 22916 0 _0972_
rlabel metal1 39146 17612 39146 17612 0 _0973_
rlabel metal1 20700 25670 20700 25670 0 _0974_
rlabel metal1 19642 26962 19642 26962 0 _0975_
rlabel metal2 20562 29886 20562 29886 0 _0976_
rlabel metal1 28152 9894 28152 9894 0 _0977_
rlabel metal1 34868 7378 34868 7378 0 _0978_
rlabel metal1 34224 16490 34224 16490 0 _0979_
rlabel metal1 27600 21522 27600 21522 0 _0980_
rlabel metal2 27830 23358 27830 23358 0 _0981_
rlabel metal1 23828 19346 23828 19346 0 _0982_
rlabel metal1 19780 21114 19780 21114 0 _0983_
rlabel metal1 18538 25942 18538 25942 0 _0984_
rlabel metal1 19918 16626 19918 16626 0 _0985_
rlabel metal1 28474 9010 28474 9010 0 _0986_
rlabel metal1 25162 24242 25162 24242 0 _0987_
rlabel metal1 26036 14518 26036 14518 0 _0988_
rlabel metal1 26818 14382 26818 14382 0 _0989_
rlabel metal2 26266 26775 26266 26775 0 _0990_
rlabel metal1 26634 26758 26634 26758 0 _0991_
rlabel metal2 26956 23868 26956 23868 0 _0992_
rlabel metal1 30268 15470 30268 15470 0 _0993_
rlabel metal1 26864 13430 26864 13430 0 _0994_
rlabel metal1 26588 15470 26588 15470 0 _0995_
rlabel metal1 26358 15504 26358 15504 0 _0996_
rlabel metal1 27048 13362 27048 13362 0 _0997_
rlabel metal1 27186 14416 27186 14416 0 _0998_
rlabel metal2 27738 5253 27738 5253 0 _0999_
rlabel metal2 27922 15079 27922 15079 0 _1000_
rlabel metal1 25208 20434 25208 20434 0 _1001_
rlabel metal1 21298 29138 21298 29138 0 _1002_
rlabel metal2 28152 20502 28152 20502 0 _1003_
rlabel metal2 29486 16728 29486 16728 0 _1004_
rlabel via2 30038 17323 30038 17323 0 _1005_
rlabel metal1 20884 18598 20884 18598 0 _1006_
rlabel metal1 28106 36210 28106 36210 0 _1007_
rlabel metal2 28474 36788 28474 36788 0 _1008_
rlabel metal2 18906 22304 18906 22304 0 _1009_
rlabel metal3 19251 18292 19251 18292 0 _1010_
rlabel via2 28474 15147 28474 15147 0 _1011_
rlabel metal1 27462 36720 27462 36720 0 _1012_
rlabel metal2 18538 29478 18538 29478 0 _1013_
rlabel metal1 26174 28560 26174 28560 0 _1014_
rlabel metal2 21206 18972 21206 18972 0 _1015_
rlabel via1 26084 18734 26084 18734 0 _1016_
rlabel metal1 23460 7854 23460 7854 0 _1017_
rlabel metal1 21942 7446 21942 7446 0 _1018_
rlabel metal1 32384 12614 32384 12614 0 _1019_
rlabel metal1 35972 7174 35972 7174 0 _1020_
rlabel metal2 18446 8007 18446 8007 0 _1021_
rlabel metal1 32338 9588 32338 9588 0 _1022_
rlabel metal1 32522 10710 32522 10710 0 _1023_
rlabel metal1 33994 20842 33994 20842 0 _1024_
rlabel via1 28566 8891 28566 8891 0 _1025_
rlabel metal1 29394 7718 29394 7718 0 _1026_
rlabel metal1 30222 9962 30222 9962 0 _1027_
rlabel metal1 26910 10132 26910 10132 0 _1028_
rlabel metal1 25070 9044 25070 9044 0 _1029_
rlabel metal1 30360 11798 30360 11798 0 _1030_
rlabel via1 36123 13906 36123 13906 0 _1031_
rlabel metal1 35282 19822 35282 19822 0 _1032_
rlabel metal1 39146 13328 39146 13328 0 _1033_
rlabel metal1 39514 21658 39514 21658 0 _1034_
rlabel metal1 30038 10642 30038 10642 0 _1035_
rlabel metal1 32890 12750 32890 12750 0 _1036_
rlabel metal1 35742 13226 35742 13226 0 _1037_
rlabel metal2 36708 12818 36708 12818 0 _1038_
rlabel metal1 33028 10778 33028 10778 0 _1039_
rlabel metal1 32108 8398 32108 8398 0 _1040_
rlabel metal1 29578 11696 29578 11696 0 _1041_
rlabel metal1 34546 7344 34546 7344 0 _1042_
rlabel metal2 28658 7038 28658 7038 0 _1043_
rlabel metal1 28934 7412 28934 7412 0 _1044_
rlabel metal1 28898 6630 28898 6630 0 _1045_
rlabel metal1 26542 6256 26542 6256 0 _1046_
rlabel metal1 28198 9044 28198 9044 0 _1047_
rlabel metal1 27646 8534 27646 8534 0 _1048_
rlabel metal1 34822 8466 34822 8466 0 _1049_
rlabel metal1 31280 7378 31280 7378 0 _1050_
rlabel metal1 37260 7854 37260 7854 0 _1051_
rlabel metal1 35926 13872 35926 13872 0 _1052_
rlabel metal1 36340 7514 36340 7514 0 _1053_
rlabel metal1 32798 12104 32798 12104 0 _1054_
rlabel metal1 33442 6800 33442 6800 0 _1055_
rlabel metal1 36938 7820 36938 7820 0 _1056_
rlabel metal1 35558 15402 35558 15402 0 _1057_
rlabel metal1 31786 7208 31786 7208 0 _1058_
rlabel metal1 33626 6868 33626 6868 0 _1059_
rlabel metal1 33672 6698 33672 6698 0 _1060_
rlabel metal1 30038 6698 30038 6698 0 _1061_
rlabel metal2 26818 7072 26818 7072 0 _1062_
rlabel metal1 33764 6766 33764 6766 0 _1063_
rlabel metal1 33442 9928 33442 9928 0 _1064_
rlabel metal1 31280 6290 31280 6290 0 _1065_
rlabel metal1 30590 5712 30590 5712 0 _1066_
rlabel metal1 32338 6766 32338 6766 0 _1067_
rlabel metal1 32522 5338 32522 5338 0 _1068_
rlabel metal1 27876 8602 27876 8602 0 _1069_
rlabel metal1 35052 6766 35052 6766 0 _1070_
rlabel metal1 36386 6970 36386 6970 0 _1071_
rlabel metal1 27002 7446 27002 7446 0 _1072_
rlabel metal1 30222 12138 30222 12138 0 _1073_
rlabel metal1 32499 7378 32499 7378 0 _1074_
rlabel metal1 32108 6834 32108 6834 0 _1075_
rlabel metal1 31510 5338 31510 5338 0 _1076_
rlabel metal1 30866 4114 30866 4114 0 _1077_
rlabel metal1 24610 26418 24610 26418 0 _1078_
rlabel metal2 14766 3553 14766 3553 0 _1079_
rlabel metal2 33718 8704 33718 8704 0 _1080_
rlabel metal1 37536 16082 37536 16082 0 _1081_
rlabel metal2 33810 16864 33810 16864 0 _1082_
rlabel metal1 37490 16728 37490 16728 0 _1083_
rlabel metal1 30544 19754 30544 19754 0 _1084_
rlabel metal1 35880 22610 35880 22610 0 _1085_
rlabel metal1 33120 14314 33120 14314 0 _1086_
rlabel metal1 32016 19822 32016 19822 0 _1087_
rlabel metal1 37582 20468 37582 20468 0 _1088_
rlabel metal1 38364 17646 38364 17646 0 _1089_
rlabel metal2 36110 11220 36110 11220 0 _1090_
rlabel metal2 37674 14144 37674 14144 0 _1091_
rlabel metal2 38962 22610 38962 22610 0 _1092_
rlabel metal1 33534 14382 33534 14382 0 _1093_
rlabel metal2 35282 10506 35282 10506 0 _1094_
rlabel metal2 38870 16116 38870 16116 0 _1095_
rlabel metal1 35006 19856 35006 19856 0 _1096_
rlabel metal2 33534 9826 33534 9826 0 _1097_
rlabel metal1 38916 13226 38916 13226 0 _1098_
rlabel metal1 34638 19822 34638 19822 0 _1099_
rlabel metal1 37996 18734 37996 18734 0 _1100_
rlabel metal1 37260 21114 37260 21114 0 _1101_
rlabel metal1 30544 14382 30544 14382 0 _1102_
rlabel metal1 35052 8874 35052 8874 0 _1103_
rlabel metal1 38686 13192 38686 13192 0 _1104_
rlabel metal2 35834 15504 35834 15504 0 _1105_
rlabel metal1 36754 18190 36754 18190 0 _1106_
rlabel via1 38870 13379 38870 13379 0 _1107_
rlabel metal1 32798 12818 32798 12818 0 _1108_
rlabel metal1 36478 18666 36478 18666 0 _1109_
rlabel metal1 32798 20842 32798 20842 0 _1110_
rlabel metal1 32706 21114 32706 21114 0 _1111_
rlabel metal1 36708 20230 36708 20230 0 _1112_
rlabel metal1 32203 16558 32203 16558 0 _1113_
rlabel metal1 33212 12818 33212 12818 0 _1114_
rlabel metal1 33166 11152 33166 11152 0 _1115_
rlabel metal1 33166 12682 33166 12682 0 _1116_
rlabel metal1 32890 12954 32890 12954 0 _1117_
rlabel metal1 38870 17578 38870 17578 0 _1118_
rlabel metal2 40158 17986 40158 17986 0 _1119_
rlabel metal3 37743 18564 37743 18564 0 _1120_
rlabel metal1 31096 22950 31096 22950 0 _1121_
rlabel metal1 38870 21386 38870 21386 0 _1122_
rlabel metal1 38824 15130 38824 15130 0 _1123_
rlabel metal1 37122 21522 37122 21522 0 _1124_
rlabel metal1 38272 18938 38272 18938 0 _1125_
rlabel metal1 36708 18938 36708 18938 0 _1126_
rlabel metal2 37858 20332 37858 20332 0 _1127_
rlabel metal1 36662 18734 36662 18734 0 _1128_
rlabel metal1 37674 18802 37674 18802 0 _1129_
rlabel via1 35742 7259 35742 7259 0 _1130_
rlabel metal1 35834 16048 35834 16048 0 _1131_
rlabel metal2 35558 21114 35558 21114 0 _1132_
rlabel metal1 38502 18802 38502 18802 0 _1133_
rlabel metal1 40066 18768 40066 18768 0 _1134_
rlabel metal1 34178 13294 34178 13294 0 _1135_
rlabel metal1 33120 9962 33120 9962 0 _1136_
rlabel metal1 33948 8942 33948 8942 0 _1137_
rlabel metal1 34224 9146 34224 9146 0 _1138_
rlabel metal1 35788 9554 35788 9554 0 _1139_
rlabel metal1 34638 9588 34638 9588 0 _1140_
rlabel metal2 33994 11458 33994 11458 0 _1141_
rlabel metal1 39974 13396 39974 13396 0 _1142_
rlabel metal1 39652 12954 39652 12954 0 _1143_
rlabel metal1 39606 13294 39606 13294 0 _1144_
rlabel metal1 40112 14382 40112 14382 0 _1145_
rlabel via3 35995 12036 35995 12036 0 _1146_
rlabel metal1 35466 9690 35466 9690 0 _1147_
rlabel metal3 34799 22508 34799 22508 0 _1148_
rlabel metal1 35650 11696 35650 11696 0 _1149_
rlabel metal2 36570 14450 36570 14450 0 _1150_
rlabel metal1 29440 32402 29440 32402 0 _1151_
rlabel metal1 30958 11764 30958 11764 0 _1152_
rlabel metal1 30820 12750 30820 12750 0 _1153_
rlabel metal1 29716 12954 29716 12954 0 _1154_
rlabel metal1 32568 13906 32568 13906 0 _1155_
rlabel metal1 36018 12818 36018 12818 0 _1156_
rlabel metal1 39882 14552 39882 14552 0 _1157_
rlabel via1 31694 14858 31694 14858 0 _1158_
rlabel metal1 31694 14246 31694 14246 0 _1159_
rlabel via2 39974 14467 39974 14467 0 _1160_
rlabel metal1 37306 14246 37306 14246 0 _1161_
rlabel metal2 40342 16422 40342 16422 0 _1162_
rlabel metal1 41078 18122 41078 18122 0 _1163_
rlabel metal1 37490 11084 37490 11084 0 _1164_
rlabel metal2 34914 18530 34914 18530 0 _1165_
rlabel metal1 39790 18224 39790 18224 0 _1166_
rlabel metal1 33580 14586 33580 14586 0 _1167_
rlabel metal1 36294 18666 36294 18666 0 _1168_
rlabel metal1 37076 14382 37076 14382 0 _1169_
rlabel metal1 39284 16082 39284 16082 0 _1170_
rlabel metal2 39698 18598 39698 18598 0 _1171_
rlabel metal1 38870 23630 38870 23630 0 _1172_
rlabel metal1 40434 16558 40434 16558 0 _1173_
rlabel metal1 38042 21454 38042 21454 0 _1174_
rlabel metal2 32062 14841 32062 14841 0 _1175_
rlabel metal2 30084 9010 30084 9010 0 _1176_
rlabel metal1 31694 13838 31694 13838 0 _1177_
rlabel metal1 38962 15878 38962 15878 0 _1178_
rlabel metal2 39882 14348 39882 14348 0 _1179_
rlabel via3 37099 24956 37099 24956 0 _1180_
rlabel metal1 38364 11118 38364 11118 0 _1181_
rlabel metal1 39606 16490 39606 16490 0 _1182_
rlabel metal1 40158 16762 40158 16762 0 _1183_
rlabel metal2 30498 35088 30498 35088 0 _1184_
rlabel metal1 39376 20910 39376 20910 0 _1185_
rlabel metal1 30038 20876 30038 20876 0 _1186_
rlabel metal1 32154 14008 32154 14008 0 _1187_
rlabel metal1 31188 16150 31188 16150 0 _1188_
rlabel metal1 38410 16014 38410 16014 0 _1189_
rlabel metal1 40066 17238 40066 17238 0 _1190_
rlabel metal1 40296 17306 40296 17306 0 _1191_
rlabel metal1 41124 18394 41124 18394 0 _1192_
rlabel metal1 38180 21590 38180 21590 0 _1193_
rlabel metal1 38410 21318 38410 21318 0 _1194_
rlabel metal2 37352 16116 37352 16116 0 _1195_
rlabel metal1 37904 8602 37904 8602 0 _1196_
rlabel via2 33626 19397 33626 19397 0 _1197_
rlabel metal1 37996 10234 37996 10234 0 _1198_
rlabel via3 38893 20740 38893 20740 0 _1199_
rlabel metal1 39376 19142 39376 19142 0 _1200_
rlabel metal1 39928 20978 39928 20978 0 _1201_
rlabel metal1 37444 20434 37444 20434 0 _1202_
rlabel metal1 39146 20434 39146 20434 0 _1203_
rlabel metal2 39606 19788 39606 19788 0 _1204_
rlabel metal1 39284 19414 39284 19414 0 _1205_
rlabel viali 39884 18734 39884 18734 0 _1206_
rlabel metal1 40066 23290 40066 23290 0 _1207_
rlabel metal2 37950 18054 37950 18054 0 _1208_
rlabel via2 19826 13923 19826 13923 0 _1209_
rlabel metal1 37904 14382 37904 14382 0 _1210_
rlabel metal1 36892 14586 36892 14586 0 _1211_
rlabel metal1 37582 13260 37582 13260 0 _1212_
rlabel metal1 37904 13498 37904 13498 0 _1213_
rlabel via1 31799 18734 31799 18734 0 _1214_
rlabel metal1 37628 18734 37628 18734 0 _1215_
rlabel metal1 37858 18666 37858 18666 0 _1216_
rlabel metal1 37858 18326 37858 18326 0 _1217_
rlabel metal2 37674 19822 37674 19822 0 _1218_
rlabel metal2 38134 18156 38134 18156 0 _1219_
rlabel metal1 39974 18360 39974 18360 0 _1220_
rlabel metal1 34730 13804 34730 13804 0 _1221_
rlabel metal2 39882 15810 39882 15810 0 _1222_
rlabel metal1 39422 14586 39422 14586 0 _1223_
rlabel metal1 39790 15470 39790 15470 0 _1224_
rlabel metal1 40480 15674 40480 15674 0 _1225_
rlabel metal1 36248 26486 36248 26486 0 _1226_
rlabel metal1 39330 22406 39330 22406 0 _1227_
rlabel metal1 39238 20978 39238 20978 0 _1228_
rlabel metal1 34799 22066 34799 22066 0 _1229_
rlabel metal1 39928 22746 39928 22746 0 _1230_
rlabel metal2 40342 23732 40342 23732 0 _1231_
rlabel via2 40066 11645 40066 11645 0 _1232_
rlabel metal1 35926 7922 35926 7922 0 _1233_
rlabel metal1 37536 8058 37536 8058 0 _1234_
rlabel metal1 38088 8398 38088 8398 0 _1235_
rlabel metal3 32821 13804 32821 13804 0 _1236_
rlabel metal1 39238 10234 39238 10234 0 _1237_
rlabel metal1 40710 20434 40710 20434 0 _1238_
rlabel metal1 40434 20808 40434 20808 0 _1239_
rlabel metal1 40158 20264 40158 20264 0 _1240_
rlabel metal2 36662 19822 36662 19822 0 _1241_
rlabel metal1 39974 20468 39974 20468 0 _1242_
rlabel metal1 40204 20570 40204 20570 0 _1243_
rlabel metal1 21850 39066 21850 39066 0 _1244_
rlabel metal1 17664 29002 17664 29002 0 _1245_
rlabel metal1 18676 18190 18676 18190 0 _1246_
rlabel metal1 17894 19414 17894 19414 0 _1247_
rlabel metal1 17480 14382 17480 14382 0 _1248_
rlabel metal1 19182 14382 19182 14382 0 _1249_
rlabel metal1 29118 28152 29118 28152 0 _1250_
rlabel metal1 20102 17136 20102 17136 0 _1251_
rlabel metal1 21390 17646 21390 17646 0 _1252_
rlabel metal1 22402 17170 22402 17170 0 _1253_
rlabel metal1 29762 16626 29762 16626 0 _1254_
rlabel metal2 21942 16422 21942 16422 0 _1255_
rlabel metal2 23598 14654 23598 14654 0 _1256_
rlabel metal1 19918 17646 19918 17646 0 _1257_
rlabel via2 27830 14331 27830 14331 0 _1258_
rlabel metal1 17710 13362 17710 13362 0 _1259_
rlabel metal1 20838 13872 20838 13872 0 _1260_
rlabel metal1 15180 7378 15180 7378 0 _1261_
rlabel metal1 25783 25874 25783 25874 0 _1262_
rlabel metal1 25024 14246 25024 14246 0 _1263_
rlabel metal2 24886 19805 24886 19805 0 _1264_
rlabel metal1 24472 12886 24472 12886 0 _1265_
rlabel metal1 25576 18938 25576 18938 0 _1266_
rlabel metal1 25530 24072 25530 24072 0 _1267_
rlabel metal1 25622 18700 25622 18700 0 _1268_
rlabel metal1 25070 18598 25070 18598 0 _1269_
rlabel metal2 21666 15725 21666 15725 0 _1270_
rlabel metal2 20838 27863 20838 27863 0 _1271_
rlabel metal1 23184 18734 23184 18734 0 _1272_
rlabel metal2 24058 23647 24058 23647 0 _1273_
rlabel metal1 23276 21998 23276 21998 0 _1274_
rlabel metal1 26496 30634 26496 30634 0 _1275_
rlabel metal2 23690 18054 23690 18054 0 _1276_
rlabel metal1 23092 18938 23092 18938 0 _1277_
rlabel metal1 18538 22508 18538 22508 0 _1278_
rlabel metal1 24058 21454 24058 21454 0 _1279_
rlabel metal1 23000 22134 23000 22134 0 _1280_
rlabel metal2 29992 19822 29992 19822 0 _1281_
rlabel metal1 28290 19346 28290 19346 0 _1282_
rlabel metal1 23690 18768 23690 18768 0 _1283_
rlabel metal1 23368 17170 23368 17170 0 _1284_
rlabel metal1 18354 28492 18354 28492 0 _1285_
rlabel metal2 22310 15742 22310 15742 0 _1286_
rlabel metal1 21620 21114 21620 21114 0 _1287_
rlabel metal2 21850 21250 21850 21250 0 _1288_
rlabel metal2 20746 22406 20746 22406 0 _1289_
rlabel metal1 21804 17102 21804 17102 0 _1290_
rlabel metal1 23046 20332 23046 20332 0 _1291_
rlabel metal1 23368 16966 23368 16966 0 _1292_
rlabel metal1 21528 16966 21528 16966 0 _1293_
rlabel metal2 31786 31008 31786 31008 0 _1294_
rlabel metal1 33442 27064 33442 27064 0 _1295_
rlabel metal4 21068 19584 21068 19584 0 _1296_
rlabel metal1 21712 19278 21712 19278 0 _1297_
rlabel metal1 21298 15436 21298 15436 0 _1298_
rlabel metal2 21298 17340 21298 17340 0 _1299_
rlabel metal1 22678 17306 22678 17306 0 _1300_
rlabel metal2 23276 20774 23276 20774 0 _1301_
rlabel metal2 26082 14450 26082 14450 0 _1302_
rlabel metal1 26128 16762 26128 16762 0 _1303_
rlabel metal2 23966 16422 23966 16422 0 _1304_
rlabel metal2 16238 14149 16238 14149 0 _1305_
rlabel metal2 18170 29070 18170 29070 0 _1306_
rlabel metal1 16514 28662 16514 28662 0 _1307_
rlabel metal1 28198 24752 28198 24752 0 _1308_
rlabel metal2 28658 26146 28658 26146 0 _1309_
rlabel metal1 28658 24378 28658 24378 0 _1310_
rlabel metal1 21068 24786 21068 24786 0 _1311_
rlabel metal1 20746 27880 20746 27880 0 _1312_
rlabel metal1 26082 21556 26082 21556 0 _1313_
rlabel metal1 26956 13974 26956 13974 0 _1314_
rlabel metal1 27186 21964 27186 21964 0 _1315_
rlabel metal1 28198 32368 28198 32368 0 _1316_
rlabel metal1 27462 14960 27462 14960 0 _1317_
rlabel metal1 29716 22202 29716 22202 0 _1318_
rlabel metal1 29210 21998 29210 21998 0 _1319_
rlabel metal1 28566 20026 28566 20026 0 _1320_
rlabel metal2 32338 34969 32338 34969 0 _1321_
rlabel metal1 28658 21386 28658 21386 0 _1322_
rlabel metal1 28336 21522 28336 21522 0 _1323_
rlabel metal2 27830 18938 27830 18938 0 _1324_
rlabel metal1 34178 26792 34178 26792 0 _1325_
rlabel metal2 28106 21692 28106 21692 0 _1326_
rlabel metal2 32062 32572 32062 32572 0 _1327_
rlabel metal1 28106 21998 28106 21998 0 _1328_
rlabel metal1 28520 21658 28520 21658 0 _1329_
rlabel metal1 28290 22066 28290 22066 0 _1330_
rlabel via2 21666 22219 21666 22219 0 _1331_
rlabel metal1 14030 25194 14030 25194 0 _1332_
rlabel metal1 7222 26894 7222 26894 0 _1333_
rlabel via1 17526 29206 17526 29206 0 _1334_
rlabel metal1 23276 20910 23276 20910 0 _1335_
rlabel metal1 21574 30056 21574 30056 0 _1336_
rlabel metal1 25668 15674 25668 15674 0 _1337_
rlabel metal1 21850 26248 21850 26248 0 _1338_
rlabel metal1 20700 26554 20700 26554 0 _1339_
rlabel metal1 17342 28526 17342 28526 0 _1340_
rlabel metal1 17296 29274 17296 29274 0 _1341_
rlabel metal3 5750 28900 5750 28900 0 _1342_
rlabel metal1 14306 29274 14306 29274 0 _1343_
rlabel metal1 28014 19448 28014 19448 0 _1344_
rlabel metal2 20746 19516 20746 19516 0 _1345_
rlabel via2 21482 34051 21482 34051 0 _1346_
rlabel metal1 26588 31246 26588 31246 0 _1347_
rlabel metal2 28934 28288 28934 28288 0 _1348_
rlabel metal1 29578 34000 29578 34000 0 _1349_
rlabel metal2 28750 28237 28750 28237 0 _1350_
rlabel metal1 29302 28016 29302 28016 0 _1351_
rlabel metal1 28520 28118 28520 28118 0 _1352_
rlabel metal1 25852 22134 25852 22134 0 _1353_
rlabel metal1 25714 21930 25714 21930 0 _1354_
rlabel metal1 25622 21318 25622 21318 0 _1355_
rlabel metal2 25346 22882 25346 22882 0 _1356_
rlabel metal1 24288 14994 24288 14994 0 _1357_
rlabel metal1 28336 23086 28336 23086 0 _1358_
rlabel metal1 27968 23290 27968 23290 0 _1359_
rlabel via1 26910 23290 26910 23290 0 _1360_
rlabel metal1 20286 20910 20286 20910 0 _1361_
rlabel metal1 26726 15436 26726 15436 0 _1362_
rlabel metal1 26910 15130 26910 15130 0 _1363_
rlabel metal1 27186 11866 27186 11866 0 _1364_
rlabel metal1 26910 12172 26910 12172 0 _1365_
rlabel metal2 26956 14042 26956 14042 0 _1366_
rlabel metal3 20677 18972 20677 18972 0 _1367_
rlabel metal1 16100 20842 16100 20842 0 _1368_
rlabel metal1 28842 21046 28842 21046 0 _1369_
rlabel metal2 26634 12631 26634 12631 0 _1370_
rlabel metal1 27646 20978 27646 20978 0 _1371_
rlabel metal1 18998 21080 18998 21080 0 _1372_
rlabel metal1 16974 20944 16974 20944 0 _1373_
rlabel metal1 27140 24038 27140 24038 0 _1374_
rlabel metal1 26726 23120 26726 23120 0 _1375_
rlabel metal1 16836 13294 16836 13294 0 _1376_
rlabel metal2 25806 14875 25806 14875 0 _1377_
rlabel metal1 16836 20910 16836 20910 0 _1378_
rlabel metal1 16744 20502 16744 20502 0 _1379_
rlabel metal1 12765 18734 12765 18734 0 _1380_
rlabel metal2 16192 22406 16192 22406 0 _1381_
rlabel metal1 15594 21658 15594 21658 0 _1382_
rlabel metal2 16514 22882 16514 22882 0 _1383_
rlabel via1 8236 24786 8236 24786 0 _1384_
rlabel metal1 15134 20910 15134 20910 0 _1385_
rlabel metal1 5474 24174 5474 24174 0 _1386_
rlabel metal1 15226 19788 15226 19788 0 _1387_
rlabel metal2 14582 19550 14582 19550 0 _1388_
rlabel metal2 16146 20876 16146 20876 0 _1389_
rlabel metal1 15640 20570 15640 20570 0 _1390_
rlabel metal1 15410 20366 15410 20366 0 _1391_
rlabel metal2 4738 20876 4738 20876 0 _1392_
rlabel metal1 5336 20026 5336 20026 0 _1393_
rlabel metal1 4784 24718 4784 24718 0 _1394_
rlabel metal2 14674 23596 14674 23596 0 _1395_
rlabel metal1 5796 27438 5796 27438 0 _1396_
rlabel metal1 29854 29648 29854 29648 0 _1397_
rlabel metal1 30498 27642 30498 27642 0 _1398_
rlabel metal2 27278 31943 27278 31943 0 _1399_
rlabel via1 23856 31314 23856 31314 0 _1400_
rlabel metal1 33488 29750 33488 29750 0 _1401_
rlabel metal2 30130 30736 30130 30736 0 _1402_
rlabel metal1 33350 31382 33350 31382 0 _1403_
rlabel metal2 33810 31518 33810 31518 0 _1404_
rlabel metal1 29946 31348 29946 31348 0 _1405_
rlabel metal1 30406 31212 30406 31212 0 _1406_
rlabel metal1 24748 31790 24748 31790 0 _1407_
rlabel metal1 24656 31450 24656 31450 0 _1408_
rlabel metal1 24932 32198 24932 32198 0 _1409_
rlabel metal1 28520 32266 28520 32266 0 _1410_
rlabel metal1 23092 20502 23092 20502 0 _1411_
rlabel metal1 27278 31926 27278 31926 0 _1412_
rlabel metal2 24702 32895 24702 32895 0 _1413_
rlabel metal1 26404 35122 26404 35122 0 _1414_
rlabel metal1 26956 34578 26956 34578 0 _1415_
rlabel via2 27646 34731 27646 34731 0 _1416_
rlabel metal1 24564 32878 24564 32878 0 _1417_
rlabel metal1 23966 33014 23966 33014 0 _1418_
rlabel metal1 21850 26452 21850 26452 0 _1419_
rlabel metal1 24334 26758 24334 26758 0 _1420_
rlabel metal2 21758 26537 21758 26537 0 _1421_
rlabel metal2 24702 17782 24702 17782 0 _1422_
rlabel metal1 24196 26282 24196 26282 0 _1423_
rlabel metal1 21965 26894 21965 26894 0 _1424_
rlabel metal2 19458 27642 19458 27642 0 _1425_
rlabel metal1 23138 33626 23138 33626 0 _1426_
rlabel metal1 22310 31382 22310 31382 0 _1427_
rlabel metal1 23736 26962 23736 26962 0 _1428_
rlabel metal1 24196 26554 24196 26554 0 _1429_
rlabel metal1 24426 26010 24426 26010 0 _1430_
rlabel metal1 23966 26486 23966 26486 0 _1431_
rlabel metal1 20332 29070 20332 29070 0 _1432_
rlabel metal1 19642 28594 19642 28594 0 _1433_
rlabel metal1 16606 29002 16606 29002 0 _1434_
rlabel metal2 8234 29376 8234 29376 0 _1435_
rlabel metal1 20608 28730 20608 28730 0 _1436_
rlabel metal1 19918 28594 19918 28594 0 _1437_
rlabel metal1 16238 28560 16238 28560 0 _1438_
rlabel metal2 15594 28288 15594 28288 0 _1439_
rlabel metal1 15318 29070 15318 29070 0 _1440_
rlabel metal1 5796 28526 5796 28526 0 _1441_
rlabel metal1 5888 27030 5888 27030 0 _1442_
rlabel metal1 25622 28492 25622 28492 0 _1443_
rlabel metal1 26266 28084 26266 28084 0 _1444_
rlabel metal1 25484 25466 25484 25466 0 _1445_
rlabel metal1 23460 12342 23460 12342 0 _1446_
rlabel metal1 24012 12614 24012 12614 0 _1447_
rlabel metal1 24840 12818 24840 12818 0 _1448_
rlabel metal1 23966 11696 23966 11696 0 _1449_
rlabel metal1 24112 12886 24112 12886 0 _1450_
rlabel metal2 24334 13311 24334 13311 0 _1451_
rlabel metal1 29164 23834 29164 23834 0 _1452_
rlabel metal1 27692 24378 27692 24378 0 _1453_
rlabel metal1 27876 25466 27876 25466 0 _1454_
rlabel metal1 27554 25874 27554 25874 0 _1455_
rlabel metal1 27232 24786 27232 24786 0 _1456_
rlabel metal1 25254 25194 25254 25194 0 _1457_
rlabel metal1 18998 26962 18998 26962 0 _1458_
rlabel metal1 21022 28084 21022 28084 0 _1459_
rlabel metal2 19550 27744 19550 27744 0 _1460_
rlabel metal1 26680 27642 26680 27642 0 _1461_
rlabel metal1 25990 26418 25990 26418 0 _1462_
rlabel metal1 26818 14586 26818 14586 0 _1463_
rlabel metal1 26220 23562 26220 23562 0 _1464_
rlabel metal2 18906 27030 18906 27030 0 _1465_
rlabel metal1 18217 26350 18217 26350 0 _1466_
rlabel metal1 18124 27438 18124 27438 0 _1467_
rlabel metal1 7774 27472 7774 27472 0 _1468_
rlabel metal1 9522 26928 9522 26928 0 _1469_
rlabel metal1 21758 23698 21758 23698 0 _1470_
rlabel metal1 20562 23766 20562 23766 0 _1471_
rlabel metal1 18676 26826 18676 26826 0 _1472_
rlabel metal1 18734 27030 18734 27030 0 _1473_
rlabel metal1 16698 26894 16698 26894 0 _1474_
rlabel metal1 8050 27404 8050 27404 0 _1475_
rlabel metal1 9246 26248 9246 26248 0 _1476_
rlabel metal1 16790 27472 16790 27472 0 _1477_
rlabel metal2 9614 25534 9614 25534 0 _1478_
rlabel metal1 8694 26010 8694 26010 0 _1479_
rlabel metal1 9614 26520 9614 26520 0 _1480_
rlabel metal1 5796 27098 5796 27098 0 _1481_
rlabel metal1 3634 15334 3634 15334 0 _1482_
rlabel metal1 8878 13838 8878 13838 0 _1483_
rlabel metal2 15318 15283 15318 15283 0 _1484_
rlabel metal1 22954 13260 22954 13260 0 _1485_
rlabel metal1 23138 20570 23138 20570 0 _1486_
rlabel metal1 22494 22134 22494 22134 0 _1487_
rlabel metal1 22494 20876 22494 20876 0 _1488_
rlabel metal1 22448 12886 22448 12886 0 _1489_
rlabel metal1 23736 11866 23736 11866 0 _1490_
rlabel metal1 22816 12818 22816 12818 0 _1491_
rlabel metal2 21942 12517 21942 12517 0 _1492_
rlabel metal1 7958 24276 7958 24276 0 _1493_
rlabel metal2 15134 37536 15134 37536 0 _1494_
rlabel metal1 10672 14382 10672 14382 0 _1495_
rlabel metal2 21850 28815 21850 28815 0 _1496_
rlabel metal1 18400 25194 18400 25194 0 _1497_
rlabel metal1 25530 31246 25530 31246 0 _1498_
rlabel metal1 24610 24276 24610 24276 0 _1499_
rlabel metal1 24472 17850 24472 17850 0 _1500_
rlabel metal1 19780 24582 19780 24582 0 _1501_
rlabel metal2 21482 31994 21482 31994 0 _1502_
rlabel metal2 22126 31382 22126 31382 0 _1503_
rlabel metal1 21850 31246 21850 31246 0 _1504_
rlabel metal1 19136 24786 19136 24786 0 _1505_
rlabel metal1 18676 25262 18676 25262 0 _1506_
rlabel metal1 22954 26928 22954 26928 0 _1507_
rlabel metal1 23046 27098 23046 27098 0 _1508_
rlabel via2 21298 23035 21298 23035 0 clk
rlabel metal1 16744 13906 16744 13906 0 clknet_0_clk
rlabel metal2 2714 20910 2714 20910 0 clknet_4_0_0_clk
rlabel metal1 33350 5270 33350 5270 0 clknet_4_10_0_clk
rlabel metal2 21850 7378 21850 7378 0 clknet_4_11_0_clk
rlabel metal1 17434 19890 17434 19890 0 clknet_4_12_0_clk
rlabel metal1 27876 36686 27876 36686 0 clknet_4_13_0_clk
rlabel metal1 37904 24718 37904 24718 0 clknet_4_14_0_clk
rlabel metal1 38870 32436 38870 32436 0 clknet_4_15_0_clk
rlabel metal2 2438 24786 2438 24786 0 clknet_4_1_0_clk
rlabel metal1 1794 16694 1794 16694 0 clknet_4_2_0_clk
rlabel metal2 13110 20196 13110 20196 0 clknet_4_3_0_clk
rlabel metal1 2254 31382 2254 31382 0 clknet_4_4_0_clk
rlabel metal1 2070 38862 2070 38862 0 clknet_4_5_0_clk
rlabel metal1 16652 34034 16652 34034 0 clknet_4_6_0_clk
rlabel metal1 18124 41650 18124 41650 0 clknet_4_7_0_clk
rlabel metal1 21804 9010 21804 9010 0 clknet_4_8_0_clk
rlabel metal1 14122 16660 14122 16660 0 clknet_4_9_0_clk
rlabel metal3 820 7548 820 7548 0 dataBusIn[0]
rlabel metal2 29026 1588 29026 1588 0 dataBusIn[1]
rlabel metal1 38732 42194 38732 42194 0 dataBusIn[2]
rlabel metal2 40618 959 40618 959 0 dataBusIn[3]
rlabel metal1 31004 42194 31004 42194 0 dataBusIn[4]
rlabel metal1 9154 42262 9154 42262 0 dataBusIn[5]
rlabel metal3 820 11628 820 11628 0 dataBusIn[6]
rlabel metal1 41078 5678 41078 5678 0 dataBusIn[7]
rlabel metal2 40986 36941 40986 36941 0 dataBusOut[0]
rlabel metal2 21942 1571 21942 1571 0 dataBusOut[1]
rlabel metal3 751 15028 751 15028 0 dataBusOut[2]
rlabel metal2 40986 32623 40986 32623 0 dataBusOut[3]
rlabel metal2 32890 1095 32890 1095 0 dataBusOut[4]
rlabel metal2 7130 1520 7130 1520 0 dataBusOut[5]
rlabel via2 40986 40885 40986 40885 0 dataBusOut[6]
rlabel metal1 1472 42330 1472 42330 0 dataBusOut[7]
rlabel metal2 35098 43163 35098 43163 0 dataBusSelect
rlabel metal2 23874 42510 23874 42510 0 gpio[0]
rlabel metal2 3634 25823 3634 25823 0 gpio[10]
rlabel metal1 20700 41650 20700 41650 0 gpio[11]
rlabel metal2 3818 37825 3818 37825 0 gpio[12]
rlabel metal2 2806 30515 2806 30515 0 gpio[13]
rlabel metal2 5297 43996 5297 43996 0 gpio[14]
rlabel metal2 46 2132 46 2132 0 gpio[15]
rlabel metal3 820 3468 820 3468 0 gpio[16]
rlabel metal3 40856 29308 40856 29308 0 gpio[17]
rlabel metal1 14536 3434 14536 3434 0 gpio[18]
rlabel metal1 21850 25398 21850 25398 0 gpio[19]
rlabel metal2 36754 2098 36754 2098 0 gpio[1]
rlabel metal2 27685 43996 27685 43996 0 gpio[20]
rlabel metal3 39031 13396 39031 13396 0 gpio[21]
rlabel metal2 3266 1792 3266 1792 0 gpio[22]
rlabel metal2 10994 2336 10994 2336 0 gpio[23]
rlabel metal1 1564 34714 1564 34714 0 gpio[24]
rlabel metal1 18124 5610 18124 5610 0 gpio[2]
rlabel metal1 12742 30668 12742 30668 0 gpio[3]
rlabel metal2 41906 42612 41906 42612 0 gpio[4]
rlabel metal1 13616 41514 13616 41514 0 gpio[5]
rlabel metal2 16146 42782 16146 42782 0 gpio[6]
rlabel metal1 24840 6698 24840 6698 0 gpio[7]
rlabel metal3 2016 19108 2016 19108 0 gpio[8]
rlabel metal3 2062 42908 2062 42908 0 gpio[9]
rlabel viali 14214 21998 14214 21998 0 net1
rlabel metal2 40802 36788 40802 36788 0 net10
rlabel metal2 21114 6324 21114 6324 0 net11
rlabel metal1 3266 13906 3266 13906 0 net12
rlabel metal2 21390 32861 21390 32861 0 net13
rlabel metal1 31372 2414 31372 2414 0 net14
rlabel metal1 7222 6766 7222 6766 0 net15
rlabel metal2 40802 40630 40802 40630 0 net16
rlabel metal2 1518 40834 1518 40834 0 net17
rlabel metal1 34776 42194 34776 42194 0 net18
rlabel metal1 8004 29614 8004 29614 0 net19
rlabel metal2 16974 12716 16974 12716 0 net2
rlabel metal1 9890 24684 9890 24684 0 net20
rlabel metal2 12834 24327 12834 24327 0 net21
rlabel metal2 9890 23120 9890 23120 0 net22
rlabel metal1 21022 13362 21022 13362 0 net23
rlabel metal1 9499 21522 9499 21522 0 net24
rlabel metal1 13501 26962 13501 26962 0 net25
rlabel metal1 38456 13294 38456 13294 0 net26
rlabel metal1 22218 26962 22218 26962 0 net27
rlabel metal1 22310 27472 22310 27472 0 net28
rlabel metal1 29348 17578 29348 17578 0 net29
rlabel metal1 38088 42126 38088 42126 0 net3
rlabel metal1 21022 13158 21022 13158 0 net30
rlabel metal1 22402 14926 22402 14926 0 net31
rlabel metal1 22540 13158 22540 13158 0 net32
rlabel metal1 28474 5644 28474 5644 0 net33
rlabel metal2 5842 22440 5842 22440 0 net34
rlabel metal1 11454 20230 11454 20230 0 net35
rlabel metal1 9108 19686 9108 19686 0 net36
rlabel metal1 8786 19754 8786 19754 0 net37
rlabel metal1 18959 10710 18959 10710 0 net38
rlabel metal2 13938 20128 13938 20128 0 net39
rlabel metal2 40802 5168 40802 5168 0 net4
rlabel metal1 2951 30702 2951 30702 0 net40
rlabel metal2 10626 41457 10626 41457 0 net41
rlabel metal1 20891 41514 20891 41514 0 net42
rlabel metal1 18545 41582 18545 41582 0 net43
rlabel metal2 16928 21284 16928 21284 0 net44
rlabel metal2 22586 6188 22586 6188 0 net45
rlabel metal1 27791 4522 27791 4522 0 net46
rlabel metal1 32561 4522 32561 4522 0 net47
rlabel metal1 23835 41514 23835 41514 0 net48
rlabel metal2 40066 30838 40066 30838 0 net49
rlabel via3 31349 41412 31349 41412 0 net5
rlabel metal2 18262 19601 18262 19601 0 net50
rlabel metal2 41078 33252 41078 33252 0 net51
rlabel metal1 14398 5066 14398 5066 0 net52
rlabel metal1 19274 8534 19274 8534 0 net53
rlabel metal1 36202 5542 36202 5542 0 net54
rlabel metal1 22310 10064 22310 10064 0 net55
rlabel metal1 20286 30736 20286 30736 0 net56
rlabel metal1 19044 30770 19044 30770 0 net57
rlabel metal2 28382 8313 28382 8313 0 net58
rlabel metal1 32982 5202 32982 5202 0 net59
rlabel metal1 13846 16184 13846 16184 0 net6
rlabel metal2 26726 6528 26726 6528 0 net60
rlabel metal1 27876 9622 27876 9622 0 net61
rlabel metal2 21482 10370 21482 10370 0 net62
rlabel metal1 5014 13328 5014 13328 0 net63
rlabel metal1 22402 38828 22402 38828 0 net64
rlabel metal1 5934 18258 5934 18258 0 net65
rlabel metal2 2622 19958 2622 19958 0 net66
rlabel metal1 21298 7310 21298 7310 0 net67
rlabel metal1 8464 18938 8464 18938 0 net68
rlabel metal1 5750 9622 5750 9622 0 net69
rlabel metal2 1702 11492 1702 11492 0 net7
rlabel metal1 12466 17170 12466 17170 0 net70
rlabel metal1 4738 18666 4738 18666 0 net71
rlabel metal1 12834 17612 12834 17612 0 net72
rlabel metal1 26772 38998 26772 38998 0 net73
rlabel metal1 14306 11696 14306 11696 0 net74
rlabel metal1 10948 40426 10948 40426 0 net75
rlabel viali 7412 31790 7412 31790 0 net76
rlabel metal1 27784 7446 27784 7446 0 net77
rlabel metal1 7176 13974 7176 13974 0 net78
rlabel metal1 3864 14314 3864 14314 0 net79
rlabel metal1 18170 6766 18170 6766 0 net8
rlabel metal2 9338 16269 9338 16269 0 net80
rlabel metal1 3450 18258 3450 18258 0 net81
rlabel metal1 22862 35666 22862 35666 0 net82
rlabel metal1 8004 17306 8004 17306 0 net83
rlabel metal1 4416 38318 4416 38318 0 net84
rlabel metal1 20516 6426 20516 6426 0 net85
rlabel metal1 7222 6426 7222 6426 0 net86
rlabel metal1 6440 16082 6440 16082 0 net87
rlabel metal1 14858 34646 14858 34646 0 net88
rlabel metal1 3726 17170 3726 17170 0 net89
rlabel metal2 40802 26282 40802 26282 0 net9
rlabel metal2 15410 38488 15410 38488 0 net90
rlabel metal1 34960 6426 34960 6426 0 net91
rlabel metal1 5290 16490 5290 16490 0 net92
rlabel metal1 14674 23290 14674 23290 0 net93
rlabel metal1 15548 27370 15548 27370 0 net94
rlabel metal1 41262 21522 41262 21522 0 nrst
rlabel metal1 19504 17238 19504 17238 0 top8227.PSRCurrentValue\[0\]
rlabel metal2 33350 24463 33350 24463 0 top8227.PSRCurrentValue\[1\]
rlabel metal1 20976 9010 20976 9010 0 top8227.PSRCurrentValue\[2\]
rlabel metal1 13110 13702 13110 13702 0 top8227.PSRCurrentValue\[3\]
rlabel viali 19734 15062 19734 15062 0 top8227.PSRCurrentValue\[6\]
rlabel metal2 17342 20247 17342 20247 0 top8227.PSRCurrentValue\[7\]
rlabel metal1 20516 30158 20516 30158 0 top8227.branchBackward
rlabel metal1 20516 31110 20516 31110 0 top8227.branchForward
rlabel metal1 28244 5678 28244 5678 0 top8227.demux.isAddressing
rlabel metal1 18906 21590 18906 21590 0 top8227.demux.nmi
rlabel metal3 20769 19108 20769 19108 0 top8227.demux.reset
rlabel metal1 20654 20502 20654 20502 0 top8227.demux.setInterruptFlag
rlabel metal1 33442 5678 33442 5678 0 top8227.demux.state_machine.currentAddress\[0\]
rlabel metal1 27140 12818 27140 12818 0 top8227.demux.state_machine.currentAddress\[10\]
rlabel metal1 27876 9486 27876 9486 0 top8227.demux.state_machine.currentAddress\[11\]
rlabel metal1 25668 21590 25668 21590 0 top8227.demux.state_machine.currentAddress\[12\]
rlabel metal1 27232 14858 27232 14858 0 top8227.demux.state_machine.currentAddress\[1\]
rlabel metal2 34822 5678 34822 5678 0 top8227.demux.state_machine.currentAddress\[2\]
rlabel metal2 27002 8228 27002 8228 0 top8227.demux.state_machine.currentAddress\[3\]
rlabel metal1 26312 12818 26312 12818 0 top8227.demux.state_machine.currentAddress\[4\]
rlabel metal1 27232 13294 27232 13294 0 top8227.demux.state_machine.currentAddress\[5\]
rlabel metal2 25162 18853 25162 18853 0 top8227.demux.state_machine.currentAddress\[6\]
rlabel metal1 26312 11050 26312 11050 0 top8227.demux.state_machine.currentAddress\[7\]
rlabel metal1 36616 5678 36616 5678 0 top8227.demux.state_machine.currentAddress\[8\]
rlabel metal1 33810 5678 33810 5678 0 top8227.demux.state_machine.currentAddress\[9\]
rlabel metal1 39100 29614 39100 29614 0 top8227.demux.state_machine.currentInstruction\[0\]
rlabel metal1 39054 30736 39054 30736 0 top8227.demux.state_machine.currentInstruction\[1\]
rlabel metal2 38870 29512 38870 29512 0 top8227.demux.state_machine.currentInstruction\[2\]
rlabel metal1 38916 29818 38916 29818 0 top8227.demux.state_machine.currentInstruction\[3\]
rlabel metal1 39330 26248 39330 26248 0 top8227.demux.state_machine.currentInstruction\[4\]
rlabel metal1 39652 26282 39652 26282 0 top8227.demux.state_machine.currentInstruction\[5\]
rlabel metal1 31418 31790 31418 31790 0 top8227.demux.state_machine.timeState\[0\]
rlabel metal1 24932 33966 24932 33966 0 top8227.demux.state_machine.timeState\[1\]
rlabel metal2 30038 37468 30038 37468 0 top8227.demux.state_machine.timeState\[2\]
rlabel metal1 27462 38930 27462 38930 0 top8227.demux.state_machine.timeState\[3\]
rlabel metal1 28796 31790 28796 31790 0 top8227.demux.state_machine.timeState\[4\]
rlabel metal1 26220 37910 26220 37910 0 top8227.demux.state_machine.timeState\[5\]
rlabel metal1 29486 36142 29486 36142 0 top8227.demux.state_machine.timeState\[6\]
rlabel metal2 21344 12988 21344 12988 0 top8227.freeCarry
rlabel metal1 39376 32334 39376 32334 0 top8227.instructionLoader.interruptInjector.interruptRequest
rlabel metal1 20654 10030 20654 10030 0 top8227.instructionLoader.interruptInjector.irqGenerated
rlabel metal2 41032 32844 41032 32844 0 top8227.instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ
rlabel metal1 40572 32538 40572 32538 0 top8227.instructionLoader.interruptInjector.irqSync.nextQ2
rlabel metal1 19044 8806 19044 8806 0 top8227.instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning
rlabel metal2 17802 6324 17802 6324 0 top8227.instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI
rlabel metal1 2070 4250 2070 4250 0 top8227.instructionLoader.interruptInjector.nmiSync.in
rlabel metal1 6808 4794 6808 4794 0 top8227.instructionLoader.interruptInjector.nmiSync.nextQ2
rlabel via1 24127 9486 24127 9486 0 top8227.instructionLoader.interruptInjector.resetDetected
rlabel metal1 9844 20502 9844 20502 0 top8227.internalDataflow.accRegToDB\[0\]
rlabel metal1 14720 19822 14720 19822 0 top8227.internalDataflow.accRegToDB\[1\]
rlabel metal1 7820 24922 7820 24922 0 top8227.internalDataflow.accRegToDB\[2\]
rlabel metal2 13386 19516 13386 19516 0 top8227.internalDataflow.accRegToDB\[3\]
rlabel metal2 8326 25874 8326 25874 0 top8227.internalDataflow.accRegToDB\[4\]
rlabel metal1 3542 26350 3542 26350 0 top8227.internalDataflow.accRegToDB\[5\]
rlabel metal1 6394 24038 6394 24038 0 top8227.internalDataflow.accRegToDB\[6\]
rlabel metal1 5612 24038 5612 24038 0 top8227.internalDataflow.accRegToDB\[7\]
rlabel metal1 11592 41446 11592 41446 0 top8227.internalDataflow.addressHighBusModule.busInputs\[16\]
rlabel metal1 15180 38862 15180 38862 0 top8227.internalDataflow.addressHighBusModule.busInputs\[17\]
rlabel metal1 9200 38998 9200 38998 0 top8227.internalDataflow.addressHighBusModule.busInputs\[18\]
rlabel metal1 6348 38862 6348 38862 0 top8227.internalDataflow.addressHighBusModule.busInputs\[19\]
rlabel metal1 8004 36074 8004 36074 0 top8227.internalDataflow.addressHighBusModule.busInputs\[20\]
rlabel metal1 7544 34578 7544 34578 0 top8227.internalDataflow.addressHighBusModule.busInputs\[21\]
rlabel metal2 9200 27438 9200 27438 0 top8227.internalDataflow.addressHighBusModule.busInputs\[22\]
rlabel metal3 9798 26996 9798 26996 0 top8227.internalDataflow.addressHighBusModule.busInputs\[23\]
rlabel via1 20102 40358 20102 40358 0 top8227.internalDataflow.addressLowBusModule.busInputs\[16\]
rlabel metal1 20056 33966 20056 33966 0 top8227.internalDataflow.addressLowBusModule.busInputs\[17\]
rlabel metal1 16576 35666 16576 35666 0 top8227.internalDataflow.addressLowBusModule.busInputs\[18\]
rlabel metal1 16054 38998 16054 38998 0 top8227.internalDataflow.addressLowBusModule.busInputs\[19\]
rlabel metal1 7590 26894 7590 26894 0 top8227.internalDataflow.addressLowBusModule.busInputs\[20\]
rlabel metal1 13938 37196 13938 37196 0 top8227.internalDataflow.addressLowBusModule.busInputs\[21\]
rlabel metal1 13202 39304 13202 39304 0 top8227.internalDataflow.addressLowBusModule.busInputs\[22\]
rlabel metal1 18952 41582 18952 41582 0 top8227.internalDataflow.addressLowBusModule.busInputs\[23\]
rlabel metal2 14490 21624 14490 21624 0 top8227.internalDataflow.addressLowBusModule.busInputs\[24\]
rlabel metal2 16836 12818 16836 12818 0 top8227.internalDataflow.addressLowBusModule.busInputs\[25\]
rlabel metal2 7682 19907 7682 19907 0 top8227.internalDataflow.addressLowBusModule.busInputs\[26\]
rlabel metal2 13110 21216 13110 21216 0 top8227.internalDataflow.addressLowBusModule.busInputs\[27\]
rlabel metal1 8188 7310 8188 7310 0 top8227.internalDataflow.addressLowBusModule.busInputs\[28\]
rlabel metal1 5152 20434 5152 20434 0 top8227.internalDataflow.addressLowBusModule.busInputs\[29\]
rlabel metal2 5382 14535 5382 14535 0 top8227.internalDataflow.addressLowBusModule.busInputs\[30\]
rlabel metal1 5290 20944 5290 20944 0 top8227.internalDataflow.addressLowBusModule.busInputs\[31\]
rlabel metal1 12627 22678 12627 22678 0 top8227.internalDataflow.addressLowBusModule.busInputs\[32\]
rlabel metal1 15640 24854 15640 24854 0 top8227.internalDataflow.addressLowBusModule.busInputs\[33\]
rlabel metal1 7728 21658 7728 21658 0 top8227.internalDataflow.addressLowBusModule.busInputs\[34\]
rlabel metal2 12190 19686 12190 19686 0 top8227.internalDataflow.addressLowBusModule.busInputs\[35\]
rlabel metal1 5612 21998 5612 21998 0 top8227.internalDataflow.addressLowBusModule.busInputs\[36\]
rlabel metal1 5566 20400 5566 20400 0 top8227.internalDataflow.addressLowBusModule.busInputs\[37\]
rlabel metal1 5382 23052 5382 23052 0 top8227.internalDataflow.addressLowBusModule.busInputs\[38\]
rlabel metal1 5566 20944 5566 20944 0 top8227.internalDataflow.addressLowBusModule.busInputs\[39\]
rlabel metal1 18078 17102 18078 17102 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[0\]
rlabel metal1 16185 17850 16185 17850 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[1\]
rlabel metal1 17480 12818 17480 12818 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[2\]
rlabel metal1 16928 15062 16928 15062 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[3\]
rlabel metal1 18722 11832 18722 11832 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[6\]
rlabel metal1 9614 19788 9614 19788 0 top8227.internalDataflow.stackBusModule.busInputs\[32\]
rlabel metal1 14582 16218 14582 16218 0 top8227.internalDataflow.stackBusModule.busInputs\[33\]
rlabel metal1 8050 17646 8050 17646 0 top8227.internalDataflow.stackBusModule.busInputs\[34\]
rlabel metal1 12466 18632 12466 18632 0 top8227.internalDataflow.stackBusModule.busInputs\[35\]
rlabel metal1 6302 16014 6302 16014 0 top8227.internalDataflow.stackBusModule.busInputs\[36\]
rlabel metal1 5336 16626 5336 16626 0 top8227.internalDataflow.stackBusModule.busInputs\[37\]
rlabel metal1 3404 15470 3404 15470 0 top8227.internalDataflow.stackBusModule.busInputs\[38\]
rlabel metal1 3818 17102 3818 17102 0 top8227.internalDataflow.stackBusModule.busInputs\[39\]
rlabel via1 9798 18394 9798 18394 0 top8227.internalDataflow.stackBusModule.busInputs\[40\]
rlabel metal2 14490 18836 14490 18836 0 top8227.internalDataflow.stackBusModule.busInputs\[41\]
rlabel metal2 7866 19380 7866 19380 0 top8227.internalDataflow.stackBusModule.busInputs\[42\]
rlabel metal1 12650 17748 12650 17748 0 top8227.internalDataflow.stackBusModule.busInputs\[43\]
rlabel metal1 6026 18190 6026 18190 0 top8227.internalDataflow.stackBusModule.busInputs\[44\]
rlabel metal1 4968 19482 4968 19482 0 top8227.internalDataflow.stackBusModule.busInputs\[45\]
rlabel metal1 3680 20366 3680 20366 0 top8227.internalDataflow.stackBusModule.busInputs\[46\]
rlabel metal1 3772 18190 3772 18190 0 top8227.internalDataflow.stackBusModule.busInputs\[47\]
rlabel metal1 20240 14994 20240 14994 0 top8227.negEdgeDetector.q1
rlabel metal2 22034 38726 22034 38726 0 top8227.pulse_slower.currentEnableState\[0\]
rlabel metal1 22954 38998 22954 38998 0 top8227.pulse_slower.currentEnableState\[1\]
rlabel metal1 20240 35054 20240 35054 0 top8227.pulse_slower.nextEnableState\[0\]
rlabel metal1 21666 39474 21666 39474 0 top8227.pulse_slower.nextEnableState\[1\]
<< properties >>
string FIXED_BBOX 0 0 42549 44693
<< end >>
