// This is the unpowered netlist.
module top_asic (clk,
    reset,
    sigout,
    mode_out,
    pb);
 input clk;
 input reset;
 output sigout;
 output [1:0] mode_out;
 input [14:0] pb;

 wire \FSM.next_mode[0] ;
 wire \FSM.next_mode[1] ;
 wire \PWM.counter[0] ;
 wire \PWM.counter[1] ;
 wire \PWM.counter[2] ;
 wire \PWM.counter[3] ;
 wire \PWM.counter[4] ;
 wire \PWM.counter[5] ;
 wire \PWM.counter[6] ;
 wire \PWM.counter[7] ;
 wire \PWM.final_in[0] ;
 wire \PWM.final_in[1] ;
 wire \PWM.final_in[2] ;
 wire \PWM.final_in[3] ;
 wire \PWM.final_in[4] ;
 wire \PWM.final_in[5] ;
 wire \PWM.final_in[6] ;
 wire \PWM.final_in[7] ;
 wire \PWM.final_sample_in[0] ;
 wire \PWM.final_sample_in[1] ;
 wire \PWM.final_sample_in[2] ;
 wire \PWM.final_sample_in[3] ;
 wire \PWM.final_sample_in[4] ;
 wire \PWM.final_sample_in[5] ;
 wire \PWM.final_sample_in[6] ;
 wire \PWM.final_sample_in[7] ;
 wire \PWM.next_counter[0] ;
 wire \PWM.next_counter[1] ;
 wire \PWM.next_counter[2] ;
 wire \PWM.next_counter[3] ;
 wire \PWM.next_counter[4] ;
 wire \PWM.next_counter[5] ;
 wire \PWM.next_counter[6] ;
 wire \PWM.next_counter[7] ;
 wire \PWM.next_pwm_out ;
 wire \PWM.pwm_out ;
 wire \PWM.start ;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_9_clk;
 wire \freq_div.state[0] ;
 wire \freq_div.state[1] ;
 wire \freq_div.state[2] ;
 wire \genblk1[0].osc.clkdiv_C.cnt[0] ;
 wire \genblk1[0].osc.clkdiv_C.cnt[10] ;
 wire \genblk1[0].osc.clkdiv_C.cnt[11] ;
 wire \genblk1[0].osc.clkdiv_C.cnt[12] ;
 wire \genblk1[0].osc.clkdiv_C.cnt[13] ;
 wire \genblk1[0].osc.clkdiv_C.cnt[14] ;
 wire \genblk1[0].osc.clkdiv_C.cnt[15] ;
 wire \genblk1[0].osc.clkdiv_C.cnt[16] ;
 wire \genblk1[0].osc.clkdiv_C.cnt[17] ;
 wire \genblk1[0].osc.clkdiv_C.cnt[1] ;
 wire \genblk1[0].osc.clkdiv_C.cnt[2] ;
 wire \genblk1[0].osc.clkdiv_C.cnt[3] ;
 wire \genblk1[0].osc.clkdiv_C.cnt[4] ;
 wire \genblk1[0].osc.clkdiv_C.cnt[5] ;
 wire \genblk1[0].osc.clkdiv_C.cnt[6] ;
 wire \genblk1[0].osc.clkdiv_C.cnt[7] ;
 wire \genblk1[0].osc.clkdiv_C.cnt[8] ;
 wire \genblk1[0].osc.clkdiv_C.cnt[9] ;
 wire \genblk1[0].osc.clkdiv_C.next_cnt[0] ;
 wire \genblk1[0].osc.clkdiv_C.next_cnt[10] ;
 wire \genblk1[0].osc.clkdiv_C.next_cnt[11] ;
 wire \genblk1[0].osc.clkdiv_C.next_cnt[12] ;
 wire \genblk1[0].osc.clkdiv_C.next_cnt[13] ;
 wire \genblk1[0].osc.clkdiv_C.next_cnt[14] ;
 wire \genblk1[0].osc.clkdiv_C.next_cnt[15] ;
 wire \genblk1[0].osc.clkdiv_C.next_cnt[16] ;
 wire \genblk1[0].osc.clkdiv_C.next_cnt[17] ;
 wire \genblk1[0].osc.clkdiv_C.next_cnt[1] ;
 wire \genblk1[0].osc.clkdiv_C.next_cnt[2] ;
 wire \genblk1[0].osc.clkdiv_C.next_cnt[3] ;
 wire \genblk1[0].osc.clkdiv_C.next_cnt[4] ;
 wire \genblk1[0].osc.clkdiv_C.next_cnt[5] ;
 wire \genblk1[0].osc.clkdiv_C.next_cnt[6] ;
 wire \genblk1[0].osc.clkdiv_C.next_cnt[7] ;
 wire \genblk1[0].osc.clkdiv_C.next_cnt[8] ;
 wire \genblk1[0].osc.clkdiv_C.next_cnt[9] ;
 wire \genblk1[10].osc.clkdiv_C.cnt[0] ;
 wire \genblk1[10].osc.clkdiv_C.cnt[10] ;
 wire \genblk1[10].osc.clkdiv_C.cnt[11] ;
 wire \genblk1[10].osc.clkdiv_C.cnt[12] ;
 wire \genblk1[10].osc.clkdiv_C.cnt[13] ;
 wire \genblk1[10].osc.clkdiv_C.cnt[14] ;
 wire \genblk1[10].osc.clkdiv_C.cnt[15] ;
 wire \genblk1[10].osc.clkdiv_C.cnt[16] ;
 wire \genblk1[10].osc.clkdiv_C.cnt[17] ;
 wire \genblk1[10].osc.clkdiv_C.cnt[1] ;
 wire \genblk1[10].osc.clkdiv_C.cnt[2] ;
 wire \genblk1[10].osc.clkdiv_C.cnt[3] ;
 wire \genblk1[10].osc.clkdiv_C.cnt[4] ;
 wire \genblk1[10].osc.clkdiv_C.cnt[5] ;
 wire \genblk1[10].osc.clkdiv_C.cnt[6] ;
 wire \genblk1[10].osc.clkdiv_C.cnt[7] ;
 wire \genblk1[10].osc.clkdiv_C.cnt[8] ;
 wire \genblk1[10].osc.clkdiv_C.cnt[9] ;
 wire \genblk1[10].osc.clkdiv_C.next_cnt[0] ;
 wire \genblk1[10].osc.clkdiv_C.next_cnt[10] ;
 wire \genblk1[10].osc.clkdiv_C.next_cnt[11] ;
 wire \genblk1[10].osc.clkdiv_C.next_cnt[12] ;
 wire \genblk1[10].osc.clkdiv_C.next_cnt[13] ;
 wire \genblk1[10].osc.clkdiv_C.next_cnt[14] ;
 wire \genblk1[10].osc.clkdiv_C.next_cnt[15] ;
 wire \genblk1[10].osc.clkdiv_C.next_cnt[16] ;
 wire \genblk1[10].osc.clkdiv_C.next_cnt[17] ;
 wire \genblk1[10].osc.clkdiv_C.next_cnt[1] ;
 wire \genblk1[10].osc.clkdiv_C.next_cnt[2] ;
 wire \genblk1[10].osc.clkdiv_C.next_cnt[3] ;
 wire \genblk1[10].osc.clkdiv_C.next_cnt[4] ;
 wire \genblk1[10].osc.clkdiv_C.next_cnt[5] ;
 wire \genblk1[10].osc.clkdiv_C.next_cnt[6] ;
 wire \genblk1[10].osc.clkdiv_C.next_cnt[7] ;
 wire \genblk1[10].osc.clkdiv_C.next_cnt[8] ;
 wire \genblk1[10].osc.clkdiv_C.next_cnt[9] ;
 wire \genblk1[11].osc.clkdiv_C.cnt[0] ;
 wire \genblk1[11].osc.clkdiv_C.cnt[10] ;
 wire \genblk1[11].osc.clkdiv_C.cnt[11] ;
 wire \genblk1[11].osc.clkdiv_C.cnt[12] ;
 wire \genblk1[11].osc.clkdiv_C.cnt[13] ;
 wire \genblk1[11].osc.clkdiv_C.cnt[14] ;
 wire \genblk1[11].osc.clkdiv_C.cnt[15] ;
 wire \genblk1[11].osc.clkdiv_C.cnt[16] ;
 wire \genblk1[11].osc.clkdiv_C.cnt[17] ;
 wire \genblk1[11].osc.clkdiv_C.cnt[1] ;
 wire \genblk1[11].osc.clkdiv_C.cnt[2] ;
 wire \genblk1[11].osc.clkdiv_C.cnt[3] ;
 wire \genblk1[11].osc.clkdiv_C.cnt[4] ;
 wire \genblk1[11].osc.clkdiv_C.cnt[5] ;
 wire \genblk1[11].osc.clkdiv_C.cnt[6] ;
 wire \genblk1[11].osc.clkdiv_C.cnt[7] ;
 wire \genblk1[11].osc.clkdiv_C.cnt[8] ;
 wire \genblk1[11].osc.clkdiv_C.cnt[9] ;
 wire \genblk1[11].osc.clkdiv_C.next_cnt[0] ;
 wire \genblk1[11].osc.clkdiv_C.next_cnt[10] ;
 wire \genblk1[11].osc.clkdiv_C.next_cnt[11] ;
 wire \genblk1[11].osc.clkdiv_C.next_cnt[12] ;
 wire \genblk1[11].osc.clkdiv_C.next_cnt[13] ;
 wire \genblk1[11].osc.clkdiv_C.next_cnt[14] ;
 wire \genblk1[11].osc.clkdiv_C.next_cnt[15] ;
 wire \genblk1[11].osc.clkdiv_C.next_cnt[16] ;
 wire \genblk1[11].osc.clkdiv_C.next_cnt[17] ;
 wire \genblk1[11].osc.clkdiv_C.next_cnt[1] ;
 wire \genblk1[11].osc.clkdiv_C.next_cnt[2] ;
 wire \genblk1[11].osc.clkdiv_C.next_cnt[3] ;
 wire \genblk1[11].osc.clkdiv_C.next_cnt[4] ;
 wire \genblk1[11].osc.clkdiv_C.next_cnt[5] ;
 wire \genblk1[11].osc.clkdiv_C.next_cnt[6] ;
 wire \genblk1[11].osc.clkdiv_C.next_cnt[7] ;
 wire \genblk1[11].osc.clkdiv_C.next_cnt[8] ;
 wire \genblk1[11].osc.clkdiv_C.next_cnt[9] ;
 wire \genblk1[1].osc.clkdiv_C.cnt[0] ;
 wire \genblk1[1].osc.clkdiv_C.cnt[10] ;
 wire \genblk1[1].osc.clkdiv_C.cnt[11] ;
 wire \genblk1[1].osc.clkdiv_C.cnt[12] ;
 wire \genblk1[1].osc.clkdiv_C.cnt[13] ;
 wire \genblk1[1].osc.clkdiv_C.cnt[14] ;
 wire \genblk1[1].osc.clkdiv_C.cnt[15] ;
 wire \genblk1[1].osc.clkdiv_C.cnt[16] ;
 wire \genblk1[1].osc.clkdiv_C.cnt[17] ;
 wire \genblk1[1].osc.clkdiv_C.cnt[1] ;
 wire \genblk1[1].osc.clkdiv_C.cnt[2] ;
 wire \genblk1[1].osc.clkdiv_C.cnt[3] ;
 wire \genblk1[1].osc.clkdiv_C.cnt[4] ;
 wire \genblk1[1].osc.clkdiv_C.cnt[5] ;
 wire \genblk1[1].osc.clkdiv_C.cnt[6] ;
 wire \genblk1[1].osc.clkdiv_C.cnt[7] ;
 wire \genblk1[1].osc.clkdiv_C.cnt[8] ;
 wire \genblk1[1].osc.clkdiv_C.cnt[9] ;
 wire \genblk1[1].osc.clkdiv_C.next_cnt[0] ;
 wire \genblk1[1].osc.clkdiv_C.next_cnt[10] ;
 wire \genblk1[1].osc.clkdiv_C.next_cnt[11] ;
 wire \genblk1[1].osc.clkdiv_C.next_cnt[12] ;
 wire \genblk1[1].osc.clkdiv_C.next_cnt[13] ;
 wire \genblk1[1].osc.clkdiv_C.next_cnt[14] ;
 wire \genblk1[1].osc.clkdiv_C.next_cnt[15] ;
 wire \genblk1[1].osc.clkdiv_C.next_cnt[16] ;
 wire \genblk1[1].osc.clkdiv_C.next_cnt[17] ;
 wire \genblk1[1].osc.clkdiv_C.next_cnt[1] ;
 wire \genblk1[1].osc.clkdiv_C.next_cnt[2] ;
 wire \genblk1[1].osc.clkdiv_C.next_cnt[3] ;
 wire \genblk1[1].osc.clkdiv_C.next_cnt[4] ;
 wire \genblk1[1].osc.clkdiv_C.next_cnt[5] ;
 wire \genblk1[1].osc.clkdiv_C.next_cnt[6] ;
 wire \genblk1[1].osc.clkdiv_C.next_cnt[7] ;
 wire \genblk1[1].osc.clkdiv_C.next_cnt[8] ;
 wire \genblk1[1].osc.clkdiv_C.next_cnt[9] ;
 wire \genblk1[2].osc.clkdiv_C.cnt[0] ;
 wire \genblk1[2].osc.clkdiv_C.cnt[10] ;
 wire \genblk1[2].osc.clkdiv_C.cnt[11] ;
 wire \genblk1[2].osc.clkdiv_C.cnt[12] ;
 wire \genblk1[2].osc.clkdiv_C.cnt[13] ;
 wire \genblk1[2].osc.clkdiv_C.cnt[14] ;
 wire \genblk1[2].osc.clkdiv_C.cnt[15] ;
 wire \genblk1[2].osc.clkdiv_C.cnt[16] ;
 wire \genblk1[2].osc.clkdiv_C.cnt[17] ;
 wire \genblk1[2].osc.clkdiv_C.cnt[1] ;
 wire \genblk1[2].osc.clkdiv_C.cnt[2] ;
 wire \genblk1[2].osc.clkdiv_C.cnt[3] ;
 wire \genblk1[2].osc.clkdiv_C.cnt[4] ;
 wire \genblk1[2].osc.clkdiv_C.cnt[5] ;
 wire \genblk1[2].osc.clkdiv_C.cnt[6] ;
 wire \genblk1[2].osc.clkdiv_C.cnt[7] ;
 wire \genblk1[2].osc.clkdiv_C.cnt[8] ;
 wire \genblk1[2].osc.clkdiv_C.cnt[9] ;
 wire \genblk1[2].osc.clkdiv_C.next_cnt[0] ;
 wire \genblk1[2].osc.clkdiv_C.next_cnt[10] ;
 wire \genblk1[2].osc.clkdiv_C.next_cnt[11] ;
 wire \genblk1[2].osc.clkdiv_C.next_cnt[12] ;
 wire \genblk1[2].osc.clkdiv_C.next_cnt[13] ;
 wire \genblk1[2].osc.clkdiv_C.next_cnt[14] ;
 wire \genblk1[2].osc.clkdiv_C.next_cnt[15] ;
 wire \genblk1[2].osc.clkdiv_C.next_cnt[16] ;
 wire \genblk1[2].osc.clkdiv_C.next_cnt[17] ;
 wire \genblk1[2].osc.clkdiv_C.next_cnt[1] ;
 wire \genblk1[2].osc.clkdiv_C.next_cnt[2] ;
 wire \genblk1[2].osc.clkdiv_C.next_cnt[3] ;
 wire \genblk1[2].osc.clkdiv_C.next_cnt[4] ;
 wire \genblk1[2].osc.clkdiv_C.next_cnt[5] ;
 wire \genblk1[2].osc.clkdiv_C.next_cnt[6] ;
 wire \genblk1[2].osc.clkdiv_C.next_cnt[7] ;
 wire \genblk1[2].osc.clkdiv_C.next_cnt[8] ;
 wire \genblk1[2].osc.clkdiv_C.next_cnt[9] ;
 wire \genblk1[3].osc.clkdiv_C.cnt[0] ;
 wire \genblk1[3].osc.clkdiv_C.cnt[10] ;
 wire \genblk1[3].osc.clkdiv_C.cnt[11] ;
 wire \genblk1[3].osc.clkdiv_C.cnt[12] ;
 wire \genblk1[3].osc.clkdiv_C.cnt[13] ;
 wire \genblk1[3].osc.clkdiv_C.cnt[14] ;
 wire \genblk1[3].osc.clkdiv_C.cnt[15] ;
 wire \genblk1[3].osc.clkdiv_C.cnt[16] ;
 wire \genblk1[3].osc.clkdiv_C.cnt[17] ;
 wire \genblk1[3].osc.clkdiv_C.cnt[1] ;
 wire \genblk1[3].osc.clkdiv_C.cnt[2] ;
 wire \genblk1[3].osc.clkdiv_C.cnt[3] ;
 wire \genblk1[3].osc.clkdiv_C.cnt[4] ;
 wire \genblk1[3].osc.clkdiv_C.cnt[5] ;
 wire \genblk1[3].osc.clkdiv_C.cnt[6] ;
 wire \genblk1[3].osc.clkdiv_C.cnt[7] ;
 wire \genblk1[3].osc.clkdiv_C.cnt[8] ;
 wire \genblk1[3].osc.clkdiv_C.cnt[9] ;
 wire \genblk1[3].osc.clkdiv_C.next_cnt[0] ;
 wire \genblk1[3].osc.clkdiv_C.next_cnt[10] ;
 wire \genblk1[3].osc.clkdiv_C.next_cnt[11] ;
 wire \genblk1[3].osc.clkdiv_C.next_cnt[12] ;
 wire \genblk1[3].osc.clkdiv_C.next_cnt[13] ;
 wire \genblk1[3].osc.clkdiv_C.next_cnt[14] ;
 wire \genblk1[3].osc.clkdiv_C.next_cnt[15] ;
 wire \genblk1[3].osc.clkdiv_C.next_cnt[16] ;
 wire \genblk1[3].osc.clkdiv_C.next_cnt[17] ;
 wire \genblk1[3].osc.clkdiv_C.next_cnt[1] ;
 wire \genblk1[3].osc.clkdiv_C.next_cnt[2] ;
 wire \genblk1[3].osc.clkdiv_C.next_cnt[3] ;
 wire \genblk1[3].osc.clkdiv_C.next_cnt[4] ;
 wire \genblk1[3].osc.clkdiv_C.next_cnt[5] ;
 wire \genblk1[3].osc.clkdiv_C.next_cnt[6] ;
 wire \genblk1[3].osc.clkdiv_C.next_cnt[7] ;
 wire \genblk1[3].osc.clkdiv_C.next_cnt[8] ;
 wire \genblk1[3].osc.clkdiv_C.next_cnt[9] ;
 wire \genblk1[4].osc.clkdiv_C.cnt[0] ;
 wire \genblk1[4].osc.clkdiv_C.cnt[10] ;
 wire \genblk1[4].osc.clkdiv_C.cnt[11] ;
 wire \genblk1[4].osc.clkdiv_C.cnt[12] ;
 wire \genblk1[4].osc.clkdiv_C.cnt[13] ;
 wire \genblk1[4].osc.clkdiv_C.cnt[14] ;
 wire \genblk1[4].osc.clkdiv_C.cnt[15] ;
 wire \genblk1[4].osc.clkdiv_C.cnt[16] ;
 wire \genblk1[4].osc.clkdiv_C.cnt[17] ;
 wire \genblk1[4].osc.clkdiv_C.cnt[1] ;
 wire \genblk1[4].osc.clkdiv_C.cnt[2] ;
 wire \genblk1[4].osc.clkdiv_C.cnt[3] ;
 wire \genblk1[4].osc.clkdiv_C.cnt[4] ;
 wire \genblk1[4].osc.clkdiv_C.cnt[5] ;
 wire \genblk1[4].osc.clkdiv_C.cnt[6] ;
 wire \genblk1[4].osc.clkdiv_C.cnt[7] ;
 wire \genblk1[4].osc.clkdiv_C.cnt[8] ;
 wire \genblk1[4].osc.clkdiv_C.cnt[9] ;
 wire \genblk1[4].osc.clkdiv_C.next_cnt[0] ;
 wire \genblk1[4].osc.clkdiv_C.next_cnt[10] ;
 wire \genblk1[4].osc.clkdiv_C.next_cnt[11] ;
 wire \genblk1[4].osc.clkdiv_C.next_cnt[12] ;
 wire \genblk1[4].osc.clkdiv_C.next_cnt[13] ;
 wire \genblk1[4].osc.clkdiv_C.next_cnt[14] ;
 wire \genblk1[4].osc.clkdiv_C.next_cnt[15] ;
 wire \genblk1[4].osc.clkdiv_C.next_cnt[16] ;
 wire \genblk1[4].osc.clkdiv_C.next_cnt[17] ;
 wire \genblk1[4].osc.clkdiv_C.next_cnt[1] ;
 wire \genblk1[4].osc.clkdiv_C.next_cnt[2] ;
 wire \genblk1[4].osc.clkdiv_C.next_cnt[3] ;
 wire \genblk1[4].osc.clkdiv_C.next_cnt[4] ;
 wire \genblk1[4].osc.clkdiv_C.next_cnt[5] ;
 wire \genblk1[4].osc.clkdiv_C.next_cnt[6] ;
 wire \genblk1[4].osc.clkdiv_C.next_cnt[7] ;
 wire \genblk1[4].osc.clkdiv_C.next_cnt[8] ;
 wire \genblk1[4].osc.clkdiv_C.next_cnt[9] ;
 wire \genblk1[5].osc.clkdiv_C.cnt[0] ;
 wire \genblk1[5].osc.clkdiv_C.cnt[10] ;
 wire \genblk1[5].osc.clkdiv_C.cnt[11] ;
 wire \genblk1[5].osc.clkdiv_C.cnt[12] ;
 wire \genblk1[5].osc.clkdiv_C.cnt[13] ;
 wire \genblk1[5].osc.clkdiv_C.cnt[14] ;
 wire \genblk1[5].osc.clkdiv_C.cnt[15] ;
 wire \genblk1[5].osc.clkdiv_C.cnt[16] ;
 wire \genblk1[5].osc.clkdiv_C.cnt[17] ;
 wire \genblk1[5].osc.clkdiv_C.cnt[1] ;
 wire \genblk1[5].osc.clkdiv_C.cnt[2] ;
 wire \genblk1[5].osc.clkdiv_C.cnt[3] ;
 wire \genblk1[5].osc.clkdiv_C.cnt[4] ;
 wire \genblk1[5].osc.clkdiv_C.cnt[5] ;
 wire \genblk1[5].osc.clkdiv_C.cnt[6] ;
 wire \genblk1[5].osc.clkdiv_C.cnt[7] ;
 wire \genblk1[5].osc.clkdiv_C.cnt[8] ;
 wire \genblk1[5].osc.clkdiv_C.cnt[9] ;
 wire \genblk1[5].osc.clkdiv_C.next_cnt[0] ;
 wire \genblk1[5].osc.clkdiv_C.next_cnt[10] ;
 wire \genblk1[5].osc.clkdiv_C.next_cnt[11] ;
 wire \genblk1[5].osc.clkdiv_C.next_cnt[12] ;
 wire \genblk1[5].osc.clkdiv_C.next_cnt[13] ;
 wire \genblk1[5].osc.clkdiv_C.next_cnt[14] ;
 wire \genblk1[5].osc.clkdiv_C.next_cnt[15] ;
 wire \genblk1[5].osc.clkdiv_C.next_cnt[16] ;
 wire \genblk1[5].osc.clkdiv_C.next_cnt[17] ;
 wire \genblk1[5].osc.clkdiv_C.next_cnt[1] ;
 wire \genblk1[5].osc.clkdiv_C.next_cnt[2] ;
 wire \genblk1[5].osc.clkdiv_C.next_cnt[3] ;
 wire \genblk1[5].osc.clkdiv_C.next_cnt[4] ;
 wire \genblk1[5].osc.clkdiv_C.next_cnt[5] ;
 wire \genblk1[5].osc.clkdiv_C.next_cnt[6] ;
 wire \genblk1[5].osc.clkdiv_C.next_cnt[7] ;
 wire \genblk1[5].osc.clkdiv_C.next_cnt[8] ;
 wire \genblk1[5].osc.clkdiv_C.next_cnt[9] ;
 wire \genblk1[6].osc.clkdiv_C.cnt[0] ;
 wire \genblk1[6].osc.clkdiv_C.cnt[10] ;
 wire \genblk1[6].osc.clkdiv_C.cnt[11] ;
 wire \genblk1[6].osc.clkdiv_C.cnt[12] ;
 wire \genblk1[6].osc.clkdiv_C.cnt[13] ;
 wire \genblk1[6].osc.clkdiv_C.cnt[14] ;
 wire \genblk1[6].osc.clkdiv_C.cnt[15] ;
 wire \genblk1[6].osc.clkdiv_C.cnt[16] ;
 wire \genblk1[6].osc.clkdiv_C.cnt[17] ;
 wire \genblk1[6].osc.clkdiv_C.cnt[1] ;
 wire \genblk1[6].osc.clkdiv_C.cnt[2] ;
 wire \genblk1[6].osc.clkdiv_C.cnt[3] ;
 wire \genblk1[6].osc.clkdiv_C.cnt[4] ;
 wire \genblk1[6].osc.clkdiv_C.cnt[5] ;
 wire \genblk1[6].osc.clkdiv_C.cnt[6] ;
 wire \genblk1[6].osc.clkdiv_C.cnt[7] ;
 wire \genblk1[6].osc.clkdiv_C.cnt[8] ;
 wire \genblk1[6].osc.clkdiv_C.cnt[9] ;
 wire \genblk1[6].osc.clkdiv_C.next_cnt[0] ;
 wire \genblk1[6].osc.clkdiv_C.next_cnt[10] ;
 wire \genblk1[6].osc.clkdiv_C.next_cnt[11] ;
 wire \genblk1[6].osc.clkdiv_C.next_cnt[12] ;
 wire \genblk1[6].osc.clkdiv_C.next_cnt[13] ;
 wire \genblk1[6].osc.clkdiv_C.next_cnt[14] ;
 wire \genblk1[6].osc.clkdiv_C.next_cnt[15] ;
 wire \genblk1[6].osc.clkdiv_C.next_cnt[16] ;
 wire \genblk1[6].osc.clkdiv_C.next_cnt[17] ;
 wire \genblk1[6].osc.clkdiv_C.next_cnt[1] ;
 wire \genblk1[6].osc.clkdiv_C.next_cnt[2] ;
 wire \genblk1[6].osc.clkdiv_C.next_cnt[3] ;
 wire \genblk1[6].osc.clkdiv_C.next_cnt[4] ;
 wire \genblk1[6].osc.clkdiv_C.next_cnt[5] ;
 wire \genblk1[6].osc.clkdiv_C.next_cnt[6] ;
 wire \genblk1[6].osc.clkdiv_C.next_cnt[7] ;
 wire \genblk1[6].osc.clkdiv_C.next_cnt[8] ;
 wire \genblk1[6].osc.clkdiv_C.next_cnt[9] ;
 wire \genblk1[7].osc.clkdiv_C.cnt[0] ;
 wire \genblk1[7].osc.clkdiv_C.cnt[10] ;
 wire \genblk1[7].osc.clkdiv_C.cnt[11] ;
 wire \genblk1[7].osc.clkdiv_C.cnt[12] ;
 wire \genblk1[7].osc.clkdiv_C.cnt[13] ;
 wire \genblk1[7].osc.clkdiv_C.cnt[14] ;
 wire \genblk1[7].osc.clkdiv_C.cnt[15] ;
 wire \genblk1[7].osc.clkdiv_C.cnt[16] ;
 wire \genblk1[7].osc.clkdiv_C.cnt[17] ;
 wire \genblk1[7].osc.clkdiv_C.cnt[1] ;
 wire \genblk1[7].osc.clkdiv_C.cnt[2] ;
 wire \genblk1[7].osc.clkdiv_C.cnt[3] ;
 wire \genblk1[7].osc.clkdiv_C.cnt[4] ;
 wire \genblk1[7].osc.clkdiv_C.cnt[5] ;
 wire \genblk1[7].osc.clkdiv_C.cnt[6] ;
 wire \genblk1[7].osc.clkdiv_C.cnt[7] ;
 wire \genblk1[7].osc.clkdiv_C.cnt[8] ;
 wire \genblk1[7].osc.clkdiv_C.cnt[9] ;
 wire \genblk1[7].osc.clkdiv_C.next_cnt[0] ;
 wire \genblk1[7].osc.clkdiv_C.next_cnt[10] ;
 wire \genblk1[7].osc.clkdiv_C.next_cnt[11] ;
 wire \genblk1[7].osc.clkdiv_C.next_cnt[12] ;
 wire \genblk1[7].osc.clkdiv_C.next_cnt[13] ;
 wire \genblk1[7].osc.clkdiv_C.next_cnt[14] ;
 wire \genblk1[7].osc.clkdiv_C.next_cnt[15] ;
 wire \genblk1[7].osc.clkdiv_C.next_cnt[16] ;
 wire \genblk1[7].osc.clkdiv_C.next_cnt[17] ;
 wire \genblk1[7].osc.clkdiv_C.next_cnt[1] ;
 wire \genblk1[7].osc.clkdiv_C.next_cnt[2] ;
 wire \genblk1[7].osc.clkdiv_C.next_cnt[3] ;
 wire \genblk1[7].osc.clkdiv_C.next_cnt[4] ;
 wire \genblk1[7].osc.clkdiv_C.next_cnt[5] ;
 wire \genblk1[7].osc.clkdiv_C.next_cnt[6] ;
 wire \genblk1[7].osc.clkdiv_C.next_cnt[7] ;
 wire \genblk1[7].osc.clkdiv_C.next_cnt[8] ;
 wire \genblk1[7].osc.clkdiv_C.next_cnt[9] ;
 wire \genblk1[8].osc.clkdiv_C.cnt[0] ;
 wire \genblk1[8].osc.clkdiv_C.cnt[10] ;
 wire \genblk1[8].osc.clkdiv_C.cnt[11] ;
 wire \genblk1[8].osc.clkdiv_C.cnt[12] ;
 wire \genblk1[8].osc.clkdiv_C.cnt[13] ;
 wire \genblk1[8].osc.clkdiv_C.cnt[14] ;
 wire \genblk1[8].osc.clkdiv_C.cnt[15] ;
 wire \genblk1[8].osc.clkdiv_C.cnt[16] ;
 wire \genblk1[8].osc.clkdiv_C.cnt[17] ;
 wire \genblk1[8].osc.clkdiv_C.cnt[1] ;
 wire \genblk1[8].osc.clkdiv_C.cnt[2] ;
 wire \genblk1[8].osc.clkdiv_C.cnt[3] ;
 wire \genblk1[8].osc.clkdiv_C.cnt[4] ;
 wire \genblk1[8].osc.clkdiv_C.cnt[5] ;
 wire \genblk1[8].osc.clkdiv_C.cnt[6] ;
 wire \genblk1[8].osc.clkdiv_C.cnt[7] ;
 wire \genblk1[8].osc.clkdiv_C.cnt[8] ;
 wire \genblk1[8].osc.clkdiv_C.cnt[9] ;
 wire \genblk1[8].osc.clkdiv_C.next_cnt[0] ;
 wire \genblk1[8].osc.clkdiv_C.next_cnt[10] ;
 wire \genblk1[8].osc.clkdiv_C.next_cnt[11] ;
 wire \genblk1[8].osc.clkdiv_C.next_cnt[12] ;
 wire \genblk1[8].osc.clkdiv_C.next_cnt[13] ;
 wire \genblk1[8].osc.clkdiv_C.next_cnt[14] ;
 wire \genblk1[8].osc.clkdiv_C.next_cnt[15] ;
 wire \genblk1[8].osc.clkdiv_C.next_cnt[16] ;
 wire \genblk1[8].osc.clkdiv_C.next_cnt[17] ;
 wire \genblk1[8].osc.clkdiv_C.next_cnt[1] ;
 wire \genblk1[8].osc.clkdiv_C.next_cnt[2] ;
 wire \genblk1[8].osc.clkdiv_C.next_cnt[3] ;
 wire \genblk1[8].osc.clkdiv_C.next_cnt[4] ;
 wire \genblk1[8].osc.clkdiv_C.next_cnt[5] ;
 wire \genblk1[8].osc.clkdiv_C.next_cnt[6] ;
 wire \genblk1[8].osc.clkdiv_C.next_cnt[7] ;
 wire \genblk1[8].osc.clkdiv_C.next_cnt[8] ;
 wire \genblk1[8].osc.clkdiv_C.next_cnt[9] ;
 wire \genblk1[9].osc.clkdiv_C.cnt[0] ;
 wire \genblk1[9].osc.clkdiv_C.cnt[10] ;
 wire \genblk1[9].osc.clkdiv_C.cnt[11] ;
 wire \genblk1[9].osc.clkdiv_C.cnt[12] ;
 wire \genblk1[9].osc.clkdiv_C.cnt[13] ;
 wire \genblk1[9].osc.clkdiv_C.cnt[14] ;
 wire \genblk1[9].osc.clkdiv_C.cnt[15] ;
 wire \genblk1[9].osc.clkdiv_C.cnt[16] ;
 wire \genblk1[9].osc.clkdiv_C.cnt[17] ;
 wire \genblk1[9].osc.clkdiv_C.cnt[1] ;
 wire \genblk1[9].osc.clkdiv_C.cnt[2] ;
 wire \genblk1[9].osc.clkdiv_C.cnt[3] ;
 wire \genblk1[9].osc.clkdiv_C.cnt[4] ;
 wire \genblk1[9].osc.clkdiv_C.cnt[5] ;
 wire \genblk1[9].osc.clkdiv_C.cnt[6] ;
 wire \genblk1[9].osc.clkdiv_C.cnt[7] ;
 wire \genblk1[9].osc.clkdiv_C.cnt[8] ;
 wire \genblk1[9].osc.clkdiv_C.cnt[9] ;
 wire \genblk1[9].osc.clkdiv_C.next_cnt[0] ;
 wire \genblk1[9].osc.clkdiv_C.next_cnt[10] ;
 wire \genblk1[9].osc.clkdiv_C.next_cnt[11] ;
 wire \genblk1[9].osc.clkdiv_C.next_cnt[12] ;
 wire \genblk1[9].osc.clkdiv_C.next_cnt[13] ;
 wire \genblk1[9].osc.clkdiv_C.next_cnt[14] ;
 wire \genblk1[9].osc.clkdiv_C.next_cnt[15] ;
 wire \genblk1[9].osc.clkdiv_C.next_cnt[16] ;
 wire \genblk1[9].osc.clkdiv_C.next_cnt[17] ;
 wire \genblk1[9].osc.clkdiv_C.next_cnt[1] ;
 wire \genblk1[9].osc.clkdiv_C.next_cnt[2] ;
 wire \genblk1[9].osc.clkdiv_C.next_cnt[3] ;
 wire \genblk1[9].osc.clkdiv_C.next_cnt[4] ;
 wire \genblk1[9].osc.clkdiv_C.next_cnt[5] ;
 wire \genblk1[9].osc.clkdiv_C.next_cnt[6] ;
 wire \genblk1[9].osc.clkdiv_C.next_cnt[7] ;
 wire \genblk1[9].osc.clkdiv_C.next_cnt[8] ;
 wire \genblk1[9].osc.clkdiv_C.next_cnt[9] ;
 wire \genblk2[0].wave_shpr.div.acc[0] ;
 wire \genblk2[0].wave_shpr.div.acc[10] ;
 wire \genblk2[0].wave_shpr.div.acc[11] ;
 wire \genblk2[0].wave_shpr.div.acc[12] ;
 wire \genblk2[0].wave_shpr.div.acc[13] ;
 wire \genblk2[0].wave_shpr.div.acc[14] ;
 wire \genblk2[0].wave_shpr.div.acc[15] ;
 wire \genblk2[0].wave_shpr.div.acc[16] ;
 wire \genblk2[0].wave_shpr.div.acc[17] ;
 wire \genblk2[0].wave_shpr.div.acc[18] ;
 wire \genblk2[0].wave_shpr.div.acc[19] ;
 wire \genblk2[0].wave_shpr.div.acc[1] ;
 wire \genblk2[0].wave_shpr.div.acc[20] ;
 wire \genblk2[0].wave_shpr.div.acc[21] ;
 wire \genblk2[0].wave_shpr.div.acc[22] ;
 wire \genblk2[0].wave_shpr.div.acc[23] ;
 wire \genblk2[0].wave_shpr.div.acc[24] ;
 wire \genblk2[0].wave_shpr.div.acc[25] ;
 wire \genblk2[0].wave_shpr.div.acc[26] ;
 wire \genblk2[0].wave_shpr.div.acc[2] ;
 wire \genblk2[0].wave_shpr.div.acc[3] ;
 wire \genblk2[0].wave_shpr.div.acc[4] ;
 wire \genblk2[0].wave_shpr.div.acc[5] ;
 wire \genblk2[0].wave_shpr.div.acc[6] ;
 wire \genblk2[0].wave_shpr.div.acc[7] ;
 wire \genblk2[0].wave_shpr.div.acc[8] ;
 wire \genblk2[0].wave_shpr.div.acc[9] ;
 wire \genblk2[0].wave_shpr.div.acc_next[0] ;
 wire \genblk2[0].wave_shpr.div.b1[0] ;
 wire \genblk2[0].wave_shpr.div.b1[10] ;
 wire \genblk2[0].wave_shpr.div.b1[11] ;
 wire \genblk2[0].wave_shpr.div.b1[12] ;
 wire \genblk2[0].wave_shpr.div.b1[13] ;
 wire \genblk2[0].wave_shpr.div.b1[14] ;
 wire \genblk2[0].wave_shpr.div.b1[15] ;
 wire \genblk2[0].wave_shpr.div.b1[16] ;
 wire \genblk2[0].wave_shpr.div.b1[17] ;
 wire \genblk2[0].wave_shpr.div.b1[1] ;
 wire \genblk2[0].wave_shpr.div.b1[2] ;
 wire \genblk2[0].wave_shpr.div.b1[3] ;
 wire \genblk2[0].wave_shpr.div.b1[4] ;
 wire \genblk2[0].wave_shpr.div.b1[5] ;
 wire \genblk2[0].wave_shpr.div.b1[6] ;
 wire \genblk2[0].wave_shpr.div.b1[7] ;
 wire \genblk2[0].wave_shpr.div.b1[8] ;
 wire \genblk2[0].wave_shpr.div.b1[9] ;
 wire \genblk2[0].wave_shpr.div.busy ;
 wire \genblk2[0].wave_shpr.div.done ;
 wire \genblk2[0].wave_shpr.div.fin_quo[0] ;
 wire \genblk2[0].wave_shpr.div.fin_quo[1] ;
 wire \genblk2[0].wave_shpr.div.fin_quo[2] ;
 wire \genblk2[0].wave_shpr.div.fin_quo[3] ;
 wire \genblk2[0].wave_shpr.div.fin_quo[4] ;
 wire \genblk2[0].wave_shpr.div.fin_quo[5] ;
 wire \genblk2[0].wave_shpr.div.fin_quo[6] ;
 wire \genblk2[0].wave_shpr.div.fin_quo[7] ;
 wire \genblk2[0].wave_shpr.div.i[0] ;
 wire \genblk2[0].wave_shpr.div.i[1] ;
 wire \genblk2[0].wave_shpr.div.i[2] ;
 wire \genblk2[0].wave_shpr.div.i[3] ;
 wire \genblk2[0].wave_shpr.div.i[4] ;
 wire \genblk2[0].wave_shpr.div.quo[0] ;
 wire \genblk2[0].wave_shpr.div.quo[10] ;
 wire \genblk2[0].wave_shpr.div.quo[11] ;
 wire \genblk2[0].wave_shpr.div.quo[12] ;
 wire \genblk2[0].wave_shpr.div.quo[13] ;
 wire \genblk2[0].wave_shpr.div.quo[14] ;
 wire \genblk2[0].wave_shpr.div.quo[15] ;
 wire \genblk2[0].wave_shpr.div.quo[16] ;
 wire \genblk2[0].wave_shpr.div.quo[17] ;
 wire \genblk2[0].wave_shpr.div.quo[18] ;
 wire \genblk2[0].wave_shpr.div.quo[19] ;
 wire \genblk2[0].wave_shpr.div.quo[1] ;
 wire \genblk2[0].wave_shpr.div.quo[20] ;
 wire \genblk2[0].wave_shpr.div.quo[21] ;
 wire \genblk2[0].wave_shpr.div.quo[22] ;
 wire \genblk2[0].wave_shpr.div.quo[23] ;
 wire \genblk2[0].wave_shpr.div.quo[24] ;
 wire \genblk2[0].wave_shpr.div.quo[2] ;
 wire \genblk2[0].wave_shpr.div.quo[3] ;
 wire \genblk2[0].wave_shpr.div.quo[4] ;
 wire \genblk2[0].wave_shpr.div.quo[5] ;
 wire \genblk2[0].wave_shpr.div.quo[6] ;
 wire \genblk2[0].wave_shpr.div.quo[7] ;
 wire \genblk2[0].wave_shpr.div.quo[8] ;
 wire \genblk2[0].wave_shpr.div.quo[9] ;
 wire \genblk2[0].wave_shpr.div.start ;
 wire \genblk2[10].wave_shpr.div.acc[0] ;
 wire \genblk2[10].wave_shpr.div.acc[10] ;
 wire \genblk2[10].wave_shpr.div.acc[11] ;
 wire \genblk2[10].wave_shpr.div.acc[12] ;
 wire \genblk2[10].wave_shpr.div.acc[13] ;
 wire \genblk2[10].wave_shpr.div.acc[14] ;
 wire \genblk2[10].wave_shpr.div.acc[15] ;
 wire \genblk2[10].wave_shpr.div.acc[16] ;
 wire \genblk2[10].wave_shpr.div.acc[17] ;
 wire \genblk2[10].wave_shpr.div.acc[18] ;
 wire \genblk2[10].wave_shpr.div.acc[19] ;
 wire \genblk2[10].wave_shpr.div.acc[1] ;
 wire \genblk2[10].wave_shpr.div.acc[20] ;
 wire \genblk2[10].wave_shpr.div.acc[21] ;
 wire \genblk2[10].wave_shpr.div.acc[22] ;
 wire \genblk2[10].wave_shpr.div.acc[23] ;
 wire \genblk2[10].wave_shpr.div.acc[24] ;
 wire \genblk2[10].wave_shpr.div.acc[25] ;
 wire \genblk2[10].wave_shpr.div.acc[26] ;
 wire \genblk2[10].wave_shpr.div.acc[2] ;
 wire \genblk2[10].wave_shpr.div.acc[3] ;
 wire \genblk2[10].wave_shpr.div.acc[4] ;
 wire \genblk2[10].wave_shpr.div.acc[5] ;
 wire \genblk2[10].wave_shpr.div.acc[6] ;
 wire \genblk2[10].wave_shpr.div.acc[7] ;
 wire \genblk2[10].wave_shpr.div.acc[8] ;
 wire \genblk2[10].wave_shpr.div.acc[9] ;
 wire \genblk2[10].wave_shpr.div.acc_next[0] ;
 wire \genblk2[10].wave_shpr.div.b1[0] ;
 wire \genblk2[10].wave_shpr.div.b1[10] ;
 wire \genblk2[10].wave_shpr.div.b1[11] ;
 wire \genblk2[10].wave_shpr.div.b1[12] ;
 wire \genblk2[10].wave_shpr.div.b1[13] ;
 wire \genblk2[10].wave_shpr.div.b1[14] ;
 wire \genblk2[10].wave_shpr.div.b1[15] ;
 wire \genblk2[10].wave_shpr.div.b1[16] ;
 wire \genblk2[10].wave_shpr.div.b1[17] ;
 wire \genblk2[10].wave_shpr.div.b1[1] ;
 wire \genblk2[10].wave_shpr.div.b1[2] ;
 wire \genblk2[10].wave_shpr.div.b1[3] ;
 wire \genblk2[10].wave_shpr.div.b1[4] ;
 wire \genblk2[10].wave_shpr.div.b1[5] ;
 wire \genblk2[10].wave_shpr.div.b1[6] ;
 wire \genblk2[10].wave_shpr.div.b1[7] ;
 wire \genblk2[10].wave_shpr.div.b1[8] ;
 wire \genblk2[10].wave_shpr.div.b1[9] ;
 wire \genblk2[10].wave_shpr.div.busy ;
 wire \genblk2[10].wave_shpr.div.done ;
 wire \genblk2[10].wave_shpr.div.fin_quo[0] ;
 wire \genblk2[10].wave_shpr.div.fin_quo[1] ;
 wire \genblk2[10].wave_shpr.div.fin_quo[2] ;
 wire \genblk2[10].wave_shpr.div.fin_quo[3] ;
 wire \genblk2[10].wave_shpr.div.fin_quo[4] ;
 wire \genblk2[10].wave_shpr.div.fin_quo[5] ;
 wire \genblk2[10].wave_shpr.div.fin_quo[6] ;
 wire \genblk2[10].wave_shpr.div.fin_quo[7] ;
 wire \genblk2[10].wave_shpr.div.i[0] ;
 wire \genblk2[10].wave_shpr.div.i[1] ;
 wire \genblk2[10].wave_shpr.div.i[2] ;
 wire \genblk2[10].wave_shpr.div.i[3] ;
 wire \genblk2[10].wave_shpr.div.i[4] ;
 wire \genblk2[10].wave_shpr.div.quo[0] ;
 wire \genblk2[10].wave_shpr.div.quo[10] ;
 wire \genblk2[10].wave_shpr.div.quo[11] ;
 wire \genblk2[10].wave_shpr.div.quo[12] ;
 wire \genblk2[10].wave_shpr.div.quo[13] ;
 wire \genblk2[10].wave_shpr.div.quo[14] ;
 wire \genblk2[10].wave_shpr.div.quo[15] ;
 wire \genblk2[10].wave_shpr.div.quo[16] ;
 wire \genblk2[10].wave_shpr.div.quo[17] ;
 wire \genblk2[10].wave_shpr.div.quo[18] ;
 wire \genblk2[10].wave_shpr.div.quo[19] ;
 wire \genblk2[10].wave_shpr.div.quo[1] ;
 wire \genblk2[10].wave_shpr.div.quo[20] ;
 wire \genblk2[10].wave_shpr.div.quo[21] ;
 wire \genblk2[10].wave_shpr.div.quo[22] ;
 wire \genblk2[10].wave_shpr.div.quo[23] ;
 wire \genblk2[10].wave_shpr.div.quo[24] ;
 wire \genblk2[10].wave_shpr.div.quo[2] ;
 wire \genblk2[10].wave_shpr.div.quo[3] ;
 wire \genblk2[10].wave_shpr.div.quo[4] ;
 wire \genblk2[10].wave_shpr.div.quo[5] ;
 wire \genblk2[10].wave_shpr.div.quo[6] ;
 wire \genblk2[10].wave_shpr.div.quo[7] ;
 wire \genblk2[10].wave_shpr.div.quo[8] ;
 wire \genblk2[10].wave_shpr.div.quo[9] ;
 wire \genblk2[11].wave_shpr.div.acc[0] ;
 wire \genblk2[11].wave_shpr.div.acc[10] ;
 wire \genblk2[11].wave_shpr.div.acc[11] ;
 wire \genblk2[11].wave_shpr.div.acc[12] ;
 wire \genblk2[11].wave_shpr.div.acc[13] ;
 wire \genblk2[11].wave_shpr.div.acc[14] ;
 wire \genblk2[11].wave_shpr.div.acc[15] ;
 wire \genblk2[11].wave_shpr.div.acc[16] ;
 wire \genblk2[11].wave_shpr.div.acc[17] ;
 wire \genblk2[11].wave_shpr.div.acc[18] ;
 wire \genblk2[11].wave_shpr.div.acc[19] ;
 wire \genblk2[11].wave_shpr.div.acc[1] ;
 wire \genblk2[11].wave_shpr.div.acc[20] ;
 wire \genblk2[11].wave_shpr.div.acc[21] ;
 wire \genblk2[11].wave_shpr.div.acc[22] ;
 wire \genblk2[11].wave_shpr.div.acc[23] ;
 wire \genblk2[11].wave_shpr.div.acc[24] ;
 wire \genblk2[11].wave_shpr.div.acc[25] ;
 wire \genblk2[11].wave_shpr.div.acc[26] ;
 wire \genblk2[11].wave_shpr.div.acc[2] ;
 wire \genblk2[11].wave_shpr.div.acc[3] ;
 wire \genblk2[11].wave_shpr.div.acc[4] ;
 wire \genblk2[11].wave_shpr.div.acc[5] ;
 wire \genblk2[11].wave_shpr.div.acc[6] ;
 wire \genblk2[11].wave_shpr.div.acc[7] ;
 wire \genblk2[11].wave_shpr.div.acc[8] ;
 wire \genblk2[11].wave_shpr.div.acc[9] ;
 wire \genblk2[11].wave_shpr.div.acc_next[0] ;
 wire \genblk2[11].wave_shpr.div.b1[0] ;
 wire \genblk2[11].wave_shpr.div.b1[10] ;
 wire \genblk2[11].wave_shpr.div.b1[11] ;
 wire \genblk2[11].wave_shpr.div.b1[12] ;
 wire \genblk2[11].wave_shpr.div.b1[13] ;
 wire \genblk2[11].wave_shpr.div.b1[14] ;
 wire \genblk2[11].wave_shpr.div.b1[15] ;
 wire \genblk2[11].wave_shpr.div.b1[16] ;
 wire \genblk2[11].wave_shpr.div.b1[17] ;
 wire \genblk2[11].wave_shpr.div.b1[1] ;
 wire \genblk2[11].wave_shpr.div.b1[2] ;
 wire \genblk2[11].wave_shpr.div.b1[3] ;
 wire \genblk2[11].wave_shpr.div.b1[4] ;
 wire \genblk2[11].wave_shpr.div.b1[5] ;
 wire \genblk2[11].wave_shpr.div.b1[6] ;
 wire \genblk2[11].wave_shpr.div.b1[7] ;
 wire \genblk2[11].wave_shpr.div.b1[8] ;
 wire \genblk2[11].wave_shpr.div.b1[9] ;
 wire \genblk2[11].wave_shpr.div.busy ;
 wire \genblk2[11].wave_shpr.div.done ;
 wire \genblk2[11].wave_shpr.div.fin_quo[0] ;
 wire \genblk2[11].wave_shpr.div.fin_quo[1] ;
 wire \genblk2[11].wave_shpr.div.fin_quo[2] ;
 wire \genblk2[11].wave_shpr.div.fin_quo[3] ;
 wire \genblk2[11].wave_shpr.div.fin_quo[4] ;
 wire \genblk2[11].wave_shpr.div.fin_quo[5] ;
 wire \genblk2[11].wave_shpr.div.fin_quo[6] ;
 wire \genblk2[11].wave_shpr.div.fin_quo[7] ;
 wire \genblk2[11].wave_shpr.div.i[0] ;
 wire \genblk2[11].wave_shpr.div.i[1] ;
 wire \genblk2[11].wave_shpr.div.i[2] ;
 wire \genblk2[11].wave_shpr.div.i[3] ;
 wire \genblk2[11].wave_shpr.div.i[4] ;
 wire \genblk2[11].wave_shpr.div.quo[0] ;
 wire \genblk2[11].wave_shpr.div.quo[10] ;
 wire \genblk2[11].wave_shpr.div.quo[11] ;
 wire \genblk2[11].wave_shpr.div.quo[12] ;
 wire \genblk2[11].wave_shpr.div.quo[13] ;
 wire \genblk2[11].wave_shpr.div.quo[14] ;
 wire \genblk2[11].wave_shpr.div.quo[15] ;
 wire \genblk2[11].wave_shpr.div.quo[16] ;
 wire \genblk2[11].wave_shpr.div.quo[17] ;
 wire \genblk2[11].wave_shpr.div.quo[18] ;
 wire \genblk2[11].wave_shpr.div.quo[19] ;
 wire \genblk2[11].wave_shpr.div.quo[1] ;
 wire \genblk2[11].wave_shpr.div.quo[20] ;
 wire \genblk2[11].wave_shpr.div.quo[21] ;
 wire \genblk2[11].wave_shpr.div.quo[22] ;
 wire \genblk2[11].wave_shpr.div.quo[23] ;
 wire \genblk2[11].wave_shpr.div.quo[24] ;
 wire \genblk2[11].wave_shpr.div.quo[2] ;
 wire \genblk2[11].wave_shpr.div.quo[3] ;
 wire \genblk2[11].wave_shpr.div.quo[4] ;
 wire \genblk2[11].wave_shpr.div.quo[5] ;
 wire \genblk2[11].wave_shpr.div.quo[6] ;
 wire \genblk2[11].wave_shpr.div.quo[7] ;
 wire \genblk2[11].wave_shpr.div.quo[8] ;
 wire \genblk2[11].wave_shpr.div.quo[9] ;
 wire \genblk2[1].wave_shpr.div.acc[0] ;
 wire \genblk2[1].wave_shpr.div.acc[10] ;
 wire \genblk2[1].wave_shpr.div.acc[11] ;
 wire \genblk2[1].wave_shpr.div.acc[12] ;
 wire \genblk2[1].wave_shpr.div.acc[13] ;
 wire \genblk2[1].wave_shpr.div.acc[14] ;
 wire \genblk2[1].wave_shpr.div.acc[15] ;
 wire \genblk2[1].wave_shpr.div.acc[16] ;
 wire \genblk2[1].wave_shpr.div.acc[17] ;
 wire \genblk2[1].wave_shpr.div.acc[18] ;
 wire \genblk2[1].wave_shpr.div.acc[19] ;
 wire \genblk2[1].wave_shpr.div.acc[1] ;
 wire \genblk2[1].wave_shpr.div.acc[20] ;
 wire \genblk2[1].wave_shpr.div.acc[21] ;
 wire \genblk2[1].wave_shpr.div.acc[22] ;
 wire \genblk2[1].wave_shpr.div.acc[23] ;
 wire \genblk2[1].wave_shpr.div.acc[24] ;
 wire \genblk2[1].wave_shpr.div.acc[25] ;
 wire \genblk2[1].wave_shpr.div.acc[26] ;
 wire \genblk2[1].wave_shpr.div.acc[2] ;
 wire \genblk2[1].wave_shpr.div.acc[3] ;
 wire \genblk2[1].wave_shpr.div.acc[4] ;
 wire \genblk2[1].wave_shpr.div.acc[5] ;
 wire \genblk2[1].wave_shpr.div.acc[6] ;
 wire \genblk2[1].wave_shpr.div.acc[7] ;
 wire \genblk2[1].wave_shpr.div.acc[8] ;
 wire \genblk2[1].wave_shpr.div.acc[9] ;
 wire \genblk2[1].wave_shpr.div.acc_next[0] ;
 wire \genblk2[1].wave_shpr.div.b1[0] ;
 wire \genblk2[1].wave_shpr.div.b1[10] ;
 wire \genblk2[1].wave_shpr.div.b1[11] ;
 wire \genblk2[1].wave_shpr.div.b1[12] ;
 wire \genblk2[1].wave_shpr.div.b1[13] ;
 wire \genblk2[1].wave_shpr.div.b1[14] ;
 wire \genblk2[1].wave_shpr.div.b1[15] ;
 wire \genblk2[1].wave_shpr.div.b1[16] ;
 wire \genblk2[1].wave_shpr.div.b1[17] ;
 wire \genblk2[1].wave_shpr.div.b1[1] ;
 wire \genblk2[1].wave_shpr.div.b1[2] ;
 wire \genblk2[1].wave_shpr.div.b1[3] ;
 wire \genblk2[1].wave_shpr.div.b1[4] ;
 wire \genblk2[1].wave_shpr.div.b1[5] ;
 wire \genblk2[1].wave_shpr.div.b1[6] ;
 wire \genblk2[1].wave_shpr.div.b1[7] ;
 wire \genblk2[1].wave_shpr.div.b1[8] ;
 wire \genblk2[1].wave_shpr.div.b1[9] ;
 wire \genblk2[1].wave_shpr.div.busy ;
 wire \genblk2[1].wave_shpr.div.done ;
 wire \genblk2[1].wave_shpr.div.fin_quo[0] ;
 wire \genblk2[1].wave_shpr.div.fin_quo[1] ;
 wire \genblk2[1].wave_shpr.div.fin_quo[2] ;
 wire \genblk2[1].wave_shpr.div.fin_quo[3] ;
 wire \genblk2[1].wave_shpr.div.fin_quo[4] ;
 wire \genblk2[1].wave_shpr.div.fin_quo[5] ;
 wire \genblk2[1].wave_shpr.div.fin_quo[6] ;
 wire \genblk2[1].wave_shpr.div.fin_quo[7] ;
 wire \genblk2[1].wave_shpr.div.i[0] ;
 wire \genblk2[1].wave_shpr.div.i[1] ;
 wire \genblk2[1].wave_shpr.div.i[2] ;
 wire \genblk2[1].wave_shpr.div.i[3] ;
 wire \genblk2[1].wave_shpr.div.i[4] ;
 wire \genblk2[1].wave_shpr.div.quo[0] ;
 wire \genblk2[1].wave_shpr.div.quo[10] ;
 wire \genblk2[1].wave_shpr.div.quo[11] ;
 wire \genblk2[1].wave_shpr.div.quo[12] ;
 wire \genblk2[1].wave_shpr.div.quo[13] ;
 wire \genblk2[1].wave_shpr.div.quo[14] ;
 wire \genblk2[1].wave_shpr.div.quo[15] ;
 wire \genblk2[1].wave_shpr.div.quo[16] ;
 wire \genblk2[1].wave_shpr.div.quo[17] ;
 wire \genblk2[1].wave_shpr.div.quo[18] ;
 wire \genblk2[1].wave_shpr.div.quo[19] ;
 wire \genblk2[1].wave_shpr.div.quo[1] ;
 wire \genblk2[1].wave_shpr.div.quo[20] ;
 wire \genblk2[1].wave_shpr.div.quo[21] ;
 wire \genblk2[1].wave_shpr.div.quo[22] ;
 wire \genblk2[1].wave_shpr.div.quo[23] ;
 wire \genblk2[1].wave_shpr.div.quo[24] ;
 wire \genblk2[1].wave_shpr.div.quo[2] ;
 wire \genblk2[1].wave_shpr.div.quo[3] ;
 wire \genblk2[1].wave_shpr.div.quo[4] ;
 wire \genblk2[1].wave_shpr.div.quo[5] ;
 wire \genblk2[1].wave_shpr.div.quo[6] ;
 wire \genblk2[1].wave_shpr.div.quo[7] ;
 wire \genblk2[1].wave_shpr.div.quo[8] ;
 wire \genblk2[1].wave_shpr.div.quo[9] ;
 wire \genblk2[2].wave_shpr.div.acc[0] ;
 wire \genblk2[2].wave_shpr.div.acc[10] ;
 wire \genblk2[2].wave_shpr.div.acc[11] ;
 wire \genblk2[2].wave_shpr.div.acc[12] ;
 wire \genblk2[2].wave_shpr.div.acc[13] ;
 wire \genblk2[2].wave_shpr.div.acc[14] ;
 wire \genblk2[2].wave_shpr.div.acc[15] ;
 wire \genblk2[2].wave_shpr.div.acc[16] ;
 wire \genblk2[2].wave_shpr.div.acc[17] ;
 wire \genblk2[2].wave_shpr.div.acc[18] ;
 wire \genblk2[2].wave_shpr.div.acc[19] ;
 wire \genblk2[2].wave_shpr.div.acc[1] ;
 wire \genblk2[2].wave_shpr.div.acc[20] ;
 wire \genblk2[2].wave_shpr.div.acc[21] ;
 wire \genblk2[2].wave_shpr.div.acc[22] ;
 wire \genblk2[2].wave_shpr.div.acc[23] ;
 wire \genblk2[2].wave_shpr.div.acc[24] ;
 wire \genblk2[2].wave_shpr.div.acc[25] ;
 wire \genblk2[2].wave_shpr.div.acc[26] ;
 wire \genblk2[2].wave_shpr.div.acc[2] ;
 wire \genblk2[2].wave_shpr.div.acc[3] ;
 wire \genblk2[2].wave_shpr.div.acc[4] ;
 wire \genblk2[2].wave_shpr.div.acc[5] ;
 wire \genblk2[2].wave_shpr.div.acc[6] ;
 wire \genblk2[2].wave_shpr.div.acc[7] ;
 wire \genblk2[2].wave_shpr.div.acc[8] ;
 wire \genblk2[2].wave_shpr.div.acc[9] ;
 wire \genblk2[2].wave_shpr.div.acc_next[0] ;
 wire \genblk2[2].wave_shpr.div.b1[0] ;
 wire \genblk2[2].wave_shpr.div.b1[10] ;
 wire \genblk2[2].wave_shpr.div.b1[11] ;
 wire \genblk2[2].wave_shpr.div.b1[12] ;
 wire \genblk2[2].wave_shpr.div.b1[13] ;
 wire \genblk2[2].wave_shpr.div.b1[14] ;
 wire \genblk2[2].wave_shpr.div.b1[15] ;
 wire \genblk2[2].wave_shpr.div.b1[16] ;
 wire \genblk2[2].wave_shpr.div.b1[17] ;
 wire \genblk2[2].wave_shpr.div.b1[1] ;
 wire \genblk2[2].wave_shpr.div.b1[2] ;
 wire \genblk2[2].wave_shpr.div.b1[3] ;
 wire \genblk2[2].wave_shpr.div.b1[4] ;
 wire \genblk2[2].wave_shpr.div.b1[5] ;
 wire \genblk2[2].wave_shpr.div.b1[6] ;
 wire \genblk2[2].wave_shpr.div.b1[7] ;
 wire \genblk2[2].wave_shpr.div.b1[8] ;
 wire \genblk2[2].wave_shpr.div.b1[9] ;
 wire \genblk2[2].wave_shpr.div.busy ;
 wire \genblk2[2].wave_shpr.div.done ;
 wire \genblk2[2].wave_shpr.div.fin_quo[0] ;
 wire \genblk2[2].wave_shpr.div.fin_quo[1] ;
 wire \genblk2[2].wave_shpr.div.fin_quo[2] ;
 wire \genblk2[2].wave_shpr.div.fin_quo[3] ;
 wire \genblk2[2].wave_shpr.div.fin_quo[4] ;
 wire \genblk2[2].wave_shpr.div.fin_quo[5] ;
 wire \genblk2[2].wave_shpr.div.fin_quo[6] ;
 wire \genblk2[2].wave_shpr.div.fin_quo[7] ;
 wire \genblk2[2].wave_shpr.div.i[0] ;
 wire \genblk2[2].wave_shpr.div.i[1] ;
 wire \genblk2[2].wave_shpr.div.i[2] ;
 wire \genblk2[2].wave_shpr.div.i[3] ;
 wire \genblk2[2].wave_shpr.div.i[4] ;
 wire \genblk2[2].wave_shpr.div.quo[0] ;
 wire \genblk2[2].wave_shpr.div.quo[10] ;
 wire \genblk2[2].wave_shpr.div.quo[11] ;
 wire \genblk2[2].wave_shpr.div.quo[12] ;
 wire \genblk2[2].wave_shpr.div.quo[13] ;
 wire \genblk2[2].wave_shpr.div.quo[14] ;
 wire \genblk2[2].wave_shpr.div.quo[15] ;
 wire \genblk2[2].wave_shpr.div.quo[16] ;
 wire \genblk2[2].wave_shpr.div.quo[17] ;
 wire \genblk2[2].wave_shpr.div.quo[18] ;
 wire \genblk2[2].wave_shpr.div.quo[19] ;
 wire \genblk2[2].wave_shpr.div.quo[1] ;
 wire \genblk2[2].wave_shpr.div.quo[20] ;
 wire \genblk2[2].wave_shpr.div.quo[21] ;
 wire \genblk2[2].wave_shpr.div.quo[22] ;
 wire \genblk2[2].wave_shpr.div.quo[23] ;
 wire \genblk2[2].wave_shpr.div.quo[24] ;
 wire \genblk2[2].wave_shpr.div.quo[2] ;
 wire \genblk2[2].wave_shpr.div.quo[3] ;
 wire \genblk2[2].wave_shpr.div.quo[4] ;
 wire \genblk2[2].wave_shpr.div.quo[5] ;
 wire \genblk2[2].wave_shpr.div.quo[6] ;
 wire \genblk2[2].wave_shpr.div.quo[7] ;
 wire \genblk2[2].wave_shpr.div.quo[8] ;
 wire \genblk2[2].wave_shpr.div.quo[9] ;
 wire \genblk2[3].wave_shpr.div.acc[0] ;
 wire \genblk2[3].wave_shpr.div.acc[10] ;
 wire \genblk2[3].wave_shpr.div.acc[11] ;
 wire \genblk2[3].wave_shpr.div.acc[12] ;
 wire \genblk2[3].wave_shpr.div.acc[13] ;
 wire \genblk2[3].wave_shpr.div.acc[14] ;
 wire \genblk2[3].wave_shpr.div.acc[15] ;
 wire \genblk2[3].wave_shpr.div.acc[16] ;
 wire \genblk2[3].wave_shpr.div.acc[17] ;
 wire \genblk2[3].wave_shpr.div.acc[18] ;
 wire \genblk2[3].wave_shpr.div.acc[19] ;
 wire \genblk2[3].wave_shpr.div.acc[1] ;
 wire \genblk2[3].wave_shpr.div.acc[20] ;
 wire \genblk2[3].wave_shpr.div.acc[21] ;
 wire \genblk2[3].wave_shpr.div.acc[22] ;
 wire \genblk2[3].wave_shpr.div.acc[23] ;
 wire \genblk2[3].wave_shpr.div.acc[24] ;
 wire \genblk2[3].wave_shpr.div.acc[25] ;
 wire \genblk2[3].wave_shpr.div.acc[26] ;
 wire \genblk2[3].wave_shpr.div.acc[2] ;
 wire \genblk2[3].wave_shpr.div.acc[3] ;
 wire \genblk2[3].wave_shpr.div.acc[4] ;
 wire \genblk2[3].wave_shpr.div.acc[5] ;
 wire \genblk2[3].wave_shpr.div.acc[6] ;
 wire \genblk2[3].wave_shpr.div.acc[7] ;
 wire \genblk2[3].wave_shpr.div.acc[8] ;
 wire \genblk2[3].wave_shpr.div.acc[9] ;
 wire \genblk2[3].wave_shpr.div.acc_next[0] ;
 wire \genblk2[3].wave_shpr.div.b1[0] ;
 wire \genblk2[3].wave_shpr.div.b1[10] ;
 wire \genblk2[3].wave_shpr.div.b1[11] ;
 wire \genblk2[3].wave_shpr.div.b1[12] ;
 wire \genblk2[3].wave_shpr.div.b1[13] ;
 wire \genblk2[3].wave_shpr.div.b1[14] ;
 wire \genblk2[3].wave_shpr.div.b1[15] ;
 wire \genblk2[3].wave_shpr.div.b1[16] ;
 wire \genblk2[3].wave_shpr.div.b1[17] ;
 wire \genblk2[3].wave_shpr.div.b1[1] ;
 wire \genblk2[3].wave_shpr.div.b1[2] ;
 wire \genblk2[3].wave_shpr.div.b1[3] ;
 wire \genblk2[3].wave_shpr.div.b1[4] ;
 wire \genblk2[3].wave_shpr.div.b1[5] ;
 wire \genblk2[3].wave_shpr.div.b1[6] ;
 wire \genblk2[3].wave_shpr.div.b1[7] ;
 wire \genblk2[3].wave_shpr.div.b1[8] ;
 wire \genblk2[3].wave_shpr.div.b1[9] ;
 wire \genblk2[3].wave_shpr.div.busy ;
 wire \genblk2[3].wave_shpr.div.done ;
 wire \genblk2[3].wave_shpr.div.fin_quo[0] ;
 wire \genblk2[3].wave_shpr.div.fin_quo[1] ;
 wire \genblk2[3].wave_shpr.div.fin_quo[2] ;
 wire \genblk2[3].wave_shpr.div.fin_quo[3] ;
 wire \genblk2[3].wave_shpr.div.fin_quo[4] ;
 wire \genblk2[3].wave_shpr.div.fin_quo[5] ;
 wire \genblk2[3].wave_shpr.div.fin_quo[6] ;
 wire \genblk2[3].wave_shpr.div.fin_quo[7] ;
 wire \genblk2[3].wave_shpr.div.i[0] ;
 wire \genblk2[3].wave_shpr.div.i[1] ;
 wire \genblk2[3].wave_shpr.div.i[2] ;
 wire \genblk2[3].wave_shpr.div.i[3] ;
 wire \genblk2[3].wave_shpr.div.i[4] ;
 wire \genblk2[3].wave_shpr.div.quo[0] ;
 wire \genblk2[3].wave_shpr.div.quo[10] ;
 wire \genblk2[3].wave_shpr.div.quo[11] ;
 wire \genblk2[3].wave_shpr.div.quo[12] ;
 wire \genblk2[3].wave_shpr.div.quo[13] ;
 wire \genblk2[3].wave_shpr.div.quo[14] ;
 wire \genblk2[3].wave_shpr.div.quo[15] ;
 wire \genblk2[3].wave_shpr.div.quo[16] ;
 wire \genblk2[3].wave_shpr.div.quo[17] ;
 wire \genblk2[3].wave_shpr.div.quo[18] ;
 wire \genblk2[3].wave_shpr.div.quo[19] ;
 wire \genblk2[3].wave_shpr.div.quo[1] ;
 wire \genblk2[3].wave_shpr.div.quo[20] ;
 wire \genblk2[3].wave_shpr.div.quo[21] ;
 wire \genblk2[3].wave_shpr.div.quo[22] ;
 wire \genblk2[3].wave_shpr.div.quo[23] ;
 wire \genblk2[3].wave_shpr.div.quo[24] ;
 wire \genblk2[3].wave_shpr.div.quo[2] ;
 wire \genblk2[3].wave_shpr.div.quo[3] ;
 wire \genblk2[3].wave_shpr.div.quo[4] ;
 wire \genblk2[3].wave_shpr.div.quo[5] ;
 wire \genblk2[3].wave_shpr.div.quo[6] ;
 wire \genblk2[3].wave_shpr.div.quo[7] ;
 wire \genblk2[3].wave_shpr.div.quo[8] ;
 wire \genblk2[3].wave_shpr.div.quo[9] ;
 wire \genblk2[4].wave_shpr.div.acc[0] ;
 wire \genblk2[4].wave_shpr.div.acc[10] ;
 wire \genblk2[4].wave_shpr.div.acc[11] ;
 wire \genblk2[4].wave_shpr.div.acc[12] ;
 wire \genblk2[4].wave_shpr.div.acc[13] ;
 wire \genblk2[4].wave_shpr.div.acc[14] ;
 wire \genblk2[4].wave_shpr.div.acc[15] ;
 wire \genblk2[4].wave_shpr.div.acc[16] ;
 wire \genblk2[4].wave_shpr.div.acc[17] ;
 wire \genblk2[4].wave_shpr.div.acc[18] ;
 wire \genblk2[4].wave_shpr.div.acc[19] ;
 wire \genblk2[4].wave_shpr.div.acc[1] ;
 wire \genblk2[4].wave_shpr.div.acc[20] ;
 wire \genblk2[4].wave_shpr.div.acc[21] ;
 wire \genblk2[4].wave_shpr.div.acc[22] ;
 wire \genblk2[4].wave_shpr.div.acc[23] ;
 wire \genblk2[4].wave_shpr.div.acc[24] ;
 wire \genblk2[4].wave_shpr.div.acc[25] ;
 wire \genblk2[4].wave_shpr.div.acc[26] ;
 wire \genblk2[4].wave_shpr.div.acc[2] ;
 wire \genblk2[4].wave_shpr.div.acc[3] ;
 wire \genblk2[4].wave_shpr.div.acc[4] ;
 wire \genblk2[4].wave_shpr.div.acc[5] ;
 wire \genblk2[4].wave_shpr.div.acc[6] ;
 wire \genblk2[4].wave_shpr.div.acc[7] ;
 wire \genblk2[4].wave_shpr.div.acc[8] ;
 wire \genblk2[4].wave_shpr.div.acc[9] ;
 wire \genblk2[4].wave_shpr.div.acc_next[0] ;
 wire \genblk2[4].wave_shpr.div.b1[0] ;
 wire \genblk2[4].wave_shpr.div.b1[10] ;
 wire \genblk2[4].wave_shpr.div.b1[11] ;
 wire \genblk2[4].wave_shpr.div.b1[12] ;
 wire \genblk2[4].wave_shpr.div.b1[13] ;
 wire \genblk2[4].wave_shpr.div.b1[14] ;
 wire \genblk2[4].wave_shpr.div.b1[15] ;
 wire \genblk2[4].wave_shpr.div.b1[16] ;
 wire \genblk2[4].wave_shpr.div.b1[17] ;
 wire \genblk2[4].wave_shpr.div.b1[1] ;
 wire \genblk2[4].wave_shpr.div.b1[2] ;
 wire \genblk2[4].wave_shpr.div.b1[3] ;
 wire \genblk2[4].wave_shpr.div.b1[4] ;
 wire \genblk2[4].wave_shpr.div.b1[5] ;
 wire \genblk2[4].wave_shpr.div.b1[6] ;
 wire \genblk2[4].wave_shpr.div.b1[7] ;
 wire \genblk2[4].wave_shpr.div.b1[8] ;
 wire \genblk2[4].wave_shpr.div.b1[9] ;
 wire \genblk2[4].wave_shpr.div.busy ;
 wire \genblk2[4].wave_shpr.div.done ;
 wire \genblk2[4].wave_shpr.div.fin_quo[0] ;
 wire \genblk2[4].wave_shpr.div.fin_quo[1] ;
 wire \genblk2[4].wave_shpr.div.fin_quo[2] ;
 wire \genblk2[4].wave_shpr.div.fin_quo[3] ;
 wire \genblk2[4].wave_shpr.div.fin_quo[4] ;
 wire \genblk2[4].wave_shpr.div.fin_quo[5] ;
 wire \genblk2[4].wave_shpr.div.fin_quo[6] ;
 wire \genblk2[4].wave_shpr.div.fin_quo[7] ;
 wire \genblk2[4].wave_shpr.div.i[0] ;
 wire \genblk2[4].wave_shpr.div.i[1] ;
 wire \genblk2[4].wave_shpr.div.i[2] ;
 wire \genblk2[4].wave_shpr.div.i[3] ;
 wire \genblk2[4].wave_shpr.div.i[4] ;
 wire \genblk2[4].wave_shpr.div.quo[0] ;
 wire \genblk2[4].wave_shpr.div.quo[10] ;
 wire \genblk2[4].wave_shpr.div.quo[11] ;
 wire \genblk2[4].wave_shpr.div.quo[12] ;
 wire \genblk2[4].wave_shpr.div.quo[13] ;
 wire \genblk2[4].wave_shpr.div.quo[14] ;
 wire \genblk2[4].wave_shpr.div.quo[15] ;
 wire \genblk2[4].wave_shpr.div.quo[16] ;
 wire \genblk2[4].wave_shpr.div.quo[17] ;
 wire \genblk2[4].wave_shpr.div.quo[18] ;
 wire \genblk2[4].wave_shpr.div.quo[19] ;
 wire \genblk2[4].wave_shpr.div.quo[1] ;
 wire \genblk2[4].wave_shpr.div.quo[20] ;
 wire \genblk2[4].wave_shpr.div.quo[21] ;
 wire \genblk2[4].wave_shpr.div.quo[22] ;
 wire \genblk2[4].wave_shpr.div.quo[23] ;
 wire \genblk2[4].wave_shpr.div.quo[24] ;
 wire \genblk2[4].wave_shpr.div.quo[2] ;
 wire \genblk2[4].wave_shpr.div.quo[3] ;
 wire \genblk2[4].wave_shpr.div.quo[4] ;
 wire \genblk2[4].wave_shpr.div.quo[5] ;
 wire \genblk2[4].wave_shpr.div.quo[6] ;
 wire \genblk2[4].wave_shpr.div.quo[7] ;
 wire \genblk2[4].wave_shpr.div.quo[8] ;
 wire \genblk2[4].wave_shpr.div.quo[9] ;
 wire \genblk2[5].wave_shpr.div.acc[0] ;
 wire \genblk2[5].wave_shpr.div.acc[10] ;
 wire \genblk2[5].wave_shpr.div.acc[11] ;
 wire \genblk2[5].wave_shpr.div.acc[12] ;
 wire \genblk2[5].wave_shpr.div.acc[13] ;
 wire \genblk2[5].wave_shpr.div.acc[14] ;
 wire \genblk2[5].wave_shpr.div.acc[15] ;
 wire \genblk2[5].wave_shpr.div.acc[16] ;
 wire \genblk2[5].wave_shpr.div.acc[17] ;
 wire \genblk2[5].wave_shpr.div.acc[18] ;
 wire \genblk2[5].wave_shpr.div.acc[19] ;
 wire \genblk2[5].wave_shpr.div.acc[1] ;
 wire \genblk2[5].wave_shpr.div.acc[20] ;
 wire \genblk2[5].wave_shpr.div.acc[21] ;
 wire \genblk2[5].wave_shpr.div.acc[22] ;
 wire \genblk2[5].wave_shpr.div.acc[23] ;
 wire \genblk2[5].wave_shpr.div.acc[24] ;
 wire \genblk2[5].wave_shpr.div.acc[25] ;
 wire \genblk2[5].wave_shpr.div.acc[26] ;
 wire \genblk2[5].wave_shpr.div.acc[2] ;
 wire \genblk2[5].wave_shpr.div.acc[3] ;
 wire \genblk2[5].wave_shpr.div.acc[4] ;
 wire \genblk2[5].wave_shpr.div.acc[5] ;
 wire \genblk2[5].wave_shpr.div.acc[6] ;
 wire \genblk2[5].wave_shpr.div.acc[7] ;
 wire \genblk2[5].wave_shpr.div.acc[8] ;
 wire \genblk2[5].wave_shpr.div.acc[9] ;
 wire \genblk2[5].wave_shpr.div.acc_next[0] ;
 wire \genblk2[5].wave_shpr.div.b1[0] ;
 wire \genblk2[5].wave_shpr.div.b1[10] ;
 wire \genblk2[5].wave_shpr.div.b1[11] ;
 wire \genblk2[5].wave_shpr.div.b1[12] ;
 wire \genblk2[5].wave_shpr.div.b1[13] ;
 wire \genblk2[5].wave_shpr.div.b1[14] ;
 wire \genblk2[5].wave_shpr.div.b1[15] ;
 wire \genblk2[5].wave_shpr.div.b1[16] ;
 wire \genblk2[5].wave_shpr.div.b1[17] ;
 wire \genblk2[5].wave_shpr.div.b1[1] ;
 wire \genblk2[5].wave_shpr.div.b1[2] ;
 wire \genblk2[5].wave_shpr.div.b1[3] ;
 wire \genblk2[5].wave_shpr.div.b1[4] ;
 wire \genblk2[5].wave_shpr.div.b1[5] ;
 wire \genblk2[5].wave_shpr.div.b1[6] ;
 wire \genblk2[5].wave_shpr.div.b1[7] ;
 wire \genblk2[5].wave_shpr.div.b1[8] ;
 wire \genblk2[5].wave_shpr.div.b1[9] ;
 wire \genblk2[5].wave_shpr.div.busy ;
 wire \genblk2[5].wave_shpr.div.done ;
 wire \genblk2[5].wave_shpr.div.fin_quo[0] ;
 wire \genblk2[5].wave_shpr.div.fin_quo[1] ;
 wire \genblk2[5].wave_shpr.div.fin_quo[2] ;
 wire \genblk2[5].wave_shpr.div.fin_quo[3] ;
 wire \genblk2[5].wave_shpr.div.fin_quo[4] ;
 wire \genblk2[5].wave_shpr.div.fin_quo[5] ;
 wire \genblk2[5].wave_shpr.div.fin_quo[6] ;
 wire \genblk2[5].wave_shpr.div.fin_quo[7] ;
 wire \genblk2[5].wave_shpr.div.i[0] ;
 wire \genblk2[5].wave_shpr.div.i[1] ;
 wire \genblk2[5].wave_shpr.div.i[2] ;
 wire \genblk2[5].wave_shpr.div.i[3] ;
 wire \genblk2[5].wave_shpr.div.i[4] ;
 wire \genblk2[5].wave_shpr.div.quo[0] ;
 wire \genblk2[5].wave_shpr.div.quo[10] ;
 wire \genblk2[5].wave_shpr.div.quo[11] ;
 wire \genblk2[5].wave_shpr.div.quo[12] ;
 wire \genblk2[5].wave_shpr.div.quo[13] ;
 wire \genblk2[5].wave_shpr.div.quo[14] ;
 wire \genblk2[5].wave_shpr.div.quo[15] ;
 wire \genblk2[5].wave_shpr.div.quo[16] ;
 wire \genblk2[5].wave_shpr.div.quo[17] ;
 wire \genblk2[5].wave_shpr.div.quo[18] ;
 wire \genblk2[5].wave_shpr.div.quo[19] ;
 wire \genblk2[5].wave_shpr.div.quo[1] ;
 wire \genblk2[5].wave_shpr.div.quo[20] ;
 wire \genblk2[5].wave_shpr.div.quo[21] ;
 wire \genblk2[5].wave_shpr.div.quo[22] ;
 wire \genblk2[5].wave_shpr.div.quo[23] ;
 wire \genblk2[5].wave_shpr.div.quo[24] ;
 wire \genblk2[5].wave_shpr.div.quo[2] ;
 wire \genblk2[5].wave_shpr.div.quo[3] ;
 wire \genblk2[5].wave_shpr.div.quo[4] ;
 wire \genblk2[5].wave_shpr.div.quo[5] ;
 wire \genblk2[5].wave_shpr.div.quo[6] ;
 wire \genblk2[5].wave_shpr.div.quo[7] ;
 wire \genblk2[5].wave_shpr.div.quo[8] ;
 wire \genblk2[5].wave_shpr.div.quo[9] ;
 wire \genblk2[6].wave_shpr.div.acc[0] ;
 wire \genblk2[6].wave_shpr.div.acc[10] ;
 wire \genblk2[6].wave_shpr.div.acc[11] ;
 wire \genblk2[6].wave_shpr.div.acc[12] ;
 wire \genblk2[6].wave_shpr.div.acc[13] ;
 wire \genblk2[6].wave_shpr.div.acc[14] ;
 wire \genblk2[6].wave_shpr.div.acc[15] ;
 wire \genblk2[6].wave_shpr.div.acc[16] ;
 wire \genblk2[6].wave_shpr.div.acc[17] ;
 wire \genblk2[6].wave_shpr.div.acc[18] ;
 wire \genblk2[6].wave_shpr.div.acc[19] ;
 wire \genblk2[6].wave_shpr.div.acc[1] ;
 wire \genblk2[6].wave_shpr.div.acc[20] ;
 wire \genblk2[6].wave_shpr.div.acc[21] ;
 wire \genblk2[6].wave_shpr.div.acc[22] ;
 wire \genblk2[6].wave_shpr.div.acc[23] ;
 wire \genblk2[6].wave_shpr.div.acc[24] ;
 wire \genblk2[6].wave_shpr.div.acc[25] ;
 wire \genblk2[6].wave_shpr.div.acc[26] ;
 wire \genblk2[6].wave_shpr.div.acc[2] ;
 wire \genblk2[6].wave_shpr.div.acc[3] ;
 wire \genblk2[6].wave_shpr.div.acc[4] ;
 wire \genblk2[6].wave_shpr.div.acc[5] ;
 wire \genblk2[6].wave_shpr.div.acc[6] ;
 wire \genblk2[6].wave_shpr.div.acc[7] ;
 wire \genblk2[6].wave_shpr.div.acc[8] ;
 wire \genblk2[6].wave_shpr.div.acc[9] ;
 wire \genblk2[6].wave_shpr.div.acc_next[0] ;
 wire \genblk2[6].wave_shpr.div.b1[0] ;
 wire \genblk2[6].wave_shpr.div.b1[10] ;
 wire \genblk2[6].wave_shpr.div.b1[11] ;
 wire \genblk2[6].wave_shpr.div.b1[12] ;
 wire \genblk2[6].wave_shpr.div.b1[13] ;
 wire \genblk2[6].wave_shpr.div.b1[14] ;
 wire \genblk2[6].wave_shpr.div.b1[15] ;
 wire \genblk2[6].wave_shpr.div.b1[16] ;
 wire \genblk2[6].wave_shpr.div.b1[17] ;
 wire \genblk2[6].wave_shpr.div.b1[1] ;
 wire \genblk2[6].wave_shpr.div.b1[2] ;
 wire \genblk2[6].wave_shpr.div.b1[3] ;
 wire \genblk2[6].wave_shpr.div.b1[4] ;
 wire \genblk2[6].wave_shpr.div.b1[5] ;
 wire \genblk2[6].wave_shpr.div.b1[6] ;
 wire \genblk2[6].wave_shpr.div.b1[7] ;
 wire \genblk2[6].wave_shpr.div.b1[8] ;
 wire \genblk2[6].wave_shpr.div.b1[9] ;
 wire \genblk2[6].wave_shpr.div.busy ;
 wire \genblk2[6].wave_shpr.div.done ;
 wire \genblk2[6].wave_shpr.div.fin_quo[0] ;
 wire \genblk2[6].wave_shpr.div.fin_quo[1] ;
 wire \genblk2[6].wave_shpr.div.fin_quo[2] ;
 wire \genblk2[6].wave_shpr.div.fin_quo[3] ;
 wire \genblk2[6].wave_shpr.div.fin_quo[4] ;
 wire \genblk2[6].wave_shpr.div.fin_quo[5] ;
 wire \genblk2[6].wave_shpr.div.fin_quo[6] ;
 wire \genblk2[6].wave_shpr.div.fin_quo[7] ;
 wire \genblk2[6].wave_shpr.div.i[0] ;
 wire \genblk2[6].wave_shpr.div.i[1] ;
 wire \genblk2[6].wave_shpr.div.i[2] ;
 wire \genblk2[6].wave_shpr.div.i[3] ;
 wire \genblk2[6].wave_shpr.div.i[4] ;
 wire \genblk2[6].wave_shpr.div.quo[0] ;
 wire \genblk2[6].wave_shpr.div.quo[10] ;
 wire \genblk2[6].wave_shpr.div.quo[11] ;
 wire \genblk2[6].wave_shpr.div.quo[12] ;
 wire \genblk2[6].wave_shpr.div.quo[13] ;
 wire \genblk2[6].wave_shpr.div.quo[14] ;
 wire \genblk2[6].wave_shpr.div.quo[15] ;
 wire \genblk2[6].wave_shpr.div.quo[16] ;
 wire \genblk2[6].wave_shpr.div.quo[17] ;
 wire \genblk2[6].wave_shpr.div.quo[18] ;
 wire \genblk2[6].wave_shpr.div.quo[19] ;
 wire \genblk2[6].wave_shpr.div.quo[1] ;
 wire \genblk2[6].wave_shpr.div.quo[20] ;
 wire \genblk2[6].wave_shpr.div.quo[21] ;
 wire \genblk2[6].wave_shpr.div.quo[22] ;
 wire \genblk2[6].wave_shpr.div.quo[23] ;
 wire \genblk2[6].wave_shpr.div.quo[24] ;
 wire \genblk2[6].wave_shpr.div.quo[2] ;
 wire \genblk2[6].wave_shpr.div.quo[3] ;
 wire \genblk2[6].wave_shpr.div.quo[4] ;
 wire \genblk2[6].wave_shpr.div.quo[5] ;
 wire \genblk2[6].wave_shpr.div.quo[6] ;
 wire \genblk2[6].wave_shpr.div.quo[7] ;
 wire \genblk2[6].wave_shpr.div.quo[8] ;
 wire \genblk2[6].wave_shpr.div.quo[9] ;
 wire \genblk2[7].wave_shpr.div.acc[0] ;
 wire \genblk2[7].wave_shpr.div.acc[10] ;
 wire \genblk2[7].wave_shpr.div.acc[11] ;
 wire \genblk2[7].wave_shpr.div.acc[12] ;
 wire \genblk2[7].wave_shpr.div.acc[13] ;
 wire \genblk2[7].wave_shpr.div.acc[14] ;
 wire \genblk2[7].wave_shpr.div.acc[15] ;
 wire \genblk2[7].wave_shpr.div.acc[16] ;
 wire \genblk2[7].wave_shpr.div.acc[17] ;
 wire \genblk2[7].wave_shpr.div.acc[18] ;
 wire \genblk2[7].wave_shpr.div.acc[19] ;
 wire \genblk2[7].wave_shpr.div.acc[1] ;
 wire \genblk2[7].wave_shpr.div.acc[20] ;
 wire \genblk2[7].wave_shpr.div.acc[21] ;
 wire \genblk2[7].wave_shpr.div.acc[22] ;
 wire \genblk2[7].wave_shpr.div.acc[23] ;
 wire \genblk2[7].wave_shpr.div.acc[24] ;
 wire \genblk2[7].wave_shpr.div.acc[25] ;
 wire \genblk2[7].wave_shpr.div.acc[26] ;
 wire \genblk2[7].wave_shpr.div.acc[2] ;
 wire \genblk2[7].wave_shpr.div.acc[3] ;
 wire \genblk2[7].wave_shpr.div.acc[4] ;
 wire \genblk2[7].wave_shpr.div.acc[5] ;
 wire \genblk2[7].wave_shpr.div.acc[6] ;
 wire \genblk2[7].wave_shpr.div.acc[7] ;
 wire \genblk2[7].wave_shpr.div.acc[8] ;
 wire \genblk2[7].wave_shpr.div.acc[9] ;
 wire \genblk2[7].wave_shpr.div.acc_next[0] ;
 wire \genblk2[7].wave_shpr.div.b1[0] ;
 wire \genblk2[7].wave_shpr.div.b1[10] ;
 wire \genblk2[7].wave_shpr.div.b1[11] ;
 wire \genblk2[7].wave_shpr.div.b1[12] ;
 wire \genblk2[7].wave_shpr.div.b1[13] ;
 wire \genblk2[7].wave_shpr.div.b1[14] ;
 wire \genblk2[7].wave_shpr.div.b1[15] ;
 wire \genblk2[7].wave_shpr.div.b1[16] ;
 wire \genblk2[7].wave_shpr.div.b1[17] ;
 wire \genblk2[7].wave_shpr.div.b1[1] ;
 wire \genblk2[7].wave_shpr.div.b1[2] ;
 wire \genblk2[7].wave_shpr.div.b1[3] ;
 wire \genblk2[7].wave_shpr.div.b1[4] ;
 wire \genblk2[7].wave_shpr.div.b1[5] ;
 wire \genblk2[7].wave_shpr.div.b1[6] ;
 wire \genblk2[7].wave_shpr.div.b1[7] ;
 wire \genblk2[7].wave_shpr.div.b1[8] ;
 wire \genblk2[7].wave_shpr.div.b1[9] ;
 wire \genblk2[7].wave_shpr.div.busy ;
 wire \genblk2[7].wave_shpr.div.done ;
 wire \genblk2[7].wave_shpr.div.fin_quo[0] ;
 wire \genblk2[7].wave_shpr.div.fin_quo[1] ;
 wire \genblk2[7].wave_shpr.div.fin_quo[2] ;
 wire \genblk2[7].wave_shpr.div.fin_quo[3] ;
 wire \genblk2[7].wave_shpr.div.fin_quo[4] ;
 wire \genblk2[7].wave_shpr.div.fin_quo[5] ;
 wire \genblk2[7].wave_shpr.div.fin_quo[6] ;
 wire \genblk2[7].wave_shpr.div.fin_quo[7] ;
 wire \genblk2[7].wave_shpr.div.i[0] ;
 wire \genblk2[7].wave_shpr.div.i[1] ;
 wire \genblk2[7].wave_shpr.div.i[2] ;
 wire \genblk2[7].wave_shpr.div.i[3] ;
 wire \genblk2[7].wave_shpr.div.i[4] ;
 wire \genblk2[7].wave_shpr.div.quo[0] ;
 wire \genblk2[7].wave_shpr.div.quo[10] ;
 wire \genblk2[7].wave_shpr.div.quo[11] ;
 wire \genblk2[7].wave_shpr.div.quo[12] ;
 wire \genblk2[7].wave_shpr.div.quo[13] ;
 wire \genblk2[7].wave_shpr.div.quo[14] ;
 wire \genblk2[7].wave_shpr.div.quo[15] ;
 wire \genblk2[7].wave_shpr.div.quo[16] ;
 wire \genblk2[7].wave_shpr.div.quo[17] ;
 wire \genblk2[7].wave_shpr.div.quo[18] ;
 wire \genblk2[7].wave_shpr.div.quo[19] ;
 wire \genblk2[7].wave_shpr.div.quo[1] ;
 wire \genblk2[7].wave_shpr.div.quo[20] ;
 wire \genblk2[7].wave_shpr.div.quo[21] ;
 wire \genblk2[7].wave_shpr.div.quo[22] ;
 wire \genblk2[7].wave_shpr.div.quo[23] ;
 wire \genblk2[7].wave_shpr.div.quo[24] ;
 wire \genblk2[7].wave_shpr.div.quo[2] ;
 wire \genblk2[7].wave_shpr.div.quo[3] ;
 wire \genblk2[7].wave_shpr.div.quo[4] ;
 wire \genblk2[7].wave_shpr.div.quo[5] ;
 wire \genblk2[7].wave_shpr.div.quo[6] ;
 wire \genblk2[7].wave_shpr.div.quo[7] ;
 wire \genblk2[7].wave_shpr.div.quo[8] ;
 wire \genblk2[7].wave_shpr.div.quo[9] ;
 wire \genblk2[8].wave_shpr.div.acc[0] ;
 wire \genblk2[8].wave_shpr.div.acc[10] ;
 wire \genblk2[8].wave_shpr.div.acc[11] ;
 wire \genblk2[8].wave_shpr.div.acc[12] ;
 wire \genblk2[8].wave_shpr.div.acc[13] ;
 wire \genblk2[8].wave_shpr.div.acc[14] ;
 wire \genblk2[8].wave_shpr.div.acc[15] ;
 wire \genblk2[8].wave_shpr.div.acc[16] ;
 wire \genblk2[8].wave_shpr.div.acc[17] ;
 wire \genblk2[8].wave_shpr.div.acc[18] ;
 wire \genblk2[8].wave_shpr.div.acc[19] ;
 wire \genblk2[8].wave_shpr.div.acc[1] ;
 wire \genblk2[8].wave_shpr.div.acc[20] ;
 wire \genblk2[8].wave_shpr.div.acc[21] ;
 wire \genblk2[8].wave_shpr.div.acc[22] ;
 wire \genblk2[8].wave_shpr.div.acc[23] ;
 wire \genblk2[8].wave_shpr.div.acc[24] ;
 wire \genblk2[8].wave_shpr.div.acc[25] ;
 wire \genblk2[8].wave_shpr.div.acc[26] ;
 wire \genblk2[8].wave_shpr.div.acc[2] ;
 wire \genblk2[8].wave_shpr.div.acc[3] ;
 wire \genblk2[8].wave_shpr.div.acc[4] ;
 wire \genblk2[8].wave_shpr.div.acc[5] ;
 wire \genblk2[8].wave_shpr.div.acc[6] ;
 wire \genblk2[8].wave_shpr.div.acc[7] ;
 wire \genblk2[8].wave_shpr.div.acc[8] ;
 wire \genblk2[8].wave_shpr.div.acc[9] ;
 wire \genblk2[8].wave_shpr.div.acc_next[0] ;
 wire \genblk2[8].wave_shpr.div.b1[0] ;
 wire \genblk2[8].wave_shpr.div.b1[10] ;
 wire \genblk2[8].wave_shpr.div.b1[11] ;
 wire \genblk2[8].wave_shpr.div.b1[12] ;
 wire \genblk2[8].wave_shpr.div.b1[13] ;
 wire \genblk2[8].wave_shpr.div.b1[14] ;
 wire \genblk2[8].wave_shpr.div.b1[15] ;
 wire \genblk2[8].wave_shpr.div.b1[16] ;
 wire \genblk2[8].wave_shpr.div.b1[17] ;
 wire \genblk2[8].wave_shpr.div.b1[1] ;
 wire \genblk2[8].wave_shpr.div.b1[2] ;
 wire \genblk2[8].wave_shpr.div.b1[3] ;
 wire \genblk2[8].wave_shpr.div.b1[4] ;
 wire \genblk2[8].wave_shpr.div.b1[5] ;
 wire \genblk2[8].wave_shpr.div.b1[6] ;
 wire \genblk2[8].wave_shpr.div.b1[7] ;
 wire \genblk2[8].wave_shpr.div.b1[8] ;
 wire \genblk2[8].wave_shpr.div.b1[9] ;
 wire \genblk2[8].wave_shpr.div.busy ;
 wire \genblk2[8].wave_shpr.div.done ;
 wire \genblk2[8].wave_shpr.div.fin_quo[0] ;
 wire \genblk2[8].wave_shpr.div.fin_quo[1] ;
 wire \genblk2[8].wave_shpr.div.fin_quo[2] ;
 wire \genblk2[8].wave_shpr.div.fin_quo[3] ;
 wire \genblk2[8].wave_shpr.div.fin_quo[4] ;
 wire \genblk2[8].wave_shpr.div.fin_quo[5] ;
 wire \genblk2[8].wave_shpr.div.fin_quo[6] ;
 wire \genblk2[8].wave_shpr.div.fin_quo[7] ;
 wire \genblk2[8].wave_shpr.div.i[0] ;
 wire \genblk2[8].wave_shpr.div.i[1] ;
 wire \genblk2[8].wave_shpr.div.i[2] ;
 wire \genblk2[8].wave_shpr.div.i[3] ;
 wire \genblk2[8].wave_shpr.div.i[4] ;
 wire \genblk2[8].wave_shpr.div.quo[0] ;
 wire \genblk2[8].wave_shpr.div.quo[10] ;
 wire \genblk2[8].wave_shpr.div.quo[11] ;
 wire \genblk2[8].wave_shpr.div.quo[12] ;
 wire \genblk2[8].wave_shpr.div.quo[13] ;
 wire \genblk2[8].wave_shpr.div.quo[14] ;
 wire \genblk2[8].wave_shpr.div.quo[15] ;
 wire \genblk2[8].wave_shpr.div.quo[16] ;
 wire \genblk2[8].wave_shpr.div.quo[17] ;
 wire \genblk2[8].wave_shpr.div.quo[18] ;
 wire \genblk2[8].wave_shpr.div.quo[19] ;
 wire \genblk2[8].wave_shpr.div.quo[1] ;
 wire \genblk2[8].wave_shpr.div.quo[20] ;
 wire \genblk2[8].wave_shpr.div.quo[21] ;
 wire \genblk2[8].wave_shpr.div.quo[22] ;
 wire \genblk2[8].wave_shpr.div.quo[23] ;
 wire \genblk2[8].wave_shpr.div.quo[24] ;
 wire \genblk2[8].wave_shpr.div.quo[2] ;
 wire \genblk2[8].wave_shpr.div.quo[3] ;
 wire \genblk2[8].wave_shpr.div.quo[4] ;
 wire \genblk2[8].wave_shpr.div.quo[5] ;
 wire \genblk2[8].wave_shpr.div.quo[6] ;
 wire \genblk2[8].wave_shpr.div.quo[7] ;
 wire \genblk2[8].wave_shpr.div.quo[8] ;
 wire \genblk2[8].wave_shpr.div.quo[9] ;
 wire \genblk2[9].wave_shpr.div.acc[0] ;
 wire \genblk2[9].wave_shpr.div.acc[10] ;
 wire \genblk2[9].wave_shpr.div.acc[11] ;
 wire \genblk2[9].wave_shpr.div.acc[12] ;
 wire \genblk2[9].wave_shpr.div.acc[13] ;
 wire \genblk2[9].wave_shpr.div.acc[14] ;
 wire \genblk2[9].wave_shpr.div.acc[15] ;
 wire \genblk2[9].wave_shpr.div.acc[16] ;
 wire \genblk2[9].wave_shpr.div.acc[17] ;
 wire \genblk2[9].wave_shpr.div.acc[18] ;
 wire \genblk2[9].wave_shpr.div.acc[19] ;
 wire \genblk2[9].wave_shpr.div.acc[1] ;
 wire \genblk2[9].wave_shpr.div.acc[20] ;
 wire \genblk2[9].wave_shpr.div.acc[21] ;
 wire \genblk2[9].wave_shpr.div.acc[22] ;
 wire \genblk2[9].wave_shpr.div.acc[23] ;
 wire \genblk2[9].wave_shpr.div.acc[24] ;
 wire \genblk2[9].wave_shpr.div.acc[25] ;
 wire \genblk2[9].wave_shpr.div.acc[26] ;
 wire \genblk2[9].wave_shpr.div.acc[2] ;
 wire \genblk2[9].wave_shpr.div.acc[3] ;
 wire \genblk2[9].wave_shpr.div.acc[4] ;
 wire \genblk2[9].wave_shpr.div.acc[5] ;
 wire \genblk2[9].wave_shpr.div.acc[6] ;
 wire \genblk2[9].wave_shpr.div.acc[7] ;
 wire \genblk2[9].wave_shpr.div.acc[8] ;
 wire \genblk2[9].wave_shpr.div.acc[9] ;
 wire \genblk2[9].wave_shpr.div.acc_next[0] ;
 wire \genblk2[9].wave_shpr.div.b1[0] ;
 wire \genblk2[9].wave_shpr.div.b1[10] ;
 wire \genblk2[9].wave_shpr.div.b1[11] ;
 wire \genblk2[9].wave_shpr.div.b1[12] ;
 wire \genblk2[9].wave_shpr.div.b1[13] ;
 wire \genblk2[9].wave_shpr.div.b1[14] ;
 wire \genblk2[9].wave_shpr.div.b1[15] ;
 wire \genblk2[9].wave_shpr.div.b1[16] ;
 wire \genblk2[9].wave_shpr.div.b1[17] ;
 wire \genblk2[9].wave_shpr.div.b1[1] ;
 wire \genblk2[9].wave_shpr.div.b1[2] ;
 wire \genblk2[9].wave_shpr.div.b1[3] ;
 wire \genblk2[9].wave_shpr.div.b1[4] ;
 wire \genblk2[9].wave_shpr.div.b1[5] ;
 wire \genblk2[9].wave_shpr.div.b1[6] ;
 wire \genblk2[9].wave_shpr.div.b1[7] ;
 wire \genblk2[9].wave_shpr.div.b1[8] ;
 wire \genblk2[9].wave_shpr.div.b1[9] ;
 wire \genblk2[9].wave_shpr.div.busy ;
 wire \genblk2[9].wave_shpr.div.done ;
 wire \genblk2[9].wave_shpr.div.fin_quo[0] ;
 wire \genblk2[9].wave_shpr.div.fin_quo[1] ;
 wire \genblk2[9].wave_shpr.div.fin_quo[2] ;
 wire \genblk2[9].wave_shpr.div.fin_quo[3] ;
 wire \genblk2[9].wave_shpr.div.fin_quo[4] ;
 wire \genblk2[9].wave_shpr.div.fin_quo[5] ;
 wire \genblk2[9].wave_shpr.div.fin_quo[6] ;
 wire \genblk2[9].wave_shpr.div.fin_quo[7] ;
 wire \genblk2[9].wave_shpr.div.i[0] ;
 wire \genblk2[9].wave_shpr.div.i[1] ;
 wire \genblk2[9].wave_shpr.div.i[2] ;
 wire \genblk2[9].wave_shpr.div.i[3] ;
 wire \genblk2[9].wave_shpr.div.i[4] ;
 wire \genblk2[9].wave_shpr.div.quo[0] ;
 wire \genblk2[9].wave_shpr.div.quo[10] ;
 wire \genblk2[9].wave_shpr.div.quo[11] ;
 wire \genblk2[9].wave_shpr.div.quo[12] ;
 wire \genblk2[9].wave_shpr.div.quo[13] ;
 wire \genblk2[9].wave_shpr.div.quo[14] ;
 wire \genblk2[9].wave_shpr.div.quo[15] ;
 wire \genblk2[9].wave_shpr.div.quo[16] ;
 wire \genblk2[9].wave_shpr.div.quo[17] ;
 wire \genblk2[9].wave_shpr.div.quo[18] ;
 wire \genblk2[9].wave_shpr.div.quo[19] ;
 wire \genblk2[9].wave_shpr.div.quo[1] ;
 wire \genblk2[9].wave_shpr.div.quo[20] ;
 wire \genblk2[9].wave_shpr.div.quo[21] ;
 wire \genblk2[9].wave_shpr.div.quo[22] ;
 wire \genblk2[9].wave_shpr.div.quo[23] ;
 wire \genblk2[9].wave_shpr.div.quo[24] ;
 wire \genblk2[9].wave_shpr.div.quo[2] ;
 wire \genblk2[9].wave_shpr.div.quo[3] ;
 wire \genblk2[9].wave_shpr.div.quo[4] ;
 wire \genblk2[9].wave_shpr.div.quo[5] ;
 wire \genblk2[9].wave_shpr.div.quo[6] ;
 wire \genblk2[9].wave_shpr.div.quo[7] ;
 wire \genblk2[9].wave_shpr.div.quo[8] ;
 wire \genblk2[9].wave_shpr.div.quo[9] ;
 wire \modein.delay_in[0] ;
 wire \modein.delay_in[1] ;
 wire \modein.delay_octave_down_in[0] ;
 wire \modein.delay_octave_down_in[1] ;
 wire \modein.delay_octave_up_in[0] ;
 wire \modein.delay_octave_up_in[1] ;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire \sig_norm.acc[0] ;
 wire \sig_norm.acc[10] ;
 wire \sig_norm.acc[11] ;
 wire \sig_norm.acc[12] ;
 wire \sig_norm.acc[1] ;
 wire \sig_norm.acc[2] ;
 wire \sig_norm.acc[3] ;
 wire \sig_norm.acc[4] ;
 wire \sig_norm.acc[5] ;
 wire \sig_norm.acc[6] ;
 wire \sig_norm.acc[7] ;
 wire \sig_norm.acc[8] ;
 wire \sig_norm.acc[9] ;
 wire \sig_norm.acc_next[0] ;
 wire \sig_norm.b1[0] ;
 wire \sig_norm.b1[1] ;
 wire \sig_norm.b1[2] ;
 wire \sig_norm.b1[3] ;
 wire \sig_norm.busy ;
 wire \sig_norm.i[0] ;
 wire \sig_norm.i[1] ;
 wire \sig_norm.i[2] ;
 wire \sig_norm.i[3] ;
 wire \sig_norm.quo[0] ;
 wire \sig_norm.quo[10] ;
 wire \sig_norm.quo[1] ;
 wire \sig_norm.quo[2] ;
 wire \sig_norm.quo[3] ;
 wire \sig_norm.quo[4] ;
 wire \sig_norm.quo[5] ;
 wire \sig_norm.quo[6] ;
 wire \sig_norm.quo[7] ;
 wire \sig_norm.quo[8] ;
 wire \sig_norm.quo[9] ;
 wire \smpl_rt_clkdiv.clkDiv_inst.cnt[0] ;
 wire \smpl_rt_clkdiv.clkDiv_inst.cnt[1] ;
 wire \smpl_rt_clkdiv.clkDiv_inst.cnt[2] ;
 wire \smpl_rt_clkdiv.clkDiv_inst.cnt[3] ;
 wire \smpl_rt_clkdiv.clkDiv_inst.cnt[4] ;
 wire \smpl_rt_clkdiv.clkDiv_inst.cnt[5] ;
 wire \smpl_rt_clkdiv.clkDiv_inst.cnt[6] ;
 wire \smpl_rt_clkdiv.clkDiv_inst.cnt[7] ;
 wire \smpl_rt_clkdiv.clkDiv_inst.next_cnt[0] ;
 wire \smpl_rt_clkdiv.clkDiv_inst.next_cnt[1] ;
 wire \smpl_rt_clkdiv.clkDiv_inst.next_cnt[2] ;
 wire \smpl_rt_clkdiv.clkDiv_inst.next_cnt[3] ;
 wire \smpl_rt_clkdiv.clkDiv_inst.next_cnt[4] ;
 wire \smpl_rt_clkdiv.clkDiv_inst.next_cnt[5] ;
 wire \smpl_rt_clkdiv.clkDiv_inst.next_cnt[6] ;
 wire \smpl_rt_clkdiv.clkDiv_inst.next_cnt[7] ;
 wire \smpl_rt_clkdiv.clkDiv_inst.next_hzX ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06125__B (.DIODE(_01095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06125__C (.DIODE(_01096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06126__A (.DIODE(_01097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06128__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__06128__B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__06129__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__06129__B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__06131__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__06132__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__06132__B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__06133__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__06133__B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__06135__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__06136__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06136__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__06137__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06137__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__06141__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__06142__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__06143__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__06145__A (.DIODE(_01114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06146__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__06147__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06147__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__06153__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__06158__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__06159__A (.DIODE(_01114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06162__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__06183__A1 (.DIODE(_01099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06184__B (.DIODE(_01095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06184__C (.DIODE(_01096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06185__B (.DIODE(_01097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06186__A1 (.DIODE(_01155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06187__A (.DIODE(_01157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06210__A (.DIODE(_01171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06218__A1 (.DIODE(_01174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06218__B1 (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06219__A (.DIODE(_01174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06221__A (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06221__B (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06222__A1 (.DIODE(_01172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06222__A2 (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06222__B1 (.DIODE(_01183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06224__A (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06227__A1 (.DIODE(_01174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06227__B1_N (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06228__B (.DIODE(_01189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06231__A (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06231__B (.DIODE(_01192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06235__A (.DIODE(_01196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06236__A (.DIODE(_01174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06237__A1 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06237__A2 (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06238__A (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06239__A (.DIODE(_01200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06240__A1 (.DIODE(_01201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06241__A1 (.DIODE(_01201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06243__A1 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06243__A2 (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06244__A2 (.DIODE(_01190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06247__A (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06248__A (.DIODE(_01209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06249__A (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06250__A2 (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06250__B1 (.DIODE(_01210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06250__B2 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06251__A (.DIODE(_01174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06252__B (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06253__A (.DIODE(_01213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06253__B (.DIODE(_01214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06254__A1_N (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06254__A2_N (.DIODE(_01215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06255__A2 (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06255__B1 (.DIODE(_01215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06255__B2 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06256__A1 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06256__A2 (.DIODE(_01210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06262__A2 (.DIODE(_01221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06262__B1 (.DIODE(_01223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06265__A (.DIODE(_01224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06265__B (.DIODE(_01226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06269__A (.DIODE(_01229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06272__A1 (.DIODE(_01229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06273__A (.DIODE(_01231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06273__B (.DIODE(_01234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06274__A2 (.DIODE(_01227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06274__B1 (.DIODE(_01235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06277__B (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06278__A (.DIODE(_01238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06280__A (.DIODE(_01241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06281__B (.DIODE(_01242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06282__B (.DIODE(_01242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06287__B (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06288__A (.DIODE(_01248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06288__B (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06289__A (.DIODE(_01246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06289__B (.DIODE(_01250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06291__A2 (.DIODE(_01240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06293__A (.DIODE(_01196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06294__A (.DIODE(_01255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06295__A1 (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06296__A (.DIODE(_01238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06297__A2_N (.DIODE(_01190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06298__A1 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06298__A2 (.DIODE(_01256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06298__B1 (.DIODE(_01240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06301__A (.DIODE(_01238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06301__B (.DIODE(_01262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06302__B (.DIODE(_01263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06303__A1 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06303__A2 (.DIODE(_01256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06304__A2 (.DIODE(_01235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06305__A2 (.DIODE(_01227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06320__A1 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06322__B (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06323__A1 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06346__B1 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06347__A (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06349__A (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06351__A1 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06352__B (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06355__A (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06356__A1 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06359__A (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06359__C (.DIODE(_01302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06361__A (.DIODE(_01223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06361__B (.DIODE(_01226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06365__A (.DIODE(_01171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06366__A (.DIODE(_01308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06366__B (.DIODE(_01309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06368__A (.DIODE(_01309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06368__B (.DIODE(_01221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06369__A (.DIODE(_01192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06369__B (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06370__B (.DIODE(_01313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06371__A2 (.DIODE(_01311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06371__B2 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06373__B (.DIODE(_01240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06374__A2 (.DIODE(_01311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06374__B2 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06377__A_N (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06378__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__06382__A (.DIODE(_01229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06384__B (.DIODE(_01327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06385__A (.DIODE(_01326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06385__B (.DIODE(_01328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06387__A2 (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06387__B1 (.DIODE(_01329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06389__A (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06391__A (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06391__B (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06392__A (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06393__A (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06393__B (.DIODE(_01226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06394__A2 (.DIODE(_01210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06394__B1 (.DIODE(_01337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06394__B2 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06395__A2 (.DIODE(_01210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06395__B1 (.DIODE(_01337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06395__B2 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06396__A (.DIODE(_01238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06396__B (.DIODE(_01262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06398__A (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06401__A1 (.DIODE(_01342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06401__A2 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06401__B1 (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06401__B2 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06402__A2 (.DIODE(_01340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06402__B1 (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06403__A (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06403__B (.DIODE(_01327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06404__A (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06404__B (.DIODE(_01327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06405__A (.DIODE(_01172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06406__A1 (.DIODE(_01201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06406__A2 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06406__B1 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06407__A2_N (.DIODE(_01349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06407__B2 (.DIODE(_01342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06408__A2 (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06412__A (.DIODE(_01226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06412__B (.DIODE(_01355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06413__A (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06413__B (.DIODE(_01356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06416__A (.DIODE(_01359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06417__A (.DIODE(_01360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06418__A (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06419__A (.DIODE(_01362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06420__A2 (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06421__A (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06422__B (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06424__A (.DIODE(_01365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06424__B (.DIODE(_01367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06425__A1_N (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06425__A2_N (.DIODE(_01368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06425__B1 (.DIODE(_01340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06426__A1 (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06426__B1 (.DIODE(_01368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06426__B2 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06428__A2 (.DIODE(_01304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06452__A (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06453__A (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06456__A (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06456__B (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06457__A1 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06457__B1 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06459__A (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06460__A (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06462__A (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06463__A1 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06464__A1 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06464__B1 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06465__A (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06465__B (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06467__A (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06469__A1 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06470__A (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06470__B (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06472__A1 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06473__A (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06475__A1 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06476__B (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06485__A (.DIODE(_01241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06485__B (.DIODE(_01337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06487__A2_N (.DIODE(_01411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06487__B2 (.DIODE(_01183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06489__S (.DIODE(_01210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06491__A2 (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06492__A (.DIODE(_01229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06492__B (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06493__A1 (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06493__B1 (.DIODE(_01418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06494__A (.DIODE(_01242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06494__B (.DIODE(_01223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06495__C (.DIODE(_01327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06496__C (.DIODE(_01327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06498__B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__06499__C (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__06500__C (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__06503__A2 (.DIODE(_01411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06504__A (.DIODE(_01224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06505__A1 (.DIODE(_01362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06505__A2 (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06505__B1 (.DIODE(_01196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06507__A (.DIODE(_01200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06507__B (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06508__A1 (.DIODE(_01201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06508__B1 (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06509__A2 (.DIODE(_01365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06509__B1 (.DIODE(_01326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06510__A (.DIODE(_01349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06512__B (.DIODE(_01437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06513__A (.DIODE(_01213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06515__A (.DIODE(_01440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06516__A (.DIODE(_01200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06516__B (.DIODE(_01441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06517__A2_N (.DIODE(_01439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06517__B1 (.DIODE(_01442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06518__A2_N (.DIODE(_01442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06518__B1 (.DIODE(_01439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06519__B1 (.DIODE(_01418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06521__B2 (.DIODE(_01436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06524__A2 (.DIODE(_01231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06575__A (.DIODE(_01196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06575__B (.DIODE(_01327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06576__A (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06576__B (.DIODE(_01302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06579__A (.DIODE(_01172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06579__B (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06580__A2 (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06582__A (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06583__B (.DIODE(_01250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06584__A2 (.DIODE(_01231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06584__B2 (.DIODE(_01490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06585__A1_N (.DIODE(_01490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06585__B1 (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06586__A (.DIODE(_01342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06586__B (.DIODE(_01248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06587__B (.DIODE(_01494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06588__A (.DIODE(_01437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06591__B1 (.DIODE(_01498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06592__B (.DIODE(_01437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06593__A2_N (.DIODE(_01498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06593__B1 (.DIODE(_01500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06594__A2_N (.DIODE(_01500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06595__A2 (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06597__B (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06598__B (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06599__A (.DIODE(_01441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06599__B (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06600__A (.DIODE(_01241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06600__B (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06601__A2_N (.DIODE(_01507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06601__B1 (.DIODE(_01508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06602__A2 (.DIODE(_01484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06603__A2 (.DIODE(_01487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06604__A (.DIODE(_01171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06604__B (.DIODE(_01192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06604__C (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06606__A (.DIODE(_01234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06607__A2_N (.DIODE(_01513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06607__B1 (.DIODE(_01514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06608__B (.DIODE(_01210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06609__A2_N (.DIODE(_01514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06609__B1 (.DIODE(_01513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06610__A2 (.DIODE(_01231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06611__B1 (.DIODE(_01171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06612__B (.DIODE(_01519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06613__A2 (.DIODE(_01256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06614__A2 (.DIODE(_01483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06614__B1 (.DIODE(_01484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06666__A2 (.DIODE(_01221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06666__B1 (.DIODE(_01223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06667__A (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06667__B (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06669__A (.DIODE(_01349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06669__B (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06672__A2_N (.DIODE(_01326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06672__B1 (.DIODE(_01498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06675__B (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06676__B (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06677__B (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06679__A2 (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06679__B1 (.DIODE(_01242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06681__A2 (.DIODE(_01362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06681__B1 (.DIODE(_01248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06682__A2 (.DIODE(_01439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06682__B1 (.DIODE(_01340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06684__S (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06687__A (.DIODE(_01576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06688__A (.DIODE(_01577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06689__A2_N (.DIODE(_01574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06689__B1 (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06690__A2_N (.DIODE(_01209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06690__B1 (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06691__A2 (.DIODE(_01210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06691__B1 (.DIODE(_01498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06693__A2_N (.DIODE(_01313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06693__B1 (.DIODE(_01340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06694__A2 (.DIODE(_01313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06695__B (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06696__A2 (.DIODE(_01326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06696__B1 (.DIODE(_01574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06697__A2 (.DIODE(_01436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06697__B1 (.DIODE(_01304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06700__B (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06702__A (.DIODE(_01171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06702__B (.DIODE(_01591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06703__B (.DIODE(_01592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06704__B (.DIODE(_01592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06705__A (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06705__B (.DIODE(_01196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06706__B (.DIODE(_01595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06707__A2 (.DIODE(_01304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06784__A1 (.DIODE(_01436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06784__A2 (.DIODE(_01304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06785__B (.DIODE(_01483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06786__A (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06786__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__06787__B (.DIODE(_01658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06788__A (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06788__B (.DIODE(_01262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06790__B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__06791__B (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06793__B (.DIODE(_01592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06794__A (.DIODE(_01440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06794__B (.DIODE(_01171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06796__A2_N (.DIODE(_01666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06799__A2 (.DIODE(_01210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06799__B1 (.DIODE(_01304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06800__B1 (.DIODE(_01666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06801__B2 (.DIODE(_01436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06802__A (.DIODE(_01238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06802__B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__06804__A2 (.DIODE(_01362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06805__B (.DIODE(_01362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06805__C (.DIODE(_01226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06806__A (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06806__B (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06807__B (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06808__B (.DIODE(_01359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06810__B (.DIODE(_01326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06811__B (.DIODE(_01326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06812__A (.DIODE(_01189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06812__B (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06813__A (.DIODE(\genblk1[5].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06813__B (.DIODE(_01684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06814__A2 (.DIODE(_01242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06815__B (.DIODE(_01355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06816__B (.DIODE(_01355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06818__B1 (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06824__B (.DIODE(\genblk1[5].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06825__B (.DIODE(\genblk1[5].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06828__C (.DIODE(\genblk1[5].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06829__A2 (.DIODE(\genblk1[5].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06872__A (.DIODE(_01441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06873__A2 (.DIODE(_01726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06874__B (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06876__A (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06876__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__06877__B (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06879__B1 (.DIODE(_01732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06880__A2 (.DIODE(_01684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06881__A (.DIODE(_01189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06881__B (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06882__A2_N (.DIODE(_01732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06882__B1 (.DIODE(_01735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06883__A2 (.DIODE(_01484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06884__A (.DIODE(_01241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06885__A (.DIODE(_01349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06885__B (.DIODE(_01209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06885__C (.DIODE(_01439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06886__A2 (.DIODE(_01738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06886__B1 (.DIODE(_01739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06887__A2 (.DIODE(_01738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06888__A (.DIODE(_01658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06888__B (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06889__A2_N (.DIODE(_01519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06890__A2 (.DIODE(_01519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06890__B1 (.DIODE(_01739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06891__A2_N (.DIODE(_01666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06891__B1 (.DIODE(_01484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06892__A2 (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06892__B1 (.DIODE(_01666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06893__A (.DIODE(_01308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06893__B (.DIODE(_01577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06895__B (.DIODE(_01362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06896__A (.DIODE(_01342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06896__B (.DIODE(_01439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06897__A2 (.DIODE(_01367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06898__A2 (.DIODE(_01367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06900__B1 (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06903__B (.DIODE(_01327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06904__A (.DIODE(_01576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06904__B (.DIODE(_01757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06906__A1 (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06956__A2 (.DIODE(_01311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06956__B1 (.DIODE(_01732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__A2 (.DIODE(_01227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__B1 (.DIODE(_01732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06959__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__C (.DIODE(_01514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__A (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__B (.DIODE(_01221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06962__B (.DIODE(_01797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__A1 (.DIODE(_01229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__B1 (.DIODE(_01238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06964__B (.DIODE(_01799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__A (.DIODE(_01213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__B (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06966__A (.DIODE(_01192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06967__A2 (.DIODE(_01574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06968__A2 (.DIODE(_01801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06969__A (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06970__A2_N (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06970__B1 (.DIODE(_01801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06971__B1 (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06972__B (.DIODE(_01214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06973__A2 (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06973__B1 (.DIODE(_01311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06974__B (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06975__A (.DIODE(_01365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06975__B (.DIODE(_01355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06976__B (.DIODE(_01811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06979__A2 (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06979__B1 (.DIODE(_01196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06980__A2 (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06980__B1 (.DIODE(_01574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06983__A (.DIODE(_01436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06983__B (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06984__B (.DIODE(_01819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__A2 (.DIODE(_01227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07034__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07034__B (.DIODE(_01359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07035__B1 (.DIODE(_01248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__B1 (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07037__B (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07038__A1 (.DIODE(_01436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07038__A2 (.DIODE(_01855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07039__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07039__B (.DIODE(_01487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07040__A (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07040__B (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07041__A (.DIODE(_01439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07041__B (.DIODE(_01576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07042__A2 (.DIODE(_01436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07042__A3 (.DIODE(_01855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__A2 (.DIODE(_01487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__B1 (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__B2 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__B (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07046__B (.DIODE(_01328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07047__A (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07047__B (.DIODE(_01223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07048__A1 (.DIODE(_01174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07048__A2 (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07048__B1 (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07049__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07051__A (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07051__B (.DIODE(_01183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__A (.DIODE(_01441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__B (.DIODE(_01226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__A1_N (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__A2_N (.DIODE(_01869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__B1 (.DIODE(_01870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__B2 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07054__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07054__A2 (.DIODE(_01436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07055__B (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07056__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07056__B (.DIODE(_01498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07057__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07057__A2 (.DIODE(_01246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07058__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07058__A2 (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07058__B1 (.DIODE(_01246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07058__B2 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07059__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07059__B1 (.DIODE(_01869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07059__B2 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07062__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07062__A2 (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07062__C1 (.DIODE(_01490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07062__D1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07063__A1 (.DIODE(_01441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07065__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07065__A2 (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07066__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07066__A2 (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07066__B1 (.DIODE(_01870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07066__B2 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07071__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07072__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07077__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07078__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07080__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07082__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07082__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07083__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07083__B1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07085__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07086__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07088__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07090__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07099__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07101__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07102__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07102__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07104__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07105__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07111__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07111__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07113__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07114__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07115__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07119__B (.DIODE(_01227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__A (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__B (.DIODE(_01221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07121__A1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07121__B1 (.DIODE(_01855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07121__B2 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__A2 (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__B1 (.DIODE(_01328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__B2 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07123__A (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07123__B (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__A (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__B (.DIODE(_01355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07126__A1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07126__A2 (.DIODE(_01925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07126__B1 (.DIODE(_01855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07126__B2 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07127__A1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07127__B1 (.DIODE(_01923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07129__B (.DIODE(_01801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07131__B (.DIODE(_01250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07132__A1_N (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07132__A2_N (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07132__B1 (.DIODE(_01349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07132__B2 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07133__A2 (.DIODE(_01513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07134__A1_N (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07134__A2_N (.DIODE(_01311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07134__B1 (.DIODE(_01923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__A1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__A2 (.DIODE(_01311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__B1 (.DIODE(_01925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__B2 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07136__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07136__B (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07137__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07138__A1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07138__A2 (.DIODE(_01246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07138__B1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07139__A1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07139__A2 (.DIODE(_01246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07139__B1 (.DIODE(_01196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__A2 (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__B1 (.DIODE(_01328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__B2 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07142__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07142__B (.DIODE(_01514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07143__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07143__B (.DIODE(_01514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07145__A2 (.DIODE(_01514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07145__B1 (.DIODE(_01513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__A (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__A (.DIODE(_01241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__B (.DIODE(_01946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07148__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__A2_N (.DIODE(_01799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__B2 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__A2 (.DIODE(_01799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07151__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07156__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07156__B (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__B (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07160__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07160__B (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07160__C (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__A1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__A2 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__B1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07164__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07166__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07167__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07170__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07170__B (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__A1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__B1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07194__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__A1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07197__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07199__A1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07200__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07200__B (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07202__A1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07209__A (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07209__B (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07210__A1 (.DIODE(_01359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07210__A2 (.DIODE(_01224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07210__B1 (.DIODE(_01241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07212__A1 (.DIODE(_01308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07212__B1 (.DIODE(_01214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07214__A (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07215__A1 (.DIODE(_01490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07216__B (.DIODE(_01442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07217__A2 (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07217__B2 (.DIODE(_01342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__A2 (.DIODE(_01246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__B1 (.DIODE(_01442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__A (.DIODE(_01365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__B (.DIODE(_01189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__A2_N (.DIODE(_02001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__B1 (.DIODE(_02002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07223__A1 (.DIODE(_01174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07223__B1 (.DIODE(_01196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__A2_N (.DIODE(_01235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__B1 (.DIODE(_01227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07229__A (.DIODE(_01229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07230__B (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07232__B1 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07233__A2 (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__B (.DIODE(_01359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07236__A2_N (.DIODE(_02001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07236__B1 (.DIODE(_02002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07237__A1 (.DIODE(_01242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07237__B2 (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07238__A2 (.DIODE(_02011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07239__B (.DIODE(_01215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07240__A2 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07242__B1 (.DIODE(_01183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__A2 (.DIODE(_01235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__A2 (.DIODE(_01991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07299__B (.DIODE(_01235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07300__A (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07300__B (.DIODE(_01226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__B (.DIODE(_01595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__A2 (.DIODE(_01256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__B1 (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__A2_N (.DIODE(_01256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__B1 (.DIODE(_01595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__A2_N (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__B1 (.DIODE(_01925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__A1 (.DIODE(_01223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__A2 (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07307__B (.DIODE(_01223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07307__C (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07308__A2 (.DIODE(_01513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07309__B (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07310__B (.DIODE(_02002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__A2_N (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__B1 (.DIODE(_01262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__A2 (.DIODE(_01210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__B1 (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__A (.DIODE(_01308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__B (.DIODE(_01439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__A2 (.DIODE(_02077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__B1 (.DIODE(\genblk1[11].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07315__A2 (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07315__B1 (.DIODE(_02077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07318__B (.DIODE(_01262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__A2 (.DIODE(_01242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__A2 (.DIODE(_01513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07321__B (.DIODE(_01359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__A2_N (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07324__A2 (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07324__B2 (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07325__B1 (.DIODE(_01925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__A (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__A (.DIODE(_02147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07408__A (.DIODE(_02152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07409__B (.DIODE(_02153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__A (.DIODE(_02154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07415__A (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07417__B (.DIODE(_02153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__A (.DIODE(_02160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07422__A (.DIODE(_02147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07424__B (.DIODE(_02153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__A (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__A (.DIODE(_02152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07432__A (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07434__A (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07439__A (.DIODE(_02147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07441__B (.DIODE(_02153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__A (.DIODE(_02147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07448__A (.DIODE(_02183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07449__B (.DIODE(_02153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07450__A (.DIODE(_02184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07454__A (.DIODE(_02147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__B (.DIODE(_02153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__A (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__A (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07463__B (.DIODE(_02153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07468__A (.DIODE(_02147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07470__B (.DIODE(_02153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07475__A (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07476__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07477__B (.DIODE(_02153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07478__A (.DIODE(_02204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07482__A (.DIODE(_02147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07484__B (.DIODE(_02153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07485__A (.DIODE(_02209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07489__A (.DIODE(_02147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__B (.DIODE(_02152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07492__A (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__A (.DIODE(\modein.delay_in[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07494__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__A (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07499__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__07499__B_N (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__07501__A_N (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__07501__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__07502__A (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__A (.DIODE(_02223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07504__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__07504__B_N (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__07505__B1 (.DIODE(_02225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__A2 (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__A3 (.DIODE(_02224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__B1 (.DIODE(_01099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07529__A (.DIODE(_01099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07531__A (.DIODE(_01155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__A (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__B1 (.DIODE(_01099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07553__A (.DIODE(_01157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__A (.DIODE(_02223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__A1 (.DIODE(_01200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__A2 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__B1 (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__C1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07560__A1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07560__B1 (.DIODE(_01328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07562__A2_N (.DIODE(_01799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07563__A2 (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07563__A3 (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07563__B1 (.DIODE(_01801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07564__A2 (.DIODE(_01227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07564__B1 (.DIODE(_01732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07565__A2 (.DIODE(_01328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07565__B1 (.DIODE(_01799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07567__A1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07567__B1 (.DIODE(_01349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__A1_N (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__A2_N (.DIODE(_01349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__B1 (.DIODE(_01246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__B2 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07569__A1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07569__A2 (.DIODE(_01577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07571__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07571__C (.DIODE(_01355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07572__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07572__C (.DIODE(_01437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07574__A1 (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07574__A2 (.DIODE(_01437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07574__A3 (.DIODE(_01226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07574__B1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__A1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__A2 (.DIODE(_01925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07576__B1 (.DIODE(_01234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__B (.DIODE(_01234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07580__A1 (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07580__A2 (.DIODE(_01221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07580__B1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__A2 (.DIODE(_01437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__A3 (.DIODE(_01226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__B1 (.DIODE(_01171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__C1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__C (.DIODE(_01221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07583__A1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07583__A2 (.DIODE(_01234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07584__A1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07584__A2 (.DIODE(_01234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07584__B2 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07585__A1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07585__A2 (.DIODE(_01311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07587__A2 (.DIODE(_01234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07587__B1 (.DIODE(_01513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07590__A2 (.DIODE(_01991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07590__B1 (.DIODE(_01923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__B (.DIODE(_01801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07595__B1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07595__C1 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07596__A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__07599__A (.DIODE(_02261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__07602__A (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__A (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__A2 (.DIODE(_02309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__07606__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__07606__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__07609__A (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07610__B (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__A2 (.DIODE(_01437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__A1 (.DIODE(_01171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__A2 (.DIODE(_01192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__A3 (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07615__C (.DIODE(_01437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__A2 (.DIODE(_01513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__B1 (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07618__B (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07619__A2 (.DIODE(_01595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07620__A2 (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07620__B1 (.DIODE(_01595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__A2 (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07622__B (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07624__B1 (.DIODE(_01172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__A2 (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__B1 (.DIODE(_01576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07626__A2 (.DIODE(_01241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__A2 (.DIODE(_01209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__B1 (.DIODE(_01256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07628__A2 (.DIODE(_01256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__A (.DIODE(_01174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07630__B (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07630__C (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__B (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__C (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07632__A2 (.DIODE(_01262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07633__A2_N (.DIODE(_01262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07633__B1 (.DIODE(_01494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07634__A2 (.DIODE(_01190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__A2 (.DIODE(_01190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__B1 (.DIODE(_01235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07638__A1 (.DIODE(_01229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07642__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07643__B (.DIODE(\genblk1[11].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07644__A (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07652__A (.DIODE(_02316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07653__B1 (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07655__A (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07656__B (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07657__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07659__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__07659__B (.DIODE(_02364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07659__C (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07661__A2 (.DIODE(_01190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07661__B1 (.DIODE(_01235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07662__B (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__A1 (.DIODE(_01360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__A2 (.DIODE(_01224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__B1 (.DIODE(_01241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07664__A2 (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07664__A3 (.DIODE(_01794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07664__B2 (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07666__B2 (.DIODE(_01190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07667__A (.DIODE(_01308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07668__A2 (.DIODE(_02374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07668__B1 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07669__A (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07669__B (.DIODE(_01440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07671__A (.DIODE(_01308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07672__A (.DIODE(_01308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__A2 (.DIODE(_02001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__B1 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07676__A2 (.DIODE(_01190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__A2_N (.DIODE(_01215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__B1 (.DIODE(_01991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07679__A (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07680__A (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__A2 (.DIODE(_01246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__A (.DIODE(_01174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__A0 (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07687__A2 (.DIODE(_02011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__A2 (.DIODE(_01215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__B1 (.DIODE(_02011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07690__A2 (.DIODE(_01991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07692__B (.DIODE(_02011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07697__A (.DIODE(_02403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07707__A (.DIODE(_02316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__A (.DIODE(_02225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__B (.DIODE(_02403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07710__A2 (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07711__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__07711__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__07717__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__07717__B (.DIODE(_02364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07717__C (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07718__A (.DIODE(_01360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07718__B (.DIODE(_01302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07719__A2 (.DIODE(_01309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07719__B1 (.DIODE(_01209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07719__B2 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__A2 (.DIODE(_01309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__B1 (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__B2 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07721__A1 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07721__A2 (.DIODE(_02425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07722__A2 (.DIODE(_01262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07722__B1 (.DIODE(_01591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07722__C1 (.DIODE(_01172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__A2 (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__A2 (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__B1 (.DIODE(_01313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__B1 (.DIODE(_01313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07726__A (.DIODE(_01342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07726__B (.DIODE(_01241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07727__A2 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__A (.DIODE(_01342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__B (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__A1 (.DIODE(_01360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07730__A (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07730__B (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__A2 (.DIODE(_01360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__A3 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07732__A2 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07735__A2 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__A (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07738__B (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07739__A1 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07739__A2 (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07739__B2 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07740__A1 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07740__A2 (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07740__B1 (.DIODE(_01356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07740__B2 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07741__A1 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07741__A2 (.DIODE(_01337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07741__B2 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07744__A1 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07744__A2 (.DIODE(_02425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07744__B1 (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07744__B2 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07745__A1 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07745__A2 (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07745__B1 (.DIODE(_01337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07745__B2 (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__B (.DIODE(_01172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07748__B (.DIODE(_01576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07752__A2 (.DIODE(_01577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07753__A (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07753__B (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__B1 (.DIODE(_02224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__A (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__A (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__A1 (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__A2 (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__A2 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__A1 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__A2 (.DIODE(_01309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__B1 (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__B2 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07766__B (.DIODE(_01255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07767__A1 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07767__A2 (.DIODE(_01309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07767__B1 (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07767__B2 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__A2 (.DIODE(_01256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__B1 (.DIODE(_01240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07770__A2 (.DIODE(_01240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07772__A2 (.DIODE(_01190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07772__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07772__D1 (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__A2 (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__A3 (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__B1 (.DIODE(_01190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07774__B (.DIODE(_01215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07775__A2 (.DIODE(_01227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07776__A (.DIODE(_01229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07776__B (.DIODE(_01359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07777__A (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07778__A1 (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__A1 (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07780__B1 (.DIODE(_01215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07782__A1 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07782__A2 (.DIODE(_01241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07783__A1 (.DIODE(_01200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07789__B (.DIODE(_01263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07790__B (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07790__C (.DIODE(_01801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__B (.DIODE(_01263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07792__A1 (.DIODE(_01246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07792__A2 (.DIODE(_01439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07792__A3 (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07798__A (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07798__B (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07798__C (.DIODE(_01209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__A1 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__A2 (.DIODE(_01349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__B1 (.DIODE(_01577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__A2 (.DIODE(_01577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__C1 (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07802__A (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07802__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07803__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07808__B1 (.DIODE(_02224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07809__B2 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07810__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07810__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07814__A (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07817__A_N (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__07817__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__A (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07820__A (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__A2 (.DIODE(_02521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__B2 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07822__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__07822__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07825__B1 (.DIODE(_02223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07827__A2 (.DIODE(_02309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__B1 (.DIODE(_02224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__A (.DIODE(_02309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__A2 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07836__B1 (.DIODE(_02261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07838__A2 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__B1 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07845__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__07850__B1 (.DIODE(_02316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07852__A2 (.DIODE(_02309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__B1 (.DIODE(_02316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__A (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07860__C (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07860__D (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07861__A2 (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07861__A3 (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07862__A1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07862__B1 (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07865__A (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07866__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__A1 (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07885__A (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07886__A2 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07886__B2 (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__A2 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__B2 (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__C (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__A1_N (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__A2_N (.DIODE(_01309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__B1 (.DIODE(_01576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__B2 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__A1_N (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07900__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07900__A2 (.DIODE(_01172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__A2 (.DIODE(_01246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__B1 (.DIODE(_01328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__B2 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__A2 (.DIODE(_01328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__B (.DIODE(_01360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__C (.DIODE(_02011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__B (.DIODE(_01869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07905__B (.DIODE(_01870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07908__B (.DIODE(_01870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07909__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07909__A2 (.DIODE(_01869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__A2 (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__C1 (.DIODE(_01238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__A2 (.DIODE(_01308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__A3 (.DIODE(_01440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__A2 (.DIODE(_01309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__A3 (.DIODE(_01855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__B2 (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07915__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07915__B1 (.DIODE(_01487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07915__B2 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__B (.DIODE(_01487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__A2 (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__A (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__A2 (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__B1 (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__B2 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A2 (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__B1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__C1 (.DIODE(_01441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__B (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07927__A1 (.DIODE(_01200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07927__A2 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07927__B1 (.DIODE(_01362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07927__C1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__C1 (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07929__A (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07929__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__A (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__B (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__C (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07933__A (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07935__B1 (.DIODE(_02223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07938__A2 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07940__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__07940__B (.DIODE(_02364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07942__A2 (.DIODE(_01311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07942__B1 (.DIODE(_01925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07943__A2 (.DIODE(_01925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__B1 (.DIODE(_01514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07945__B1 (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__A2 (.DIODE(_01574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07947__B (.DIODE(_01574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__A (.DIODE(_01172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__B (.DIODE(_02011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__A1 (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__A2 (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07951__A2 (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07951__A3 (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07951__B1 (.DIODE(_01732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07952__A2 (.DIODE(_01801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__A2 (.DIODE(_01732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__B1 (.DIODE(_02656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07954__B (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07956__A2 (.DIODE(_02656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07959__A2 (.DIODE(_01311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07959__B1 (.DIODE(_01925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__A2 (.DIODE(_01514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07961__B (.DIODE(_01360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07962__B (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07963__A1 (.DIODE(_01200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07963__A3 (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07965__A2 (.DIODE(_01577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07965__B1 (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__A2 (.DIODE(_01214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__B1 (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07967__A2 (.DIODE(_01214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07970__A2 (.DIODE(_01577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__A1 (.DIODE(_01201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__A3 (.DIODE(_01362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__A (.DIODE(\genblk2[7].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__B1 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07987__A (.DIODE(_02225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07993__A2 (.DIODE(_01484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07993__B1 (.DIODE(_01519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__A2 (.DIODE(_01732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07995__A2 (.DIODE(_01484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07997__B (.DIODE(_01360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07998__B (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__A1 (.DIODE(_01200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__A3 (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08001__A2 (.DIODE(_01577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08001__B1 (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__A2 (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__B1 (.DIODE(_01666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08003__A2 (.DIODE(_01666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__A2 (.DIODE(_01519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08006__A2 (.DIODE(_01735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08006__B1 (.DIODE(_01738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08007__B1 (.DIODE(_01735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08010__A2 (.DIODE(_01365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08011__A2 (.DIODE(_01367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08013__A2 (.DIODE(_01367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__B (.DIODE(_01367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__B1 (.DIODE(_01739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08018__A (.DIODE(_01739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08019__A2_N (.DIODE(_01732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08021__A2 (.DIODE(_01577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08023__A1 (.DIODE(_01229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08027__A (.DIODE(_02733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08028__A (.DIODE(\genblk2[6].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08028__B (.DIODE(\genblk2[6].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08032__B1 (.DIODE(_02261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08035__A (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08035__B (.DIODE(_02733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__A1 (.DIODE(\genblk2[6].wave_shpr.div.fin_quo[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__A2 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08037__A (.DIODE(_02364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08038__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__08038__C (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__B (.DIODE(_01576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08042__B (.DIODE(_01359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08043__B (.DIODE(_01360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08044__A1 (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08045__A2 (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__B1 (.DIODE(_01666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__A2 (.DIODE(_01666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08049__B (.DIODE(_01355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08050__B (.DIODE(_01355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__A1 (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__A3 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__08054__B (.DIODE(_01223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08055__A1 (.DIODE(_01309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08055__A2 (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08057__B (.DIODE(_01223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08058__A2 (.DIODE(_01172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08058__A3 (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__A2 (.DIODE(_01238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__B (.DIODE(_01238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__B (.DIODE(_01238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__C (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__08066__A1 (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08066__B1 (.DIODE(_01171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08066__C1 (.DIODE(\genblk1[5].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08068__A1 (.DIODE(_01196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08069__A2 (.DIODE(_01592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__A2 (.DIODE(_01309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__A3 (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__A2 (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__B1 (.DIODE(_01726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__A2 (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08079__A2 (.DIODE(_01355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08080__A1 (.DIODE(_01200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__A (.DIODE(_02225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__B (.DIODE(_02789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08087__B (.DIODE(_02789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08089__A2 (.DIODE(_02309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08089__B2 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__B (.DIODE(_02364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__C (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08093__B (.DIODE(_01360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__A2 (.DIODE(_01359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__B1 (.DIODE(_01498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08095__B (.DIODE(_01196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__A (.DIODE(_01174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__C (.DIODE(_01359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__A (.DIODE(_01440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__B (.DIODE(_01576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__A2 (.DIODE(_01498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__B1 (.DIODE(_02805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08100__A2 (.DIODE(_02805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08102__B (.DIODE(_01574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__B (.DIODE(_01574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__A2 (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__B1 (.DIODE(_01592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08105__B (.DIODE(_01192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08105__C (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08106__B (.DIODE(_01574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__A1 (.DIODE(_01192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__A2 (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08109__A2 (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08110__A2 (.DIODE(_01313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__A2 (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__A2 (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__B1 (.DIODE(_01592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08115__A1 (.DIODE(_01172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08115__A2 (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__B (.DIODE(_01326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08118__A2 (.DIODE(_01326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08118__B1 (.DIODE(_01213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08120__A1 (.DIODE(_01224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08120__A2 (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08121__A2 (.DIODE(_01439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__A2 (.DIODE(_01340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__B1 (.DIODE(_01304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__A2 (.DIODE(_01224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__A3 (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__B1 (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__A2 (.DIODE(_01340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__B1 (.DIODE(_01304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08125__A2 (.DIODE(_01870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__A2 (.DIODE(_01340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08131__A (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08131__B (.DIODE(_02837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__C_N (.DIODE(_02837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__A2 (.DIODE(_02309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__B2 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__B (.DIODE(_02364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__C (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__B (.DIODE(_01576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08145__A1 (.DIODE(_01201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08145__C1 (.DIODE(_01362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08147__B1 (.DIODE(_01519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08148__B1 (.DIODE(_01513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08149__B (.DIODE(_01513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08150__A2 (.DIODE(_01234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08151__A2 (.DIODE(_01250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08151__B1 (.DIODE(_01514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08152__A2 (.DIODE(_01500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08152__B1 (.DIODE(_01250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08153__A2 (.DIODE(_01500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08153__B1 (.DIODE(_01494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08155__A2 (.DIODE(_01483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08155__B1 (.DIODE(_01494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08156__A2_N (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08156__B1 (.DIODE(_01576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08157__A2 (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08158__A2 (.DIODE(_01483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08158__B1 (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08159__A (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08160__A (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08161__B (.DIODE(_01498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08163__A2 (.DIODE(_01498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08164__A (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08164__C (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08165__B (.DIODE(_01508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08167__B (.DIODE(_01231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__A2 (.DIODE(_01508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__B1 (.DIODE(_01507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__A2 (.DIODE(_01498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__B (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08181__B (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__B1 (.DIODE(_02224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08184__A (.DIODE(_02225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08184__B (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08185__B (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08186__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__08186__C (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__08196__A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__08196__A3 (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08196__B1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08197__B (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08200__A2 (.DIODE(_02403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08201__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__08205__B1 (.DIODE(_02316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08206__B2 (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__B (.DIODE(_02789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08222__A1 (.DIODE(_02789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__A2 (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__A1 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__A (.DIODE(_02837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08227__B1 (.DIODE(_02316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__B2 (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08232__A (.DIODE(_02225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08232__B (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__B (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08234__A1 (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08235__A1 (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08235__B1 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__C (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__B1 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08242__B (.DIODE(_02309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08243__A (.DIODE(_02225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08247__B1 (.DIODE(_02223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__A2 (.DIODE(_02309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08254__A2 (.DIODE(_02733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08254__B1 (.DIODE(_02261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08255__B2 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__A3 (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__B1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08268__B (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__B1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08275__A2 (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08279__B1 (.DIODE(_02223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08281__A2 (.DIODE(_02521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08308__B1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08309__B (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08313__B1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08314__A (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08319__B1 (.DIODE(_02316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__B2 (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08325__B1 (.DIODE(_02223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08327__A2 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08331__B1 (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08337__B1 (.DIODE(_02261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__A2 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__A_N (.DIODE(_02789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08350__B1 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08352__A2 (.DIODE(_02521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08355__B1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__A2 (.DIODE(_02521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08360__A (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08362__A2 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08362__B2 (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08380__A2 (.DIODE(_01209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08380__B1 (.DIODE(_02425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__A2 (.DIODE(_01209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__B1 (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08382__A2 (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08382__B1 (.DIODE(_01418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08384__A_N (.DIODE(_01437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08385__A2 (.DIODE(_01439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08385__B1 (.DIODE(_01418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08386__A1 (.DIODE(_01200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08386__C1 (.DIODE(_01441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__B2 (.DIODE(_02011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08390__A2 (.DIODE(_01442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08390__B1 (.DIODE(_02011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__B (.DIODE(_01302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08394__B (.DIODE(_01411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08396__A2 (.DIODE(_01349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08396__B1 (.DIODE(_01209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08397__A2 (.DIODE(_01209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08397__B1 (.DIODE(_02425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08398__B (.DIODE(_01349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08400__A2 (.DIODE(_02425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08400__B1 (.DIODE(_01591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__A2 (.DIODE(_01591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08402__A2 (.DIODE(_01411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08404__A1 (.DIODE(_01201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08404__A3 (.DIODE(_01362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08405__A2 (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08406__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__08407__A (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08412__C_N (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__08414__A2 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08414__B2 (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08415__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__08415__C (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08431__A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__08431__B1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08432__B2 (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08434__B1 (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__A2 (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__A1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__B1 (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__B (.DIODE(_02403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__A1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__B1 (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__B1 (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08449__A1 (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08449__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__08449__B1 (.DIODE(_02316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__B2 (.DIODE(_02521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__B1 (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08454__A (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08459__B1 (.DIODE(_02261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08471__B1 (.DIODE(_02789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__B1 (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08474__A2 (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__B1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__B2 (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08484__B1 (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08486__A2 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08486__B2 (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08505__B1 (.DIODE(_02224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08506__B2 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08519__A (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08520__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__08520__C1 (.DIODE(_02364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__A (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__B1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__C1 (.DIODE(_02364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__A (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__C1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__A2 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__B1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__C1 (.DIODE(_02364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__A2 (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__B1 (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08541__A1 (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08541__A2 (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08541__B1 (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08541__B2 (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__A1 (.DIODE(\genblk2[7].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__A2 (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__B1 (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08543__A1 (.DIODE(_02225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08547__A1 (.DIODE(\genblk2[6].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08547__A2 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08547__B1 (.DIODE(_02309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08547__B2 (.DIODE(\genblk2[6].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08552__A1 (.DIODE(\genblk2[6].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08552__B1 (.DIODE(\genblk2[6].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08553__A1 (.DIODE(\genblk2[6].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08553__A2 (.DIODE(\genblk2[6].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08553__B1 (.DIODE(_02261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08557__A1 (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08557__B1 (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08558__A1 (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08558__A2 (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08558__B1 (.DIODE(_02223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08560__A1 (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08560__A2 (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08562__C1 (.DIODE(\genblk2[7].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08564__B (.DIODE(_02521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08565__A1 (.DIODE(_02261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__B1 (.DIODE(_02316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__B2 (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08574__A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__08574__A3 (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08576__A1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08576__B1 (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__B1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08583__A2 (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08592__A2 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08592__B1 (.DIODE(_02521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__A2 (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__B1 (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08594__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__08594__B (.DIODE(_02364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__A2 (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__B1 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__C (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08603__A2 (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08604__A (.DIODE(_02261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08605__B (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08609__A2 (.DIODE(_02789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08610__C (.DIODE(_02789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08611__B (.DIODE(_02223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08612__A2 (.DIODE(_02521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08615__B1 (.DIODE(_02223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08617__A2 (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__A2 (.DIODE(_02733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__B1 (.DIODE(_02261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08634__A1 (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08634__A2 (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__A (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08636__A (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08636__C (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08637__A1 (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08639__B1 (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08640__A (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08656__B1 (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08658__A2 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08658__B2 (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08660__A (.DIODE(_02789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__A2 (.DIODE(_02789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__B1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__A2 (.DIODE(_02521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08666__B1 (.DIODE(_02316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08667__B2 (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08682__B1 (.DIODE(_02224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08683__B2 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08707__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__08707__B1 (.DIODE(_02224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08708__B2 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08728__B1 (.DIODE(_02224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08729__B2 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08746__C (.DIODE(\genblk2[6].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__C (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08749__A1 (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08749__A2 (.DIODE(_02309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08751__A (.DIODE(\genblk2[7].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08751__B (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08759__A2 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08760__A2 (.DIODE(_02521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08761__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__08762__A2 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08763__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__08786__B1 (.DIODE(_02224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08787__B2 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08827__A2 (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08827__B1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08828__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__08834__A2 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__08838__B (.DIODE(_03544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__B (.DIODE(_03544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08865__B1 (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08866__A2 (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08893__A (.DIODE(_01099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08899__B1 (.DIODE(_01157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08903__B1 (.DIODE(_01157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__B1 (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__S (.DIODE(_01157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08927__A (.DIODE(_01099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08933__B (.DIODE(_01157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08934__A1 (.DIODE(_01099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08943__C1 (.DIODE(_01155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08954__S (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08959__S (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08966__S (.DIODE(_01155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08978__S (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08979__B (.DIODE(_01157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08980__A1 (.DIODE(_01157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08982__A (.DIODE(_01097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08989__S (.DIODE(_01155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08994__A2 (.DIODE(_01099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08994__B1 (.DIODE(_01157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09013__A (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09014__C1 (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09016__A (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09017__A (.DIODE(_03689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09018__C1 (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09020__A (.DIODE(_02152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09022__A (.DIODE(_03693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09024__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09025__A2 (.DIODE(_03694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09025__B1 (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09029__A1 (.DIODE(_03694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09029__B1 (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09031__A (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09032__A (.DIODE(_03701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__B1 (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09035__A (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09036__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09036__B (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09037__A1 (.DIODE(_03704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09037__B1_N (.DIODE(_03705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09038__A (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09038__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09039__A (.DIODE(_02147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09040__A (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09041__A1 (.DIODE(_03706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09041__S (.DIODE(_03708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__A1 (.DIODE(_02002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__S (.DIODE(_03708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09045__A1 (.DIODE(_01991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09045__S (.DIODE(_03708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09047__A (.DIODE(_01248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09047__B (.DIODE(_02374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09048__A1 (.DIODE(_03712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09048__S (.DIODE(_03708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09050__A (.DIODE(_03708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09052__A (.DIODE(_03689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09052__B (.DIODE(_01242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09054__A1 (.DIODE(_03714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09054__C1 (.DIODE(_03717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09055__A1 (.DIODE(_03704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09056__A1 (.DIODE(_01201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09056__S (.DIODE(_03708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09058__A (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09059__A0 (.DIODE(_01229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09059__S (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09062__A (.DIODE(_03701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09063__S (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09065__S (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09067__A (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09069__A (.DIODE(_03701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09069__B (.DIODE(_01221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__B (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09071__A1 (.DIODE(_03726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09071__B1 (.DIODE(_01302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09071__B2 (.DIODE(_03727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09071__C1 (.DIODE(_03728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__A1 (.DIODE(_01340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__S (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__A1 (.DIODE(_01592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__S (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09076__A1 (.DIODE(_01483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09076__S (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09078__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__A (.DIODE(_03708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__B (.DIODE(_01210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__A1 (.DIODE(_03732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__B1 (.DIODE(_03733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09081__A1 (.DIODE(_03704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09081__B1_N (.DIODE(_03717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09083__A (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09083__B (.DIODE(_01201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09083__C (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09084__A (.DIODE(_03735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09085__A1 (.DIODE(_03714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09085__B1 (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__A (.DIODE(\modein.delay_octave_down_in[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09088__B1 (.DIODE(_01591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09088__C1 (.DIODE(_03738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__C (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__D (.DIODE(_03738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09091__A (.DIODE(_01201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__A (.DIODE(_01367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__A1 (.DIODE(_01367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__B2 (.DIODE(_01342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09094__A (.DIODE(_01367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09095__A0 (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09095__A1 (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__A1 (.DIODE(_01490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09157__A1 (.DIODE(_03804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09159__A1 (.DIODE(\genblk2[0].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09173__A (.DIODE(_01342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09173__B (.DIODE(_01441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__A1 (.DIODE(_03813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__S (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09176__A1 (.DIODE(_01368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09176__S (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09178__A1 (.DIODE(_01342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09178__S (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__A1 (.DIODE(_01356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__S (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__A1 (.DIODE(_01214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__S (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09184__A (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__A1 (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__A2 (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__B1 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09186__A1 (.DIODE(_03704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__A1 (.DIODE(_03714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__B1 (.DIODE(_03705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09189__A (.DIODE(_03701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09190__A1 (.DIODE(_03706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09190__S (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09192__A1 (.DIODE(_02002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09192__S (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09194__A1 (.DIODE(_01991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09194__S (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__A1 (.DIODE(_03712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__S (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09199__S (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__A1 (.DIODE(_01183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__S (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09203__A1 (.DIODE(_01302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09203__S (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09205__A1 (.DIODE(_03704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09205__B1_N (.DIODE(_03728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09206__A (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09207__A1 (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09207__B1_N (.DIODE(_03717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09209__A1 (.DIODE(_03714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09209__B1 (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09210__A (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09211__A (.DIODE(_03833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09215__A (.DIODE(_02152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__A (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__A2 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__B1 (.DIODE(_03804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__B2 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__A (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09220__A2 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09220__B1 (.DIODE(_03840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09220__B2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__A2 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__B1 (.DIODE(_03840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09222__A2 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09222__B1 (.DIODE(_03840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09223__A2 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09223__B1 (.DIODE(_03840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09224__A2 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09224__B1 (.DIODE(_03840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09225__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__09225__A2 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09225__B1 (.DIODE(_03840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__A2 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__B1 (.DIODE(_03840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__A2 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__B1 (.DIODE(_03840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09230__A2 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09230__B1 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09232__A2 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09232__B1 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09234__A2 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09234__B1 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09237__B1 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09238__A (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09239__B (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09249__A (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09252__A (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__A (.DIODE(_03855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09255__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09259__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09261__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09261__B (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09262__B1 (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09263__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09263__B (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__B1 (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09266__B1 (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__A (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09268__A (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09268__B (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09270__A2 (.DIODE(_03804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__A3 (.DIODE(_03804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__B2 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__A (.DIODE(_03804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__A1 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__B1 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09280__S (.DIODE(_03804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__B1 (.DIODE(_03840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09284__S (.DIODE(_03804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__B1 (.DIODE(_03840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09286__A (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__S (.DIODE(_03804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09293__S (.DIODE(_03804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__S (.DIODE(_03804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__A (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__A2 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09364__A2 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__A2 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__B1 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__A2 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__B1 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__A (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__A0 (.DIODE(_03941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__A1 (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09379__A (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__A1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__B1 (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09384__A1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09384__B1 (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__A (.DIODE(_03726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09388__B1 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__B_N (.DIODE(\genblk2[1].wave_shpr.div.b1[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__A_N (.DIODE(\genblk2[1].wave_shpr.div.b1[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__A1 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__S (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__A1 (.DIODE(\genblk2[1].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__S (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09452__S (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__S (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__S (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__S (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09460__S (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09462__S (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09464__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09464__S (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__A1 (.DIODE(_01327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__S (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__A1 (.DIODE(_03732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__B1 (.DIODE(_03733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09469__A1 (.DIODE(_01231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09469__S (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09471__A (.DIODE(_01418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09472__A (.DIODE(_03701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__A1 (.DIODE(_04023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09475__A1 (.DIODE(_01248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09477__A1 (.DIODE(_01437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09480__A1 (.DIODE(_04028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09482__A1 (.DIODE(_01183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09484__A1 (.DIODE(_01302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__A1 (.DIODE(_04032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09490__A1 (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09492__A (.DIODE(_01411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09493__A1 (.DIODE(_04036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09495__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09497__A (.DIODE(_03701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09498__A1 (.DIODE(_01327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09498__S (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09500__A1 (.DIODE(_03732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09500__B1 (.DIODE(_03733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09501__A1 (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09501__B1_N (.DIODE(_03717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__A1 (.DIODE(_03714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__B1 (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09505__A (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09506__A (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__A1 (.DIODE(\genblk2[1].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__A2 (.DIODE(_04043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__B1 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__B2 (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__A (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__A2 (.DIODE(_04043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__B1 (.DIODE(_04047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__B2 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA__09512__A2 (.DIODE(_04043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09512__B1 (.DIODE(_04047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09513__A2 (.DIODE(_04043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09513__B1 (.DIODE(_04047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09514__A2 (.DIODE(_04043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09514__B1 (.DIODE(_04047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__A2 (.DIODE(_04043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__B1 (.DIODE(_04047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09516__A1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__09516__A2 (.DIODE(_04043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09516__B1 (.DIODE(_04047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__A1 (.DIODE(\genblk2[1].wave_shpr.div.quo[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__A2 (.DIODE(_04043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__B1 (.DIODE(_04047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__B2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__09518__A2 (.DIODE(_04043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09518__B1 (.DIODE(_04047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09518__B2 (.DIODE(\genblk2[1].wave_shpr.div.quo[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09519__A (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__A (.DIODE(_03855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__A2 (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__B1 (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09522__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__A2 (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__B1 (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09524__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__A2 (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__B1 (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09526__A (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09527__A (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09528__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09530__A (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09535__A (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09536__A (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09538__B (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__A (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__B (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09544__B (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09546__B (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__B (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__B (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__A2 (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__B1 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__B (.DIODE(\genblk1[1].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09553__A2 (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09553__B1 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09555__A2 (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09555__B1 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09556__A (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09557__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09558__A2 (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09558__B1 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09559__B_N (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__A1 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09561__C (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__A2 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__A1 (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__B1 (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09565__S (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__A2 (.DIODE(_04043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__B1 (.DIODE(_04047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09567__A (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09570__S (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__B1 (.DIODE(_04047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09572__A (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09575__S (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09579__S (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09583__S (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09587__S (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__S (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09596__S (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__S (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09604__S (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09608__S (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__A (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__S (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__A (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09618__S (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09622__S (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09626__S (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09630__S (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09652__A2 (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09655__A1 (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09655__B1 (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__A2 (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__B1 (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__A2 (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__B1 (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09662__A0 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09662__A1 (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09666__A1 (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09666__B1 (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09670__A1 (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09670__B1 (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__A (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09674__B1 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09735__A1 (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09735__S (.DIODE(_00009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09737__S (.DIODE(_00009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__S (.DIODE(_00009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__S (.DIODE(_00009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09743__S (.DIODE(_00009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09745__S (.DIODE(_00009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09747__S (.DIODE(_00009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__S (.DIODE(_00009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09751__A (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09751__B (.DIODE(_01302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09752__A1 (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09752__S (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09754__A (.DIODE(_01436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09754__B (.DIODE(_01925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09755__A1 (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09755__S (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09758__A1 (.DIODE(_04227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09758__S (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09761__A (.DIODE(_01436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09761__B (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09762__A1 (.DIODE(_04230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09762__S (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09764__A1 (.DIODE(_01794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09764__S (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09766__A (.DIODE(_01302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09766__B (.DIODE(_03727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09767__A1 (.DIODE(_03704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09767__B1 (.DIODE(_04233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09768__A1 (.DIODE(_01262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09768__S (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__A1 (.DIODE(_02077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__S (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09772__A1 (.DIODE(_01256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09772__S (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09774__A1 (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09774__B1_N (.DIODE(_03733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09775__A1 (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09775__S (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09777__A (.DIODE(_03701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__A1 (.DIODE(_01487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__S (.DIODE(_04238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09780__A1 (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09780__S (.DIODE(_04238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09782__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09782__B (.DIODE(_01490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09783__A1 (.DIODE(_03732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09783__B1 (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09784__A (.DIODE(_01490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__A1 (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__S (.DIODE(_04238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09787__A1 (.DIODE(_01365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09787__S (.DIODE(_04238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09790__A1 (.DIODE(_03714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09790__B1 (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__A (.DIODE(_03833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09794__A (.DIODE(_04247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__A (.DIODE(_02152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09797__A (.DIODE(_04250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09798__A2 (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09798__B1 (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09798__B2 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09799__A (.DIODE(_04250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09800__A2 (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09800__B1 (.DIODE(_04252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__A2 (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__B1 (.DIODE(_04252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09802__A2 (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09802__B1 (.DIODE(_04252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09803__A2 (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09803__B1 (.DIODE(_04252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__A2 (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__B1 (.DIODE(_04252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__A2 (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__B1 (.DIODE(_04252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09806__A2 (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09806__B1 (.DIODE(_04252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09807__A1 (.DIODE(\genblk2[2].wave_shpr.div.quo[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09807__A2 (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09807__B1 (.DIODE(_04252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__A (.DIODE(_04247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09809__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09810__A2 (.DIODE(_04253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09810__B1 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09811__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09812__A2 (.DIODE(_04253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09812__B1 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09813__A (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09814__A2 (.DIODE(_04253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09814__B1 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09815__A (.DIODE(_04247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09816__A (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__B1 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09818__A (.DIODE(_04250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09819__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09821__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09823__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__A (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09829__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09831__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09835__A (.DIODE(_02147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09836__A (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09837__A (.DIODE(_04269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09839__A (.DIODE(_04269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09840__A2 (.DIODE(_04247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09841__A (.DIODE(_04269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09842__A2 (.DIODE(_04247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09842__B1 (.DIODE(_04250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__A (.DIODE(_04269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09844__A2 (.DIODE(_04247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09844__B1 (.DIODE(_04250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__A (.DIODE(_04269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09846__A2 (.DIODE(_04247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09846__B1 (.DIODE(_04250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09847__A (.DIODE(_04250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09848__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09850__A2 (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09851__A3 (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09852__B2 (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09855__A (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09856__A1 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09856__B1 (.DIODE(_04253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09857__A (.DIODE(_04247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__S (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09861__B1 (.DIODE(_04252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__S (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__B1 (.DIODE(_04252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__A (.DIODE(_04250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09869__S (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__S (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09877__S (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__A (.DIODE(_04247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09909__A (.DIODE(_04250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__A2 (.DIODE(_04253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09944__A2 (.DIODE(_04253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09946__A2 (.DIODE(_04253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09946__B1 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09950__A2 (.DIODE(_04253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09950__B1 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__A0 (.DIODE(_04250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__A1 (.DIODE(_04247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__A1 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__B1 (.DIODE(_04253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__A1 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__B1 (.DIODE(_04253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09962__A (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__B1 (.DIODE(_03855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09969__B_N (.DIODE(\genblk2[3].wave_shpr.div.b1[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10009__A_N (.DIODE(\genblk2[3].wave_shpr.div.b1[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10025__A (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10026__A (.DIODE(_04421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10027__A1 (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10029__A1 (.DIODE(\genblk2[3].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__A1 (.DIODE(_03732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__B1 (.DIODE(_03733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10045__A1 (.DIODE(_03714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10045__B1 (.DIODE(_03717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10046__B (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10047__A1_N (.DIODE(_03727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10047__A2_N (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10047__B2 (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10048__A1 (.DIODE(_01223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10048__S (.DIODE(_04238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10050__A1 (.DIODE(_01248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10050__S (.DIODE(_04238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10052__A1 (.DIODE(_01870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10052__S (.DIODE(_04238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10055__A1 (.DIODE(_04436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10055__S (.DIODE(_04238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__A1 (.DIODE(_01329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__S (.DIODE(_04238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10059__A1 (.DIODE(_01263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10059__S (.DIODE(_04238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__A (.DIODE(_03701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10062__A1 (.DIODE(_01240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10062__S (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10064__A1 (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10064__S (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__A1 (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__S (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10068__B (.DIODE(_01226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10069__A1 (.DIODE(_04444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10069__S (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10071__A1 (.DIODE(_01595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10071__S (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10073__A1 (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10073__S (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10075__A1 (.DIODE(_01365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10075__S (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10078__A1 (.DIODE(_03714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10078__B1 (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10079__A (.DIODE(_03833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10082__A (.DIODE(_04451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__A (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10085__A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__10085__A2 (.DIODE(_04452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10085__B1 (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10085__B2 (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10087__A (.DIODE(_04455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10088__A2 (.DIODE(_04452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10088__B1 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10088__B2 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__10089__A2 (.DIODE(_04452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10089__B1 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10090__A2 (.DIODE(_04452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10090__B1 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__A2 (.DIODE(_04452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__B1 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10092__A2 (.DIODE(_04452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10092__B1 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10093__A2 (.DIODE(_04452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10093__B1 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__A1 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__A2 (.DIODE(_04452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__B1 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10095__A1 (.DIODE(\genblk2[3].wave_shpr.div.quo[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10095__A2 (.DIODE(_04452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10095__B1 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10095__B2 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__A (.DIODE(_04451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10097__A (.DIODE(_04269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__B1 (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__B2 (.DIODE(\genblk2[3].wave_shpr.div.quo[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10099__A (.DIODE(_04269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10100__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10100__B1 (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10101__A (.DIODE(_04269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10102__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10102__B1 (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10103__A (.DIODE(_04451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__A (.DIODE(_04455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10105__A (.DIODE(_04269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10107__A (.DIODE(_04269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10109__A (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10122__A (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__A2 (.DIODE(_04451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__B1 (.DIODE(_04455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10129__A2 (.DIODE(_04451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10129__B1 (.DIODE(_04455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10131__A2 (.DIODE(_04451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10131__B1 (.DIODE(_04455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10132__A (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10133__A (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10134__A2 (.DIODE(_04451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10134__B1 (.DIODE(_04455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10135__B_N (.DIODE(_04455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__A1 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10138__A (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10139__A2 (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__A1 (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__B1 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__S (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__A2 (.DIODE(_04452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__B1 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__A (.DIODE(_04451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__S (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10149__B1 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__A (.DIODE(_04455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10153__S (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__S (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10160__S (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10164__S (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__S (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10173__S (.DIODE(_04507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10177__S (.DIODE(_04507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10181__S (.DIODE(_04507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__S (.DIODE(_04507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10187__A (.DIODE(_04451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10190__S (.DIODE(_04507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10192__A (.DIODE(_04455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__S (.DIODE(_04507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__S (.DIODE(_04507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10203__S (.DIODE(_04507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10207__S (.DIODE(_04507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10211__S (.DIODE(_04507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10213__B (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__A2 (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10224__A2_N (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10232__A2 (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10232__B1 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__B (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__B1 (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10238__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10238__B1 (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__A0 (.DIODE(_04455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__A1 (.DIODE(_04451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10243__A1 (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10243__B1 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__A1 (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__B1 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10250__A (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10251__B1 (.DIODE(_03855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__A1 (.DIODE(_01735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__S (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10331__A1 (.DIODE(_01304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10331__S (.DIODE(_03689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10332__A (.DIODE(_03717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10333__A1 (.DIODE(_03714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10333__B1 (.DIODE(_01262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10333__B2 (.DIODE(_03705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10334__A1 (.DIODE(_01240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10334__S (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__A1 (.DIODE(_01256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__S (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__A1 (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__B1_N (.DIODE(_03733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__A1 (.DIODE(_03732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__B1 (.DIODE(_03717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10340__A1 (.DIODE(_03714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10340__B1 (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10340__B2 (.DIODE(_03727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10341__A (.DIODE(_03701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10342__A1 (.DIODE(_01326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10342__S (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10344__A (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10345__S (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10347__A1 (.DIODE(_01658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10347__S (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10349__A1 (.DIODE(_01757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10349__S (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10351__A (.DIODE(_01355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10352__A1 (.DIODE(_04643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10352__S (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__A (.DIODE(_01490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__B (.DIODE(_01242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10355__A1 (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10355__S (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__A (.DIODE(_03708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__B (.DIODE(_01441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__C (.DIODE(_01367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__A1 (.DIODE(_03704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__B1 (.DIODE(_04647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__A1 (.DIODE(_01365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__S (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__A1 (.DIODE(_03726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__B1 (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10363__A (.DIODE(_03833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10366__A (.DIODE(_04651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10367__A (.DIODE(_02152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10369__A (.DIODE(_04654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10370__B2 (.DIODE(_04655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10371__A (.DIODE(_04654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10380__A (.DIODE(_04651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10381__A (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10382__A2 (.DIODE(_04657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10382__B1 (.DIODE(_04655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10383__A (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10384__A2 (.DIODE(_04657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10384__B1 (.DIODE(_04655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__A (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10386__A2 (.DIODE(_04657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10386__B1 (.DIODE(_04655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10387__A (.DIODE(_04651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10388__A (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10389__B1 (.DIODE(_04655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10390__A (.DIODE(_04654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__A (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10393__A (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10395__A (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10397__A (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10399__A (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10401__A (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10403__A (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10405__A (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10407__A (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10408__A (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__A (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10411__A2 (.DIODE(_04651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10412__A (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10413__A2 (.DIODE(_04651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10413__B1 (.DIODE(_04654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10414__A (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10415__A (.DIODE(_04676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10416__A2 (.DIODE(_04651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10416__B1 (.DIODE(_04654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__A (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__A2 (.DIODE(_04651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__B1 (.DIODE(_04654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10419__A (.DIODE(_04654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10420__A (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__A (.DIODE(_04651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__A (.DIODE(_04654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10453__S (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__S (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10461__S (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10465__S (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10467__A (.DIODE(_04651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10470__S (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10471__A2 (.DIODE(_04715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10474__S (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10475__A2 (.DIODE(_04715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10476__A (.DIODE(_04654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__S (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__A2 (.DIODE(_04715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10483__S (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10484__A2 (.DIODE(_04715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__S (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__A2 (.DIODE(_04715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10491__S (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__A2 (.DIODE(_04715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__A2 (.DIODE(_04715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10499__A2 (.DIODE(_04715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10503__A2 (.DIODE(_04715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10505__A2 (.DIODE(_04715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10509__A2 (.DIODE(_04657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10511__A2 (.DIODE(_04657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10514__A2 (.DIODE(_04657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10514__B1 (.DIODE(_04655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__A2 (.DIODE(_04657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__B1 (.DIODE(_04655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10520__A2 (.DIODE(_04657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10520__B1 (.DIODE(_04655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10521__A0 (.DIODE(_04654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10521__A1 (.DIODE(_04651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__A1 (.DIODE(_04655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__B1 (.DIODE(_04657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__A1 (.DIODE(_04655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__B1 (.DIODE(_04657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10532__A (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10533__B1 (.DIODE(_03855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10545__B_N (.DIODE(\genblk2[5].wave_shpr.div.b1[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10566__A_N (.DIODE(\genblk2[5].wave_shpr.div.b1[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10594__A1 (.DIODE(_04821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10594__S (.DIODE(_00015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10596__A1 (.DIODE(\genblk2[5].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10596__S (.DIODE(_00015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10598__S (.DIODE(_00015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10600__S (.DIODE(_00015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10602__S (.DIODE(_00015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10604__S (.DIODE(_00015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10606__S (.DIODE(_00015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__S (.DIODE(_00015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10610__A1 (.DIODE(_01189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10610__S (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10612__A (.DIODE(_01738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10613__S (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10615__A1 (.DIODE(_01684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10615__S (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10617__A (.DIODE(_03701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__S (.DIODE(_04834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10621__S (.DIODE(_04834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10624__S (.DIODE(_04834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10626__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10626__S (.DIODE(_04834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__A1 (.DIODE(_01189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__S (.DIODE(_04834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10630__S (.DIODE(_04834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10632__A1 (.DIODE(_01923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10632__S (.DIODE(_04834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10635__S (.DIODE(_04834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10637__A1 (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10637__S (.DIODE(_04834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10639__A1 (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10639__S (.DIODE(_04834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10641__A (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10642__A1 (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10642__S (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__A1 (.DIODE(_03704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__B1 (.DIODE(_04647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10645__A1 (.DIODE(_01365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10645__S (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__A1 (.DIODE(_03726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__B1 (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__A (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10651__A (.DIODE(_02183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10652__A (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__A2 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__B1 (.DIODE(_04821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__B2 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10656__A (.DIODE(_04856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__A2 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__B1 (.DIODE(_04857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10658__A2 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10658__B1 (.DIODE(_04857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10659__A2 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10659__B1 (.DIODE(_04857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10660__A2 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10660__B1 (.DIODE(_04857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10661__A2 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10661__B1 (.DIODE(_04857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10662__A2 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10662__B1 (.DIODE(_04857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10663__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__10663__A2 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10663__B1 (.DIODE(_04857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10664__A2 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10664__B1 (.DIODE(_04857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10664__B2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__A (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__B (.DIODE(\genblk1[5].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__A2 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__B1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10668__A (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10669__A2 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10669__B1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10672__A (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__A (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10676__A (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__A (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__A (.DIODE(_04676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10682__A (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__A (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10694__A2 (.DIODE(_02183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10694__B1 (.DIODE(_04856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10696__A2 (.DIODE(_02183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10696__B1 (.DIODE(_04856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10698__A2 (.DIODE(_02183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10698__B1 (.DIODE(_04856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__A2 (.DIODE(_02183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__B1 (.DIODE(_04856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10702__A2 (.DIODE(_02183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10702__B1 (.DIODE(_04856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10703__B_N (.DIODE(_04856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10704__A1 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__A (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10707__A2 (.DIODE(_04821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__B1 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10711__S (.DIODE(_04821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10712__A2 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10712__B1 (.DIODE(_04857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10713__A (.DIODE(_02183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__S (.DIODE(_04821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10717__B1 (.DIODE(_04857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10718__A (.DIODE(_04856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10721__S (.DIODE(_04821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10724__S (.DIODE(_04821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10728__S (.DIODE(_04821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10732__S (.DIODE(_04821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10736__S (.DIODE(_04821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10755__A (.DIODE(_02183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10760__A (.DIODE(_04856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10781__B (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10782__A2 (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10792__A2_N (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10796__A2 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10800__A2 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10800__B1 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10802__B (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10804__A2 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10804__B1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10806__A2 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10806__B1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__A0 (.DIODE(_04856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__A1 (.DIODE(_02183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__B1 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10814__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10814__B1 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10818__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10818__B1 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10820__B1 (.DIODE(_03708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10880__A0 (.DIODE(\genblk2[6].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10880__A1 (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10882__A0 (.DIODE(\genblk2[6].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10882__A1 (.DIODE(\genblk2[6].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10894__A0 (.DIODE(\genblk2[6].wave_shpr.div.fin_quo[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10896__A1 (.DIODE(_01514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10896__S (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__A1 (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__B1 (.DIODE(_04233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10900__A1 (.DIODE(_01991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10900__S (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10902__A1 (.DIODE(_01923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10902__S (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10904__A1 (.DIODE(_01799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10904__S (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10906__A (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10907__S (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10909__A1 (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10909__S (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__A0 (.DIODE(\genblk2[7].wave_shpr.div.b1[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__A1 (.DIODE(_04444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__S (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10913__A1 (.DIODE(_01819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10913__S (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10915__A (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10916__A1 (.DIODE(_01797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10916__S (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__S (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10920__A1 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10920__S (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10922__A1 (.DIODE(_01811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10922__S (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10924__A1 (.DIODE(_02374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10924__S (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10926__A1 (.DIODE(_03704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10926__B1 (.DIODE(_04647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__A1 (.DIODE(_01365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__S (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__A1 (.DIODE(_03726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__B1 (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10931__A (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10934__A (.DIODE(_05051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10935__A (.DIODE(_02152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10937__A (.DIODE(_05054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10938__A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__10938__A2 (.DIODE(_05052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10938__B1 (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10938__B2 (.DIODE(_05055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10939__A (.DIODE(_05054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__A2 (.DIODE(_05052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__B1 (.DIODE(_05056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__B2 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__10941__A2 (.DIODE(_05052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10941__B1 (.DIODE(_05056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__A2 (.DIODE(_05052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__B1 (.DIODE(_05056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__A2 (.DIODE(_05052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__B1 (.DIODE(_05056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__A2 (.DIODE(_05052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__B1 (.DIODE(_05056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10945__A2 (.DIODE(_05052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10945__B1 (.DIODE(_05056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10946__A2 (.DIODE(_05052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10946__B1 (.DIODE(_05056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__A2 (.DIODE(_05052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__B1 (.DIODE(_05056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10948__A (.DIODE(_05051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__A2 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__B1 (.DIODE(_05055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__A (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10953__A2 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10953__B1 (.DIODE(_05055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10954__A (.DIODE(_04676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__A2 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__B1 (.DIODE(_05055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10956__A (.DIODE(_05051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10958__B1 (.DIODE(_05055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10959__A (.DIODE(_05054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10966__A (.DIODE(_04676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10978__A (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__A (.DIODE(_05074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__A2 (.DIODE(_05051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10981__A (.DIODE(_05074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10982__A2 (.DIODE(_05051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10982__B1 (.DIODE(_05054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10983__A (.DIODE(_05074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__A2 (.DIODE(_05051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__B1 (.DIODE(_05054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10985__A (.DIODE(_05074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10986__A2 (.DIODE(_05051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10986__B1 (.DIODE(_05054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10987__A (.DIODE(_05054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10988__A (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10990__A2 (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10991__A3 (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10992__B2 (.DIODE(_05052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10995__A (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10996__A1 (.DIODE(_05055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10996__B1 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10997__A (.DIODE(_05051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11000__S (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11001__B1 (.DIODE(_05056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11004__S (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11005__B1 (.DIODE(_05056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11006__A (.DIODE(_05054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11009__S (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11013__S (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11017__S (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__A (.DIODE(_05051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11049__A (.DIODE(_05054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11080__A2 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11083__A2 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11085__A2 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11085__B1 (.DIODE(_05055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11089__A2 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11089__B1 (.DIODE(_05055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11090__A0 (.DIODE(_05054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11090__A1 (.DIODE(_05051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11094__A1 (.DIODE(_05055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11094__B1 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11098__A1 (.DIODE(_05055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11098__B1 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11101__A (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11102__B1 (.DIODE(_03855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11114__B_N (.DIODE(\genblk2[7].wave_shpr.div.b1[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11135__A_N (.DIODE(\genblk2[7].wave_shpr.div.b1[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11163__A0 (.DIODE(\genblk2[7].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11163__A1 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11179__A1 (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11179__B1_N (.DIODE(_03705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11180__A (.DIODE(_03708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11180__B (.DIODE(\genblk2[8].wave_shpr.div.b1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11181__A1 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11181__A2 (.DIODE(_01242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11181__A3 (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__A1 (.DIODE(_03732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__B1 (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11183__A1 (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11183__S (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11185__A1_N (.DIODE(_03727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11185__A2_N (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11185__B2 (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__A1 (.DIODE(_01508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__S (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__A1 (.DIODE(_01507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__S (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11190__A1 (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11190__B1_N (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__A1 (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__S (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11194__A (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11195__A1 (.DIODE(_05236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11198__A1 (.DIODE(_05239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11200__A1 (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11202__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11203__A1 (.DIODE(_03726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11203__A2 (.DIODE(_01869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11204__A1_N (.DIODE(_03727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11204__A2_N (.DIODE(_01490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11204__B1 (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11205__A1 (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11205__B1_N (.DIODE(_03728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11206__A1 (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11206__B1_N (.DIODE(_03717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11208__A1 (.DIODE(_03726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11208__B1 (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11209__A (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11212__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11213__A (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__A2 (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__B1 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__B2 (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11217__A (.DIODE(_05249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11218__A2 (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11218__B1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__A2 (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__B1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11220__A2 (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11220__B1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11221__A2 (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11221__B1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11222__A2 (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11222__B1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11223__A2 (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11223__B1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11224__A2 (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11224__B1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__A2 (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__B1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11226__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__A (.DIODE(_05074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11228__B1 (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11229__A (.DIODE(_05074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11230__B1 (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11231__A (.DIODE(_05074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__B1 (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11233__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11234__A (.DIODE(_05249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__A (.DIODE(_05074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__A (.DIODE(_05074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11239__A (.DIODE(_05074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11241__A (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11257__A2 (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11257__B1 (.DIODE(_05249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11259__A2 (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11259__B1 (.DIODE(_05249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__A2 (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__B1 (.DIODE(_05249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11262__A (.DIODE(_04676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11263__A2 (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11263__B1 (.DIODE(_05249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11264__B_N (.DIODE(_05249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11265__A1 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__A2 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11269__A1 (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__S (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11273__A2 (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11273__B1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11274__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11277__S (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__A2 (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__B1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11279__A (.DIODE(_05249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11282__S (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__A2 (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__B1 (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11285__S (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__A2 (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__B1 (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11289__S (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11290__A2 (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11290__B1 (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11293__S (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11294__A2 (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11294__B1 (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11297__S (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11298__A2 (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11298__B1 (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11303__A2 (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11303__B1 (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11307__A2 (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11307__B1 (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11311__A2 (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11311__B1 (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11315__A2 (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11315__B1 (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11316__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11320__B1 (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11321__A (.DIODE(_05249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11361__A2 (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__B1 (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11367__B1 (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11368__A0 (.DIODE(_05249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11368__A1 (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__A1 (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11376__A1 (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__A (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11380__B1 (.DIODE(_03855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11387__B_N (.DIODE(\genblk2[8].wave_shpr.div.b1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11398__B (.DIODE(\genblk2[8].wave_shpr.div.b1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11400__A (.DIODE(\genblk2[8].wave_shpr.div.b1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11422__A_N (.DIODE(\genblk2[8].wave_shpr.div.b1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11442__A0 (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11442__A1 (.DIODE(_05417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11444__A0 (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11446__A0 (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11448__A0 (.DIODE(\genblk2[8].wave_shpr.div.fin_quo[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11458__A1 (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11460__A1 (.DIODE(_01819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__A1 (.DIODE(_01797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11464__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11466__A1 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11468__A1 (.DIODE(_01811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11470__A1 (.DIODE(_01946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11472__A (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11473__A1 (.DIODE(_04230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11477__A1 (.DIODE(_03704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11477__B1 (.DIODE(_04233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11478__A1 (.DIODE(_01227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11480__A1 (.DIODE(_01732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__A1 (.DIODE(_02656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__A1_N (.DIODE(_03727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__A2_N (.DIODE(_01490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__B1 (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__A1 (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__B1_N (.DIODE(_03728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11486__A1 (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11486__B1_N (.DIODE(_03717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__A1 (.DIODE(_03726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__B1 (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11489__A (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11492__A (.DIODE(_05441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11493__A (.DIODE(_02152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11495__A (.DIODE(_05444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__B1 (.DIODE(_05417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11497__A (.DIODE(_05444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11498__B1 (.DIODE(_05446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11499__B1 (.DIODE(_05446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11500__B1 (.DIODE(_05446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11501__B1 (.DIODE(_05446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11502__B1 (.DIODE(_05446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11503__B1 (.DIODE(_05446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11504__B1 (.DIODE(_05446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11505__A (.DIODE(_05441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11506__B1 (.DIODE(_05446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11507__A (.DIODE(_05441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11508__A (.DIODE(_05444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11509__A (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11510__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__A2 (.DIODE(_05448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__B1 (.DIODE(_05449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11513__A2 (.DIODE(_05448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11513__B1 (.DIODE(_05449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11514__A (.DIODE(_04676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11515__A2 (.DIODE(_05448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11515__B1 (.DIODE(_05449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11516__A (.DIODE(_05441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11518__B1 (.DIODE(_05449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11519__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11520__B1 (.DIODE(_05449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11521__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11522__B1 (.DIODE(_05449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11523__A (.DIODE(_05444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11524__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11526__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11534__A (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11535__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11540__A2 (.DIODE(_05441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11541__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11542__A2 (.DIODE(_05441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11544__A2 (.DIODE(_05441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11545__B (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11546__A2 (.DIODE(_05441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11546__B1 (.DIODE(_05444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__A (.DIODE(_05444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11548__A (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11549__C1 (.DIODE(_05472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11550__A2 (.DIODE(_05417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11551__A3 (.DIODE(_05417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__A (.DIODE(_05417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11556__A1 (.DIODE(_05449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11556__B1 (.DIODE(_05448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__S (.DIODE(_05417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11560__B1 (.DIODE(_05446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__S (.DIODE(_05417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11564__B1 (.DIODE(_05446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__A (.DIODE(_05444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__S (.DIODE(_05417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11572__S (.DIODE(_05417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11595__A (.DIODE(_05441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11636__A1 (.DIODE(_05449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11636__B1 (.DIODE(_05448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__B1 (.DIODE(_05417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11642__A2 (.DIODE(_05448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11644__A2 (.DIODE(_05448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11647__A2 (.DIODE(_05448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11648__A0 (.DIODE(_05444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11648__A1 (.DIODE(_05441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11652__A1 (.DIODE(_05449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11652__B1 (.DIODE(_05448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__A1 (.DIODE(_05449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__B1 (.DIODE(_05448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11659__A (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11660__B1 (.DIODE(_03855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11722__A1 (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11722__S (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11724__S (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__S (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__S (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__S (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11732__S (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11734__S (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11736__S (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11738__A (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__A1_N (.DIODE(_01099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__A1_N (.DIODE(_01099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11741__A1 (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11742__A1 (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11743__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11744__A (.DIODE(_03693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11745__A2 (.DIODE(_05623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11745__B1 (.DIODE(_05624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11745__B2 (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11746__A2 (.DIODE(_05623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11746__B1 (.DIODE(_05624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11747__A2 (.DIODE(_05623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11747__B1 (.DIODE(_05624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11748__A2 (.DIODE(_05623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11748__B1 (.DIODE(_05624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11749__A2 (.DIODE(_05623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11749__B1 (.DIODE(_05624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11750__A2 (.DIODE(_05623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11750__B1 (.DIODE(_05624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11751__A2 (.DIODE(_05623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11751__B1 (.DIODE(_05624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11752__A2 (.DIODE(_05623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11752__B1 (.DIODE(_05624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11753__A1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__11753__A2 (.DIODE(_05623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11753__B1 (.DIODE(_05624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11754__B (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11755__A2 (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11755__B1 (.DIODE(_03694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11755__B2 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__B (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11757__A2 (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11757__B1 (.DIODE(_03694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11758__B (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11759__A2 (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11759__B1 (.DIODE(_03694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11761__A (.DIODE(_03693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__B (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__A (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11765__B (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11767__B (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11773__A (.DIODE(_04676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11775__A (.DIODE(_04676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11777__A (.DIODE(_04676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11783__B (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11784__A2 (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11784__B1 (.DIODE(_03693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11785__B (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11786__A2 (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11786__B1 (.DIODE(_03693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11787__B (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11788__A2 (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11788__B1 (.DIODE(_03693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11789__B (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11790__A2 (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11790__B1 (.DIODE(_03693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11791__B_N (.DIODE(_03693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11792__A1 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11792__A2 (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11795__A2 (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11796__A1 (.DIODE(_03694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11796__B1 (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11799__S (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11800__A2 (.DIODE(_05623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11800__B1 (.DIODE(_05624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11801__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11802__A (.DIODE(_03693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11805__S (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11809__S (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11812__S (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11816__S (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11820__S (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11824__S (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11844__A (.DIODE(_03693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__A2 (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__B1 (.DIODE(_03694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11888__A1 (.DIODE(_03694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11888__B1 (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11892__A2 (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11892__B1 (.DIODE(_03694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11894__A2 (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11894__B1 (.DIODE(_03694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11895__A0 (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11899__A1 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11899__B1 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11903__A1 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11903__B1 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11906__A (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11907__B1 (.DIODE(_03855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11966__A1 (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11968__A1 (.DIODE(\genblk2[10].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11980__A1 (.DIODE(\genblk2[10].wave_shpr.div.quo[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11982__A1 (.DIODE(_01441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11982__B1 (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11983__A1 (.DIODE(_03732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11983__B1 (.DIODE(_05796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11984__A1 (.DIODE(_03813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11986__A1 (.DIODE(_01811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11988__A1 (.DIODE(_01946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11990__A1 (.DIODE(_04230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11992__A1 (.DIODE(_01855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11994__A (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__A1 (.DIODE(_02805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__S (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__A1 (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__S (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11999__A1 (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11999__B1_N (.DIODE(_03705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12000__A1 (.DIODE(_03706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12000__S (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__A1 (.DIODE(_02002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__S (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__A0 (.DIODE(\genblk2[11].wave_shpr.div.b1[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__A1 (.DIODE(_01500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__S (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__A1 (.DIODE(_01494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__S (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12008__A1 (.DIODE(_01483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12008__S (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12010__A1 (.DIODE(_03732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12010__B1 (.DIODE(_03733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12011__A1 (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12011__B1_N (.DIODE(_03717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12013__A1 (.DIODE(_03726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12013__B1 (.DIODE(_03735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12014__A (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__A (.DIODE(_02152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12020__A (.DIODE(_05815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12021__A1 (.DIODE(\genblk2[10].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12021__A2 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12021__B1 (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12021__B2 (.DIODE(_05816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12022__A (.DIODE(_05815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12023__A2 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12023__B1 (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12024__A2 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12024__B1 (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12025__A2 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12025__B1 (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12026__A2 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12026__B1 (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12027__A2 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12027__B1 (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12028__A1 (.DIODE(\genblk2[10].wave_shpr.div.quo[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12028__A2 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12028__B1 (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12029__A2 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12029__B1 (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12029__B2 (.DIODE(\genblk2[10].wave_shpr.div.quo[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12030__A1 (.DIODE(\genblk2[10].wave_shpr.div.quo[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12030__A2 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12030__B1 (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12032__A (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12034__A2 (.DIODE(_05818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12034__B1 (.DIODE(_05816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12034__B2 (.DIODE(\genblk2[10].wave_shpr.div.quo[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12036__A2 (.DIODE(_05818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12036__B1 (.DIODE(_05816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12038__A2 (.DIODE(_05818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12038__B1 (.DIODE(_05816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12041__B1 (.DIODE(_05816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12042__A (.DIODE(_05815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12043__A (.DIODE(_04676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12051__A (.DIODE(_03833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12059__A (.DIODE(_03833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__A (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12064__A (.DIODE(_03833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12065__B1 (.DIODE(_05815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12067__B1 (.DIODE(_05815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12069__B1 (.DIODE(_05815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12070__A (.DIODE(_05815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12071__A (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12073__A2 (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12074__A3 (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12075__B2 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12078__S (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12079__A2 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12079__B1 (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12082__S (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12083__A2 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12083__B1 (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12084__A (.DIODE(_05815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12087__S (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12088__A2 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12091__S (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12092__A2 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12095__S (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12096__A2 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12099__S (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12100__A2 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12104__S (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12105__A2 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__S (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12109__A2 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12112__S (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12113__A2 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12116__S (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__A2 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12121__S (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12125__S (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12127__A (.DIODE(_05815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12130__S (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12134__S (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12138__S (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__S (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12160__A2 (.DIODE(_05818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12163__A2 (.DIODE(_05818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12166__A1 (.DIODE(_05816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12166__B1 (.DIODE(_05818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12169__A2 (.DIODE(_05818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12169__B1 (.DIODE(_05816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12172__A2 (.DIODE(_05818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12172__B1 (.DIODE(_05816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12173__A0 (.DIODE(_05815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__A1 (.DIODE(_05816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__B1 (.DIODE(_05818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__A1 (.DIODE(_05816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__B1 (.DIODE(_05818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12184__A (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12185__B1 (.DIODE(_03855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12193__B_N (.DIODE(\genblk2[11].wave_shpr.div.b1[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12225__A_N (.DIODE(\genblk2[11].wave_shpr.div.b1[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12245__A1 (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12261__A1 (.DIODE(_01329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12261__S (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12263__A1 (.DIODE(_01263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12263__S (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12265__A1 (.DIODE(_01240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12265__S (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12267__A (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12268__A1 (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12270__A1 (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12275__A1 (.DIODE(_01311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12277__A1 (.DIODE(_02001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12279__A0 (.DIODE(_01308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12279__S (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__A1 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12283__A1 (.DIODE(_01946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12285__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12286__A1 (.DIODE(_03726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12287__A (.DIODE(_01337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12290__A1 (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__A1 (.DIODE(_01327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12294__A1 (.DIODE(_03732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12294__B1 (.DIODE(_03733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12295__A1 (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12296__A1 (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12296__B1_N (.DIODE(_03735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12297__A (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12298__A (.DIODE(_03941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__A2 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__B1 (.DIODE(_06010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__B2 (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__A2 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__B1 (.DIODE(_06010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__A2 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__B1 (.DIODE(_06010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12302__A2 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12302__B1 (.DIODE(_06010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12303__A2 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12303__B1 (.DIODE(_06010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12304__A2 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12304__B1 (.DIODE(_06010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12305__A1 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__12305__A2 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12305__B1 (.DIODE(_06010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12306__A2 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12306__B1 (.DIODE(_06010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12306__B2 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__12307__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__12307__A2 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12307__B1 (.DIODE(_06010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__A2 (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__B1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__B2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__12311__A2 (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12311__B1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12313__A2 (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12313__B1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12314__A (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12315__A (.DIODE(_03941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12324__A (.DIODE(_03689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12326__A (.DIODE(_03689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12328__A (.DIODE(_03689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12330__A (.DIODE(_03689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12332__A (.DIODE(_03833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12334__A (.DIODE(_03689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12336__A (.DIODE(_03689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12337__A2 (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12337__B1 (.DIODE(_03941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12338__A (.DIODE(_03833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__A2 (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__B1 (.DIODE(_03941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__A (.DIODE(_03833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__A2 (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__B1 (.DIODE(_03941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12342__A (.DIODE(_03689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__A1 (.DIODE(\genblk2[11].wave_shpr.div.acc_next[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__A2 (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__B1 (.DIODE(_03941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12344__A (.DIODE(\genblk2[11].wave_shpr.div.acc_next[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12344__B_N (.DIODE(_03941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12345__A1 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12345__A2 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__12346__C (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12347__A2 (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12348__A1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12348__B1 (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12351__A (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12352__A1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12352__B1 (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12355__S (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12356__A2 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12356__B1 (.DIODE(_06010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12357__A (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12358__A (.DIODE(_03941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12361__S (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12365__S (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12369__S (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12373__S (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12400__A (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12401__A (.DIODE(_03941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__A2 (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__B1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__A2 (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__B1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__A2 (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__B1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12451__CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12451__RESET_B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__12452__D (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__12452__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__12474__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__12475__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__12477__RESET_B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__12478__RESET_B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__12479__RESET_B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__12480__RESET_B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__12490__RESET_B (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__12491__RESET_B (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__12493__RESET_B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__12496__RESET_B (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__12582__RESET_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__12586__RESET_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__12614__RESET_B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__12623__RESET_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__12624__RESET_B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__RESET_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__12626__RESET_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__12631__RESET_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__12632__RESET_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__12633__RESET_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__12634__RESET_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__12635__RESET_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__12636__RESET_B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__12638__RESET_B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__RESET_B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__12663__RESET_B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__RESET_B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__12666__RESET_B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__12667__RESET_B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__12688__RESET_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__12762__SET_B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__12844__D (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12844__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__12886__RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__12890__RESET_B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__12891__RESET_B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__12892__RESET_B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__12893__RESET_B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__12911__RESET_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__12912__RESET_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__12930__D (.DIODE(_00009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12930__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__12938__RESET_B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__12939__RESET_B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__12940__RESET_B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__12941__RESET_B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__12981__RESET_B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__13000__RESET_B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__13056__RESET_B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__13073__RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__13080__RESET_B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__13081__RESET_B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__13094__RESET_B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__13165__RESET_B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__13170__RESET_B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__13180__RESET_B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__13181__RESET_B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__13188__D (.DIODE(_00015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13206__RESET_B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__13208__RESET_B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__13236__RESET_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__13260__RESET_B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__13261__RESET_B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__13262__RESET_B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__13263__RESET_B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__13264__RESET_B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__13265__RESET_B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__13266__RESET_B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__13267__RESET_B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__13268__RESET_B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__13295__RESET_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__13316__RESET_B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__13317__RESET_B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__13329__RESET_B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__13330__RESET_B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__13338__RESET_B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__13388__RESET_B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__13394__RESET_B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__13516__RESET_B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__13517__RESET_B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__13532__D (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13546__RESET_B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__13547__RESET_B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__13548__RESET_B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__13549__RESET_B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__13550__RESET_B (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__13558__RESET_B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__13596__RESET_B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__13597__RESET_B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__13598__RESET_B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__13599__RESET_B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__13600__RESET_B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__13632__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__13633__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__13648__RESET_B (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__13649__RESET_B (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__13757__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__13759__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__13760__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__13765__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__13766__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__13768__RESET_B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__13769__RESET_B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__13773__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__13774__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_100_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_101_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_102_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_103_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_104_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_105_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_106_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_107_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_108_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_109_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_110_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_111_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_112_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_113_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_114_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_115_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_116_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_117_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_118_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_119_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_120_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_121_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_122_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_123_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_124_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_125_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_126_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_127_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_128_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_129_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_130_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_131_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_132_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_133_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_134_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_135_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_136_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_137_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_138_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_139_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_78_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_79_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_80_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_81_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_82_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_83_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_84_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_85_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_86_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_87_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_88_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_89_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_90_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_91_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_92_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_93_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_94_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_95_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_96_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_97_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_98_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_99_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout38_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout39_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout40_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout43_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout44_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout47_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout48_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout49_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout57_A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout65_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout67_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout69_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1002_A (.DIODE(\genblk1[11].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1124_A (.DIODE(\genblk2[5].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4_A (.DIODE(\modein.delay_in[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold522_A (.DIODE(\genblk2[10].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold546_A (.DIODE(\genblk2[1].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold574_A (.DIODE(\genblk2[6].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold576_A (.DIODE(\genblk2[3].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold586_A (.DIODE(\genblk2[0].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold7_A (.DIODE(\modein.delay_octave_down_in[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold82_A (.DIODE(\genblk2[2].wave_shpr.div.quo[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold838_A (.DIODE(\genblk2[5].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold874_A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold879_A (.DIODE(\genblk2[5].wave_shpr.div.b1[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold902_A (.DIODE(\genblk1[5].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold903_A (.DIODE(\genblk2[1].wave_shpr.div.b1[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold915_A (.DIODE(\genblk1[0].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold918_A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold929_A (.DIODE(\genblk2[8].wave_shpr.div.b1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold934_A (.DIODE(\genblk2[3].wave_shpr.div.b1[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold944_A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold967_A (.DIODE(\genblk1[8].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold976_A (.DIODE(\genblk1[9].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap34_A (.DIODE(_01794_));
 sky130_fd_sc_hd__diode_2 ANTENNA_output17_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_output18_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire32_A (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire33_A (.DIODE(_02348_));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_812 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_871 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__and3_1 _06105_ (.A(\smpl_rt_clkdiv.clkDiv_inst.cnt[1] ),
    .B(\smpl_rt_clkdiv.clkDiv_inst.cnt[0] ),
    .C(\smpl_rt_clkdiv.clkDiv_inst.cnt[2] ),
    .X(_01086_));
 sky130_fd_sc_hd__and2_1 _06106_ (.A(\smpl_rt_clkdiv.clkDiv_inst.cnt[3] ),
    .B(_01086_),
    .X(_01087_));
 sky130_fd_sc_hd__and3_1 _06107_ (.A(\smpl_rt_clkdiv.clkDiv_inst.cnt[5] ),
    .B(\smpl_rt_clkdiv.clkDiv_inst.cnt[4] ),
    .C(_01087_),
    .X(_01088_));
 sky130_fd_sc_hd__and3_1 _06108_ (.A(net1179),
    .B(net395),
    .C(_01088_),
    .X(_01089_));
 sky130_fd_sc_hd__clkbuf_1 _06109_ (.A(_01089_),
    .X(\smpl_rt_clkdiv.clkDiv_inst.next_hzX ));
 sky130_fd_sc_hd__inv_2 _06110_ (.A(net338),
    .Y(\smpl_rt_clkdiv.clkDiv_inst.next_cnt[0] ));
 sky130_fd_sc_hd__xor2_1 _06111_ (.A(net364),
    .B(net338),
    .X(\smpl_rt_clkdiv.clkDiv_inst.next_cnt[1] ));
 sky130_fd_sc_hd__a21oi_1 _06112_ (.A1(\smpl_rt_clkdiv.clkDiv_inst.cnt[1] ),
    .A2(net338),
    .B1(net359),
    .Y(_01090_));
 sky130_fd_sc_hd__nor2_1 _06113_ (.A(_01086_),
    .B(net360),
    .Y(\smpl_rt_clkdiv.clkDiv_inst.next_cnt[2] ));
 sky130_fd_sc_hd__nor2_1 _06114_ (.A(net368),
    .B(_01086_),
    .Y(_01091_));
 sky130_fd_sc_hd__nor2_1 _06115_ (.A(_01087_),
    .B(_01091_),
    .Y(\smpl_rt_clkdiv.clkDiv_inst.next_cnt[3] ));
 sky130_fd_sc_hd__xor2_1 _06116_ (.A(net380),
    .B(_01087_),
    .X(\smpl_rt_clkdiv.clkDiv_inst.next_cnt[4] ));
 sky130_fd_sc_hd__a21oi_1 _06117_ (.A1(net380),
    .A2(_01087_),
    .B1(net407),
    .Y(_01092_));
 sky130_fd_sc_hd__nor2_1 _06118_ (.A(_01088_),
    .B(_01092_),
    .Y(\smpl_rt_clkdiv.clkDiv_inst.next_cnt[5] ));
 sky130_fd_sc_hd__xor2_1 _06119_ (.A(net365),
    .B(_01088_),
    .X(\smpl_rt_clkdiv.clkDiv_inst.next_cnt[6] ));
 sky130_fd_sc_hd__a21oi_1 _06120_ (.A1(net365),
    .A2(_01088_),
    .B1(net395),
    .Y(_01093_));
 sky130_fd_sc_hd__nor2_1 _06121_ (.A(\smpl_rt_clkdiv.clkDiv_inst.next_hzX ),
    .B(_01093_),
    .Y(\smpl_rt_clkdiv.clkDiv_inst.next_cnt[7] ));
 sky130_fd_sc_hd__or4_2 _06122_ (.A(\genblk2[9].wave_shpr.div.done ),
    .B(\genblk2[8].wave_shpr.div.done ),
    .C(\genblk2[11].wave_shpr.div.done ),
    .D(\genblk2[10].wave_shpr.div.done ),
    .X(_01094_));
 sky130_fd_sc_hd__or4_4 _06123_ (.A(\genblk2[5].wave_shpr.div.done ),
    .B(\genblk2[4].wave_shpr.div.done ),
    .C(\genblk2[7].wave_shpr.div.done ),
    .D(\genblk2[6].wave_shpr.div.done ),
    .X(_01095_));
 sky130_fd_sc_hd__or4_2 _06124_ (.A(\genblk2[1].wave_shpr.div.done ),
    .B(\genblk2[0].wave_shpr.div.done ),
    .C(\genblk2[3].wave_shpr.div.done ),
    .D(\genblk2[2].wave_shpr.div.done ),
    .X(_01096_));
 sky130_fd_sc_hd__nor3_2 _06125_ (.A(_01094_),
    .B(_01095_),
    .C(_01096_),
    .Y(_01097_));
 sky130_fd_sc_hd__clkbuf_4 _06126_ (.A(_01097_),
    .X(_01098_));
 sky130_fd_sc_hd__buf_2 _06127_ (.A(_01098_),
    .X(_01099_));
 sky130_fd_sc_hd__or2_1 _06128_ (.A(net13),
    .B(net15),
    .X(_01100_));
 sky130_fd_sc_hd__nand2_1 _06129_ (.A(net13),
    .B(net15),
    .Y(_01101_));
 sky130_fd_sc_hd__nand2_1 _06130_ (.A(_01100_),
    .B(_01101_),
    .Y(_01102_));
 sky130_fd_sc_hd__xor2_1 _06131_ (.A(net3),
    .B(_01102_),
    .X(_01103_));
 sky130_fd_sc_hd__nand2_1 _06132_ (.A(net8),
    .B(net9),
    .Y(_01104_));
 sky130_fd_sc_hd__or2_1 _06133_ (.A(net8),
    .B(net9),
    .X(_01105_));
 sky130_fd_sc_hd__nand2_1 _06134_ (.A(_01104_),
    .B(_01105_),
    .Y(_01106_));
 sky130_fd_sc_hd__xor2_1 _06135_ (.A(net11),
    .B(_01106_),
    .X(_01107_));
 sky130_fd_sc_hd__nand2_1 _06136_ (.A(net1),
    .B(net7),
    .Y(_01108_));
 sky130_fd_sc_hd__or2_1 _06137_ (.A(net1),
    .B(net7),
    .X(_01109_));
 sky130_fd_sc_hd__nand2_1 _06138_ (.A(_01108_),
    .B(_01109_),
    .Y(_01110_));
 sky130_fd_sc_hd__xor2_1 _06139_ (.A(_01107_),
    .B(_01110_),
    .X(_01111_));
 sky130_fd_sc_hd__xnor2_1 _06140_ (.A(_01103_),
    .B(_01111_),
    .Y(_01112_));
 sky130_fd_sc_hd__nand2_1 _06141_ (.A(net14),
    .B(_01112_),
    .Y(_01113_));
 sky130_fd_sc_hd__inv_2 _06142_ (.A(net2),
    .Y(_01114_));
 sky130_fd_sc_hd__or2_1 _06143_ (.A(net14),
    .B(_01112_),
    .X(_01115_));
 sky130_fd_sc_hd__nand2_1 _06144_ (.A(_01113_),
    .B(_01115_),
    .Y(_01116_));
 sky130_fd_sc_hd__or2_1 _06145_ (.A(_01114_),
    .B(_01116_),
    .X(_01117_));
 sky130_fd_sc_hd__a21bo_1 _06146_ (.A1(net11),
    .A2(_01105_),
    .B1_N(_01104_),
    .X(_01118_));
 sky130_fd_sc_hd__and3_1 _06147_ (.A(net1),
    .B(net7),
    .C(_01118_),
    .X(_01119_));
 sky130_fd_sc_hd__and2b_1 _06148_ (.A_N(_01118_),
    .B(_01108_),
    .X(_01120_));
 sky130_fd_sc_hd__nor2_1 _06149_ (.A(_01119_),
    .B(_01120_),
    .Y(_01121_));
 sky130_fd_sc_hd__and2b_1 _06150_ (.A_N(_01103_),
    .B(_01111_),
    .X(_01122_));
 sky130_fd_sc_hd__o21bai_1 _06151_ (.A1(_01107_),
    .A2(_01110_),
    .B1_N(_01122_),
    .Y(_01123_));
 sky130_fd_sc_hd__xnor2_1 _06152_ (.A(_01121_),
    .B(_01123_),
    .Y(_01124_));
 sky130_fd_sc_hd__a21boi_1 _06153_ (.A1(net3),
    .A2(_01100_),
    .B1_N(_01101_),
    .Y(_01125_));
 sky130_fd_sc_hd__nor2_1 _06154_ (.A(_01124_),
    .B(_01125_),
    .Y(_01126_));
 sky130_fd_sc_hd__and2_1 _06155_ (.A(_01124_),
    .B(_01125_),
    .X(_01127_));
 sky130_fd_sc_hd__or2_1 _06156_ (.A(_01126_),
    .B(_01127_),
    .X(_01128_));
 sky130_fd_sc_hd__a21oi_1 _06157_ (.A1(_01113_),
    .A2(_01117_),
    .B1(_01128_),
    .Y(_01129_));
 sky130_fd_sc_hd__inv_2 _06158_ (.A(net12),
    .Y(_01130_));
 sky130_fd_sc_hd__nand2_1 _06159_ (.A(_01114_),
    .B(_01116_),
    .Y(_01131_));
 sky130_fd_sc_hd__nand2_1 _06160_ (.A(_01117_),
    .B(_01131_),
    .Y(_01132_));
 sky130_fd_sc_hd__or2_1 _06161_ (.A(_01130_),
    .B(_01132_),
    .X(_01133_));
 sky130_fd_sc_hd__inv_2 _06162_ (.A(net10),
    .Y(_01134_));
 sky130_fd_sc_hd__nand2_1 _06163_ (.A(_01130_),
    .B(_01132_),
    .Y(_01135_));
 sky130_fd_sc_hd__nand2_1 _06164_ (.A(_01133_),
    .B(_01135_),
    .Y(_01136_));
 sky130_fd_sc_hd__or2_1 _06165_ (.A(_01134_),
    .B(_01136_),
    .X(_01137_));
 sky130_fd_sc_hd__and3_1 _06166_ (.A(_01128_),
    .B(_01113_),
    .C(_01117_),
    .X(_01138_));
 sky130_fd_sc_hd__or2_1 _06167_ (.A(_01129_),
    .B(_01138_),
    .X(_01139_));
 sky130_fd_sc_hd__a21oi_1 _06168_ (.A1(_01133_),
    .A2(_01137_),
    .B1(_01139_),
    .Y(_01140_));
 sky130_fd_sc_hd__nor2_1 _06169_ (.A(_01129_),
    .B(_01140_),
    .Y(_01141_));
 sky130_fd_sc_hd__xor2_1 _06170_ (.A(_01119_),
    .B(_01126_),
    .X(_01142_));
 sky130_fd_sc_hd__a21oi_1 _06171_ (.A1(_01121_),
    .A2(_01123_),
    .B1(_01142_),
    .Y(_01143_));
 sky130_fd_sc_hd__a2bb2o_1 _06172_ (.A1_N(_01141_),
    .A2_N(_01143_),
    .B1(_01119_),
    .B2(_01126_),
    .X(_01144_));
 sky130_fd_sc_hd__xor2_1 _06173_ (.A(_01141_),
    .B(_01143_),
    .X(_01145_));
 sky130_fd_sc_hd__nand2_1 _06174_ (.A(_01134_),
    .B(_01136_),
    .Y(_01146_));
 sky130_fd_sc_hd__nand2_1 _06175_ (.A(_01137_),
    .B(_01146_),
    .Y(_01147_));
 sky130_fd_sc_hd__and3_1 _06176_ (.A(_01139_),
    .B(_01133_),
    .C(_01137_),
    .X(_01148_));
 sky130_fd_sc_hd__or2_1 _06177_ (.A(_01140_),
    .B(_01148_),
    .X(_01149_));
 sky130_fd_sc_hd__or4bb_4 _06178_ (.A(_01144_),
    .B(_01145_),
    .C_N(_01147_),
    .D_N(_01149_),
    .X(_01150_));
 sky130_fd_sc_hd__inv_2 _06179_ (.A(net765),
    .Y(_01151_));
 sky130_fd_sc_hd__and4_1 _06180_ (.A(\sig_norm.i[1] ),
    .B(\sig_norm.i[0] ),
    .C(\sig_norm.i[3] ),
    .D(_01151_),
    .X(_01152_));
 sky130_fd_sc_hd__and3_1 _06181_ (.A(\sig_norm.busy ),
    .B(_01152_),
    .C(_01098_),
    .X(_01153_));
 sky130_fd_sc_hd__clkbuf_4 _06182_ (.A(_01153_),
    .X(_01154_));
 sky130_fd_sc_hd__o21bai_1 _06183_ (.A1(_01099_),
    .A2(_01150_),
    .B1_N(_01154_),
    .Y(_00025_));
 sky130_fd_sc_hd__or3_4 _06184_ (.A(_01094_),
    .B(_01095_),
    .C(_01096_),
    .X(_01155_));
 sky130_fd_sc_hd__and3b_1 _06185_ (.A_N(_01152_),
    .B(_01097_),
    .C(\sig_norm.busy ),
    .X(_01156_));
 sky130_fd_sc_hd__a21oi_4 _06186_ (.A1(_01155_),
    .A2(_01150_),
    .B1(_01156_),
    .Y(_01157_));
 sky130_fd_sc_hd__inv_2 _06187_ (.A(_01157_),
    .Y(_01158_));
 sky130_fd_sc_hd__clkbuf_4 _06188_ (.A(_01158_),
    .X(_00024_));
 sky130_fd_sc_hd__inv_2 _06189_ (.A(net361),
    .Y(\PWM.next_counter[0] ));
 sky130_fd_sc_hd__xor2_1 _06190_ (.A(net642),
    .B(net361),
    .X(\PWM.next_counter[1] ));
 sky130_fd_sc_hd__and3_1 _06191_ (.A(\PWM.counter[1] ),
    .B(\PWM.counter[0] ),
    .C(\PWM.counter[2] ),
    .X(_01159_));
 sky130_fd_sc_hd__a21oi_1 _06192_ (.A1(net642),
    .A2(\PWM.counter[0] ),
    .B1(net831),
    .Y(_01160_));
 sky130_fd_sc_hd__nor2_1 _06193_ (.A(_01159_),
    .B(net832),
    .Y(\PWM.next_counter[2] ));
 sky130_fd_sc_hd__and2_1 _06194_ (.A(\PWM.counter[3] ),
    .B(_01159_),
    .X(_01161_));
 sky130_fd_sc_hd__nor2_1 _06195_ (.A(net996),
    .B(_01159_),
    .Y(_01162_));
 sky130_fd_sc_hd__nor2_1 _06196_ (.A(_01161_),
    .B(_01162_),
    .Y(\PWM.next_counter[3] ));
 sky130_fd_sc_hd__inv_2 _06197_ (.A(net1307),
    .Y(_01163_));
 sky130_fd_sc_hd__xnor2_1 _06198_ (.A(_01163_),
    .B(_01161_),
    .Y(\PWM.next_counter[4] ));
 sky130_fd_sc_hd__and3_1 _06199_ (.A(\PWM.counter[5] ),
    .B(\PWM.counter[4] ),
    .C(_01161_),
    .X(_01164_));
 sky130_fd_sc_hd__a21oi_1 _06200_ (.A1(\PWM.counter[4] ),
    .A2(_01161_),
    .B1(net810),
    .Y(_01165_));
 sky130_fd_sc_hd__nor2_1 _06201_ (.A(_01164_),
    .B(net811),
    .Y(\PWM.next_counter[5] ));
 sky130_fd_sc_hd__nand2_1 _06202_ (.A(\PWM.counter[6] ),
    .B(_01164_),
    .Y(_01166_));
 sky130_fd_sc_hd__or2_1 _06203_ (.A(\PWM.counter[6] ),
    .B(_01164_),
    .X(_01167_));
 sky130_fd_sc_hd__and2_1 _06204_ (.A(_01166_),
    .B(_01167_),
    .X(_01168_));
 sky130_fd_sc_hd__clkbuf_1 _06205_ (.A(_01168_),
    .X(\PWM.next_counter[6] ));
 sky130_fd_sc_hd__xnor2_1 _06206_ (.A(net399),
    .B(_01166_),
    .Y(\PWM.next_counter[7] ));
 sky130_fd_sc_hd__inv_2 _06207_ (.A(\genblk1[0].osc.clkdiv_C.cnt[10] ),
    .Y(_01169_));
 sky130_fd_sc_hd__or3b_1 _06208_ (.A(\freq_div.state[1] ),
    .B(\freq_div.state[2] ),
    .C_N(\freq_div.state[0] ),
    .X(_01170_));
 sky130_fd_sc_hd__buf_4 _06209_ (.A(_01170_),
    .X(_01171_));
 sky130_fd_sc_hd__clkbuf_8 _06210_ (.A(_01171_),
    .X(_01172_));
 sky130_fd_sc_hd__clkbuf_4 _06211_ (.A(\freq_div.state[0] ),
    .X(_01173_));
 sky130_fd_sc_hd__clkbuf_8 _06212_ (.A(_01173_),
    .X(_01174_));
 sky130_fd_sc_hd__buf_4 _06213_ (.A(\freq_div.state[1] ),
    .X(_01175_));
 sky130_fd_sc_hd__buf_4 _06214_ (.A(\freq_div.state[2] ),
    .X(_01176_));
 sky130_fd_sc_hd__xnor2_4 _06215_ (.A(_01175_),
    .B(_01176_),
    .Y(_01177_));
 sky130_fd_sc_hd__buf_4 _06216_ (.A(\freq_div.state[1] ),
    .X(_01178_));
 sky130_fd_sc_hd__nor2_4 _06217_ (.A(_01178_),
    .B(_01176_),
    .Y(_01179_));
 sky130_fd_sc_hd__a21o_2 _06218_ (.A1(_01174_),
    .A2(_01177_),
    .B1(_01179_),
    .X(_01180_));
 sky130_fd_sc_hd__buf_6 _06219_ (.A(_01174_),
    .X(_01181_));
 sky130_fd_sc_hd__clkbuf_8 _06220_ (.A(_01177_),
    .X(_01182_));
 sky130_fd_sc_hd__nor2_8 _06221_ (.A(_01181_),
    .B(_01182_),
    .Y(_01183_));
 sky130_fd_sc_hd__a21oi_4 _06222_ (.A1(_01172_),
    .A2(_01180_),
    .B1(_01183_),
    .Y(_01184_));
 sky130_fd_sc_hd__inv_2 _06223_ (.A(_01184_),
    .Y(_01185_));
 sky130_fd_sc_hd__clkbuf_4 _06224_ (.A(_01179_),
    .X(_01186_));
 sky130_fd_sc_hd__buf_4 _06225_ (.A(_01176_),
    .X(_01187_));
 sky130_fd_sc_hd__buf_4 _06226_ (.A(_01178_),
    .X(_01188_));
 sky130_fd_sc_hd__a21boi_4 _06227_ (.A1(_01174_),
    .A2(_01187_),
    .B1_N(_01188_),
    .Y(_01189_));
 sky130_fd_sc_hd__nor2_4 _06228_ (.A(_01186_),
    .B(_01189_),
    .Y(_01190_));
 sky130_fd_sc_hd__buf_4 _06229_ (.A(\freq_div.state[2] ),
    .X(_01191_));
 sky130_fd_sc_hd__nand2_4 _06230_ (.A(_01175_),
    .B(_01191_),
    .Y(_01192_));
 sky130_fd_sc_hd__nand2_2 _06231_ (.A(_01181_),
    .B(_01192_),
    .Y(_01193_));
 sky130_fd_sc_hd__buf_2 _06232_ (.A(\freq_div.state[0] ),
    .X(_01194_));
 sky130_fd_sc_hd__nor3_1 _06233_ (.A(_01194_),
    .B(_01175_),
    .C(_01191_),
    .Y(_01195_));
 sky130_fd_sc_hd__clkbuf_8 _06234_ (.A(_01195_),
    .X(_01196_));
 sky130_fd_sc_hd__buf_4 _06235_ (.A(_01196_),
    .X(_01197_));
 sky130_fd_sc_hd__xor2_1 _06236_ (.A(_01174_),
    .B(\genblk1[0].osc.clkdiv_C.cnt[6] ),
    .X(_01198_));
 sky130_fd_sc_hd__a21o_1 _06237_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[17] ),
    .A2(_01197_),
    .B1(_01198_),
    .X(_01199_));
 sky130_fd_sc_hd__buf_6 _06238_ (.A(_01181_),
    .X(_01200_));
 sky130_fd_sc_hd__buf_4 _06239_ (.A(_01200_),
    .X(_01201_));
 sky130_fd_sc_hd__a21o_1 _06240_ (.A1(_01201_),
    .A2(\genblk1[0].osc.clkdiv_C.cnt[7] ),
    .B1(\genblk1[0].osc.clkdiv_C.cnt[8] ),
    .X(_01202_));
 sky130_fd_sc_hd__o21ai_1 _06241_ (.A1(_01201_),
    .A2(\genblk1[0].osc.clkdiv_C.cnt[7] ),
    .B1(\genblk1[0].osc.clkdiv_C.cnt[8] ),
    .Y(_01203_));
 sky130_fd_sc_hd__o2111a_1 _06242_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[9] ),
    .A2(_01193_),
    .B1(_01199_),
    .C1(_01202_),
    .D1(_01203_),
    .X(_01204_));
 sky130_fd_sc_hd__o21ai_1 _06243_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[17] ),
    .A2(_01197_),
    .B1(_01198_),
    .Y(_01205_));
 sky130_fd_sc_hd__o211a_1 _06244_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[2] ),
    .A2(_01190_),
    .B1(_01204_),
    .C1(_01205_),
    .X(_01206_));
 sky130_fd_sc_hd__or3b_1 _06245_ (.A(\freq_div.state[0] ),
    .B(\freq_div.state[2] ),
    .C_N(\freq_div.state[1] ),
    .X(_01207_));
 sky130_fd_sc_hd__buf_4 _06246_ (.A(_01207_),
    .X(_01208_));
 sky130_fd_sc_hd__buf_4 _06247_ (.A(_01208_),
    .X(_01209_));
 sky130_fd_sc_hd__clkbuf_8 _06248_ (.A(_01209_),
    .X(_01210_));
 sky130_fd_sc_hd__buf_4 _06249_ (.A(_01182_),
    .X(_01211_));
 sky130_fd_sc_hd__o22ai_1 _06250_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[0] ),
    .A2(_01211_),
    .B1(_01210_),
    .B2(\genblk1[0].osc.clkdiv_C.cnt[15] ),
    .Y(_01212_));
 sky130_fd_sc_hd__nand2_2 _06251_ (.A(_01174_),
    .B(_01187_),
    .Y(_01213_));
 sky130_fd_sc_hd__nand2b_4 _06252_ (.A_N(_01187_),
    .B(_01188_),
    .Y(_01214_));
 sky130_fd_sc_hd__nand2_2 _06253_ (.A(_01213_),
    .B(_01214_),
    .Y(_01215_));
 sky130_fd_sc_hd__a2bb2o_1 _06254_ (.A1_N(\genblk1[0].osc.clkdiv_C.cnt[4] ),
    .A2_N(_01215_),
    .B1(_01193_),
    .B2(\genblk1[0].osc.clkdiv_C.cnt[9] ),
    .X(_01216_));
 sky130_fd_sc_hd__a221o_1 _06255_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[0] ),
    .A2(_01211_),
    .B1(_01215_),
    .B2(\genblk1[0].osc.clkdiv_C.cnt[4] ),
    .C1(_01216_),
    .X(_01217_));
 sky130_fd_sc_hd__a211oi_1 _06256_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[15] ),
    .A2(_01210_),
    .B1(_01212_),
    .C1(_01217_),
    .Y(_01218_));
 sky130_fd_sc_hd__o211a_1 _06257_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[10] ),
    .A2(_01184_),
    .B1(_01206_),
    .C1(_01218_),
    .X(_01219_));
 sky130_fd_sc_hd__xor2_4 _06258_ (.A(\freq_div.state[1] ),
    .B(_01176_),
    .X(_01220_));
 sky130_fd_sc_hd__nand2b_4 _06259_ (.A_N(_01194_),
    .B(_01175_),
    .Y(_01221_));
 sky130_fd_sc_hd__and3b_1 _06260_ (.A_N(\freq_div.state[0] ),
    .B(\freq_div.state[1] ),
    .C(\freq_div.state[2] ),
    .X(_01222_));
 sky130_fd_sc_hd__buf_4 _06261_ (.A(_01222_),
    .X(_01223_));
 sky130_fd_sc_hd__a21oi_4 _06262_ (.A1(_01220_),
    .A2(_01221_),
    .B1(_01223_),
    .Y(_01224_));
 sky130_fd_sc_hd__nor2b_2 _06263_ (.A(_01175_),
    .B_N(_01194_),
    .Y(_01225_));
 sky130_fd_sc_hd__buf_6 _06264_ (.A(_01225_),
    .X(_01226_));
 sky130_fd_sc_hd__nor2_8 _06265_ (.A(_01224_),
    .B(_01226_),
    .Y(_01227_));
 sky130_fd_sc_hd__inv_2 _06266_ (.A(_01194_),
    .Y(_01228_));
 sky130_fd_sc_hd__buf_6 _06267_ (.A(_01228_),
    .X(_01229_));
 sky130_fd_sc_hd__clkbuf_8 _06268_ (.A(_01220_),
    .X(_01230_));
 sky130_fd_sc_hd__nor2_4 _06269_ (.A(_01229_),
    .B(_01230_),
    .Y(_01231_));
 sky130_fd_sc_hd__and2_1 _06270_ (.A(\freq_div.state[0] ),
    .B(\freq_div.state[1] ),
    .X(_01232_));
 sky130_fd_sc_hd__clkbuf_4 _06271_ (.A(_01232_),
    .X(_01233_));
 sky130_fd_sc_hd__a21o_2 _06272_ (.A1(_01229_),
    .A2(_01230_),
    .B1(_01233_),
    .X(_01234_));
 sky130_fd_sc_hd__nor2_4 _06273_ (.A(_01231_),
    .B(_01234_),
    .Y(_01235_));
 sky130_fd_sc_hd__o22ai_1 _06274_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[3] ),
    .A2(_01227_),
    .B1(_01235_),
    .B2(\genblk1[0].osc.clkdiv_C.cnt[1] ),
    .Y(_01236_));
 sky130_fd_sc_hd__nor3b_1 _06275_ (.A(_01178_),
    .B(_01176_),
    .C_N(_01194_),
    .Y(_01237_));
 sky130_fd_sc_hd__clkbuf_8 _06276_ (.A(_01237_),
    .X(_01238_));
 sky130_fd_sc_hd__nor3b_2 _06277_ (.A(_01173_),
    .B(_01188_),
    .C_N(_01191_),
    .Y(_01239_));
 sky130_fd_sc_hd__nor2_8 _06278_ (.A(_01238_),
    .B(_01239_),
    .Y(_01240_));
 sky130_fd_sc_hd__buf_4 _06279_ (.A(_01237_),
    .X(_01241_));
 sky130_fd_sc_hd__clkbuf_8 _06280_ (.A(_01241_),
    .X(_01242_));
 sky130_fd_sc_hd__or2_1 _06281_ (.A(\genblk1[0].osc.clkdiv_C.cnt[16] ),
    .B(_01242_),
    .X(_01243_));
 sky130_fd_sc_hd__nand2_1 _06282_ (.A(\genblk1[0].osc.clkdiv_C.cnt[16] ),
    .B(_01242_),
    .Y(_01244_));
 sky130_fd_sc_hd__or2_2 _06283_ (.A(_01173_),
    .B(_01187_),
    .X(_01245_));
 sky130_fd_sc_hd__buf_4 _06284_ (.A(_01245_),
    .X(_01246_));
 sky130_fd_sc_hd__and2_1 _06285_ (.A(_01173_),
    .B(_01191_),
    .X(_01247_));
 sky130_fd_sc_hd__buf_4 _06286_ (.A(_01247_),
    .X(_01248_));
 sky130_fd_sc_hd__nor2_4 _06287_ (.A(_01173_),
    .B(_01188_),
    .Y(_01249_));
 sky130_fd_sc_hd__nor2_2 _06288_ (.A(_01248_),
    .B(_01249_),
    .Y(_01250_));
 sky130_fd_sc_hd__nand2_1 _06289_ (.A(_01246_),
    .B(_01250_),
    .Y(_01251_));
 sky130_fd_sc_hd__xnor2_1 _06290_ (.A(\genblk1[0].osc.clkdiv_C.cnt[11] ),
    .B(_01251_),
    .Y(_01252_));
 sky130_fd_sc_hd__a221o_1 _06291_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[13] ),
    .A2(_01240_),
    .B1(_01243_),
    .B2(_01244_),
    .C1(_01252_),
    .X(_01253_));
 sky130_fd_sc_hd__and3b_2 _06292_ (.A_N(_01176_),
    .B(_01178_),
    .C(_01194_),
    .X(_01254_));
 sky130_fd_sc_hd__nor2_1 _06293_ (.A(_01196_),
    .B(_01254_),
    .Y(_01255_));
 sky130_fd_sc_hd__buf_4 _06294_ (.A(_01255_),
    .X(_01256_));
 sky130_fd_sc_hd__o21ba_1 _06295_ (.A1(_01188_),
    .A2(_01187_),
    .B1_N(_01173_),
    .X(_01257_));
 sky130_fd_sc_hd__or2_2 _06296_ (.A(_01238_),
    .B(_01257_),
    .X(_01258_));
 sky130_fd_sc_hd__o2bb2a_1 _06297_ (.A1_N(\genblk1[0].osc.clkdiv_C.cnt[2] ),
    .A2_N(_01190_),
    .B1(_01258_),
    .B2(\genblk1[0].osc.clkdiv_C.cnt[5] ),
    .X(_01259_));
 sky130_fd_sc_hd__o221ai_1 _06298_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[14] ),
    .A2(_01256_),
    .B1(_01240_),
    .B2(\genblk1[0].osc.clkdiv_C.cnt[13] ),
    .C1(_01259_),
    .Y(_01260_));
 sky130_fd_sc_hd__mux2_1 _06299_ (.A0(_01176_),
    .A1(_01178_),
    .S(_01194_),
    .X(_01261_));
 sky130_fd_sc_hd__buf_4 _06300_ (.A(_01261_),
    .X(_01262_));
 sky130_fd_sc_hd__or2_4 _06301_ (.A(_01238_),
    .B(_01262_),
    .X(_01263_));
 sky130_fd_sc_hd__xnor2_1 _06302_ (.A(\genblk1[0].osc.clkdiv_C.cnt[12] ),
    .B(_01263_),
    .Y(_01264_));
 sky130_fd_sc_hd__a221o_1 _06303_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[14] ),
    .A2(_01256_),
    .B1(_01258_),
    .B2(\genblk1[0].osc.clkdiv_C.cnt[5] ),
    .C1(_01264_),
    .X(_01265_));
 sky130_fd_sc_hd__a2111o_1 _06304_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[1] ),
    .A2(_01235_),
    .B1(_01253_),
    .C1(_01260_),
    .D1(_01265_),
    .X(_01266_));
 sky130_fd_sc_hd__a211oi_1 _06305_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[3] ),
    .A2(_01227_),
    .B1(_01236_),
    .C1(_01266_),
    .Y(_01267_));
 sky130_fd_sc_hd__o211a_2 _06306_ (.A1(_01169_),
    .A2(_01185_),
    .B1(_01219_),
    .C1(_01267_),
    .X(_01268_));
 sky130_fd_sc_hd__clkbuf_4 _06307_ (.A(_01268_),
    .X(_01269_));
 sky130_fd_sc_hd__nor2_1 _06308_ (.A(net1089),
    .B(_01269_),
    .Y(\genblk1[0].osc.clkdiv_C.next_cnt[0] ));
 sky130_fd_sc_hd__inv_2 _06309_ (.A(_01268_),
    .Y(_01270_));
 sky130_fd_sc_hd__or2_1 _06310_ (.A(\genblk1[0].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[0].osc.clkdiv_C.cnt[0] ),
    .X(_01271_));
 sky130_fd_sc_hd__nand2_1 _06311_ (.A(\genblk1[0].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[0].osc.clkdiv_C.cnt[0] ),
    .Y(_01272_));
 sky130_fd_sc_hd__and3_1 _06312_ (.A(_01270_),
    .B(_01271_),
    .C(_01272_),
    .X(_01273_));
 sky130_fd_sc_hd__clkbuf_1 _06313_ (.A(_01273_),
    .X(\genblk1[0].osc.clkdiv_C.next_cnt[1] ));
 sky130_fd_sc_hd__and3_1 _06314_ (.A(\genblk1[0].osc.clkdiv_C.cnt[2] ),
    .B(\genblk1[0].osc.clkdiv_C.cnt[1] ),
    .C(\genblk1[0].osc.clkdiv_C.cnt[0] ),
    .X(_01274_));
 sky130_fd_sc_hd__a21oi_1 _06315_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[1] ),
    .A2(\genblk1[0].osc.clkdiv_C.cnt[0] ),
    .B1(\genblk1[0].osc.clkdiv_C.cnt[2] ),
    .Y(_01275_));
 sky130_fd_sc_hd__nor3_1 _06316_ (.A(_01269_),
    .B(_01274_),
    .C(_01275_),
    .Y(\genblk1[0].osc.clkdiv_C.next_cnt[2] ));
 sky130_fd_sc_hd__and2_1 _06317_ (.A(\genblk1[0].osc.clkdiv_C.cnt[3] ),
    .B(_01274_),
    .X(_01276_));
 sky130_fd_sc_hd__nor2_1 _06318_ (.A(\genblk1[0].osc.clkdiv_C.cnt[3] ),
    .B(_01274_),
    .Y(_01277_));
 sky130_fd_sc_hd__nor3_1 _06319_ (.A(_01269_),
    .B(_01276_),
    .C(_01277_),
    .Y(\genblk1[0].osc.clkdiv_C.next_cnt[3] ));
 sky130_fd_sc_hd__o21ai_1 _06320_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[4] ),
    .A2(_01276_),
    .B1(_01270_),
    .Y(_01278_));
 sky130_fd_sc_hd__a21oi_1 _06321_ (.A1(net1133),
    .A2(_01276_),
    .B1(_01278_),
    .Y(\genblk1[0].osc.clkdiv_C.next_cnt[4] ));
 sky130_fd_sc_hd__and3_1 _06322_ (.A(\genblk1[0].osc.clkdiv_C.cnt[5] ),
    .B(\genblk1[0].osc.clkdiv_C.cnt[4] ),
    .C(_01276_),
    .X(_01279_));
 sky130_fd_sc_hd__a21oi_1 _06323_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[4] ),
    .A2(_01276_),
    .B1(\genblk1[0].osc.clkdiv_C.cnt[5] ),
    .Y(_01280_));
 sky130_fd_sc_hd__nor3_1 _06324_ (.A(_01269_),
    .B(_01279_),
    .C(_01280_),
    .Y(\genblk1[0].osc.clkdiv_C.next_cnt[5] ));
 sky130_fd_sc_hd__and2_1 _06325_ (.A(\genblk1[0].osc.clkdiv_C.cnt[6] ),
    .B(_01279_),
    .X(_01281_));
 sky130_fd_sc_hd__nor2_1 _06326_ (.A(\genblk1[0].osc.clkdiv_C.cnt[6] ),
    .B(_01279_),
    .Y(_01282_));
 sky130_fd_sc_hd__nor3_1 _06327_ (.A(_01269_),
    .B(_01281_),
    .C(_01282_),
    .Y(\genblk1[0].osc.clkdiv_C.next_cnt[6] ));
 sky130_fd_sc_hd__o21ai_1 _06328_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[7] ),
    .A2(_01281_),
    .B1(_01270_),
    .Y(_01283_));
 sky130_fd_sc_hd__a21oi_1 _06329_ (.A1(net592),
    .A2(_01281_),
    .B1(_01283_),
    .Y(\genblk1[0].osc.clkdiv_C.next_cnt[7] ));
 sky130_fd_sc_hd__and3_1 _06330_ (.A(\genblk1[0].osc.clkdiv_C.cnt[8] ),
    .B(\genblk1[0].osc.clkdiv_C.cnt[7] ),
    .C(_01281_),
    .X(_01284_));
 sky130_fd_sc_hd__a21oi_1 _06331_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[7] ),
    .A2(_01281_),
    .B1(\genblk1[0].osc.clkdiv_C.cnt[8] ),
    .Y(_01285_));
 sky130_fd_sc_hd__nor3_1 _06332_ (.A(_01269_),
    .B(_01284_),
    .C(_01285_),
    .Y(\genblk1[0].osc.clkdiv_C.next_cnt[8] ));
 sky130_fd_sc_hd__and2_1 _06333_ (.A(\genblk1[0].osc.clkdiv_C.cnt[9] ),
    .B(_01284_),
    .X(_01286_));
 sky130_fd_sc_hd__nor2_1 _06334_ (.A(\genblk1[0].osc.clkdiv_C.cnt[9] ),
    .B(_01284_),
    .Y(_01287_));
 sky130_fd_sc_hd__nor3_1 _06335_ (.A(_01269_),
    .B(_01286_),
    .C(_01287_),
    .Y(\genblk1[0].osc.clkdiv_C.next_cnt[9] ));
 sky130_fd_sc_hd__nand2_1 _06336_ (.A(\genblk1[0].osc.clkdiv_C.cnt[10] ),
    .B(_01286_),
    .Y(_01288_));
 sky130_fd_sc_hd__o211a_1 _06337_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[10] ),
    .A2(_01286_),
    .B1(_01288_),
    .C1(_01270_),
    .X(\genblk1[0].osc.clkdiv_C.next_cnt[10] ));
 sky130_fd_sc_hd__a21oi_1 _06338_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[10] ),
    .A2(_01286_),
    .B1(\genblk1[0].osc.clkdiv_C.cnt[11] ),
    .Y(_01289_));
 sky130_fd_sc_hd__and3_1 _06339_ (.A(\genblk1[0].osc.clkdiv_C.cnt[11] ),
    .B(\genblk1[0].osc.clkdiv_C.cnt[10] ),
    .C(_01286_),
    .X(_01290_));
 sky130_fd_sc_hd__nor3_1 _06340_ (.A(_01269_),
    .B(_01289_),
    .C(_01290_),
    .Y(\genblk1[0].osc.clkdiv_C.next_cnt[11] ));
 sky130_fd_sc_hd__and2_1 _06341_ (.A(\genblk1[0].osc.clkdiv_C.cnt[12] ),
    .B(_01290_),
    .X(_01291_));
 sky130_fd_sc_hd__nor2_1 _06342_ (.A(_01268_),
    .B(_01291_),
    .Y(_01292_));
 sky130_fd_sc_hd__o21a_1 _06343_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[12] ),
    .A2(_01290_),
    .B1(_01292_),
    .X(\genblk1[0].osc.clkdiv_C.next_cnt[12] ));
 sky130_fd_sc_hd__a21oi_1 _06344_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[13] ),
    .A2(_01291_),
    .B1(_01269_),
    .Y(_01293_));
 sky130_fd_sc_hd__o21a_1 _06345_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[13] ),
    .A2(_01291_),
    .B1(_01293_),
    .X(\genblk1[0].osc.clkdiv_C.next_cnt[13] ));
 sky130_fd_sc_hd__a21oi_1 _06346_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[13] ),
    .A2(_01291_),
    .B1(\genblk1[0].osc.clkdiv_C.cnt[14] ),
    .Y(_01294_));
 sky130_fd_sc_hd__and3_1 _06347_ (.A(\genblk1[0].osc.clkdiv_C.cnt[14] ),
    .B(\genblk1[0].osc.clkdiv_C.cnt[13] ),
    .C(_01291_),
    .X(_01295_));
 sky130_fd_sc_hd__nor3_1 _06348_ (.A(_01269_),
    .B(_01294_),
    .C(_01295_),
    .Y(\genblk1[0].osc.clkdiv_C.next_cnt[14] ));
 sky130_fd_sc_hd__and2_1 _06349_ (.A(\genblk1[0].osc.clkdiv_C.cnt[15] ),
    .B(_01295_),
    .X(_01296_));
 sky130_fd_sc_hd__nor2_1 _06350_ (.A(_01268_),
    .B(_01296_),
    .Y(_01297_));
 sky130_fd_sc_hd__o21a_1 _06351_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[15] ),
    .A2(_01295_),
    .B1(_01297_),
    .X(\genblk1[0].osc.clkdiv_C.next_cnt[15] ));
 sky130_fd_sc_hd__and3_1 _06352_ (.A(\genblk1[0].osc.clkdiv_C.cnt[16] ),
    .B(\genblk1[0].osc.clkdiv_C.cnt[15] ),
    .C(_01295_),
    .X(_01298_));
 sky130_fd_sc_hd__nor2_1 _06353_ (.A(_01268_),
    .B(_01298_),
    .Y(_01299_));
 sky130_fd_sc_hd__o21a_1 _06354_ (.A1(net1196),
    .A2(_01296_),
    .B1(_01299_),
    .X(\genblk1[0].osc.clkdiv_C.next_cnt[16] ));
 sky130_fd_sc_hd__nand2_1 _06355_ (.A(\genblk1[0].osc.clkdiv_C.cnt[17] ),
    .B(_01298_),
    .Y(_01300_));
 sky130_fd_sc_hd__o211a_1 _06356_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[17] ),
    .A2(_01298_),
    .B1(_01300_),
    .C1(_01270_),
    .X(\genblk1[0].osc.clkdiv_C.next_cnt[17] ));
 sky130_fd_sc_hd__and2b_1 _06357_ (.A_N(\freq_div.state[2] ),
    .B(\freq_div.state[0] ),
    .X(_01301_));
 sky130_fd_sc_hd__buf_6 _06358_ (.A(_01301_),
    .X(_01302_));
 sky130_fd_sc_hd__or3_1 _06359_ (.A(_01179_),
    .B(_01222_),
    .C(_01302_),
    .X(_01303_));
 sky130_fd_sc_hd__clkbuf_4 _06360_ (.A(_01303_),
    .X(_01304_));
 sky130_fd_sc_hd__or2_2 _06361_ (.A(_01223_),
    .B(_01226_),
    .X(_01305_));
 sky130_fd_sc_hd__and2_1 _06362_ (.A(\genblk1[1].osc.clkdiv_C.cnt[5] ),
    .B(_01305_),
    .X(_01306_));
 sky130_fd_sc_hd__inv_2 _06363_ (.A(\genblk1[1].osc.clkdiv_C.cnt[6] ),
    .Y(_01307_));
 sky130_fd_sc_hd__inv_4 _06364_ (.A(_01178_),
    .Y(_01308_));
 sky130_fd_sc_hd__clkbuf_4 _06365_ (.A(_01171_),
    .X(_01309_));
 sky130_fd_sc_hd__nand2_1 _06366_ (.A(_01308_),
    .B(_01309_),
    .Y(_01310_));
 sky130_fd_sc_hd__buf_4 _06367_ (.A(_01310_),
    .X(_01311_));
 sky130_fd_sc_hd__and2_2 _06368_ (.A(_01309_),
    .B(_01221_),
    .X(_01312_));
 sky130_fd_sc_hd__nand2_4 _06369_ (.A(_01192_),
    .B(_01208_),
    .Y(_01313_));
 sky130_fd_sc_hd__xnor2_1 _06370_ (.A(\genblk1[1].osc.clkdiv_C.cnt[4] ),
    .B(_01313_),
    .Y(_01314_));
 sky130_fd_sc_hd__a221o_1 _06371_ (.A1(_01307_),
    .A2(_01311_),
    .B1(_01312_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[11] ),
    .C1(_01314_),
    .X(_01315_));
 sky130_fd_sc_hd__nor2_1 _06372_ (.A(\genblk1[1].osc.clkdiv_C.cnt[5] ),
    .B(_01305_),
    .Y(_01316_));
 sky130_fd_sc_hd__xnor2_1 _06373_ (.A(\genblk1[1].osc.clkdiv_C.cnt[2] ),
    .B(_01240_),
    .Y(_01317_));
 sky130_fd_sc_hd__o221a_1 _06374_ (.A1(_01307_),
    .A2(_01311_),
    .B1(_01312_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[11] ),
    .C1(_01317_),
    .X(_01318_));
 sky130_fd_sc_hd__or4b_1 _06375_ (.A(_01306_),
    .B(_01315_),
    .C(_01316_),
    .D_N(_01318_),
    .X(_01319_));
 sky130_fd_sc_hd__xnor2_4 _06376_ (.A(\freq_div.state[0] ),
    .B(_01178_),
    .Y(_01320_));
 sky130_fd_sc_hd__nand2b_4 _06377_ (.A_N(_01188_),
    .B(_01191_),
    .Y(_01321_));
 sky130_fd_sc_hd__and2_1 _06378_ (.A(net37),
    .B(_01321_),
    .X(_01322_));
 sky130_fd_sc_hd__clkbuf_4 _06379_ (.A(_01322_),
    .X(_01323_));
 sky130_fd_sc_hd__and2_1 _06380_ (.A(_01178_),
    .B(_01176_),
    .X(_01324_));
 sky130_fd_sc_hd__clkbuf_4 _06381_ (.A(_01324_),
    .X(_01325_));
 sky130_fd_sc_hd__nand2_4 _06382_ (.A(_01229_),
    .B(_01325_),
    .Y(_01326_));
 sky130_fd_sc_hd__clkbuf_8 _06383_ (.A(_01254_),
    .X(_01327_));
 sky130_fd_sc_hd__nor2_4 _06384_ (.A(_01186_),
    .B(_01327_),
    .Y(_01328_));
 sky130_fd_sc_hd__and2_2 _06385_ (.A(_01326_),
    .B(_01328_),
    .X(_01329_));
 sky130_fd_sc_hd__inv_2 _06386_ (.A(\genblk1[1].osc.clkdiv_C.cnt[0] ),
    .Y(_01330_));
 sky130_fd_sc_hd__a22o_1 _06387_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[3] ),
    .A2(_01323_),
    .B1(_01329_),
    .B2(_01330_),
    .X(_01331_));
 sky130_fd_sc_hd__and2b_1 _06388_ (.A_N(_01194_),
    .B(_01176_),
    .X(_01332_));
 sky130_fd_sc_hd__or3_1 _06389_ (.A(_01179_),
    .B(_01332_),
    .C(_01225_),
    .X(_01333_));
 sky130_fd_sc_hd__clkbuf_4 _06390_ (.A(_01333_),
    .X(_01334_));
 sky130_fd_sc_hd__xnor2_1 _06391_ (.A(\genblk1[1].osc.clkdiv_C.cnt[10] ),
    .B(_01334_),
    .Y(_01335_));
 sky130_fd_sc_hd__clkbuf_8 _06392_ (.A(_01179_),
    .X(_01336_));
 sky130_fd_sc_hd__nor2_4 _06393_ (.A(_01336_),
    .B(_01226_),
    .Y(_01337_));
 sky130_fd_sc_hd__o22ai_1 _06394_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[15] ),
    .A2(_01210_),
    .B1(_01337_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[12] ),
    .Y(_01338_));
 sky130_fd_sc_hd__a22o_1 _06395_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[15] ),
    .A2(_01210_),
    .B1(_01337_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[12] ),
    .X(_01339_));
 sky130_fd_sc_hd__nor2_4 _06396_ (.A(_01238_),
    .B(_01262_),
    .Y(_01340_));
 sky130_fd_sc_hd__inv_2 _06397_ (.A(\genblk1[1].osc.clkdiv_C.cnt[17] ),
    .Y(_01341_));
 sky130_fd_sc_hd__clkbuf_8 _06398_ (.A(_01188_),
    .X(_01342_));
 sky130_fd_sc_hd__or2_1 _06399_ (.A(_01173_),
    .B(_01175_),
    .X(_01343_));
 sky130_fd_sc_hd__clkbuf_8 _06400_ (.A(_01343_),
    .X(_01344_));
 sky130_fd_sc_hd__a22o_1 _06401_ (.A1(_01342_),
    .A2(\genblk1[1].osc.clkdiv_C.cnt[8] ),
    .B1(_01344_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[13] ),
    .X(_01345_));
 sky130_fd_sc_hd__a221o_1 _06402_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[1] ),
    .A2(_01340_),
    .B1(_01197_),
    .B2(_01341_),
    .C1(_01345_),
    .X(_01346_));
 sky130_fd_sc_hd__nor2_1 _06403_ (.A(\genblk1[1].osc.clkdiv_C.cnt[14] ),
    .B(_01327_),
    .Y(_01347_));
 sky130_fd_sc_hd__and2_1 _06404_ (.A(\genblk1[1].osc.clkdiv_C.cnt[14] ),
    .B(_01327_),
    .X(_01348_));
 sky130_fd_sc_hd__buf_4 _06405_ (.A(_01172_),
    .X(_01349_));
 sky130_fd_sc_hd__o21a_1 _06406_ (.A1(_01201_),
    .A2(\genblk1[1].osc.clkdiv_C.cnt[13] ),
    .B1(\genblk1[1].osc.clkdiv_C.cnt[8] ),
    .X(_01350_));
 sky130_fd_sc_hd__o2bb2a_1 _06407_ (.A1_N(\genblk1[1].osc.clkdiv_C.cnt[16] ),
    .A2_N(_01349_),
    .B1(_01350_),
    .B2(_01342_),
    .X(_01351_));
 sky130_fd_sc_hd__o221a_1 _06408_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[3] ),
    .A2(_01323_),
    .B1(_01347_),
    .B2(_01348_),
    .C1(_01351_),
    .X(_01352_));
 sky130_fd_sc_hd__or4b_1 _06409_ (.A(_01338_),
    .B(_01339_),
    .C(_01346_),
    .D_N(_01352_),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_2 _06410_ (.A0(_01178_),
    .A1(_01176_),
    .S(\freq_div.state[0] ),
    .X(_01354_));
 sky130_fd_sc_hd__buf_4 _06411_ (.A(_01354_),
    .X(_01355_));
 sky130_fd_sc_hd__or2_2 _06412_ (.A(_01226_),
    .B(_01355_),
    .X(_01356_));
 sky130_fd_sc_hd__xnor2_1 _06413_ (.A(\genblk1[1].osc.clkdiv_C.cnt[9] ),
    .B(_01356_),
    .Y(_01357_));
 sky130_fd_sc_hd__or2_1 _06414_ (.A(_01178_),
    .B(\freq_div.state[2] ),
    .X(_01358_));
 sky130_fd_sc_hd__buf_4 _06415_ (.A(_01358_),
    .X(_01359_));
 sky130_fd_sc_hd__buf_4 _06416_ (.A(_01359_),
    .X(_01360_));
 sky130_fd_sc_hd__clkbuf_4 _06417_ (.A(_01360_),
    .X(_01361_));
 sky130_fd_sc_hd__buf_4 _06418_ (.A(_01361_),
    .X(_01362_));
 sky130_fd_sc_hd__buf_4 _06419_ (.A(_01362_),
    .X(_01363_));
 sky130_fd_sc_hd__o21a_1 _06420_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[16] ),
    .A2(_01363_),
    .B1(_01341_),
    .X(_01364_));
 sky130_fd_sc_hd__buf_8 _06421_ (.A(_01336_),
    .X(_01365_));
 sky130_fd_sc_hd__nor2_1 _06422_ (.A(_01233_),
    .B(_01249_),
    .Y(_01366_));
 sky130_fd_sc_hd__clkbuf_4 _06423_ (.A(_01366_),
    .X(_01367_));
 sky130_fd_sc_hd__nor2_2 _06424_ (.A(_01365_),
    .B(_01367_),
    .Y(_01368_));
 sky130_fd_sc_hd__o2bb2a_1 _06425_ (.A1_N(\genblk1[1].osc.clkdiv_C.cnt[7] ),
    .A2_N(_01368_),
    .B1(_01340_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[1] ),
    .X(_01369_));
 sky130_fd_sc_hd__o221a_1 _06426_ (.A1(_01197_),
    .A2(_01364_),
    .B1(_01368_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[7] ),
    .C1(_01369_),
    .X(_01370_));
 sky130_fd_sc_hd__or4b_1 _06427_ (.A(_01335_),
    .B(_01353_),
    .C(_01357_),
    .D_N(_01370_),
    .X(_01371_));
 sky130_fd_sc_hd__a2111oi_2 _06428_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[0] ),
    .A2(_01304_),
    .B1(_01319_),
    .C1(_01331_),
    .D1(_01371_),
    .Y(_01372_));
 sky130_fd_sc_hd__clkbuf_4 _06429_ (.A(_01372_),
    .X(_01373_));
 sky130_fd_sc_hd__nor2_1 _06430_ (.A(net718),
    .B(_01373_),
    .Y(\genblk1[1].osc.clkdiv_C.next_cnt[0] ));
 sky130_fd_sc_hd__inv_2 _06431_ (.A(net29),
    .Y(_01374_));
 sky130_fd_sc_hd__or2_1 _06432_ (.A(\genblk1[1].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[1].osc.clkdiv_C.cnt[0] ),
    .X(_01375_));
 sky130_fd_sc_hd__nand2_1 _06433_ (.A(\genblk1[1].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[1].osc.clkdiv_C.cnt[0] ),
    .Y(_01376_));
 sky130_fd_sc_hd__and3_1 _06434_ (.A(_01374_),
    .B(_01375_),
    .C(_01376_),
    .X(_01377_));
 sky130_fd_sc_hd__clkbuf_1 _06435_ (.A(_01377_),
    .X(\genblk1[1].osc.clkdiv_C.next_cnt[1] ));
 sky130_fd_sc_hd__and3_1 _06436_ (.A(\genblk1[1].osc.clkdiv_C.cnt[2] ),
    .B(\genblk1[1].osc.clkdiv_C.cnt[1] ),
    .C(\genblk1[1].osc.clkdiv_C.cnt[0] ),
    .X(_01378_));
 sky130_fd_sc_hd__a21oi_1 _06437_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[1] ),
    .A2(\genblk1[1].osc.clkdiv_C.cnt[0] ),
    .B1(\genblk1[1].osc.clkdiv_C.cnt[2] ),
    .Y(_01379_));
 sky130_fd_sc_hd__nor3_1 _06438_ (.A(_01373_),
    .B(_01378_),
    .C(_01379_),
    .Y(\genblk1[1].osc.clkdiv_C.next_cnt[2] ));
 sky130_fd_sc_hd__and2_1 _06439_ (.A(\genblk1[1].osc.clkdiv_C.cnt[3] ),
    .B(_01378_),
    .X(_01380_));
 sky130_fd_sc_hd__nor2_1 _06440_ (.A(\genblk1[1].osc.clkdiv_C.cnt[3] ),
    .B(_01378_),
    .Y(_01381_));
 sky130_fd_sc_hd__nor3_1 _06441_ (.A(_01373_),
    .B(_01380_),
    .C(_01381_),
    .Y(\genblk1[1].osc.clkdiv_C.next_cnt[3] ));
 sky130_fd_sc_hd__nand2_1 _06442_ (.A(\genblk1[1].osc.clkdiv_C.cnt[4] ),
    .B(_01380_),
    .Y(_01382_));
 sky130_fd_sc_hd__or2_1 _06443_ (.A(\genblk1[1].osc.clkdiv_C.cnt[4] ),
    .B(_01380_),
    .X(_01383_));
 sky130_fd_sc_hd__and3_1 _06444_ (.A(_01374_),
    .B(_01382_),
    .C(_01383_),
    .X(_01384_));
 sky130_fd_sc_hd__clkbuf_1 _06445_ (.A(_01384_),
    .X(\genblk1[1].osc.clkdiv_C.next_cnt[4] ));
 sky130_fd_sc_hd__and3_1 _06446_ (.A(\genblk1[1].osc.clkdiv_C.cnt[5] ),
    .B(\genblk1[1].osc.clkdiv_C.cnt[4] ),
    .C(_01380_),
    .X(_01385_));
 sky130_fd_sc_hd__a21oi_1 _06447_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[4] ),
    .A2(_01380_),
    .B1(\genblk1[1].osc.clkdiv_C.cnt[5] ),
    .Y(_01386_));
 sky130_fd_sc_hd__nor3_1 _06448_ (.A(_01373_),
    .B(_01385_),
    .C(_01386_),
    .Y(\genblk1[1].osc.clkdiv_C.next_cnt[5] ));
 sky130_fd_sc_hd__and2_1 _06449_ (.A(\genblk1[1].osc.clkdiv_C.cnt[6] ),
    .B(_01385_),
    .X(_01387_));
 sky130_fd_sc_hd__nor2_1 _06450_ (.A(\genblk1[1].osc.clkdiv_C.cnt[6] ),
    .B(_01385_),
    .Y(_01388_));
 sky130_fd_sc_hd__nor3_1 _06451_ (.A(_01373_),
    .B(_01387_),
    .C(_01388_),
    .Y(\genblk1[1].osc.clkdiv_C.next_cnt[6] ));
 sky130_fd_sc_hd__nand2_1 _06452_ (.A(\genblk1[1].osc.clkdiv_C.cnt[7] ),
    .B(_01387_),
    .Y(_01389_));
 sky130_fd_sc_hd__or2_1 _06453_ (.A(\genblk1[1].osc.clkdiv_C.cnt[7] ),
    .B(_01387_),
    .X(_01390_));
 sky130_fd_sc_hd__and3_1 _06454_ (.A(_01374_),
    .B(_01389_),
    .C(_01390_),
    .X(_01391_));
 sky130_fd_sc_hd__clkbuf_1 _06455_ (.A(_01391_),
    .X(\genblk1[1].osc.clkdiv_C.next_cnt[7] ));
 sky130_fd_sc_hd__and3_1 _06456_ (.A(\genblk1[1].osc.clkdiv_C.cnt[8] ),
    .B(\genblk1[1].osc.clkdiv_C.cnt[7] ),
    .C(_01387_),
    .X(_01392_));
 sky130_fd_sc_hd__a21oi_1 _06457_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[7] ),
    .A2(_01387_),
    .B1(\genblk1[1].osc.clkdiv_C.cnt[8] ),
    .Y(_01393_));
 sky130_fd_sc_hd__nor3_1 _06458_ (.A(_01373_),
    .B(_01392_),
    .C(_01393_),
    .Y(\genblk1[1].osc.clkdiv_C.next_cnt[8] ));
 sky130_fd_sc_hd__and2_1 _06459_ (.A(\genblk1[1].osc.clkdiv_C.cnt[9] ),
    .B(_01392_),
    .X(_01394_));
 sky130_fd_sc_hd__nor2_1 _06460_ (.A(\genblk1[1].osc.clkdiv_C.cnt[9] ),
    .B(_01392_),
    .Y(_01395_));
 sky130_fd_sc_hd__nor3_1 _06461_ (.A(_01373_),
    .B(_01394_),
    .C(_01395_),
    .Y(\genblk1[1].osc.clkdiv_C.next_cnt[9] ));
 sky130_fd_sc_hd__nand2_1 _06462_ (.A(\genblk1[1].osc.clkdiv_C.cnt[10] ),
    .B(_01394_),
    .Y(_01396_));
 sky130_fd_sc_hd__o211a_1 _06463_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[10] ),
    .A2(_01394_),
    .B1(_01396_),
    .C1(_01374_),
    .X(\genblk1[1].osc.clkdiv_C.next_cnt[10] ));
 sky130_fd_sc_hd__a21oi_1 _06464_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[10] ),
    .A2(_01394_),
    .B1(\genblk1[1].osc.clkdiv_C.cnt[11] ),
    .Y(_01397_));
 sky130_fd_sc_hd__and3_1 _06465_ (.A(\genblk1[1].osc.clkdiv_C.cnt[11] ),
    .B(\genblk1[1].osc.clkdiv_C.cnt[10] ),
    .C(_01394_),
    .X(_01398_));
 sky130_fd_sc_hd__nor3_1 _06466_ (.A(_01373_),
    .B(_01397_),
    .C(_01398_),
    .Y(\genblk1[1].osc.clkdiv_C.next_cnt[11] ));
 sky130_fd_sc_hd__and2_1 _06467_ (.A(\genblk1[1].osc.clkdiv_C.cnt[12] ),
    .B(_01398_),
    .X(_01399_));
 sky130_fd_sc_hd__nor2_1 _06468_ (.A(_01373_),
    .B(_01399_),
    .Y(_01400_));
 sky130_fd_sc_hd__o21a_1 _06469_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[12] ),
    .A2(_01398_),
    .B1(_01400_),
    .X(\genblk1[1].osc.clkdiv_C.next_cnt[12] ));
 sky130_fd_sc_hd__and3_1 _06470_ (.A(\genblk1[1].osc.clkdiv_C.cnt[13] ),
    .B(\genblk1[1].osc.clkdiv_C.cnt[12] ),
    .C(_01398_),
    .X(_01401_));
 sky130_fd_sc_hd__nor2_1 _06471_ (.A(_01373_),
    .B(_01401_),
    .Y(_01402_));
 sky130_fd_sc_hd__o21a_1 _06472_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[13] ),
    .A2(_01399_),
    .B1(_01402_),
    .X(\genblk1[1].osc.clkdiv_C.next_cnt[13] ));
 sky130_fd_sc_hd__and2_1 _06473_ (.A(\genblk1[1].osc.clkdiv_C.cnt[14] ),
    .B(_01401_),
    .X(_01403_));
 sky130_fd_sc_hd__nor2_1 _06474_ (.A(net29),
    .B(_01403_),
    .Y(_01404_));
 sky130_fd_sc_hd__o21a_1 _06475_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[14] ),
    .A2(_01401_),
    .B1(_01404_),
    .X(\genblk1[1].osc.clkdiv_C.next_cnt[14] ));
 sky130_fd_sc_hd__and3_1 _06476_ (.A(\genblk1[1].osc.clkdiv_C.cnt[15] ),
    .B(\genblk1[1].osc.clkdiv_C.cnt[14] ),
    .C(_01401_),
    .X(_01405_));
 sky130_fd_sc_hd__nor2_1 _06477_ (.A(net29),
    .B(_01405_),
    .Y(_01406_));
 sky130_fd_sc_hd__o21a_1 _06478_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[15] ),
    .A2(_01403_),
    .B1(_01406_),
    .X(\genblk1[1].osc.clkdiv_C.next_cnt[15] ));
 sky130_fd_sc_hd__and2_1 _06479_ (.A(\genblk1[1].osc.clkdiv_C.cnt[16] ),
    .B(_01405_),
    .X(_01407_));
 sky130_fd_sc_hd__nor2_1 _06480_ (.A(net29),
    .B(_01407_),
    .Y(_01408_));
 sky130_fd_sc_hd__o21a_1 _06481_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[16] ),
    .A2(_01405_),
    .B1(_01408_),
    .X(\genblk1[1].osc.clkdiv_C.next_cnt[16] ));
 sky130_fd_sc_hd__nand2_1 _06482_ (.A(\genblk1[1].osc.clkdiv_C.cnt[17] ),
    .B(_01407_),
    .Y(_01409_));
 sky130_fd_sc_hd__o211a_1 _06483_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[17] ),
    .A2(_01407_),
    .B1(_01409_),
    .C1(_01374_),
    .X(\genblk1[1].osc.clkdiv_C.next_cnt[17] ));
 sky130_fd_sc_hd__inv_2 _06484_ (.A(\genblk1[2].osc.clkdiv_C.cnt[3] ),
    .Y(_01410_));
 sky130_fd_sc_hd__or2_2 _06485_ (.A(_01241_),
    .B(_01337_),
    .X(_01411_));
 sky130_fd_sc_hd__inv_2 _06486_ (.A(\genblk1[2].osc.clkdiv_C.cnt[8] ),
    .Y(_01412_));
 sky130_fd_sc_hd__o2bb2a_1 _06487_ (.A1_N(\genblk1[2].osc.clkdiv_C.cnt[12] ),
    .A2_N(_01411_),
    .B1(_01412_),
    .B2(_01183_),
    .X(_01413_));
 sky130_fd_sc_hd__inv_2 _06488_ (.A(\genblk1[2].osc.clkdiv_C.cnt[2] ),
    .Y(_01414_));
 sky130_fd_sc_hd__mux2_1 _06489_ (.A0(\genblk1[2].osc.clkdiv_C.cnt[15] ),
    .A1(_01414_),
    .S(_01210_),
    .X(_01415_));
 sky130_fd_sc_hd__inv_2 _06490_ (.A(\genblk1[2].osc.clkdiv_C.cnt[17] ),
    .Y(_01416_));
 sky130_fd_sc_hd__o21a_1 _06491_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[16] ),
    .A2(_01363_),
    .B1(_01416_),
    .X(_01417_));
 sky130_fd_sc_hd__nand2_2 _06492_ (.A(_01229_),
    .B(_01182_),
    .Y(_01418_));
 sky130_fd_sc_hd__o22a_1 _06493_ (.A1(_01197_),
    .A2(_01417_),
    .B1(_01418_),
    .B2(\genblk1[2].osc.clkdiv_C.cnt[4] ),
    .X(_01419_));
 sky130_fd_sc_hd__nor2_2 _06494_ (.A(_01242_),
    .B(_01223_),
    .Y(_01420_));
 sky130_fd_sc_hd__nor3_1 _06495_ (.A(\genblk1[2].osc.clkdiv_C.cnt[14] ),
    .B(\genblk1[2].osc.clkdiv_C.cnt[1] ),
    .C(_01327_),
    .Y(_01421_));
 sky130_fd_sc_hd__and3_1 _06496_ (.A(\genblk1[2].osc.clkdiv_C.cnt[14] ),
    .B(\genblk1[2].osc.clkdiv_C.cnt[1] ),
    .C(_01327_),
    .X(_01422_));
 sky130_fd_sc_hd__nor3b_4 _06497_ (.A(_01173_),
    .B(_01191_),
    .C_N(_01175_),
    .Y(_01423_));
 sky130_fd_sc_hd__nand2_1 _06498_ (.A(\genblk1[2].osc.clkdiv_C.cnt[2] ),
    .B(net36),
    .Y(_01424_));
 sky130_fd_sc_hd__nor3_1 _06499_ (.A(\genblk1[2].osc.clkdiv_C.cnt[13] ),
    .B(\genblk1[2].osc.clkdiv_C.cnt[0] ),
    .C(net35),
    .Y(_01425_));
 sky130_fd_sc_hd__and3_1 _06500_ (.A(\genblk1[2].osc.clkdiv_C.cnt[13] ),
    .B(\genblk1[2].osc.clkdiv_C.cnt[0] ),
    .C(net35),
    .X(_01426_));
 sky130_fd_sc_hd__o2bb2a_1 _06501_ (.A1_N(\genblk1[2].osc.clkdiv_C.cnt[15] ),
    .A2_N(_01424_),
    .B1(_01425_),
    .B2(_01426_),
    .X(_01427_));
 sky130_fd_sc_hd__o221a_1 _06502_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[11] ),
    .A2(_01420_),
    .B1(_01421_),
    .B2(_01422_),
    .C1(_01427_),
    .X(_01428_));
 sky130_fd_sc_hd__o2111a_1 _06503_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[12] ),
    .A2(_01411_),
    .B1(_01415_),
    .C1(_01419_),
    .D1(_01428_),
    .X(_01429_));
 sky130_fd_sc_hd__clkbuf_4 _06504_ (.A(_01224_),
    .X(_01430_));
 sky130_fd_sc_hd__a21oi_4 _06505_ (.A1(_01362_),
    .A2(_01430_),
    .B1(_01196_),
    .Y(_01431_));
 sky130_fd_sc_hd__buf_8 _06506_ (.A(_01230_),
    .X(_01432_));
 sky130_fd_sc_hd__nand2_2 _06507_ (.A(_01200_),
    .B(_01432_),
    .Y(_01433_));
 sky130_fd_sc_hd__a221o_1 _06508_ (.A1(_01201_),
    .A2(_01410_),
    .B1(_01432_),
    .B2(_01412_),
    .C1(\genblk1[2].osc.clkdiv_C.cnt[7] ),
    .X(_01434_));
 sky130_fd_sc_hd__a221o_1 _06509_ (.A1(_01416_),
    .A2(_01365_),
    .B1(_01326_),
    .B2(\genblk1[2].osc.clkdiv_C.cnt[11] ),
    .C1(\genblk1[2].osc.clkdiv_C.cnt[16] ),
    .X(_01435_));
 sky130_fd_sc_hd__buf_4 _06510_ (.A(_01349_),
    .X(_01436_));
 sky130_fd_sc_hd__clkbuf_8 _06511_ (.A(_01332_),
    .X(_01437_));
 sky130_fd_sc_hd__xor2_1 _06512_ (.A(\genblk1[2].osc.clkdiv_C.cnt[6] ),
    .B(_01437_),
    .X(_01438_));
 sky130_fd_sc_hd__buf_4 _06513_ (.A(_01213_),
    .X(_01439_));
 sky130_fd_sc_hd__inv_2 _06514_ (.A(_01191_),
    .Y(_01440_));
 sky130_fd_sc_hd__buf_6 _06515_ (.A(_01440_),
    .X(_01441_));
 sky130_fd_sc_hd__nand2_4 _06516_ (.A(_01200_),
    .B(_01441_),
    .Y(_01442_));
 sky130_fd_sc_hd__a2bb2o_1 _06517_ (.A1_N(\genblk1[2].osc.clkdiv_C.cnt[5] ),
    .A2_N(_01439_),
    .B1(_01442_),
    .B2(\genblk1[2].osc.clkdiv_C.cnt[9] ),
    .X(_01443_));
 sky130_fd_sc_hd__a2bb2o_1 _06518_ (.A1_N(\genblk1[2].osc.clkdiv_C.cnt[9] ),
    .A2_N(_01442_),
    .B1(_01439_),
    .B2(\genblk1[2].osc.clkdiv_C.cnt[5] ),
    .X(_01444_));
 sky130_fd_sc_hd__a2bb2o_1 _06519_ (.A1_N(\genblk1[2].osc.clkdiv_C.cnt[7] ),
    .A2_N(_01433_),
    .B1(_01418_),
    .B2(\genblk1[2].osc.clkdiv_C.cnt[4] ),
    .X(_01445_));
 sky130_fd_sc_hd__or4_1 _06520_ (.A(_01438_),
    .B(_01443_),
    .C(_01444_),
    .D(_01445_),
    .X(_01446_));
 sky130_fd_sc_hd__a221o_1 _06521_ (.A1(_01433_),
    .A2(_01434_),
    .B1(_01435_),
    .B2(_01436_),
    .C1(_01446_),
    .X(_01447_));
 sky130_fd_sc_hd__o21bai_1 _06522_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[10] ),
    .A2(_01431_),
    .B1_N(_01447_),
    .Y(_01448_));
 sky130_fd_sc_hd__a21oi_1 _06523_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[10] ),
    .A2(_01431_),
    .B1(_01448_),
    .Y(_01449_));
 sky130_fd_sc_hd__o2111a_1 _06524_ (.A1(_01410_),
    .A2(_01231_),
    .B1(_01413_),
    .C1(_01429_),
    .D1(_01449_),
    .X(_01450_));
 sky130_fd_sc_hd__buf_2 _06525_ (.A(_01450_),
    .X(_01451_));
 sky130_fd_sc_hd__clkbuf_4 _06526_ (.A(_01451_),
    .X(_01452_));
 sky130_fd_sc_hd__nor2_1 _06527_ (.A(net1051),
    .B(_01452_),
    .Y(\genblk1[2].osc.clkdiv_C.next_cnt[0] ));
 sky130_fd_sc_hd__xnor2_1 _06528_ (.A(\genblk1[2].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[2].osc.clkdiv_C.cnt[0] ),
    .Y(_01453_));
 sky130_fd_sc_hd__nor2_1 _06529_ (.A(_01452_),
    .B(_01453_),
    .Y(\genblk1[2].osc.clkdiv_C.next_cnt[1] ));
 sky130_fd_sc_hd__and3_1 _06530_ (.A(\genblk1[2].osc.clkdiv_C.cnt[2] ),
    .B(\genblk1[2].osc.clkdiv_C.cnt[1] ),
    .C(\genblk1[2].osc.clkdiv_C.cnt[0] ),
    .X(_01454_));
 sky130_fd_sc_hd__a21oi_1 _06531_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[1] ),
    .A2(\genblk1[2].osc.clkdiv_C.cnt[0] ),
    .B1(\genblk1[2].osc.clkdiv_C.cnt[2] ),
    .Y(_01455_));
 sky130_fd_sc_hd__nor3_1 _06532_ (.A(_01452_),
    .B(_01454_),
    .C(_01455_),
    .Y(\genblk1[2].osc.clkdiv_C.next_cnt[2] ));
 sky130_fd_sc_hd__and2_1 _06533_ (.A(\genblk1[2].osc.clkdiv_C.cnt[3] ),
    .B(_01454_),
    .X(_01456_));
 sky130_fd_sc_hd__nor2_1 _06534_ (.A(\genblk1[2].osc.clkdiv_C.cnt[3] ),
    .B(_01454_),
    .Y(_01457_));
 sky130_fd_sc_hd__nor3_1 _06535_ (.A(_01452_),
    .B(_01456_),
    .C(_01457_),
    .Y(\genblk1[2].osc.clkdiv_C.next_cnt[3] ));
 sky130_fd_sc_hd__xnor2_1 _06536_ (.A(\genblk1[2].osc.clkdiv_C.cnt[4] ),
    .B(_01456_),
    .Y(_01458_));
 sky130_fd_sc_hd__nor2_1 _06537_ (.A(_01452_),
    .B(_01458_),
    .Y(\genblk1[2].osc.clkdiv_C.next_cnt[4] ));
 sky130_fd_sc_hd__and3_1 _06538_ (.A(\genblk1[2].osc.clkdiv_C.cnt[5] ),
    .B(\genblk1[2].osc.clkdiv_C.cnt[4] ),
    .C(_01456_),
    .X(_01459_));
 sky130_fd_sc_hd__a21oi_1 _06539_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[4] ),
    .A2(_01456_),
    .B1(\genblk1[2].osc.clkdiv_C.cnt[5] ),
    .Y(_01460_));
 sky130_fd_sc_hd__nor3_1 _06540_ (.A(_01452_),
    .B(_01459_),
    .C(_01460_),
    .Y(\genblk1[2].osc.clkdiv_C.next_cnt[5] ));
 sky130_fd_sc_hd__and2_1 _06541_ (.A(\genblk1[2].osc.clkdiv_C.cnt[6] ),
    .B(_01459_),
    .X(_01461_));
 sky130_fd_sc_hd__nor2_1 _06542_ (.A(\genblk1[2].osc.clkdiv_C.cnt[6] ),
    .B(_01459_),
    .Y(_01462_));
 sky130_fd_sc_hd__nor3_1 _06543_ (.A(_01452_),
    .B(_01461_),
    .C(_01462_),
    .Y(\genblk1[2].osc.clkdiv_C.next_cnt[6] ));
 sky130_fd_sc_hd__xnor2_1 _06544_ (.A(\genblk1[2].osc.clkdiv_C.cnt[7] ),
    .B(_01461_),
    .Y(_01463_));
 sky130_fd_sc_hd__nor2_1 _06545_ (.A(_01452_),
    .B(_01463_),
    .Y(\genblk1[2].osc.clkdiv_C.next_cnt[7] ));
 sky130_fd_sc_hd__and3_1 _06546_ (.A(\genblk1[2].osc.clkdiv_C.cnt[8] ),
    .B(\genblk1[2].osc.clkdiv_C.cnt[7] ),
    .C(_01461_),
    .X(_01464_));
 sky130_fd_sc_hd__a21oi_1 _06547_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[7] ),
    .A2(_01461_),
    .B1(\genblk1[2].osc.clkdiv_C.cnt[8] ),
    .Y(_01465_));
 sky130_fd_sc_hd__nor3_1 _06548_ (.A(_01452_),
    .B(_01464_),
    .C(_01465_),
    .Y(\genblk1[2].osc.clkdiv_C.next_cnt[8] ));
 sky130_fd_sc_hd__and2_1 _06549_ (.A(\genblk1[2].osc.clkdiv_C.cnt[9] ),
    .B(_01464_),
    .X(_01466_));
 sky130_fd_sc_hd__nor2_1 _06550_ (.A(\genblk1[2].osc.clkdiv_C.cnt[9] ),
    .B(_01464_),
    .Y(_01467_));
 sky130_fd_sc_hd__nor3_1 _06551_ (.A(_01451_),
    .B(_01466_),
    .C(_01467_),
    .Y(\genblk1[2].osc.clkdiv_C.next_cnt[9] ));
 sky130_fd_sc_hd__and3_1 _06552_ (.A(\genblk1[2].osc.clkdiv_C.cnt[10] ),
    .B(\genblk1[2].osc.clkdiv_C.cnt[9] ),
    .C(_01464_),
    .X(_01468_));
 sky130_fd_sc_hd__nor2_1 _06553_ (.A(_01451_),
    .B(_01468_),
    .Y(_01469_));
 sky130_fd_sc_hd__o21a_1 _06554_ (.A1(net1159),
    .A2(_01466_),
    .B1(_01469_),
    .X(\genblk1[2].osc.clkdiv_C.next_cnt[10] ));
 sky130_fd_sc_hd__and2_1 _06555_ (.A(\genblk1[2].osc.clkdiv_C.cnt[11] ),
    .B(_01468_),
    .X(_01470_));
 sky130_fd_sc_hd__nor2_1 _06556_ (.A(_01451_),
    .B(_01470_),
    .Y(_01471_));
 sky130_fd_sc_hd__o21a_1 _06557_ (.A1(net1213),
    .A2(_01468_),
    .B1(_01471_),
    .X(\genblk1[2].osc.clkdiv_C.next_cnt[11] ));
 sky130_fd_sc_hd__and3_1 _06558_ (.A(\genblk1[2].osc.clkdiv_C.cnt[12] ),
    .B(\genblk1[2].osc.clkdiv_C.cnt[11] ),
    .C(_01468_),
    .X(_01472_));
 sky130_fd_sc_hd__nor2_1 _06559_ (.A(_01451_),
    .B(_01472_),
    .Y(_01473_));
 sky130_fd_sc_hd__o21a_1 _06560_ (.A1(net1256),
    .A2(_01470_),
    .B1(_01473_),
    .X(\genblk1[2].osc.clkdiv_C.next_cnt[12] ));
 sky130_fd_sc_hd__and3_1 _06561_ (.A(\genblk1[2].osc.clkdiv_C.cnt[13] ),
    .B(\genblk1[2].osc.clkdiv_C.cnt[12] ),
    .C(_01470_),
    .X(_01474_));
 sky130_fd_sc_hd__nor2_1 _06562_ (.A(_01451_),
    .B(_01474_),
    .Y(_01475_));
 sky130_fd_sc_hd__o21a_1 _06563_ (.A1(net1166),
    .A2(_01472_),
    .B1(_01475_),
    .X(\genblk1[2].osc.clkdiv_C.next_cnt[13] ));
 sky130_fd_sc_hd__and2_1 _06564_ (.A(\genblk1[2].osc.clkdiv_C.cnt[14] ),
    .B(_01474_),
    .X(_01476_));
 sky130_fd_sc_hd__nor2_1 _06565_ (.A(_01451_),
    .B(_01476_),
    .Y(_01477_));
 sky130_fd_sc_hd__o21a_1 _06566_ (.A1(net1207),
    .A2(_01474_),
    .B1(_01477_),
    .X(\genblk1[2].osc.clkdiv_C.next_cnt[14] ));
 sky130_fd_sc_hd__and3_1 _06567_ (.A(\genblk1[2].osc.clkdiv_C.cnt[15] ),
    .B(\genblk1[2].osc.clkdiv_C.cnt[14] ),
    .C(_01474_),
    .X(_01478_));
 sky130_fd_sc_hd__nor2_1 _06568_ (.A(_01451_),
    .B(_01478_),
    .Y(_01479_));
 sky130_fd_sc_hd__o21a_1 _06569_ (.A1(net1167),
    .A2(_01476_),
    .B1(_01479_),
    .X(\genblk1[2].osc.clkdiv_C.next_cnt[15] ));
 sky130_fd_sc_hd__and2_1 _06570_ (.A(\genblk1[2].osc.clkdiv_C.cnt[16] ),
    .B(_01478_),
    .X(_01480_));
 sky130_fd_sc_hd__nor2_1 _06571_ (.A(_01451_),
    .B(_01480_),
    .Y(_01481_));
 sky130_fd_sc_hd__o21a_1 _06572_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[16] ),
    .A2(_01478_),
    .B1(_01481_),
    .X(\genblk1[2].osc.clkdiv_C.next_cnt[16] ));
 sky130_fd_sc_hd__xnor2_1 _06573_ (.A(\genblk1[2].osc.clkdiv_C.cnt[17] ),
    .B(_01480_),
    .Y(_01482_));
 sky130_fd_sc_hd__nor2_1 _06574_ (.A(_01452_),
    .B(_01482_),
    .Y(\genblk1[2].osc.clkdiv_C.next_cnt[17] ));
 sky130_fd_sc_hd__or2_4 _06575_ (.A(_01196_),
    .B(_01327_),
    .X(_01483_));
 sky130_fd_sc_hd__or2_2 _06576_ (.A(_01182_),
    .B(_01302_),
    .X(_01484_));
 sky130_fd_sc_hd__inv_2 _06577_ (.A(\genblk1[3].osc.clkdiv_C.cnt[8] ),
    .Y(_01485_));
 sky130_fd_sc_hd__inv_2 _06578_ (.A(\genblk1[3].osc.clkdiv_C.cnt[11] ),
    .Y(_01486_));
 sky130_fd_sc_hd__nand2_4 _06579_ (.A(_01172_),
    .B(_01182_),
    .Y(_01487_));
 sky130_fd_sc_hd__a21o_1 _06580_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[12] ),
    .A2(_01344_),
    .B1(\genblk1[3].osc.clkdiv_C.cnt[13] ),
    .X(_01488_));
 sky130_fd_sc_hd__clkbuf_8 _06581_ (.A(_01187_),
    .X(_01489_));
 sky130_fd_sc_hd__buf_8 _06582_ (.A(_01489_),
    .X(_01490_));
 sky130_fd_sc_hd__xnor2_1 _06583_ (.A(\genblk1[3].osc.clkdiv_C.cnt[5] ),
    .B(_01250_),
    .Y(_01491_));
 sky130_fd_sc_hd__a221o_1 _06584_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[10] ),
    .A2(_01231_),
    .B1(_01488_),
    .B2(_01490_),
    .C1(_01491_),
    .X(_01492_));
 sky130_fd_sc_hd__a2bb2o_1 _06585_ (.A1_N(_01490_),
    .A2_N(\genblk1[3].osc.clkdiv_C.cnt[13] ),
    .B1(_01363_),
    .B2(\genblk1[3].osc.clkdiv_C.cnt[15] ),
    .X(_01493_));
 sky130_fd_sc_hd__nor2_4 _06586_ (.A(_01342_),
    .B(_01248_),
    .Y(_01494_));
 sky130_fd_sc_hd__xnor2_1 _06587_ (.A(\genblk1[3].osc.clkdiv_C.cnt[7] ),
    .B(_01494_),
    .Y(_01495_));
 sky130_fd_sc_hd__or2_4 _06588_ (.A(_01437_),
    .B(_01225_),
    .X(_01496_));
 sky130_fd_sc_hd__or2_1 _06589_ (.A(_01191_),
    .B(_01233_),
    .X(_01497_));
 sky130_fd_sc_hd__clkbuf_4 _06590_ (.A(_01497_),
    .X(_01498_));
 sky130_fd_sc_hd__o2bb2a_1 _06591_ (.A1_N(\genblk1[3].osc.clkdiv_C.cnt[2] ),
    .A2_N(_01496_),
    .B1(_01498_),
    .B2(\genblk1[3].osc.clkdiv_C.cnt[14] ),
    .X(_01499_));
 sky130_fd_sc_hd__nor2_2 _06592_ (.A(_01233_),
    .B(_01437_),
    .Y(_01500_));
 sky130_fd_sc_hd__o2bb2a_1 _06593_ (.A1_N(\genblk1[3].osc.clkdiv_C.cnt[14] ),
    .A2_N(_01498_),
    .B1(_01500_),
    .B2(\genblk1[3].osc.clkdiv_C.cnt[6] ),
    .X(_01501_));
 sky130_fd_sc_hd__o2bb2a_1 _06594_ (.A1_N(\genblk1[3].osc.clkdiv_C.cnt[6] ),
    .A2_N(_01500_),
    .B1(_01496_),
    .B2(\genblk1[3].osc.clkdiv_C.cnt[2] ),
    .X(_01502_));
 sky130_fd_sc_hd__o2111a_1 _06595_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[15] ),
    .A2(_01363_),
    .B1(_01499_),
    .C1(_01501_),
    .D1(_01502_),
    .X(_01503_));
 sky130_fd_sc_hd__or4b_1 _06596_ (.A(\genblk1[3].osc.clkdiv_C.cnt[17] ),
    .B(_01493_),
    .C(_01495_),
    .D_N(_01503_),
    .X(_01504_));
 sky130_fd_sc_hd__or2_1 _06597_ (.A(\genblk1[3].osc.clkdiv_C.cnt[16] ),
    .B(_01197_),
    .X(_01505_));
 sky130_fd_sc_hd__nand2_1 _06598_ (.A(\genblk1[3].osc.clkdiv_C.cnt[16] ),
    .B(_01197_),
    .Y(_01506_));
 sky130_fd_sc_hd__nor2_2 _06599_ (.A(_01441_),
    .B(_01249_),
    .Y(_01507_));
 sky130_fd_sc_hd__nor2_2 _06600_ (.A(_01241_),
    .B(_01432_),
    .Y(_01508_));
 sky130_fd_sc_hd__a2bb2o_1 _06601_ (.A1_N(\genblk1[3].osc.clkdiv_C.cnt[12] ),
    .A2_N(_01507_),
    .B1(_01508_),
    .B2(\genblk1[3].osc.clkdiv_C.cnt[11] ),
    .X(_01509_));
 sky130_fd_sc_hd__a221o_1 _06602_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[0] ),
    .A2(_01484_),
    .B1(_01505_),
    .B2(_01506_),
    .C1(_01509_),
    .X(_01510_));
 sky130_fd_sc_hd__a2111oi_1 _06603_ (.A1(_01486_),
    .A2(_01487_),
    .B1(_01492_),
    .C1(_01504_),
    .D1(_01510_),
    .Y(_01511_));
 sky130_fd_sc_hd__and3_1 _06604_ (.A(_01171_),
    .B(_01192_),
    .C(_01208_),
    .X(_01512_));
 sky130_fd_sc_hd__clkbuf_4 _06605_ (.A(_01512_),
    .X(_01513_));
 sky130_fd_sc_hd__clkbuf_4 _06606_ (.A(_01234_),
    .X(_01514_));
 sky130_fd_sc_hd__o2bb2a_1 _06607_ (.A1_N(\genblk1[3].osc.clkdiv_C.cnt[3] ),
    .A2_N(_01513_),
    .B1(_01514_),
    .B2(\genblk1[3].osc.clkdiv_C.cnt[4] ),
    .X(_01515_));
 sky130_fd_sc_hd__xnor2_1 _06608_ (.A(\genblk1[3].osc.clkdiv_C.cnt[9] ),
    .B(_01210_),
    .Y(_01516_));
 sky130_fd_sc_hd__o2bb2a_1 _06609_ (.A1_N(\genblk1[3].osc.clkdiv_C.cnt[4] ),
    .A2_N(_01514_),
    .B1(_01513_),
    .B2(\genblk1[3].osc.clkdiv_C.cnt[3] ),
    .X(_01517_));
 sky130_fd_sc_hd__o2111a_1 _06610_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[10] ),
    .A2(_01231_),
    .B1(_01515_),
    .C1(_01516_),
    .D1(_01517_),
    .X(_01518_));
 sky130_fd_sc_hd__o21a_2 _06611_ (.A1(_01186_),
    .A2(_01354_),
    .B1(_01171_),
    .X(_01519_));
 sky130_fd_sc_hd__xor2_1 _06612_ (.A(\genblk1[3].osc.clkdiv_C.cnt[1] ),
    .B(_01519_),
    .X(_01520_));
 sky130_fd_sc_hd__o2111a_1 _06613_ (.A1(_01485_),
    .A2(_01256_),
    .B1(_01511_),
    .C1(_01518_),
    .D1(_01520_),
    .X(_01521_));
 sky130_fd_sc_hd__o221a_1 _06614_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[8] ),
    .A2(_01483_),
    .B1(_01484_),
    .B2(\genblk1[3].osc.clkdiv_C.cnt[0] ),
    .C1(_01521_),
    .X(_01522_));
 sky130_fd_sc_hd__clkbuf_4 _06615_ (.A(_01522_),
    .X(_01523_));
 sky130_fd_sc_hd__nor2_1 _06616_ (.A(net1101),
    .B(_01523_),
    .Y(\genblk1[3].osc.clkdiv_C.next_cnt[0] ));
 sky130_fd_sc_hd__inv_2 _06617_ (.A(_01522_),
    .Y(_01524_));
 sky130_fd_sc_hd__nand2_1 _06618_ (.A(\genblk1[3].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[3].osc.clkdiv_C.cnt[0] ),
    .Y(_01525_));
 sky130_fd_sc_hd__or2_1 _06619_ (.A(\genblk1[3].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[3].osc.clkdiv_C.cnt[0] ),
    .X(_01526_));
 sky130_fd_sc_hd__and3_1 _06620_ (.A(_01524_),
    .B(_01525_),
    .C(_01526_),
    .X(_01527_));
 sky130_fd_sc_hd__clkbuf_1 _06621_ (.A(_01527_),
    .X(\genblk1[3].osc.clkdiv_C.next_cnt[1] ));
 sky130_fd_sc_hd__and3_1 _06622_ (.A(\genblk1[3].osc.clkdiv_C.cnt[2] ),
    .B(\genblk1[3].osc.clkdiv_C.cnt[1] ),
    .C(\genblk1[3].osc.clkdiv_C.cnt[0] ),
    .X(_01528_));
 sky130_fd_sc_hd__a21oi_1 _06623_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[1] ),
    .A2(\genblk1[3].osc.clkdiv_C.cnt[0] ),
    .B1(\genblk1[3].osc.clkdiv_C.cnt[2] ),
    .Y(_01529_));
 sky130_fd_sc_hd__nor3_1 _06624_ (.A(_01523_),
    .B(_01528_),
    .C(_01529_),
    .Y(\genblk1[3].osc.clkdiv_C.next_cnt[2] ));
 sky130_fd_sc_hd__and2_1 _06625_ (.A(\genblk1[3].osc.clkdiv_C.cnt[3] ),
    .B(_01528_),
    .X(_01530_));
 sky130_fd_sc_hd__nor2_1 _06626_ (.A(\genblk1[3].osc.clkdiv_C.cnt[3] ),
    .B(_01528_),
    .Y(_01531_));
 sky130_fd_sc_hd__nor3_1 _06627_ (.A(_01523_),
    .B(_01530_),
    .C(_01531_),
    .Y(\genblk1[3].osc.clkdiv_C.next_cnt[3] ));
 sky130_fd_sc_hd__o21ai_1 _06628_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[4] ),
    .A2(_01530_),
    .B1(_01524_),
    .Y(_01532_));
 sky130_fd_sc_hd__a21oi_1 _06629_ (.A1(net1077),
    .A2(_01530_),
    .B1(_01532_),
    .Y(\genblk1[3].osc.clkdiv_C.next_cnt[4] ));
 sky130_fd_sc_hd__and3_1 _06630_ (.A(\genblk1[3].osc.clkdiv_C.cnt[5] ),
    .B(\genblk1[3].osc.clkdiv_C.cnt[4] ),
    .C(_01530_),
    .X(_01533_));
 sky130_fd_sc_hd__a21oi_1 _06631_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[4] ),
    .A2(_01530_),
    .B1(\genblk1[3].osc.clkdiv_C.cnt[5] ),
    .Y(_01534_));
 sky130_fd_sc_hd__nor3_1 _06632_ (.A(_01523_),
    .B(_01533_),
    .C(_01534_),
    .Y(\genblk1[3].osc.clkdiv_C.next_cnt[5] ));
 sky130_fd_sc_hd__and2_1 _06633_ (.A(\genblk1[3].osc.clkdiv_C.cnt[6] ),
    .B(_01533_),
    .X(_01535_));
 sky130_fd_sc_hd__nor2_1 _06634_ (.A(\genblk1[3].osc.clkdiv_C.cnt[6] ),
    .B(_01533_),
    .Y(_01536_));
 sky130_fd_sc_hd__nor3_1 _06635_ (.A(_01523_),
    .B(_01535_),
    .C(_01536_),
    .Y(\genblk1[3].osc.clkdiv_C.next_cnt[6] ));
 sky130_fd_sc_hd__o21ai_1 _06636_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[7] ),
    .A2(_01535_),
    .B1(_01524_),
    .Y(_01537_));
 sky130_fd_sc_hd__a21oi_1 _06637_ (.A1(net1095),
    .A2(_01535_),
    .B1(_01537_),
    .Y(\genblk1[3].osc.clkdiv_C.next_cnt[7] ));
 sky130_fd_sc_hd__and3_1 _06638_ (.A(\genblk1[3].osc.clkdiv_C.cnt[8] ),
    .B(\genblk1[3].osc.clkdiv_C.cnt[7] ),
    .C(_01535_),
    .X(_01538_));
 sky130_fd_sc_hd__a21oi_1 _06639_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[7] ),
    .A2(_01535_),
    .B1(\genblk1[3].osc.clkdiv_C.cnt[8] ),
    .Y(_01539_));
 sky130_fd_sc_hd__nor3_1 _06640_ (.A(_01523_),
    .B(_01538_),
    .C(_01539_),
    .Y(\genblk1[3].osc.clkdiv_C.next_cnt[8] ));
 sky130_fd_sc_hd__and2_1 _06641_ (.A(\genblk1[3].osc.clkdiv_C.cnt[9] ),
    .B(_01538_),
    .X(_01540_));
 sky130_fd_sc_hd__nor2_1 _06642_ (.A(_01523_),
    .B(_01540_),
    .Y(_01541_));
 sky130_fd_sc_hd__o21a_1 _06643_ (.A1(net1145),
    .A2(_01538_),
    .B1(_01541_),
    .X(\genblk1[3].osc.clkdiv_C.next_cnt[9] ));
 sky130_fd_sc_hd__nand2_1 _06644_ (.A(\genblk1[3].osc.clkdiv_C.cnt[10] ),
    .B(_01540_),
    .Y(_01542_));
 sky130_fd_sc_hd__o211a_1 _06645_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[10] ),
    .A2(_01540_),
    .B1(_01542_),
    .C1(_01524_),
    .X(\genblk1[3].osc.clkdiv_C.next_cnt[10] ));
 sky130_fd_sc_hd__nor2_1 _06646_ (.A(_01486_),
    .B(_01542_),
    .Y(_01543_));
 sky130_fd_sc_hd__or2_1 _06647_ (.A(_01522_),
    .B(_01543_),
    .X(_01544_));
 sky130_fd_sc_hd__a21oi_1 _06648_ (.A1(_01486_),
    .A2(_01542_),
    .B1(_01544_),
    .Y(\genblk1[3].osc.clkdiv_C.next_cnt[11] ));
 sky130_fd_sc_hd__and2_1 _06649_ (.A(\genblk1[3].osc.clkdiv_C.cnt[12] ),
    .B(_01543_),
    .X(_01545_));
 sky130_fd_sc_hd__nor2_1 _06650_ (.A(_01523_),
    .B(_01545_),
    .Y(_01546_));
 sky130_fd_sc_hd__o21a_1 _06651_ (.A1(net1193),
    .A2(_01543_),
    .B1(_01546_),
    .X(\genblk1[3].osc.clkdiv_C.next_cnt[12] ));
 sky130_fd_sc_hd__and3_1 _06652_ (.A(\genblk1[3].osc.clkdiv_C.cnt[13] ),
    .B(\genblk1[3].osc.clkdiv_C.cnt[12] ),
    .C(_01543_),
    .X(_01547_));
 sky130_fd_sc_hd__nor2_1 _06653_ (.A(_01523_),
    .B(_01547_),
    .Y(_01548_));
 sky130_fd_sc_hd__o21a_1 _06654_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[13] ),
    .A2(_01545_),
    .B1(_01548_),
    .X(\genblk1[3].osc.clkdiv_C.next_cnt[13] ));
 sky130_fd_sc_hd__and2_1 _06655_ (.A(\genblk1[3].osc.clkdiv_C.cnt[14] ),
    .B(_01547_),
    .X(_01549_));
 sky130_fd_sc_hd__nor2_1 _06656_ (.A(_01523_),
    .B(_01549_),
    .Y(_01550_));
 sky130_fd_sc_hd__o21a_1 _06657_ (.A1(net1195),
    .A2(_01547_),
    .B1(_01550_),
    .X(\genblk1[3].osc.clkdiv_C.next_cnt[14] ));
 sky130_fd_sc_hd__and3_1 _06658_ (.A(\genblk1[3].osc.clkdiv_C.cnt[15] ),
    .B(\genblk1[3].osc.clkdiv_C.cnt[14] ),
    .C(_01547_),
    .X(_01551_));
 sky130_fd_sc_hd__nor2_1 _06659_ (.A(_01522_),
    .B(_01551_),
    .Y(_01552_));
 sky130_fd_sc_hd__o21a_1 _06660_ (.A1(net1237),
    .A2(_01549_),
    .B1(_01552_),
    .X(\genblk1[3].osc.clkdiv_C.next_cnt[15] ));
 sky130_fd_sc_hd__or2_1 _06661_ (.A(\genblk1[3].osc.clkdiv_C.cnt[16] ),
    .B(_01551_),
    .X(_01553_));
 sky130_fd_sc_hd__nand2_1 _06662_ (.A(\genblk1[3].osc.clkdiv_C.cnt[16] ),
    .B(_01551_),
    .Y(_01554_));
 sky130_fd_sc_hd__and3_1 _06663_ (.A(_01524_),
    .B(_01553_),
    .C(_01554_),
    .X(_01555_));
 sky130_fd_sc_hd__clkbuf_1 _06664_ (.A(_01555_),
    .X(\genblk1[3].osc.clkdiv_C.next_cnt[16] ));
 sky130_fd_sc_hd__xnor2_1 _06665_ (.A(net436),
    .B(_01554_),
    .Y(\genblk1[3].osc.clkdiv_C.next_cnt[17] ));
 sky130_fd_sc_hd__a21o_4 _06666_ (.A1(_01230_),
    .A2(_01221_),
    .B1(_01223_),
    .X(_01556_));
 sky130_fd_sc_hd__nand2_1 _06667_ (.A(_01556_),
    .B(_01344_),
    .Y(_01557_));
 sky130_fd_sc_hd__nor2_1 _06668_ (.A(\genblk1[4].osc.clkdiv_C.cnt[6] ),
    .B(_01557_),
    .Y(_01558_));
 sky130_fd_sc_hd__nand2_2 _06669_ (.A(_01349_),
    .B(_01180_),
    .Y(_01559_));
 sky130_fd_sc_hd__a22o_1 _06670_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[2] ),
    .A2(_01559_),
    .B1(_01557_),
    .B2(\genblk1[4].osc.clkdiv_C.cnt[6] ),
    .X(_01560_));
 sky130_fd_sc_hd__nor2_1 _06671_ (.A(\genblk1[4].osc.clkdiv_C.cnt[2] ),
    .B(_01559_),
    .Y(_01561_));
 sky130_fd_sc_hd__a2bb2o_1 _06672_ (.A1_N(\genblk1[4].osc.clkdiv_C.cnt[3] ),
    .A2_N(_01326_),
    .B1(_01498_),
    .B2(\genblk1[4].osc.clkdiv_C.cnt[14] ),
    .X(_01562_));
 sky130_fd_sc_hd__or2b_1 _06673_ (.A(_01175_),
    .B_N(_01194_),
    .X(_01563_));
 sky130_fd_sc_hd__buf_6 _06674_ (.A(_01563_),
    .X(_01564_));
 sky130_fd_sc_hd__nand2_4 _06675_ (.A(_01187_),
    .B(_01564_),
    .Y(_01565_));
 sky130_fd_sc_hd__and2_1 _06676_ (.A(\genblk1[4].osc.clkdiv_C.cnt[5] ),
    .B(_01565_),
    .X(_01566_));
 sky130_fd_sc_hd__nor2_1 _06677_ (.A(\genblk1[4].osc.clkdiv_C.cnt[5] ),
    .B(_01565_),
    .Y(_01567_));
 sky130_fd_sc_hd__inv_2 _06678_ (.A(\genblk1[4].osc.clkdiv_C.cnt[1] ),
    .Y(_01568_));
 sky130_fd_sc_hd__a221o_1 _06679_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[15] ),
    .A2(_01363_),
    .B1(_01242_),
    .B2(_01568_),
    .C1(\genblk1[4].osc.clkdiv_C.cnt[17] ),
    .X(_01569_));
 sky130_fd_sc_hd__inv_2 _06680_ (.A(\genblk1[4].osc.clkdiv_C.cnt[4] ),
    .Y(_01570_));
 sky130_fd_sc_hd__o22a_1 _06681_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[15] ),
    .A2(_01362_),
    .B1(_01248_),
    .B2(_01570_),
    .X(_01571_));
 sky130_fd_sc_hd__o221a_1 _06682_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[4] ),
    .A2(_01439_),
    .B1(_01340_),
    .B2(\genblk1[4].osc.clkdiv_C.cnt[8] ),
    .C1(_01571_),
    .X(_01572_));
 sky130_fd_sc_hd__or4b_1 _06683_ (.A(_01566_),
    .B(_01567_),
    .C(_01569_),
    .D_N(_01572_),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_4 _06684_ (.A0(_01173_),
    .A1(_01187_),
    .S(_01188_),
    .X(_01574_));
 sky130_fd_sc_hd__or3_1 _06685_ (.A(_01194_),
    .B(_01175_),
    .C(_01191_),
    .X(_01575_));
 sky130_fd_sc_hd__buf_4 _06686_ (.A(_01575_),
    .X(_01576_));
 sky130_fd_sc_hd__clkbuf_8 _06687_ (.A(_01576_),
    .X(_01577_));
 sky130_fd_sc_hd__buf_4 _06688_ (.A(_01577_),
    .X(_01578_));
 sky130_fd_sc_hd__a2bb2o_1 _06689_ (.A1_N(\genblk1[4].osc.clkdiv_C.cnt[12] ),
    .A2_N(_01574_),
    .B1(_01578_),
    .B2(\genblk1[4].osc.clkdiv_C.cnt[16] ),
    .X(_01579_));
 sky130_fd_sc_hd__o2bb2a_1 _06690_ (.A1_N(\genblk1[4].osc.clkdiv_C.cnt[0] ),
    .A2_N(_01209_),
    .B1(_01578_),
    .B2(\genblk1[4].osc.clkdiv_C.cnt[16] ),
    .X(_01580_));
 sky130_fd_sc_hd__o221a_1 _06691_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[0] ),
    .A2(_01210_),
    .B1(_01498_),
    .B2(\genblk1[4].osc.clkdiv_C.cnt[14] ),
    .C1(_01580_),
    .X(_01581_));
 sky130_fd_sc_hd__or4b_1 _06692_ (.A(_01562_),
    .B(_01573_),
    .C(_01579_),
    .D_N(_01581_),
    .X(_01582_));
 sky130_fd_sc_hd__a2bb2o_1 _06693_ (.A1_N(\genblk1[4].osc.clkdiv_C.cnt[11] ),
    .A2_N(_01313_),
    .B1(_01340_),
    .B2(\genblk1[4].osc.clkdiv_C.cnt[8] ),
    .X(_01583_));
 sky130_fd_sc_hd__a2111o_1 _06694_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[11] ),
    .A2(_01313_),
    .B1(_01561_),
    .C1(_01582_),
    .D1(_01583_),
    .X(_01584_));
 sky130_fd_sc_hd__nor2_1 _06695_ (.A(\genblk1[4].osc.clkdiv_C.cnt[10] ),
    .B(_01323_),
    .Y(_01585_));
 sky130_fd_sc_hd__a22o_1 _06696_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[3] ),
    .A2(_01326_),
    .B1(_01574_),
    .B2(\genblk1[4].osc.clkdiv_C.cnt[12] ),
    .X(_01586_));
 sky130_fd_sc_hd__a221o_1 _06697_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[1] ),
    .A2(_01436_),
    .B1(_01304_),
    .B2(\genblk1[4].osc.clkdiv_C.cnt[7] ),
    .C1(_01586_),
    .X(_01587_));
 sky130_fd_sc_hd__inv_2 _06698_ (.A(\genblk1[4].osc.clkdiv_C.cnt[10] ),
    .Y(_01588_));
 sky130_fd_sc_hd__nand2_4 _06699_ (.A(_01320_),
    .B(_01321_),
    .Y(_01589_));
 sky130_fd_sc_hd__nor2_1 _06700_ (.A(_01588_),
    .B(_01589_),
    .Y(_01590_));
 sky130_fd_sc_hd__or3b_4 _06701_ (.A(_01173_),
    .B(_01175_),
    .C_N(_01191_),
    .X(_01591_));
 sky130_fd_sc_hd__nand2_4 _06702_ (.A(_01171_),
    .B(_01591_),
    .Y(_01592_));
 sky130_fd_sc_hd__nand2_1 _06703_ (.A(\genblk1[4].osc.clkdiv_C.cnt[9] ),
    .B(_01592_),
    .Y(_01593_));
 sky130_fd_sc_hd__or2_1 _06704_ (.A(\genblk1[4].osc.clkdiv_C.cnt[9] ),
    .B(_01592_),
    .X(_01594_));
 sky130_fd_sc_hd__nor2_4 _06705_ (.A(_01489_),
    .B(_01196_),
    .Y(_01595_));
 sky130_fd_sc_hd__xnor2_1 _06706_ (.A(\genblk1[4].osc.clkdiv_C.cnt[13] ),
    .B(_01595_),
    .Y(_01596_));
 sky130_fd_sc_hd__o2111a_1 _06707_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[7] ),
    .A2(_01304_),
    .B1(_01593_),
    .C1(_01594_),
    .D1(_01596_),
    .X(_01597_));
 sky130_fd_sc_hd__or4b_1 _06708_ (.A(_01585_),
    .B(_01587_),
    .C(_01590_),
    .D_N(_01597_),
    .X(_01598_));
 sky130_fd_sc_hd__or4_4 _06709_ (.A(_01558_),
    .B(_01560_),
    .C(_01584_),
    .D(_01598_),
    .X(_01599_));
 sky130_fd_sc_hd__buf_2 _06710_ (.A(_01599_),
    .X(_01600_));
 sky130_fd_sc_hd__and2b_1 _06711_ (.A_N(\genblk1[4].osc.clkdiv_C.cnt[0] ),
    .B(_01600_),
    .X(_01601_));
 sky130_fd_sc_hd__clkbuf_1 _06712_ (.A(_01601_),
    .X(\genblk1[4].osc.clkdiv_C.next_cnt[0] ));
 sky130_fd_sc_hd__or2_1 _06713_ (.A(\genblk1[4].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[4].osc.clkdiv_C.cnt[0] ),
    .X(_01602_));
 sky130_fd_sc_hd__nand2_1 _06714_ (.A(\genblk1[4].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[4].osc.clkdiv_C.cnt[0] ),
    .Y(_01603_));
 sky130_fd_sc_hd__and3_1 _06715_ (.A(_01600_),
    .B(_01602_),
    .C(_01603_),
    .X(_01604_));
 sky130_fd_sc_hd__clkbuf_1 _06716_ (.A(_01604_),
    .X(\genblk1[4].osc.clkdiv_C.next_cnt[1] ));
 sky130_fd_sc_hd__and3_1 _06717_ (.A(\genblk1[4].osc.clkdiv_C.cnt[2] ),
    .B(\genblk1[4].osc.clkdiv_C.cnt[1] ),
    .C(\genblk1[4].osc.clkdiv_C.cnt[0] ),
    .X(_01605_));
 sky130_fd_sc_hd__inv_2 _06718_ (.A(_01605_),
    .Y(_01606_));
 sky130_fd_sc_hd__a21o_1 _06719_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[1] ),
    .A2(\genblk1[4].osc.clkdiv_C.cnt[0] ),
    .B1(\genblk1[4].osc.clkdiv_C.cnt[2] ),
    .X(_01607_));
 sky130_fd_sc_hd__and3_1 _06720_ (.A(_01600_),
    .B(_01606_),
    .C(_01607_),
    .X(_01608_));
 sky130_fd_sc_hd__clkbuf_1 _06721_ (.A(_01608_),
    .X(\genblk1[4].osc.clkdiv_C.next_cnt[2] ));
 sky130_fd_sc_hd__and2_1 _06722_ (.A(\genblk1[4].osc.clkdiv_C.cnt[3] ),
    .B(_01605_),
    .X(_01609_));
 sky130_fd_sc_hd__inv_2 _06723_ (.A(_01609_),
    .Y(_01610_));
 sky130_fd_sc_hd__or2_1 _06724_ (.A(\genblk1[4].osc.clkdiv_C.cnt[3] ),
    .B(_01605_),
    .X(_01611_));
 sky130_fd_sc_hd__and3_1 _06725_ (.A(_01600_),
    .B(_01610_),
    .C(_01611_),
    .X(_01612_));
 sky130_fd_sc_hd__clkbuf_1 _06726_ (.A(_01612_),
    .X(\genblk1[4].osc.clkdiv_C.next_cnt[3] ));
 sky130_fd_sc_hd__nand2_1 _06727_ (.A(\genblk1[4].osc.clkdiv_C.cnt[4] ),
    .B(_01609_),
    .Y(_01613_));
 sky130_fd_sc_hd__or2_1 _06728_ (.A(\genblk1[4].osc.clkdiv_C.cnt[4] ),
    .B(_01609_),
    .X(_01614_));
 sky130_fd_sc_hd__and3_1 _06729_ (.A(_01600_),
    .B(_01613_),
    .C(_01614_),
    .X(_01615_));
 sky130_fd_sc_hd__clkbuf_1 _06730_ (.A(_01615_),
    .X(\genblk1[4].osc.clkdiv_C.next_cnt[4] ));
 sky130_fd_sc_hd__and3_1 _06731_ (.A(\genblk1[4].osc.clkdiv_C.cnt[5] ),
    .B(\genblk1[4].osc.clkdiv_C.cnt[4] ),
    .C(_01609_),
    .X(_01616_));
 sky130_fd_sc_hd__inv_2 _06732_ (.A(_01616_),
    .Y(_01617_));
 sky130_fd_sc_hd__a31o_1 _06733_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[4] ),
    .A2(\genblk1[4].osc.clkdiv_C.cnt[3] ),
    .A3(_01605_),
    .B1(\genblk1[4].osc.clkdiv_C.cnt[5] ),
    .X(_01618_));
 sky130_fd_sc_hd__and3_1 _06734_ (.A(_01600_),
    .B(_01617_),
    .C(_01618_),
    .X(_01619_));
 sky130_fd_sc_hd__clkbuf_1 _06735_ (.A(_01619_),
    .X(\genblk1[4].osc.clkdiv_C.next_cnt[5] ));
 sky130_fd_sc_hd__and2_1 _06736_ (.A(\genblk1[4].osc.clkdiv_C.cnt[6] ),
    .B(_01616_),
    .X(_01620_));
 sky130_fd_sc_hd__inv_2 _06737_ (.A(_01620_),
    .Y(_01621_));
 sky130_fd_sc_hd__or2_1 _06738_ (.A(\genblk1[4].osc.clkdiv_C.cnt[6] ),
    .B(_01616_),
    .X(_01622_));
 sky130_fd_sc_hd__and3_1 _06739_ (.A(_01600_),
    .B(_01621_),
    .C(_01622_),
    .X(_01623_));
 sky130_fd_sc_hd__clkbuf_1 _06740_ (.A(_01623_),
    .X(\genblk1[4].osc.clkdiv_C.next_cnt[6] ));
 sky130_fd_sc_hd__nand2_1 _06741_ (.A(\genblk1[4].osc.clkdiv_C.cnt[7] ),
    .B(_01620_),
    .Y(_01624_));
 sky130_fd_sc_hd__or2_1 _06742_ (.A(\genblk1[4].osc.clkdiv_C.cnt[7] ),
    .B(_01620_),
    .X(_01625_));
 sky130_fd_sc_hd__and3_1 _06743_ (.A(_01599_),
    .B(_01624_),
    .C(_01625_),
    .X(_01626_));
 sky130_fd_sc_hd__clkbuf_1 _06744_ (.A(_01626_),
    .X(\genblk1[4].osc.clkdiv_C.next_cnt[7] ));
 sky130_fd_sc_hd__and3_1 _06745_ (.A(\genblk1[4].osc.clkdiv_C.cnt[8] ),
    .B(\genblk1[4].osc.clkdiv_C.cnt[7] ),
    .C(_01620_),
    .X(_01627_));
 sky130_fd_sc_hd__inv_2 _06746_ (.A(_01627_),
    .Y(_01628_));
 sky130_fd_sc_hd__a31o_1 _06747_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[7] ),
    .A2(\genblk1[4].osc.clkdiv_C.cnt[6] ),
    .A3(_01616_),
    .B1(\genblk1[4].osc.clkdiv_C.cnt[8] ),
    .X(_01629_));
 sky130_fd_sc_hd__and3_1 _06748_ (.A(_01599_),
    .B(_01628_),
    .C(_01629_),
    .X(_01630_));
 sky130_fd_sc_hd__clkbuf_1 _06749_ (.A(_01630_),
    .X(\genblk1[4].osc.clkdiv_C.next_cnt[8] ));
 sky130_fd_sc_hd__and2_1 _06750_ (.A(\genblk1[4].osc.clkdiv_C.cnt[9] ),
    .B(_01627_),
    .X(_01631_));
 sky130_fd_sc_hd__inv_2 _06751_ (.A(_01631_),
    .Y(_01632_));
 sky130_fd_sc_hd__or2_1 _06752_ (.A(\genblk1[4].osc.clkdiv_C.cnt[9] ),
    .B(_01627_),
    .X(_01633_));
 sky130_fd_sc_hd__and3_1 _06753_ (.A(_01599_),
    .B(_01632_),
    .C(_01633_),
    .X(_01634_));
 sky130_fd_sc_hd__clkbuf_1 _06754_ (.A(_01634_),
    .X(\genblk1[4].osc.clkdiv_C.next_cnt[9] ));
 sky130_fd_sc_hd__nand2_1 _06755_ (.A(\genblk1[4].osc.clkdiv_C.cnt[10] ),
    .B(_01631_),
    .Y(_01635_));
 sky130_fd_sc_hd__o211a_1 _06756_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[10] ),
    .A2(_01631_),
    .B1(_01635_),
    .C1(_01600_),
    .X(\genblk1[4].osc.clkdiv_C.next_cnt[10] ));
 sky130_fd_sc_hd__a31o_1 _06757_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[10] ),
    .A2(\genblk1[4].osc.clkdiv_C.cnt[9] ),
    .A3(_01627_),
    .B1(\genblk1[4].osc.clkdiv_C.cnt[11] ),
    .X(_01636_));
 sky130_fd_sc_hd__and3_1 _06758_ (.A(\genblk1[4].osc.clkdiv_C.cnt[11] ),
    .B(\genblk1[4].osc.clkdiv_C.cnt[10] ),
    .C(_01631_),
    .X(_01637_));
 sky130_fd_sc_hd__inv_2 _06759_ (.A(_01637_),
    .Y(_01638_));
 sky130_fd_sc_hd__and3_1 _06760_ (.A(_01599_),
    .B(_01636_),
    .C(_01638_),
    .X(_01639_));
 sky130_fd_sc_hd__clkbuf_1 _06761_ (.A(_01639_),
    .X(\genblk1[4].osc.clkdiv_C.next_cnt[11] ));
 sky130_fd_sc_hd__or2_1 _06762_ (.A(\genblk1[4].osc.clkdiv_C.cnt[12] ),
    .B(_01637_),
    .X(_01640_));
 sky130_fd_sc_hd__and2_1 _06763_ (.A(\genblk1[4].osc.clkdiv_C.cnt[12] ),
    .B(_01637_),
    .X(_01641_));
 sky130_fd_sc_hd__inv_2 _06764_ (.A(_01641_),
    .Y(_01642_));
 sky130_fd_sc_hd__and3_1 _06765_ (.A(_01599_),
    .B(_01640_),
    .C(_01642_),
    .X(_01643_));
 sky130_fd_sc_hd__clkbuf_1 _06766_ (.A(_01643_),
    .X(\genblk1[4].osc.clkdiv_C.next_cnt[12] ));
 sky130_fd_sc_hd__inv_2 _06767_ (.A(\genblk1[4].osc.clkdiv_C.cnt[13] ),
    .Y(_01644_));
 sky130_fd_sc_hd__or2_1 _06768_ (.A(\genblk1[4].osc.clkdiv_C.cnt[13] ),
    .B(_01641_),
    .X(_01645_));
 sky130_fd_sc_hd__o211a_1 _06769_ (.A1(_01644_),
    .A2(_01642_),
    .B1(_01645_),
    .C1(_01600_),
    .X(\genblk1[4].osc.clkdiv_C.next_cnt[13] ));
 sky130_fd_sc_hd__a31o_1 _06770_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[13] ),
    .A2(\genblk1[4].osc.clkdiv_C.cnt[12] ),
    .A3(_01637_),
    .B1(\genblk1[4].osc.clkdiv_C.cnt[14] ),
    .X(_01646_));
 sky130_fd_sc_hd__and3_1 _06771_ (.A(\genblk1[4].osc.clkdiv_C.cnt[14] ),
    .B(\genblk1[4].osc.clkdiv_C.cnt[13] ),
    .C(_01641_),
    .X(_01647_));
 sky130_fd_sc_hd__inv_2 _06772_ (.A(_01647_),
    .Y(_01648_));
 sky130_fd_sc_hd__and3_1 _06773_ (.A(_01599_),
    .B(_01646_),
    .C(_01648_),
    .X(_01649_));
 sky130_fd_sc_hd__clkbuf_1 _06774_ (.A(_01649_),
    .X(\genblk1[4].osc.clkdiv_C.next_cnt[14] ));
 sky130_fd_sc_hd__inv_2 _06775_ (.A(\genblk1[4].osc.clkdiv_C.cnt[15] ),
    .Y(_01650_));
 sky130_fd_sc_hd__or2_1 _06776_ (.A(\genblk1[4].osc.clkdiv_C.cnt[15] ),
    .B(_01647_),
    .X(_01651_));
 sky130_fd_sc_hd__o211a_1 _06777_ (.A1(_01650_),
    .A2(_01648_),
    .B1(_01651_),
    .C1(_01600_),
    .X(\genblk1[4].osc.clkdiv_C.next_cnt[15] ));
 sky130_fd_sc_hd__nor2_1 _06778_ (.A(_01650_),
    .B(_01648_),
    .Y(_01652_));
 sky130_fd_sc_hd__or2_1 _06779_ (.A(\genblk1[4].osc.clkdiv_C.cnt[16] ),
    .B(_01652_),
    .X(_01653_));
 sky130_fd_sc_hd__nand2_1 _06780_ (.A(\genblk1[4].osc.clkdiv_C.cnt[16] ),
    .B(_01652_),
    .Y(_01654_));
 sky130_fd_sc_hd__and3_1 _06781_ (.A(_01599_),
    .B(_01653_),
    .C(_01654_),
    .X(_01655_));
 sky130_fd_sc_hd__clkbuf_1 _06782_ (.A(_01655_),
    .X(\genblk1[4].osc.clkdiv_C.next_cnt[16] ));
 sky130_fd_sc_hd__xnor2_1 _06783_ (.A(net851),
    .B(_01654_),
    .Y(\genblk1[4].osc.clkdiv_C.next_cnt[17] ));
 sky130_fd_sc_hd__a21oi_1 _06784_ (.A1(_01436_),
    .A2(_01304_),
    .B1(\genblk1[5].osc.clkdiv_C.cnt[1] ),
    .Y(_01656_));
 sky130_fd_sc_hd__xnor2_1 _06785_ (.A(\genblk1[5].osc.clkdiv_C.cnt[4] ),
    .B(_01483_),
    .Y(_01657_));
 sky130_fd_sc_hd__nand2_2 _06786_ (.A(_01489_),
    .B(net37),
    .Y(_01658_));
 sky130_fd_sc_hd__xor2_1 _06787_ (.A(\genblk1[5].osc.clkdiv_C.cnt[10] ),
    .B(_01658_),
    .X(_01659_));
 sky130_fd_sc_hd__nor2_1 _06788_ (.A(_01179_),
    .B(_01262_),
    .Y(_01660_));
 sky130_fd_sc_hd__xnor2_1 _06789_ (.A(\genblk1[5].osc.clkdiv_C.cnt[2] ),
    .B(_01660_),
    .Y(_01661_));
 sky130_fd_sc_hd__xnor2_1 _06790_ (.A(\genblk1[5].osc.clkdiv_C.cnt[5] ),
    .B(net36),
    .Y(_01662_));
 sky130_fd_sc_hd__xnor2_1 _06791_ (.A(\genblk1[5].osc.clkdiv_C.cnt[16] ),
    .B(_01578_),
    .Y(_01663_));
 sky130_fd_sc_hd__or4_1 _06792_ (.A(_01659_),
    .B(_01661_),
    .C(_01662_),
    .D(_01663_),
    .X(_01664_));
 sky130_fd_sc_hd__xnor2_1 _06793_ (.A(\genblk1[5].osc.clkdiv_C.cnt[3] ),
    .B(_01592_),
    .Y(_01665_));
 sky130_fd_sc_hd__nand2_4 _06794_ (.A(_01440_),
    .B(_01171_),
    .Y(_01666_));
 sky130_fd_sc_hd__or2_2 _06795_ (.A(_01325_),
    .B(_01254_),
    .X(_01667_));
 sky130_fd_sc_hd__a2bb2o_1 _06796_ (.A1_N(\genblk1[5].osc.clkdiv_C.cnt[13] ),
    .A2_N(_01666_),
    .B1(_01667_),
    .B2(\genblk1[5].osc.clkdiv_C.cnt[11] ),
    .X(_01668_));
 sky130_fd_sc_hd__inv_2 _06797_ (.A(\genblk1[5].osc.clkdiv_C.cnt[7] ),
    .Y(_01669_));
 sky130_fd_sc_hd__inv_2 _06798_ (.A(\genblk1[5].osc.clkdiv_C.cnt[6] ),
    .Y(_01670_));
 sky130_fd_sc_hd__a221o_1 _06799_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[14] ),
    .A2(_01210_),
    .B1(_01304_),
    .B2(\genblk1[5].osc.clkdiv_C.cnt[1] ),
    .C1(_01670_),
    .X(_01671_));
 sky130_fd_sc_hd__a2bb2o_1 _06800_ (.A1_N(\genblk1[5].osc.clkdiv_C.cnt[11] ),
    .A2_N(_01667_),
    .B1(_01666_),
    .B2(\genblk1[5].osc.clkdiv_C.cnt[13] ),
    .X(_01672_));
 sky130_fd_sc_hd__a221o_1 _06801_ (.A1(_01669_),
    .A2(_01559_),
    .B1(_01671_),
    .B2(_01436_),
    .C1(_01672_),
    .X(_01673_));
 sky130_fd_sc_hd__nor2_1 _06802_ (.A(_01238_),
    .B(net36),
    .Y(_01674_));
 sky130_fd_sc_hd__buf_4 _06803_ (.A(_01674_),
    .X(_01675_));
 sky130_fd_sc_hd__a21o_1 _06804_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[15] ),
    .A2(_01362_),
    .B1(\genblk1[5].osc.clkdiv_C.cnt[17] ),
    .X(_01676_));
 sky130_fd_sc_hd__and3_1 _06805_ (.A(\genblk1[5].osc.clkdiv_C.cnt[9] ),
    .B(_01362_),
    .C(_01226_),
    .X(_01677_));
 sky130_fd_sc_hd__nor2_4 _06806_ (.A(_01336_),
    .B(_01564_),
    .Y(_01678_));
 sky130_fd_sc_hd__nor2_1 _06807_ (.A(\genblk1[5].osc.clkdiv_C.cnt[9] ),
    .B(_01678_),
    .Y(_01679_));
 sky130_fd_sc_hd__or2_1 _06808_ (.A(\genblk1[5].osc.clkdiv_C.cnt[15] ),
    .B(_01359_),
    .X(_01680_));
 sky130_fd_sc_hd__or4b_1 _06809_ (.A(_01676_),
    .B(_01677_),
    .C(_01679_),
    .D_N(_01680_),
    .X(_01681_));
 sky130_fd_sc_hd__nand2_1 _06810_ (.A(\genblk1[5].osc.clkdiv_C.cnt[8] ),
    .B(_01326_),
    .Y(_01682_));
 sky130_fd_sc_hd__or2_1 _06811_ (.A(\genblk1[5].osc.clkdiv_C.cnt[8] ),
    .B(_01326_),
    .X(_01683_));
 sky130_fd_sc_hd__nor2_2 _06812_ (.A(_01189_),
    .B(_01678_),
    .Y(_01684_));
 sky130_fd_sc_hd__xnor2_1 _06813_ (.A(\genblk1[5].osc.clkdiv_C.cnt[0] ),
    .B(_01684_),
    .Y(_01685_));
 sky130_fd_sc_hd__a221o_1 _06814_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[6] ),
    .A2(_01242_),
    .B1(_01682_),
    .B2(_01683_),
    .C1(_01685_),
    .X(_01686_));
 sky130_fd_sc_hd__nand2_1 _06815_ (.A(\genblk1[5].osc.clkdiv_C.cnt[12] ),
    .B(_01355_),
    .Y(_01687_));
 sky130_fd_sc_hd__or2_1 _06816_ (.A(\genblk1[5].osc.clkdiv_C.cnt[12] ),
    .B(_01355_),
    .X(_01688_));
 sky130_fd_sc_hd__and4bb_1 _06817_ (.A_N(_01681_),
    .B_N(_01686_),
    .C(_01687_),
    .D(_01688_),
    .X(_01689_));
 sky130_fd_sc_hd__o221a_1 _06818_ (.A1(_01669_),
    .A2(_01559_),
    .B1(_01675_),
    .B2(\genblk1[5].osc.clkdiv_C.cnt[14] ),
    .C1(_01689_),
    .X(_01690_));
 sky130_fd_sc_hd__or4b_1 _06819_ (.A(_01665_),
    .B(_01668_),
    .C(_01673_),
    .D_N(_01690_),
    .X(_01691_));
 sky130_fd_sc_hd__nor4_1 _06820_ (.A(_01656_),
    .B(_01657_),
    .C(_01664_),
    .D(_01691_),
    .Y(_01692_));
 sky130_fd_sc_hd__clkbuf_4 _06821_ (.A(net27),
    .X(_01693_));
 sky130_fd_sc_hd__nor2_1 _06822_ (.A(net1120),
    .B(_01693_),
    .Y(\genblk1[5].osc.clkdiv_C.next_cnt[0] ));
 sky130_fd_sc_hd__inv_2 _06823_ (.A(net1355),
    .Y(_01694_));
 sky130_fd_sc_hd__or2_1 _06824_ (.A(\genblk1[5].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[5].osc.clkdiv_C.cnt[0] ),
    .X(_01695_));
 sky130_fd_sc_hd__nand2_1 _06825_ (.A(\genblk1[5].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[5].osc.clkdiv_C.cnt[0] ),
    .Y(_01696_));
 sky130_fd_sc_hd__and3_1 _06826_ (.A(_01694_),
    .B(_01695_),
    .C(_01696_),
    .X(_01697_));
 sky130_fd_sc_hd__clkbuf_1 _06827_ (.A(_01697_),
    .X(\genblk1[5].osc.clkdiv_C.next_cnt[1] ));
 sky130_fd_sc_hd__and3_1 _06828_ (.A(\genblk1[5].osc.clkdiv_C.cnt[2] ),
    .B(\genblk1[5].osc.clkdiv_C.cnt[1] ),
    .C(\genblk1[5].osc.clkdiv_C.cnt[0] ),
    .X(_01698_));
 sky130_fd_sc_hd__a21oi_1 _06829_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[1] ),
    .A2(\genblk1[5].osc.clkdiv_C.cnt[0] ),
    .B1(\genblk1[5].osc.clkdiv_C.cnt[2] ),
    .Y(_01699_));
 sky130_fd_sc_hd__nor3_1 _06830_ (.A(_01693_),
    .B(_01698_),
    .C(_01699_),
    .Y(\genblk1[5].osc.clkdiv_C.next_cnt[2] ));
 sky130_fd_sc_hd__and2_1 _06831_ (.A(\genblk1[5].osc.clkdiv_C.cnt[3] ),
    .B(_01698_),
    .X(_01700_));
 sky130_fd_sc_hd__nor2_1 _06832_ (.A(\genblk1[5].osc.clkdiv_C.cnt[3] ),
    .B(_01698_),
    .Y(_01701_));
 sky130_fd_sc_hd__nor3_1 _06833_ (.A(_01693_),
    .B(_01700_),
    .C(_01701_),
    .Y(\genblk1[5].osc.clkdiv_C.next_cnt[3] ));
 sky130_fd_sc_hd__o21ai_1 _06834_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[4] ),
    .A2(_01700_),
    .B1(_01694_),
    .Y(_01702_));
 sky130_fd_sc_hd__a21oi_1 _06835_ (.A1(net1105),
    .A2(_01700_),
    .B1(_01702_),
    .Y(\genblk1[5].osc.clkdiv_C.next_cnt[4] ));
 sky130_fd_sc_hd__and3_1 _06836_ (.A(\genblk1[5].osc.clkdiv_C.cnt[5] ),
    .B(\genblk1[5].osc.clkdiv_C.cnt[4] ),
    .C(_01700_),
    .X(_01703_));
 sky130_fd_sc_hd__a21oi_1 _06837_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[4] ),
    .A2(_01700_),
    .B1(\genblk1[5].osc.clkdiv_C.cnt[5] ),
    .Y(_01704_));
 sky130_fd_sc_hd__nor3_1 _06838_ (.A(_01693_),
    .B(_01703_),
    .C(_01704_),
    .Y(\genblk1[5].osc.clkdiv_C.next_cnt[5] ));
 sky130_fd_sc_hd__and2_1 _06839_ (.A(\genblk1[5].osc.clkdiv_C.cnt[6] ),
    .B(_01703_),
    .X(_01705_));
 sky130_fd_sc_hd__nor2_1 _06840_ (.A(\genblk1[5].osc.clkdiv_C.cnt[6] ),
    .B(_01703_),
    .Y(_01706_));
 sky130_fd_sc_hd__nor3_1 _06841_ (.A(_01693_),
    .B(_01705_),
    .C(_01706_),
    .Y(\genblk1[5].osc.clkdiv_C.next_cnt[6] ));
 sky130_fd_sc_hd__o21ai_1 _06842_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[7] ),
    .A2(_01705_),
    .B1(_01694_),
    .Y(_01707_));
 sky130_fd_sc_hd__a21oi_1 _06843_ (.A1(net1072),
    .A2(_01705_),
    .B1(_01707_),
    .Y(\genblk1[5].osc.clkdiv_C.next_cnt[7] ));
 sky130_fd_sc_hd__and3_1 _06844_ (.A(\genblk1[5].osc.clkdiv_C.cnt[8] ),
    .B(\genblk1[5].osc.clkdiv_C.cnt[7] ),
    .C(_01705_),
    .X(_01708_));
 sky130_fd_sc_hd__a21oi_1 _06845_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[7] ),
    .A2(_01705_),
    .B1(\genblk1[5].osc.clkdiv_C.cnt[8] ),
    .Y(_01709_));
 sky130_fd_sc_hd__nor3_1 _06846_ (.A(_01693_),
    .B(_01708_),
    .C(_01709_),
    .Y(\genblk1[5].osc.clkdiv_C.next_cnt[8] ));
 sky130_fd_sc_hd__and2_1 _06847_ (.A(\genblk1[5].osc.clkdiv_C.cnt[9] ),
    .B(_01708_),
    .X(_01710_));
 sky130_fd_sc_hd__nor2_1 _06848_ (.A(\genblk1[5].osc.clkdiv_C.cnt[9] ),
    .B(_01708_),
    .Y(_01711_));
 sky130_fd_sc_hd__nor3_1 _06849_ (.A(_01693_),
    .B(_01710_),
    .C(_01711_),
    .Y(\genblk1[5].osc.clkdiv_C.next_cnt[9] ));
 sky130_fd_sc_hd__nand2_1 _06850_ (.A(\genblk1[5].osc.clkdiv_C.cnt[10] ),
    .B(_01710_),
    .Y(_01712_));
 sky130_fd_sc_hd__o211a_1 _06851_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[10] ),
    .A2(_01710_),
    .B1(_01712_),
    .C1(_01694_),
    .X(\genblk1[5].osc.clkdiv_C.next_cnt[10] ));
 sky130_fd_sc_hd__a21oi_1 _06852_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[10] ),
    .A2(_01710_),
    .B1(\genblk1[5].osc.clkdiv_C.cnt[11] ),
    .Y(_01713_));
 sky130_fd_sc_hd__and3_1 _06853_ (.A(\genblk1[5].osc.clkdiv_C.cnt[11] ),
    .B(\genblk1[5].osc.clkdiv_C.cnt[10] ),
    .C(_01710_),
    .X(_01714_));
 sky130_fd_sc_hd__nor3_1 _06854_ (.A(_01693_),
    .B(_01713_),
    .C(_01714_),
    .Y(\genblk1[5].osc.clkdiv_C.next_cnt[11] ));
 sky130_fd_sc_hd__and2_1 _06855_ (.A(\genblk1[5].osc.clkdiv_C.cnt[12] ),
    .B(_01714_),
    .X(_01715_));
 sky130_fd_sc_hd__nor2_1 _06856_ (.A(_01693_),
    .B(_01715_),
    .Y(_01716_));
 sky130_fd_sc_hd__o21a_1 _06857_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[12] ),
    .A2(_01714_),
    .B1(_01716_),
    .X(\genblk1[5].osc.clkdiv_C.next_cnt[12] ));
 sky130_fd_sc_hd__and3_1 _06858_ (.A(\genblk1[5].osc.clkdiv_C.cnt[13] ),
    .B(\genblk1[5].osc.clkdiv_C.cnt[12] ),
    .C(_01714_),
    .X(_01717_));
 sky130_fd_sc_hd__nor2_1 _06859_ (.A(_01693_),
    .B(_01717_),
    .Y(_01718_));
 sky130_fd_sc_hd__o21a_1 _06860_ (.A1(net1229),
    .A2(_01715_),
    .B1(_01718_),
    .X(\genblk1[5].osc.clkdiv_C.next_cnt[13] ));
 sky130_fd_sc_hd__and2_1 _06861_ (.A(\genblk1[5].osc.clkdiv_C.cnt[14] ),
    .B(_01717_),
    .X(_01719_));
 sky130_fd_sc_hd__nor2_1 _06862_ (.A(net27),
    .B(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__o21a_1 _06863_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[14] ),
    .A2(_01717_),
    .B1(_01720_),
    .X(\genblk1[5].osc.clkdiv_C.next_cnt[14] ));
 sky130_fd_sc_hd__and3_1 _06864_ (.A(\genblk1[5].osc.clkdiv_C.cnt[15] ),
    .B(\genblk1[5].osc.clkdiv_C.cnt[14] ),
    .C(_01717_),
    .X(_01721_));
 sky130_fd_sc_hd__nor2_1 _06865_ (.A(net27),
    .B(_01721_),
    .Y(_01722_));
 sky130_fd_sc_hd__o21a_1 _06866_ (.A1(net1115),
    .A2(_01719_),
    .B1(_01722_),
    .X(\genblk1[5].osc.clkdiv_C.next_cnt[15] ));
 sky130_fd_sc_hd__or2_1 _06867_ (.A(\genblk1[5].osc.clkdiv_C.cnt[16] ),
    .B(_01721_),
    .X(_01723_));
 sky130_fd_sc_hd__nand2_1 _06868_ (.A(\genblk1[5].osc.clkdiv_C.cnt[16] ),
    .B(_01721_),
    .Y(_01724_));
 sky130_fd_sc_hd__and3_1 _06869_ (.A(_01694_),
    .B(_01723_),
    .C(_01724_),
    .X(_01725_));
 sky130_fd_sc_hd__clkbuf_1 _06870_ (.A(_01725_),
    .X(\genblk1[5].osc.clkdiv_C.next_cnt[16] ));
 sky130_fd_sc_hd__xnor2_1 _06871_ (.A(net493),
    .B(_01724_),
    .Y(\genblk1[5].osc.clkdiv_C.next_cnt[17] ));
 sky130_fd_sc_hd__nor2_1 _06872_ (.A(_01441_),
    .B(_01366_),
    .Y(_01726_));
 sky130_fd_sc_hd__o21bai_1 _06873_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[10] ),
    .A2(_01726_),
    .B1_N(\genblk1[6].osc.clkdiv_C.cnt[14] ),
    .Y(_01727_));
 sky130_fd_sc_hd__xnor2_1 _06874_ (.A(\genblk1[6].osc.clkdiv_C.cnt[16] ),
    .B(_01578_),
    .Y(_01728_));
 sky130_fd_sc_hd__inv_2 _06875_ (.A(\genblk1[6].osc.clkdiv_C.cnt[2] ),
    .Y(_01729_));
 sky130_fd_sc_hd__or2_1 _06876_ (.A(_01336_),
    .B(net37),
    .X(_01730_));
 sky130_fd_sc_hd__nor2_1 _06877_ (.A(_01177_),
    .B(_01249_),
    .Y(_01731_));
 sky130_fd_sc_hd__buf_4 _06878_ (.A(_01731_),
    .X(_01732_));
 sky130_fd_sc_hd__a2bb2o_1 _06879_ (.A1_N(\genblk1[6].osc.clkdiv_C.cnt[4] ),
    .A2_N(_01730_),
    .B1(_01732_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[9] ),
    .X(_01733_));
 sky130_fd_sc_hd__a221o_1 _06880_ (.A1(_01729_),
    .A2(_01684_),
    .B1(_01730_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[4] ),
    .C1(_01733_),
    .X(_01734_));
 sky130_fd_sc_hd__or2_2 _06881_ (.A(_01189_),
    .B(_01678_),
    .X(_01735_));
 sky130_fd_sc_hd__a2bb2o_1 _06882_ (.A1_N(\genblk1[6].osc.clkdiv_C.cnt[9] ),
    .A2_N(_01732_),
    .B1(_01735_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[2] ),
    .X(_01736_));
 sky130_fd_sc_hd__a2111o_1 _06883_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[11] ),
    .A2(_01484_),
    .B1(_01728_),
    .C1(_01734_),
    .D1(_01736_),
    .X(_01737_));
 sky130_fd_sc_hd__nor2_2 _06884_ (.A(_01241_),
    .B(_01660_),
    .Y(_01738_));
 sky130_fd_sc_hd__and3_2 _06885_ (.A(_01349_),
    .B(_01209_),
    .C(_01439_),
    .X(_01739_));
 sky130_fd_sc_hd__o22a_1 _06886_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[1] ),
    .A2(_01738_),
    .B1(_01739_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[8] ),
    .X(_01740_));
 sky130_fd_sc_hd__a21bo_1 _06887_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[1] ),
    .A2(_01738_),
    .B1_N(_01740_),
    .X(_01741_));
 sky130_fd_sc_hd__nand2_2 _06888_ (.A(_01658_),
    .B(_01675_),
    .Y(_01742_));
 sky130_fd_sc_hd__a2bb2o_1 _06889_ (.A1_N(\genblk1[6].osc.clkdiv_C.cnt[12] ),
    .A2_N(_01519_),
    .B1(_01742_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[10] ),
    .X(_01743_));
 sky130_fd_sc_hd__a221o_1 _06890_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[12] ),
    .A2(_01519_),
    .B1(_01739_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[8] ),
    .C1(_01743_),
    .X(_01744_));
 sky130_fd_sc_hd__o2bb2a_1 _06891_ (.A1_N(\genblk1[6].osc.clkdiv_C.cnt[13] ),
    .A2_N(_01666_),
    .B1(_01484_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[11] ),
    .X(_01745_));
 sky130_fd_sc_hd__o221ai_2 _06892_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[14] ),
    .A2(_01675_),
    .B1(_01666_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[13] ),
    .C1(_01745_),
    .Y(_01746_));
 sky130_fd_sc_hd__nand2_2 _06893_ (.A(_01308_),
    .B(_01577_),
    .Y(_01747_));
 sky130_fd_sc_hd__xnor2_1 _06894_ (.A(\genblk1[6].osc.clkdiv_C.cnt[5] ),
    .B(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__nor2_1 _06895_ (.A(\genblk1[6].osc.clkdiv_C.cnt[15] ),
    .B(_01362_),
    .Y(_01749_));
 sky130_fd_sc_hd__nand2_2 _06896_ (.A(_01342_),
    .B(_01439_),
    .Y(_01750_));
 sky130_fd_sc_hd__o22ai_1 _06897_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[6] ),
    .A2(_01367_),
    .B1(_01750_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[0] ),
    .Y(_01751_));
 sky130_fd_sc_hd__a221o_1 _06898_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[6] ),
    .A2(_01367_),
    .B1(_01750_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[7] ),
    .C1(_01751_),
    .X(_01752_));
 sky130_fd_sc_hd__inv_2 _06899_ (.A(\genblk1[6].osc.clkdiv_C.cnt[7] ),
    .Y(_01753_));
 sky130_fd_sc_hd__a221o_1 _06900_ (.A1(_01753_),
    .A2(\genblk1[6].osc.clkdiv_C.cnt[0] ),
    .B1(_01363_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[15] ),
    .C1(\genblk1[6].osc.clkdiv_C.cnt[17] ),
    .X(_01754_));
 sky130_fd_sc_hd__or4_1 _06901_ (.A(_01748_),
    .B(_01749_),
    .C(_01752_),
    .D(_01754_),
    .X(_01755_));
 sky130_fd_sc_hd__or4_1 _06902_ (.A(_01741_),
    .B(_01744_),
    .C(_01746_),
    .D(_01755_),
    .X(_01756_));
 sky130_fd_sc_hd__nor2_2 _06903_ (.A(_01325_),
    .B(_01327_),
    .Y(_01757_));
 sky130_fd_sc_hd__nand2_2 _06904_ (.A(_01576_),
    .B(_01757_),
    .Y(_01758_));
 sky130_fd_sc_hd__xor2_1 _06905_ (.A(\genblk1[6].osc.clkdiv_C.cnt[3] ),
    .B(_01758_),
    .X(_01759_));
 sky130_fd_sc_hd__a2111oi_1 _06906_ (.A1(_01675_),
    .A2(_01727_),
    .B1(_01737_),
    .C1(_01756_),
    .D1(_01759_),
    .Y(_01760_));
 sky130_fd_sc_hd__clkbuf_4 _06907_ (.A(net28),
    .X(_01761_));
 sky130_fd_sc_hd__nor2_1 _06908_ (.A(net837),
    .B(_01761_),
    .Y(\genblk1[6].osc.clkdiv_C.next_cnt[0] ));
 sky130_fd_sc_hd__xnor2_1 _06909_ (.A(\genblk1[6].osc.clkdiv_C.cnt[1] ),
    .B(net837),
    .Y(_01762_));
 sky130_fd_sc_hd__nor2_1 _06910_ (.A(_01761_),
    .B(_01762_),
    .Y(\genblk1[6].osc.clkdiv_C.next_cnt[1] ));
 sky130_fd_sc_hd__and3_1 _06911_ (.A(\genblk1[6].osc.clkdiv_C.cnt[2] ),
    .B(\genblk1[6].osc.clkdiv_C.cnt[1] ),
    .C(\genblk1[6].osc.clkdiv_C.cnt[0] ),
    .X(_01763_));
 sky130_fd_sc_hd__a21oi_1 _06912_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[1] ),
    .A2(net837),
    .B1(\genblk1[6].osc.clkdiv_C.cnt[2] ),
    .Y(_01764_));
 sky130_fd_sc_hd__nor3_1 _06913_ (.A(_01761_),
    .B(_01763_),
    .C(_01764_),
    .Y(\genblk1[6].osc.clkdiv_C.next_cnt[2] ));
 sky130_fd_sc_hd__and2_1 _06914_ (.A(\genblk1[6].osc.clkdiv_C.cnt[3] ),
    .B(_01763_),
    .X(_01765_));
 sky130_fd_sc_hd__nor2_1 _06915_ (.A(\genblk1[6].osc.clkdiv_C.cnt[3] ),
    .B(_01763_),
    .Y(_01766_));
 sky130_fd_sc_hd__nor3_1 _06916_ (.A(_01761_),
    .B(_01765_),
    .C(_01766_),
    .Y(\genblk1[6].osc.clkdiv_C.next_cnt[3] ));
 sky130_fd_sc_hd__xnor2_1 _06917_ (.A(\genblk1[6].osc.clkdiv_C.cnt[4] ),
    .B(_01765_),
    .Y(_01767_));
 sky130_fd_sc_hd__nor2_1 _06918_ (.A(_01761_),
    .B(_01767_),
    .Y(\genblk1[6].osc.clkdiv_C.next_cnt[4] ));
 sky130_fd_sc_hd__and3_1 _06919_ (.A(\genblk1[6].osc.clkdiv_C.cnt[5] ),
    .B(\genblk1[6].osc.clkdiv_C.cnt[4] ),
    .C(_01765_),
    .X(_01768_));
 sky130_fd_sc_hd__a21oi_1 _06920_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[4] ),
    .A2(_01765_),
    .B1(\genblk1[6].osc.clkdiv_C.cnt[5] ),
    .Y(_01769_));
 sky130_fd_sc_hd__nor3_1 _06921_ (.A(_01761_),
    .B(_01768_),
    .C(_01769_),
    .Y(\genblk1[6].osc.clkdiv_C.next_cnt[5] ));
 sky130_fd_sc_hd__and2_1 _06922_ (.A(\genblk1[6].osc.clkdiv_C.cnt[6] ),
    .B(_01768_),
    .X(_01770_));
 sky130_fd_sc_hd__nor2_1 _06923_ (.A(\genblk1[6].osc.clkdiv_C.cnt[6] ),
    .B(_01768_),
    .Y(_01771_));
 sky130_fd_sc_hd__nor3_1 _06924_ (.A(_01761_),
    .B(_01770_),
    .C(_01771_),
    .Y(\genblk1[6].osc.clkdiv_C.next_cnt[6] ));
 sky130_fd_sc_hd__xnor2_1 _06925_ (.A(\genblk1[6].osc.clkdiv_C.cnt[7] ),
    .B(_01770_),
    .Y(_01772_));
 sky130_fd_sc_hd__nor2_1 _06926_ (.A(_01761_),
    .B(_01772_),
    .Y(\genblk1[6].osc.clkdiv_C.next_cnt[7] ));
 sky130_fd_sc_hd__and3_1 _06927_ (.A(\genblk1[6].osc.clkdiv_C.cnt[8] ),
    .B(\genblk1[6].osc.clkdiv_C.cnt[7] ),
    .C(_01770_),
    .X(_01773_));
 sky130_fd_sc_hd__a21oi_1 _06928_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[7] ),
    .A2(_01770_),
    .B1(\genblk1[6].osc.clkdiv_C.cnt[8] ),
    .Y(_01774_));
 sky130_fd_sc_hd__nor3_1 _06929_ (.A(_01761_),
    .B(_01773_),
    .C(_01774_),
    .Y(\genblk1[6].osc.clkdiv_C.next_cnt[8] ));
 sky130_fd_sc_hd__and2_1 _06930_ (.A(\genblk1[6].osc.clkdiv_C.cnt[9] ),
    .B(_01773_),
    .X(_01775_));
 sky130_fd_sc_hd__nor2_1 _06931_ (.A(\genblk1[6].osc.clkdiv_C.cnt[9] ),
    .B(_01773_),
    .Y(_01776_));
 sky130_fd_sc_hd__nor3_1 _06932_ (.A(_01761_),
    .B(_01775_),
    .C(_01776_),
    .Y(\genblk1[6].osc.clkdiv_C.next_cnt[9] ));
 sky130_fd_sc_hd__and3_1 _06933_ (.A(\genblk1[6].osc.clkdiv_C.cnt[10] ),
    .B(\genblk1[6].osc.clkdiv_C.cnt[9] ),
    .C(_01773_),
    .X(_01777_));
 sky130_fd_sc_hd__nor2_1 _06934_ (.A(net28),
    .B(_01777_),
    .Y(_01778_));
 sky130_fd_sc_hd__o21a_1 _06935_ (.A1(net1180),
    .A2(_01775_),
    .B1(_01778_),
    .X(\genblk1[6].osc.clkdiv_C.next_cnt[10] ));
 sky130_fd_sc_hd__and2_1 _06936_ (.A(\genblk1[6].osc.clkdiv_C.cnt[11] ),
    .B(_01777_),
    .X(_01779_));
 sky130_fd_sc_hd__nor2_1 _06937_ (.A(net28),
    .B(_01779_),
    .Y(_01780_));
 sky130_fd_sc_hd__o21a_1 _06938_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[11] ),
    .A2(_01777_),
    .B1(_01780_),
    .X(\genblk1[6].osc.clkdiv_C.next_cnt[11] ));
 sky130_fd_sc_hd__and3_1 _06939_ (.A(\genblk1[6].osc.clkdiv_C.cnt[12] ),
    .B(\genblk1[6].osc.clkdiv_C.cnt[11] ),
    .C(_01777_),
    .X(_01781_));
 sky130_fd_sc_hd__nor2_1 _06940_ (.A(net28),
    .B(_01781_),
    .Y(_01782_));
 sky130_fd_sc_hd__o21a_1 _06941_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[12] ),
    .A2(_01779_),
    .B1(_01782_),
    .X(\genblk1[6].osc.clkdiv_C.next_cnt[12] ));
 sky130_fd_sc_hd__and3_1 _06942_ (.A(\genblk1[6].osc.clkdiv_C.cnt[13] ),
    .B(\genblk1[6].osc.clkdiv_C.cnt[12] ),
    .C(_01779_),
    .X(_01783_));
 sky130_fd_sc_hd__nor2_1 _06943_ (.A(net28),
    .B(_01783_),
    .Y(_01784_));
 sky130_fd_sc_hd__o21a_1 _06944_ (.A1(net1146),
    .A2(_01781_),
    .B1(_01784_),
    .X(\genblk1[6].osc.clkdiv_C.next_cnt[13] ));
 sky130_fd_sc_hd__and2_1 _06945_ (.A(\genblk1[6].osc.clkdiv_C.cnt[14] ),
    .B(_01783_),
    .X(_01785_));
 sky130_fd_sc_hd__nor2_1 _06946_ (.A(net1356),
    .B(_01785_),
    .Y(_01786_));
 sky130_fd_sc_hd__o21a_1 _06947_ (.A1(net1104),
    .A2(_01783_),
    .B1(_01786_),
    .X(\genblk1[6].osc.clkdiv_C.next_cnt[14] ));
 sky130_fd_sc_hd__and3_1 _06948_ (.A(\genblk1[6].osc.clkdiv_C.cnt[15] ),
    .B(\genblk1[6].osc.clkdiv_C.cnt[14] ),
    .C(_01783_),
    .X(_01787_));
 sky130_fd_sc_hd__nor2_1 _06949_ (.A(net1356),
    .B(_01787_),
    .Y(_01788_));
 sky130_fd_sc_hd__o21a_1 _06950_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[15] ),
    .A2(_01785_),
    .B1(_01788_),
    .X(\genblk1[6].osc.clkdiv_C.next_cnt[15] ));
 sky130_fd_sc_hd__or2_1 _06951_ (.A(\genblk1[6].osc.clkdiv_C.cnt[16] ),
    .B(_01787_),
    .X(_01789_));
 sky130_fd_sc_hd__nand2_1 _06952_ (.A(\genblk1[6].osc.clkdiv_C.cnt[16] ),
    .B(_01787_),
    .Y(_01790_));
 sky130_fd_sc_hd__and3b_1 _06953_ (.A_N(_01760_),
    .B(_01789_),
    .C(_01790_),
    .X(_01791_));
 sky130_fd_sc_hd__clkbuf_1 _06954_ (.A(_01791_),
    .X(\genblk1[6].osc.clkdiv_C.next_cnt[16] ));
 sky130_fd_sc_hd__xnor2_1 _06955_ (.A(net1063),
    .B(_01790_),
    .Y(\genblk1[6].osc.clkdiv_C.next_cnt[17] ));
 sky130_fd_sc_hd__o22ai_1 _06956_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[11] ),
    .A2(_01311_),
    .B1(_01732_),
    .B2(\genblk1[7].osc.clkdiv_C.cnt[3] ),
    .Y(_01792_));
 sky130_fd_sc_hd__a221oi_1 _06957_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[2] ),
    .A2(_01227_),
    .B1(_01732_),
    .B2(\genblk1[7].osc.clkdiv_C.cnt[3] ),
    .C1(_01792_),
    .Y(_01793_));
 sky130_fd_sc_hd__a21oi_4 _06958_ (.A1(_01228_),
    .A2(_01220_),
    .B1(_01233_),
    .Y(_01794_));
 sky130_fd_sc_hd__and3b_1 _06959_ (.A_N(\genblk1[7].osc.clkdiv_C.cnt[0] ),
    .B(net34),
    .C(\genblk1[7].osc.clkdiv_C.cnt[10] ),
    .X(_01795_));
 sky130_fd_sc_hd__and3b_1 _06960_ (.A_N(\genblk1[7].osc.clkdiv_C.cnt[10] ),
    .B(\genblk1[7].osc.clkdiv_C.cnt[0] ),
    .C(_01514_),
    .X(_01796_));
 sky130_fd_sc_hd__nand2_2 _06961_ (.A(_01432_),
    .B(_01221_),
    .Y(_01797_));
 sky130_fd_sc_hd__xnor2_1 _06962_ (.A(\genblk1[7].osc.clkdiv_C.cnt[9] ),
    .B(_01797_),
    .Y(_01798_));
 sky130_fd_sc_hd__a21oi_4 _06963_ (.A1(_01229_),
    .A2(_01230_),
    .B1(_01238_),
    .Y(_01799_));
 sky130_fd_sc_hd__xnor2_1 _06964_ (.A(\genblk1[7].osc.clkdiv_C.cnt[4] ),
    .B(_01799_),
    .Y(_01800_));
 sky130_fd_sc_hd__nand2_2 _06965_ (.A(_01213_),
    .B(_01344_),
    .Y(_01801_));
 sky130_fd_sc_hd__nand2_1 _06966_ (.A(_01192_),
    .B(_01245_),
    .Y(_01802_));
 sky130_fd_sc_hd__a22o_1 _06967_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[7] ),
    .A2(_01574_),
    .B1(_01802_),
    .B2(\genblk1[7].osc.clkdiv_C.cnt[6] ),
    .X(_01803_));
 sky130_fd_sc_hd__a21oi_1 _06968_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[1] ),
    .A2(_01801_),
    .B1(_01803_),
    .Y(_01804_));
 sky130_fd_sc_hd__or2_2 _06969_ (.A(_01179_),
    .B(_01233_),
    .X(_01805_));
 sky130_fd_sc_hd__o2bb2a_1 _06970_ (.A1_N(\genblk1[7].osc.clkdiv_C.cnt[5] ),
    .A2_N(_01805_),
    .B1(_01801_),
    .B2(\genblk1[7].osc.clkdiv_C.cnt[1] ),
    .X(_01806_));
 sky130_fd_sc_hd__o221a_1 _06971_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[6] ),
    .A2(_01802_),
    .B1(_01805_),
    .B2(\genblk1[7].osc.clkdiv_C.cnt[5] ),
    .C1(_01806_),
    .X(_01807_));
 sky130_fd_sc_hd__xnor2_1 _06972_ (.A(\genblk1[7].osc.clkdiv_C.cnt[13] ),
    .B(_01214_),
    .Y(_01808_));
 sky130_fd_sc_hd__a221o_1 _06973_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[15] ),
    .A2(_01363_),
    .B1(_01311_),
    .B2(\genblk1[7].osc.clkdiv_C.cnt[11] ),
    .C1(_01808_),
    .X(_01809_));
 sky130_fd_sc_hd__xor2_1 _06974_ (.A(\genblk1[7].osc.clkdiv_C.cnt[14] ),
    .B(_01675_),
    .X(_01810_));
 sky130_fd_sc_hd__nor2_4 _06975_ (.A(_01365_),
    .B(_01355_),
    .Y(_01811_));
 sky130_fd_sc_hd__xnor2_1 _06976_ (.A(\genblk1[7].osc.clkdiv_C.cnt[12] ),
    .B(_01811_),
    .Y(_01812_));
 sky130_fd_sc_hd__inv_2 _06977_ (.A(\genblk1[7].osc.clkdiv_C.cnt[16] ),
    .Y(_01813_));
 sky130_fd_sc_hd__inv_2 _06978_ (.A(\genblk1[7].osc.clkdiv_C.cnt[17] ),
    .Y(_01814_));
 sky130_fd_sc_hd__o221a_1 _06979_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[15] ),
    .A2(_01363_),
    .B1(_01196_),
    .B2(_01813_),
    .C1(_01814_),
    .X(_01815_));
 sky130_fd_sc_hd__o221a_1 _06980_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[16] ),
    .A2(_01578_),
    .B1(_01574_),
    .B2(\genblk1[7].osc.clkdiv_C.cnt[7] ),
    .C1(_01815_),
    .X(_01816_));
 sky130_fd_sc_hd__and4b_1 _06981_ (.A_N(_01809_),
    .B(_01810_),
    .C(_01812_),
    .D(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__and4_1 _06982_ (.A(_01800_),
    .B(_01804_),
    .C(_01807_),
    .D(_01817_),
    .X(_01818_));
 sky130_fd_sc_hd__nand2_2 _06983_ (.A(_01436_),
    .B(_01334_),
    .Y(_01819_));
 sky130_fd_sc_hd__xnor2_1 _06984_ (.A(\genblk1[7].osc.clkdiv_C.cnt[8] ),
    .B(_01819_),
    .Y(_01820_));
 sky130_fd_sc_hd__o2111a_1 _06985_ (.A1(_01795_),
    .A2(_01796_),
    .B1(_01798_),
    .C1(_01818_),
    .D1(_01820_),
    .X(_01821_));
 sky130_fd_sc_hd__o211a_2 _06986_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[2] ),
    .A2(_01227_),
    .B1(_01793_),
    .C1(_01821_),
    .X(_01822_));
 sky130_fd_sc_hd__clkbuf_4 _06987_ (.A(_01822_),
    .X(_01823_));
 sky130_fd_sc_hd__nor2_1 _06988_ (.A(net1058),
    .B(_01823_),
    .Y(\genblk1[7].osc.clkdiv_C.next_cnt[0] ));
 sky130_fd_sc_hd__xnor2_1 _06989_ (.A(\genblk1[7].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[7].osc.clkdiv_C.cnt[0] ),
    .Y(_01824_));
 sky130_fd_sc_hd__nor2_1 _06990_ (.A(_01823_),
    .B(_01824_),
    .Y(\genblk1[7].osc.clkdiv_C.next_cnt[1] ));
 sky130_fd_sc_hd__and3_1 _06991_ (.A(\genblk1[7].osc.clkdiv_C.cnt[2] ),
    .B(\genblk1[7].osc.clkdiv_C.cnt[1] ),
    .C(\genblk1[7].osc.clkdiv_C.cnt[0] ),
    .X(_01825_));
 sky130_fd_sc_hd__a21oi_1 _06992_ (.A1(net1252),
    .A2(net1058),
    .B1(\genblk1[7].osc.clkdiv_C.cnt[2] ),
    .Y(_01826_));
 sky130_fd_sc_hd__nor3_1 _06993_ (.A(_01823_),
    .B(_01825_),
    .C(_01826_),
    .Y(\genblk1[7].osc.clkdiv_C.next_cnt[2] ));
 sky130_fd_sc_hd__and2_1 _06994_ (.A(\genblk1[7].osc.clkdiv_C.cnt[3] ),
    .B(_01825_),
    .X(_01827_));
 sky130_fd_sc_hd__nor2_1 _06995_ (.A(\genblk1[7].osc.clkdiv_C.cnt[3] ),
    .B(_01825_),
    .Y(_01828_));
 sky130_fd_sc_hd__nor3_1 _06996_ (.A(_01823_),
    .B(_01827_),
    .C(_01828_),
    .Y(\genblk1[7].osc.clkdiv_C.next_cnt[3] ));
 sky130_fd_sc_hd__xnor2_1 _06997_ (.A(\genblk1[7].osc.clkdiv_C.cnt[4] ),
    .B(_01827_),
    .Y(_01829_));
 sky130_fd_sc_hd__nor2_1 _06998_ (.A(_01823_),
    .B(_01829_),
    .Y(\genblk1[7].osc.clkdiv_C.next_cnt[4] ));
 sky130_fd_sc_hd__and3_1 _06999_ (.A(\genblk1[7].osc.clkdiv_C.cnt[5] ),
    .B(\genblk1[7].osc.clkdiv_C.cnt[4] ),
    .C(_01827_),
    .X(_01830_));
 sky130_fd_sc_hd__a21oi_1 _07000_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[4] ),
    .A2(_01827_),
    .B1(\genblk1[7].osc.clkdiv_C.cnt[5] ),
    .Y(_01831_));
 sky130_fd_sc_hd__nor3_1 _07001_ (.A(_01823_),
    .B(_01830_),
    .C(_01831_),
    .Y(\genblk1[7].osc.clkdiv_C.next_cnt[5] ));
 sky130_fd_sc_hd__and2_1 _07002_ (.A(\genblk1[7].osc.clkdiv_C.cnt[6] ),
    .B(_01830_),
    .X(_01832_));
 sky130_fd_sc_hd__nor2_1 _07003_ (.A(\genblk1[7].osc.clkdiv_C.cnt[6] ),
    .B(_01830_),
    .Y(_01833_));
 sky130_fd_sc_hd__nor3_1 _07004_ (.A(_01823_),
    .B(_01832_),
    .C(_01833_),
    .Y(\genblk1[7].osc.clkdiv_C.next_cnt[6] ));
 sky130_fd_sc_hd__xnor2_1 _07005_ (.A(\genblk1[7].osc.clkdiv_C.cnt[7] ),
    .B(_01832_),
    .Y(_01834_));
 sky130_fd_sc_hd__nor2_1 _07006_ (.A(_01823_),
    .B(_01834_),
    .Y(\genblk1[7].osc.clkdiv_C.next_cnt[7] ));
 sky130_fd_sc_hd__and3_1 _07007_ (.A(\genblk1[7].osc.clkdiv_C.cnt[8] ),
    .B(\genblk1[7].osc.clkdiv_C.cnt[7] ),
    .C(_01832_),
    .X(_01835_));
 sky130_fd_sc_hd__a21oi_1 _07008_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[7] ),
    .A2(_01832_),
    .B1(\genblk1[7].osc.clkdiv_C.cnt[8] ),
    .Y(_01836_));
 sky130_fd_sc_hd__nor3_1 _07009_ (.A(_01823_),
    .B(_01835_),
    .C(_01836_),
    .Y(\genblk1[7].osc.clkdiv_C.next_cnt[8] ));
 sky130_fd_sc_hd__and2_1 _07010_ (.A(\genblk1[7].osc.clkdiv_C.cnt[9] ),
    .B(_01835_),
    .X(_01837_));
 sky130_fd_sc_hd__nor2_1 _07011_ (.A(\genblk1[7].osc.clkdiv_C.cnt[9] ),
    .B(_01835_),
    .Y(_01838_));
 sky130_fd_sc_hd__nor3_1 _07012_ (.A(_01823_),
    .B(_01837_),
    .C(_01838_),
    .Y(\genblk1[7].osc.clkdiv_C.next_cnt[9] ));
 sky130_fd_sc_hd__a21oi_1 _07013_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[10] ),
    .A2(_01837_),
    .B1(_01822_),
    .Y(_01839_));
 sky130_fd_sc_hd__o21a_1 _07014_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[10] ),
    .A2(_01837_),
    .B1(_01839_),
    .X(\genblk1[7].osc.clkdiv_C.next_cnt[10] ));
 sky130_fd_sc_hd__a21oi_1 _07015_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[10] ),
    .A2(_01837_),
    .B1(\genblk1[7].osc.clkdiv_C.cnt[11] ),
    .Y(_01840_));
 sky130_fd_sc_hd__and3_1 _07016_ (.A(\genblk1[7].osc.clkdiv_C.cnt[11] ),
    .B(\genblk1[7].osc.clkdiv_C.cnt[10] ),
    .C(_01837_),
    .X(_01841_));
 sky130_fd_sc_hd__nor3_1 _07017_ (.A(_01822_),
    .B(_01840_),
    .C(_01841_),
    .Y(\genblk1[7].osc.clkdiv_C.next_cnt[11] ));
 sky130_fd_sc_hd__and2_1 _07018_ (.A(\genblk1[7].osc.clkdiv_C.cnt[12] ),
    .B(_01841_),
    .X(_01842_));
 sky130_fd_sc_hd__nor2_1 _07019_ (.A(_01822_),
    .B(_01842_),
    .Y(_01843_));
 sky130_fd_sc_hd__o21a_1 _07020_ (.A1(net1189),
    .A2(_01841_),
    .B1(_01843_),
    .X(\genblk1[7].osc.clkdiv_C.next_cnt[12] ));
 sky130_fd_sc_hd__a21oi_1 _07021_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[13] ),
    .A2(_01842_),
    .B1(_01822_),
    .Y(_01844_));
 sky130_fd_sc_hd__o21a_1 _07022_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[13] ),
    .A2(_01842_),
    .B1(_01844_),
    .X(\genblk1[7].osc.clkdiv_C.next_cnt[13] ));
 sky130_fd_sc_hd__a21oi_1 _07023_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[13] ),
    .A2(_01842_),
    .B1(\genblk1[7].osc.clkdiv_C.cnt[14] ),
    .Y(_01845_));
 sky130_fd_sc_hd__and3_1 _07024_ (.A(\genblk1[7].osc.clkdiv_C.cnt[14] ),
    .B(\genblk1[7].osc.clkdiv_C.cnt[13] ),
    .C(_01842_),
    .X(_01846_));
 sky130_fd_sc_hd__nor3_1 _07025_ (.A(_01822_),
    .B(_01845_),
    .C(_01846_),
    .Y(\genblk1[7].osc.clkdiv_C.next_cnt[14] ));
 sky130_fd_sc_hd__and2_1 _07026_ (.A(\genblk1[7].osc.clkdiv_C.cnt[15] ),
    .B(_01846_),
    .X(_01847_));
 sky130_fd_sc_hd__nor2_1 _07027_ (.A(_01822_),
    .B(_01847_),
    .Y(_01848_));
 sky130_fd_sc_hd__o21a_1 _07028_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[15] ),
    .A2(_01846_),
    .B1(_01848_),
    .X(\genblk1[7].osc.clkdiv_C.next_cnt[15] ));
 sky130_fd_sc_hd__or2_1 _07029_ (.A(\genblk1[7].osc.clkdiv_C.cnt[16] ),
    .B(_01847_),
    .X(_01849_));
 sky130_fd_sc_hd__nand2_1 _07030_ (.A(\genblk1[7].osc.clkdiv_C.cnt[16] ),
    .B(_01847_),
    .Y(_01850_));
 sky130_fd_sc_hd__and3b_1 _07031_ (.A_N(_01822_),
    .B(_01849_),
    .C(_01850_),
    .X(_01851_));
 sky130_fd_sc_hd__clkbuf_1 _07032_ (.A(_01851_),
    .X(\genblk1[7].osc.clkdiv_C.next_cnt[16] ));
 sky130_fd_sc_hd__xnor2_1 _07033_ (.A(net848),
    .B(_01850_),
    .Y(\genblk1[7].osc.clkdiv_C.next_cnt[17] ));
 sky130_fd_sc_hd__or2_1 _07034_ (.A(\genblk1[8].osc.clkdiv_C.cnt[15] ),
    .B(_01359_),
    .X(_01852_));
 sky130_fd_sc_hd__a21oi_1 _07035_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[10] ),
    .A2(_01852_),
    .B1(_01248_),
    .Y(_01853_));
 sky130_fd_sc_hd__o21a_1 _07036_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[16] ),
    .A2(_01853_),
    .B1(_01578_),
    .X(_01854_));
 sky130_fd_sc_hd__nand2_4 _07037_ (.A(_01230_),
    .B(_01564_),
    .Y(_01855_));
 sky130_fd_sc_hd__a21oi_1 _07038_ (.A1(_01436_),
    .A2(_01855_),
    .B1(\genblk1[8].osc.clkdiv_C.cnt[1] ),
    .Y(_01856_));
 sky130_fd_sc_hd__nor2_1 _07039_ (.A(\genblk1[8].osc.clkdiv_C.cnt[5] ),
    .B(_01487_),
    .Y(_01857_));
 sky130_fd_sc_hd__nand2_4 _07040_ (.A(_01489_),
    .B(_01344_),
    .Y(_01858_));
 sky130_fd_sc_hd__nand2_2 _07041_ (.A(_01439_),
    .B(_01576_),
    .Y(_01859_));
 sky130_fd_sc_hd__a32o_1 _07042_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[1] ),
    .A2(_01436_),
    .A3(_01855_),
    .B1(_01859_),
    .B2(\genblk1[8].osc.clkdiv_C.cnt[10] ),
    .X(_01860_));
 sky130_fd_sc_hd__a221o_1 _07043_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[5] ),
    .A2(_01487_),
    .B1(_01858_),
    .B2(\genblk1[8].osc.clkdiv_C.cnt[6] ),
    .C1(_01860_),
    .X(_01861_));
 sky130_fd_sc_hd__or4_1 _07044_ (.A(_01854_),
    .B(_01856_),
    .C(_01857_),
    .D(_01861_),
    .X(_01862_));
 sky130_fd_sc_hd__and2_1 _07045_ (.A(\genblk1[8].osc.clkdiv_C.cnt[8] ),
    .B(_01430_),
    .X(_01863_));
 sky130_fd_sc_hd__xnor2_1 _07046_ (.A(\genblk1[8].osc.clkdiv_C.cnt[13] ),
    .B(_01328_),
    .Y(_01864_));
 sky130_fd_sc_hd__or2_2 _07047_ (.A(_01336_),
    .B(_01223_),
    .X(_01865_));
 sky130_fd_sc_hd__a21oi_2 _07048_ (.A1(_01174_),
    .A2(_01182_),
    .B1(_01336_),
    .Y(_01866_));
 sky130_fd_sc_hd__o22a_1 _07049_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[4] ),
    .A2(_01866_),
    .B1(_01865_),
    .B2(\genblk1[8].osc.clkdiv_C.cnt[9] ),
    .X(_01867_));
 sky130_fd_sc_hd__a21bo_1 _07050_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[9] ),
    .A2(_01865_),
    .B1_N(_01867_),
    .X(_01868_));
 sky130_fd_sc_hd__nor2_2 _07051_ (.A(_01336_),
    .B(_01183_),
    .Y(_01869_));
 sky130_fd_sc_hd__nor2_4 _07052_ (.A(_01441_),
    .B(_01226_),
    .Y(_01870_));
 sky130_fd_sc_hd__a2bb2o_1 _07053_ (.A1_N(\genblk1[8].osc.clkdiv_C.cnt[12] ),
    .A2_N(_01869_),
    .B1(_01870_),
    .B2(\genblk1[8].osc.clkdiv_C.cnt[11] ),
    .X(_01871_));
 sky130_fd_sc_hd__a2111o_1 _07054_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[15] ),
    .A2(_01436_),
    .B1(_01864_),
    .C1(_01868_),
    .D1(_01871_),
    .X(_01872_));
 sky130_fd_sc_hd__nor2_1 _07055_ (.A(\genblk1[8].osc.clkdiv_C.cnt[8] ),
    .B(_01430_),
    .Y(_01873_));
 sky130_fd_sc_hd__xnor2_1 _07056_ (.A(\genblk1[8].osc.clkdiv_C.cnt[3] ),
    .B(_01498_),
    .Y(_01874_));
 sky130_fd_sc_hd__o21bai_1 _07057_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[14] ),
    .A2(_01246_),
    .B1_N(\genblk1[8].osc.clkdiv_C.cnt[17] ),
    .Y(_01875_));
 sky130_fd_sc_hd__a221o_1 _07058_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[0] ),
    .A2(_01211_),
    .B1(_01246_),
    .B2(\genblk1[8].osc.clkdiv_C.cnt[14] ),
    .C1(_01875_),
    .X(_01876_));
 sky130_fd_sc_hd__a22o_1 _07059_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[4] ),
    .A2(_01866_),
    .B1(_01869_),
    .B2(\genblk1[8].osc.clkdiv_C.cnt[12] ),
    .X(_01877_));
 sky130_fd_sc_hd__inv_2 _07060_ (.A(\genblk1[8].osc.clkdiv_C.cnt[7] ),
    .Y(_01878_));
 sky130_fd_sc_hd__inv_2 _07061_ (.A(\genblk1[8].osc.clkdiv_C.cnt[2] ),
    .Y(_01879_));
 sky130_fd_sc_hd__o2111a_1 _07062_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[6] ),
    .A2(_01249_),
    .B1(_01879_),
    .C1(_01490_),
    .D1(\genblk1[8].osc.clkdiv_C.cnt[7] ),
    .X(_01880_));
 sky130_fd_sc_hd__a31o_1 _07063_ (.A1(_01441_),
    .A2(_01878_),
    .A3(\genblk1[8].osc.clkdiv_C.cnt[2] ),
    .B1(_01880_),
    .X(_01881_));
 sky130_fd_sc_hd__or4b_1 _07064_ (.A(_01874_),
    .B(_01876_),
    .C(_01877_),
    .D_N(_01881_),
    .X(_01882_));
 sky130_fd_sc_hd__o21ba_1 _07065_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[0] ),
    .A2(_01211_),
    .B1_N(_01882_),
    .X(_01883_));
 sky130_fd_sc_hd__o221a_1 _07066_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[16] ),
    .A2(_01578_),
    .B1(_01870_),
    .B2(\genblk1[8].osc.clkdiv_C.cnt[11] ),
    .C1(_01883_),
    .X(_01884_));
 sky130_fd_sc_hd__or4b_1 _07067_ (.A(_01863_),
    .B(_01872_),
    .C(_01873_),
    .D_N(_01884_),
    .X(_01885_));
 sky130_fd_sc_hd__nor2_2 _07068_ (.A(_01862_),
    .B(_01885_),
    .Y(_01886_));
 sky130_fd_sc_hd__clkbuf_4 _07069_ (.A(_01886_),
    .X(_01887_));
 sky130_fd_sc_hd__nor2_1 _07070_ (.A(net1092),
    .B(_01887_),
    .Y(\genblk1[8].osc.clkdiv_C.next_cnt[0] ));
 sky130_fd_sc_hd__or2_1 _07071_ (.A(\genblk1[8].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[8].osc.clkdiv_C.cnt[0] ),
    .X(_01888_));
 sky130_fd_sc_hd__nand2_2 _07072_ (.A(\genblk1[8].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[8].osc.clkdiv_C.cnt[0] ),
    .Y(_01889_));
 sky130_fd_sc_hd__o211a_1 _07073_ (.A1(_01862_),
    .A2(_01885_),
    .B1(_01888_),
    .C1(_01889_),
    .X(\genblk1[8].osc.clkdiv_C.next_cnt[1] ));
 sky130_fd_sc_hd__nor2_1 _07074_ (.A(_01879_),
    .B(_01889_),
    .Y(_01890_));
 sky130_fd_sc_hd__and2_1 _07075_ (.A(_01879_),
    .B(_01889_),
    .X(_01891_));
 sky130_fd_sc_hd__nor3_1 _07076_ (.A(_01887_),
    .B(_01890_),
    .C(_01891_),
    .Y(\genblk1[8].osc.clkdiv_C.next_cnt[2] ));
 sky130_fd_sc_hd__and2_1 _07077_ (.A(\genblk1[8].osc.clkdiv_C.cnt[3] ),
    .B(_01890_),
    .X(_01892_));
 sky130_fd_sc_hd__nor2_1 _07078_ (.A(\genblk1[8].osc.clkdiv_C.cnt[3] ),
    .B(_01890_),
    .Y(_01893_));
 sky130_fd_sc_hd__nor3_1 _07079_ (.A(_01887_),
    .B(_01892_),
    .C(_01893_),
    .Y(\genblk1[8].osc.clkdiv_C.next_cnt[3] ));
 sky130_fd_sc_hd__o21bai_1 _07080_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[4] ),
    .A2(_01892_),
    .B1_N(_01886_),
    .Y(_01894_));
 sky130_fd_sc_hd__a21oi_1 _07081_ (.A1(net1162),
    .A2(_01892_),
    .B1(_01894_),
    .Y(\genblk1[8].osc.clkdiv_C.next_cnt[4] ));
 sky130_fd_sc_hd__and3_1 _07082_ (.A(\genblk1[8].osc.clkdiv_C.cnt[5] ),
    .B(\genblk1[8].osc.clkdiv_C.cnt[4] ),
    .C(_01892_),
    .X(_01895_));
 sky130_fd_sc_hd__a21oi_1 _07083_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[4] ),
    .A2(_01892_),
    .B1(\genblk1[8].osc.clkdiv_C.cnt[5] ),
    .Y(_01896_));
 sky130_fd_sc_hd__nor3_1 _07084_ (.A(_01887_),
    .B(_01895_),
    .C(_01896_),
    .Y(\genblk1[8].osc.clkdiv_C.next_cnt[5] ));
 sky130_fd_sc_hd__and2_1 _07085_ (.A(\genblk1[8].osc.clkdiv_C.cnt[6] ),
    .B(_01895_),
    .X(_01897_));
 sky130_fd_sc_hd__nor2_1 _07086_ (.A(\genblk1[8].osc.clkdiv_C.cnt[6] ),
    .B(_01895_),
    .Y(_01898_));
 sky130_fd_sc_hd__nor3_1 _07087_ (.A(_01887_),
    .B(_01897_),
    .C(_01898_),
    .Y(\genblk1[8].osc.clkdiv_C.next_cnt[6] ));
 sky130_fd_sc_hd__o21bai_1 _07088_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[7] ),
    .A2(_01897_),
    .B1_N(_01886_),
    .Y(_01899_));
 sky130_fd_sc_hd__a21oi_1 _07089_ (.A1(net1185),
    .A2(_01897_),
    .B1(_01899_),
    .Y(\genblk1[8].osc.clkdiv_C.next_cnt[7] ));
 sky130_fd_sc_hd__and3_1 _07090_ (.A(\genblk1[8].osc.clkdiv_C.cnt[8] ),
    .B(\genblk1[8].osc.clkdiv_C.cnt[7] ),
    .C(_01897_),
    .X(_01900_));
 sky130_fd_sc_hd__a21oi_1 _07091_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[7] ),
    .A2(_01897_),
    .B1(\genblk1[8].osc.clkdiv_C.cnt[8] ),
    .Y(_01901_));
 sky130_fd_sc_hd__nor3_1 _07092_ (.A(_01887_),
    .B(_01900_),
    .C(_01901_),
    .Y(\genblk1[8].osc.clkdiv_C.next_cnt[8] ));
 sky130_fd_sc_hd__and2_1 _07093_ (.A(\genblk1[8].osc.clkdiv_C.cnt[9] ),
    .B(_01900_),
    .X(_01902_));
 sky130_fd_sc_hd__nor2_1 _07094_ (.A(\genblk1[8].osc.clkdiv_C.cnt[9] ),
    .B(_01900_),
    .Y(_01903_));
 sky130_fd_sc_hd__nor3_1 _07095_ (.A(_01887_),
    .B(_01902_),
    .C(_01903_),
    .Y(\genblk1[8].osc.clkdiv_C.next_cnt[9] ));
 sky130_fd_sc_hd__and3_1 _07096_ (.A(\genblk1[8].osc.clkdiv_C.cnt[10] ),
    .B(\genblk1[8].osc.clkdiv_C.cnt[9] ),
    .C(_01900_),
    .X(_01904_));
 sky130_fd_sc_hd__nor2_1 _07097_ (.A(_01887_),
    .B(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__o21a_1 _07098_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[10] ),
    .A2(_01902_),
    .B1(_01905_),
    .X(\genblk1[8].osc.clkdiv_C.next_cnt[10] ));
 sky130_fd_sc_hd__and2_1 _07099_ (.A(\genblk1[8].osc.clkdiv_C.cnt[11] ),
    .B(_01904_),
    .X(_01906_));
 sky130_fd_sc_hd__nor2_1 _07100_ (.A(_01887_),
    .B(_01906_),
    .Y(_01907_));
 sky130_fd_sc_hd__o21a_1 _07101_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[11] ),
    .A2(_01904_),
    .B1(_01907_),
    .X(\genblk1[8].osc.clkdiv_C.next_cnt[11] ));
 sky130_fd_sc_hd__and3_1 _07102_ (.A(\genblk1[8].osc.clkdiv_C.cnt[12] ),
    .B(\genblk1[8].osc.clkdiv_C.cnt[11] ),
    .C(_01904_),
    .X(_01908_));
 sky130_fd_sc_hd__nor2_1 _07103_ (.A(_01887_),
    .B(_01908_),
    .Y(_01909_));
 sky130_fd_sc_hd__o21a_1 _07104_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[12] ),
    .A2(_01906_),
    .B1(_01909_),
    .X(\genblk1[8].osc.clkdiv_C.next_cnt[12] ));
 sky130_fd_sc_hd__and3_1 _07105_ (.A(\genblk1[8].osc.clkdiv_C.cnt[13] ),
    .B(\genblk1[8].osc.clkdiv_C.cnt[12] ),
    .C(_01906_),
    .X(_01910_));
 sky130_fd_sc_hd__nor2_1 _07106_ (.A(_01886_),
    .B(_01910_),
    .Y(_01911_));
 sky130_fd_sc_hd__o21a_1 _07107_ (.A1(net1182),
    .A2(_01908_),
    .B1(_01911_),
    .X(\genblk1[8].osc.clkdiv_C.next_cnt[13] ));
 sky130_fd_sc_hd__and2_1 _07108_ (.A(\genblk1[8].osc.clkdiv_C.cnt[14] ),
    .B(_01910_),
    .X(_01912_));
 sky130_fd_sc_hd__nor2_1 _07109_ (.A(_01886_),
    .B(_01912_),
    .Y(_01913_));
 sky130_fd_sc_hd__o21a_1 _07110_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[14] ),
    .A2(_01910_),
    .B1(_01913_),
    .X(\genblk1[8].osc.clkdiv_C.next_cnt[14] ));
 sky130_fd_sc_hd__and3_1 _07111_ (.A(\genblk1[8].osc.clkdiv_C.cnt[15] ),
    .B(\genblk1[8].osc.clkdiv_C.cnt[14] ),
    .C(_01910_),
    .X(_01914_));
 sky130_fd_sc_hd__nor2_1 _07112_ (.A(_01886_),
    .B(_01914_),
    .Y(_01915_));
 sky130_fd_sc_hd__o21a_1 _07113_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[15] ),
    .A2(_01912_),
    .B1(_01915_),
    .X(\genblk1[8].osc.clkdiv_C.next_cnt[15] ));
 sky130_fd_sc_hd__or2_1 _07114_ (.A(\genblk1[8].osc.clkdiv_C.cnt[16] ),
    .B(_01914_),
    .X(_01916_));
 sky130_fd_sc_hd__nand2_1 _07115_ (.A(\genblk1[8].osc.clkdiv_C.cnt[16] ),
    .B(_01914_),
    .Y(_01917_));
 sky130_fd_sc_hd__and3b_1 _07116_ (.A_N(_01886_),
    .B(_01916_),
    .C(_01917_),
    .X(_01918_));
 sky130_fd_sc_hd__clkbuf_1 _07117_ (.A(_01918_),
    .X(\genblk1[8].osc.clkdiv_C.next_cnt[16] ));
 sky130_fd_sc_hd__xnor2_1 _07118_ (.A(net691),
    .B(_01917_),
    .Y(\genblk1[8].osc.clkdiv_C.next_cnt[17] ));
 sky130_fd_sc_hd__xnor2_1 _07119_ (.A(\genblk1[9].osc.clkdiv_C.cnt[10] ),
    .B(_01227_),
    .Y(_01919_));
 sky130_fd_sc_hd__and2_1 _07120_ (.A(_01432_),
    .B(_01221_),
    .X(_01920_));
 sky130_fd_sc_hd__o22a_1 _07121_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[2] ),
    .A2(_01920_),
    .B1(_01855_),
    .B2(\genblk1[9].osc.clkdiv_C.cnt[0] ),
    .X(_01921_));
 sky130_fd_sc_hd__o221a_1 _07122_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[6] ),
    .A2(_01334_),
    .B1(_01328_),
    .B2(\genblk1[9].osc.clkdiv_C.cnt[13] ),
    .C1(_01921_),
    .X(_01922_));
 sky130_fd_sc_hd__nand2_4 _07123_ (.A(_01432_),
    .B(_01344_),
    .Y(_01923_));
 sky130_fd_sc_hd__or2_1 _07124_ (.A(_01336_),
    .B(_01355_),
    .X(_01924_));
 sky130_fd_sc_hd__clkbuf_4 _07125_ (.A(_01924_),
    .X(_01925_));
 sky130_fd_sc_hd__a22o_1 _07126_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[5] ),
    .A2(_01925_),
    .B1(_01855_),
    .B2(\genblk1[9].osc.clkdiv_C.cnt[0] ),
    .X(_01926_));
 sky130_fd_sc_hd__a221oi_1 _07127_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[2] ),
    .A2(_01920_),
    .B1(_01923_),
    .B2(\genblk1[9].osc.clkdiv_C.cnt[11] ),
    .C1(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__inv_2 _07128_ (.A(\genblk1[9].osc.clkdiv_C.cnt[8] ),
    .Y(_01928_));
 sky130_fd_sc_hd__nand2_1 _07129_ (.A(\genblk1[9].osc.clkdiv_C.cnt[9] ),
    .B(_01801_),
    .Y(_01929_));
 sky130_fd_sc_hd__inv_2 _07130_ (.A(\genblk1[9].osc.clkdiv_C.cnt[9] ),
    .Y(_01930_));
 sky130_fd_sc_hd__nand2_1 _07131_ (.A(_01930_),
    .B(_01250_),
    .Y(_01931_));
 sky130_fd_sc_hd__a2bb2o_1 _07132_ (.A1_N(\genblk1[9].osc.clkdiv_C.cnt[16] ),
    .A2_N(_01578_),
    .B1(_01349_),
    .B2(\genblk1[9].osc.clkdiv_C.cnt[15] ),
    .X(_01932_));
 sky130_fd_sc_hd__a221o_1 _07133_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[7] ),
    .A2(_01513_),
    .B1(_01929_),
    .B2(_01931_),
    .C1(_01932_),
    .X(_01933_));
 sky130_fd_sc_hd__o2bb2a_1 _07134_ (.A1_N(\genblk1[9].osc.clkdiv_C.cnt[4] ),
    .A2_N(_01311_),
    .B1(_01923_),
    .B2(\genblk1[9].osc.clkdiv_C.cnt[11] ),
    .X(_01934_));
 sky130_fd_sc_hd__o221a_1 _07135_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[4] ),
    .A2(_01311_),
    .B1(_01925_),
    .B2(\genblk1[9].osc.clkdiv_C.cnt[5] ),
    .C1(_01934_),
    .X(_01935_));
 sky130_fd_sc_hd__nor2_1 _07136_ (.A(\genblk1[9].osc.clkdiv_C.cnt[15] ),
    .B(_01361_),
    .Y(_01936_));
 sky130_fd_sc_hd__nor2_1 _07137_ (.A(\genblk1[9].osc.clkdiv_C.cnt[16] ),
    .B(_01936_),
    .Y(_01937_));
 sky130_fd_sc_hd__a21oi_1 _07138_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[14] ),
    .A2(_01246_),
    .B1(\genblk1[9].osc.clkdiv_C.cnt[17] ),
    .Y(_01938_));
 sky130_fd_sc_hd__o221a_1 _07139_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[14] ),
    .A2(_01246_),
    .B1(_01196_),
    .B2(_01937_),
    .C1(_01938_),
    .X(_01939_));
 sky130_fd_sc_hd__a22oi_1 _07140_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[6] ),
    .A2(_01334_),
    .B1(_01328_),
    .B2(\genblk1[9].osc.clkdiv_C.cnt[13] ),
    .Y(_01940_));
 sky130_fd_sc_hd__and3_1 _07141_ (.A(_01935_),
    .B(_01939_),
    .C(_01940_),
    .X(_01941_));
 sky130_fd_sc_hd__or2_1 _07142_ (.A(\genblk1[9].osc.clkdiv_C.cnt[3] ),
    .B(_01514_),
    .X(_01942_));
 sky130_fd_sc_hd__nand2_1 _07143_ (.A(\genblk1[9].osc.clkdiv_C.cnt[3] ),
    .B(_01514_),
    .Y(_01943_));
 sky130_fd_sc_hd__and4b_1 _07144_ (.A_N(_01933_),
    .B(_01941_),
    .C(_01942_),
    .D(_01943_),
    .X(_01944_));
 sky130_fd_sc_hd__o22a_1 _07145_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[8] ),
    .A2(_01514_),
    .B1(_01513_),
    .B2(\genblk1[9].osc.clkdiv_C.cnt[7] ),
    .X(_01945_));
 sky130_fd_sc_hd__nor2_4 _07146_ (.A(_01336_),
    .B(_01496_),
    .Y(_01946_));
 sky130_fd_sc_hd__nor2_1 _07147_ (.A(_01241_),
    .B(_01946_),
    .Y(_01947_));
 sky130_fd_sc_hd__nand2_1 _07148_ (.A(\genblk1[9].osc.clkdiv_C.cnt[1] ),
    .B(_01947_),
    .Y(_01948_));
 sky130_fd_sc_hd__o2bb2a_1 _07149_ (.A1_N(\genblk1[9].osc.clkdiv_C.cnt[12] ),
    .A2_N(_01799_),
    .B1(_01947_),
    .B2(\genblk1[9].osc.clkdiv_C.cnt[1] ),
    .X(_01949_));
 sky130_fd_sc_hd__o211a_1 _07150_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[12] ),
    .A2(_01799_),
    .B1(_01948_),
    .C1(_01949_),
    .X(_01950_));
 sky130_fd_sc_hd__o2111a_1 _07151_ (.A1(_01928_),
    .A2(net34),
    .B1(_01944_),
    .C1(_01945_),
    .D1(_01950_),
    .X(_01951_));
 sky130_fd_sc_hd__and4_2 _07152_ (.A(_01919_),
    .B(_01922_),
    .C(_01927_),
    .D(_01951_),
    .X(_01952_));
 sky130_fd_sc_hd__clkbuf_4 _07153_ (.A(_01952_),
    .X(_01953_));
 sky130_fd_sc_hd__nor2_1 _07154_ (.A(net1136),
    .B(_01953_),
    .Y(\genblk1[9].osc.clkdiv_C.next_cnt[0] ));
 sky130_fd_sc_hd__inv_2 _07155_ (.A(_01952_),
    .Y(_01954_));
 sky130_fd_sc_hd__or2_1 _07156_ (.A(\genblk1[9].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[9].osc.clkdiv_C.cnt[0] ),
    .X(_01955_));
 sky130_fd_sc_hd__nand2_1 _07157_ (.A(\genblk1[9].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[9].osc.clkdiv_C.cnt[0] ),
    .Y(_01956_));
 sky130_fd_sc_hd__and3_1 _07158_ (.A(_01954_),
    .B(_01955_),
    .C(_01956_),
    .X(_01957_));
 sky130_fd_sc_hd__clkbuf_1 _07159_ (.A(_01957_),
    .X(\genblk1[9].osc.clkdiv_C.next_cnt[1] ));
 sky130_fd_sc_hd__and3_1 _07160_ (.A(\genblk1[9].osc.clkdiv_C.cnt[2] ),
    .B(\genblk1[9].osc.clkdiv_C.cnt[1] ),
    .C(\genblk1[9].osc.clkdiv_C.cnt[0] ),
    .X(_01958_));
 sky130_fd_sc_hd__a21oi_1 _07161_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[1] ),
    .A2(\genblk1[9].osc.clkdiv_C.cnt[0] ),
    .B1(\genblk1[9].osc.clkdiv_C.cnt[2] ),
    .Y(_01959_));
 sky130_fd_sc_hd__nor3_1 _07162_ (.A(_01953_),
    .B(_01958_),
    .C(_01959_),
    .Y(\genblk1[9].osc.clkdiv_C.next_cnt[2] ));
 sky130_fd_sc_hd__and2_1 _07163_ (.A(\genblk1[9].osc.clkdiv_C.cnt[3] ),
    .B(_01958_),
    .X(_01960_));
 sky130_fd_sc_hd__nor2_1 _07164_ (.A(\genblk1[9].osc.clkdiv_C.cnt[3] ),
    .B(_01958_),
    .Y(_01961_));
 sky130_fd_sc_hd__nor3_1 _07165_ (.A(_01953_),
    .B(_01960_),
    .C(_01961_),
    .Y(\genblk1[9].osc.clkdiv_C.next_cnt[3] ));
 sky130_fd_sc_hd__nand2_1 _07166_ (.A(\genblk1[9].osc.clkdiv_C.cnt[4] ),
    .B(_01960_),
    .Y(_01962_));
 sky130_fd_sc_hd__or2_1 _07167_ (.A(\genblk1[9].osc.clkdiv_C.cnt[4] ),
    .B(_01960_),
    .X(_01963_));
 sky130_fd_sc_hd__and3_1 _07168_ (.A(_01954_),
    .B(_01962_),
    .C(_01963_),
    .X(_01964_));
 sky130_fd_sc_hd__clkbuf_1 _07169_ (.A(_01964_),
    .X(\genblk1[9].osc.clkdiv_C.next_cnt[4] ));
 sky130_fd_sc_hd__and3_1 _07170_ (.A(\genblk1[9].osc.clkdiv_C.cnt[5] ),
    .B(\genblk1[9].osc.clkdiv_C.cnt[4] ),
    .C(_01960_),
    .X(_01965_));
 sky130_fd_sc_hd__a21oi_1 _07171_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[4] ),
    .A2(_01960_),
    .B1(\genblk1[9].osc.clkdiv_C.cnt[5] ),
    .Y(_01966_));
 sky130_fd_sc_hd__nor3_1 _07172_ (.A(_01953_),
    .B(_01965_),
    .C(_01966_),
    .Y(\genblk1[9].osc.clkdiv_C.next_cnt[5] ));
 sky130_fd_sc_hd__and2_1 _07173_ (.A(\genblk1[9].osc.clkdiv_C.cnt[6] ),
    .B(_01965_),
    .X(_01967_));
 sky130_fd_sc_hd__nor2_1 _07174_ (.A(\genblk1[9].osc.clkdiv_C.cnt[6] ),
    .B(_01965_),
    .Y(_01968_));
 sky130_fd_sc_hd__nor3_1 _07175_ (.A(_01953_),
    .B(_01967_),
    .C(_01968_),
    .Y(\genblk1[9].osc.clkdiv_C.next_cnt[6] ));
 sky130_fd_sc_hd__nand2_1 _07176_ (.A(\genblk1[9].osc.clkdiv_C.cnt[7] ),
    .B(_01967_),
    .Y(_01969_));
 sky130_fd_sc_hd__or2_1 _07177_ (.A(\genblk1[9].osc.clkdiv_C.cnt[7] ),
    .B(_01967_),
    .X(_01970_));
 sky130_fd_sc_hd__and3_1 _07178_ (.A(_01954_),
    .B(_01969_),
    .C(_01970_),
    .X(_01971_));
 sky130_fd_sc_hd__clkbuf_1 _07179_ (.A(_01971_),
    .X(\genblk1[9].osc.clkdiv_C.next_cnt[7] ));
 sky130_fd_sc_hd__and3_1 _07180_ (.A(\genblk1[9].osc.clkdiv_C.cnt[8] ),
    .B(\genblk1[9].osc.clkdiv_C.cnt[7] ),
    .C(_01967_),
    .X(_01972_));
 sky130_fd_sc_hd__a21oi_1 _07181_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[7] ),
    .A2(_01967_),
    .B1(\genblk1[9].osc.clkdiv_C.cnt[8] ),
    .Y(_01973_));
 sky130_fd_sc_hd__nor3_1 _07182_ (.A(_01953_),
    .B(_01972_),
    .C(_01973_),
    .Y(\genblk1[9].osc.clkdiv_C.next_cnt[8] ));
 sky130_fd_sc_hd__and2_1 _07183_ (.A(\genblk1[9].osc.clkdiv_C.cnt[9] ),
    .B(_01972_),
    .X(_01974_));
 sky130_fd_sc_hd__nor2_1 _07184_ (.A(\genblk1[9].osc.clkdiv_C.cnt[9] ),
    .B(_01972_),
    .Y(_01975_));
 sky130_fd_sc_hd__nor3_1 _07185_ (.A(_01953_),
    .B(_01974_),
    .C(_01975_),
    .Y(\genblk1[9].osc.clkdiv_C.next_cnt[9] ));
 sky130_fd_sc_hd__nand2_1 _07186_ (.A(\genblk1[9].osc.clkdiv_C.cnt[10] ),
    .B(_01974_),
    .Y(_01976_));
 sky130_fd_sc_hd__o211a_1 _07187_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[10] ),
    .A2(_01974_),
    .B1(_01976_),
    .C1(_01954_),
    .X(\genblk1[9].osc.clkdiv_C.next_cnt[10] ));
 sky130_fd_sc_hd__a21oi_1 _07188_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[10] ),
    .A2(_01974_),
    .B1(\genblk1[9].osc.clkdiv_C.cnt[11] ),
    .Y(_01977_));
 sky130_fd_sc_hd__and3_1 _07189_ (.A(\genblk1[9].osc.clkdiv_C.cnt[11] ),
    .B(\genblk1[9].osc.clkdiv_C.cnt[10] ),
    .C(_01974_),
    .X(_01978_));
 sky130_fd_sc_hd__nor3_1 _07190_ (.A(_01953_),
    .B(_01977_),
    .C(_01978_),
    .Y(\genblk1[9].osc.clkdiv_C.next_cnt[11] ));
 sky130_fd_sc_hd__and2_1 _07191_ (.A(\genblk1[9].osc.clkdiv_C.cnt[12] ),
    .B(_01978_),
    .X(_01979_));
 sky130_fd_sc_hd__nor2_1 _07192_ (.A(_01953_),
    .B(_01979_),
    .Y(_01980_));
 sky130_fd_sc_hd__o21a_1 _07193_ (.A1(net1296),
    .A2(_01978_),
    .B1(_01980_),
    .X(\genblk1[9].osc.clkdiv_C.next_cnt[12] ));
 sky130_fd_sc_hd__and3_1 _07194_ (.A(\genblk1[9].osc.clkdiv_C.cnt[13] ),
    .B(\genblk1[9].osc.clkdiv_C.cnt[12] ),
    .C(_01978_),
    .X(_01981_));
 sky130_fd_sc_hd__nor2_1 _07195_ (.A(_01953_),
    .B(_01981_),
    .Y(_01982_));
 sky130_fd_sc_hd__o21a_1 _07196_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[13] ),
    .A2(_01979_),
    .B1(_01982_),
    .X(\genblk1[9].osc.clkdiv_C.next_cnt[13] ));
 sky130_fd_sc_hd__and2_1 _07197_ (.A(\genblk1[9].osc.clkdiv_C.cnt[14] ),
    .B(_01981_),
    .X(_01983_));
 sky130_fd_sc_hd__nor2_1 _07198_ (.A(_01952_),
    .B(_01983_),
    .Y(_01984_));
 sky130_fd_sc_hd__o21a_1 _07199_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[14] ),
    .A2(_01981_),
    .B1(_01984_),
    .X(\genblk1[9].osc.clkdiv_C.next_cnt[14] ));
 sky130_fd_sc_hd__and3_1 _07200_ (.A(\genblk1[9].osc.clkdiv_C.cnt[15] ),
    .B(\genblk1[9].osc.clkdiv_C.cnt[14] ),
    .C(_01981_),
    .X(_01985_));
 sky130_fd_sc_hd__nor2_1 _07201_ (.A(_01952_),
    .B(_01985_),
    .Y(_01986_));
 sky130_fd_sc_hd__o21a_1 _07202_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[15] ),
    .A2(_01983_),
    .B1(_01986_),
    .X(\genblk1[9].osc.clkdiv_C.next_cnt[15] ));
 sky130_fd_sc_hd__or2_1 _07203_ (.A(\genblk1[9].osc.clkdiv_C.cnt[16] ),
    .B(_01985_),
    .X(_01987_));
 sky130_fd_sc_hd__nand2_1 _07204_ (.A(\genblk1[9].osc.clkdiv_C.cnt[16] ),
    .B(_01985_),
    .Y(_01988_));
 sky130_fd_sc_hd__and3_1 _07205_ (.A(_01954_),
    .B(_01987_),
    .C(_01988_),
    .X(_01989_));
 sky130_fd_sc_hd__clkbuf_1 _07206_ (.A(_01989_),
    .X(\genblk1[9].osc.clkdiv_C.next_cnt[16] ));
 sky130_fd_sc_hd__xnor2_1 _07207_ (.A(net1194),
    .B(_01988_),
    .Y(\genblk1[9].osc.clkdiv_C.next_cnt[17] ));
 sky130_fd_sc_hd__inv_2 _07208_ (.A(\genblk1[10].osc.clkdiv_C.cnt[9] ),
    .Y(_01990_));
 sky130_fd_sc_hd__nand2_8 _07209_ (.A(_01556_),
    .B(_01564_),
    .Y(_01991_));
 sky130_fd_sc_hd__a21o_1 _07210_ (.A1(_01359_),
    .A2(_01224_),
    .B1(_01241_),
    .X(_01992_));
 sky130_fd_sc_hd__inv_2 _07211_ (.A(\genblk1[10].osc.clkdiv_C.cnt[4] ),
    .Y(_01993_));
 sky130_fd_sc_hd__a221o_1 _07212_ (.A1(_01308_),
    .A2(\genblk1[10].osc.clkdiv_C.cnt[2] ),
    .B1(_01214_),
    .B2(_01993_),
    .C1(\genblk1[10].osc.clkdiv_C.cnt[17] ),
    .X(_01994_));
 sky130_fd_sc_hd__inv_2 _07213_ (.A(\genblk1[10].osc.clkdiv_C.cnt[14] ),
    .Y(_01995_));
 sky130_fd_sc_hd__nor2_4 _07214_ (.A(_01181_),
    .B(_01187_),
    .Y(_01996_));
 sky130_fd_sc_hd__o21ai_1 _07215_ (.A1(_01490_),
    .A2(_01993_),
    .B1(\genblk1[10].osc.clkdiv_C.cnt[2] ),
    .Y(_01997_));
 sky130_fd_sc_hd__nor2_1 _07216_ (.A(\genblk1[10].osc.clkdiv_C.cnt[13] ),
    .B(_01442_),
    .Y(_01998_));
 sky130_fd_sc_hd__a221o_1 _07217_ (.A1(_01995_),
    .A2(_01996_),
    .B1(_01997_),
    .B2(_01342_),
    .C1(_01998_),
    .X(_01999_));
 sky130_fd_sc_hd__a221o_1 _07218_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[14] ),
    .A2(_01246_),
    .B1(_01442_),
    .B2(\genblk1[10].osc.clkdiv_C.cnt[13] ),
    .C1(_01999_),
    .X(_02000_));
 sky130_fd_sc_hd__nand2_2 _07219_ (.A(_01358_),
    .B(net37),
    .Y(_02001_));
 sky130_fd_sc_hd__or2_4 _07220_ (.A(_01365_),
    .B(_01189_),
    .X(_02002_));
 sky130_fd_sc_hd__inv_2 _07221_ (.A(\genblk1[10].osc.clkdiv_C.cnt[8] ),
    .Y(_02003_));
 sky130_fd_sc_hd__a2bb2o_1 _07222_ (.A1_N(\genblk1[10].osc.clkdiv_C.cnt[1] ),
    .A2_N(_02001_),
    .B1(_02002_),
    .B2(_02003_),
    .X(_02004_));
 sky130_fd_sc_hd__a21oi_4 _07223_ (.A1(_01174_),
    .A2(_01230_),
    .B1(_01196_),
    .Y(_02005_));
 sky130_fd_sc_hd__xnor2_1 _07224_ (.A(\genblk1[10].osc.clkdiv_C.cnt[11] ),
    .B(_02005_),
    .Y(_02006_));
 sky130_fd_sc_hd__or4_1 _07225_ (.A(_01994_),
    .B(_02000_),
    .C(_02004_),
    .D(_02006_),
    .X(_02007_));
 sky130_fd_sc_hd__a21oi_1 _07226_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[5] ),
    .A2(_01992_),
    .B1(_02007_),
    .Y(_02008_));
 sky130_fd_sc_hd__o21a_1 _07227_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[5] ),
    .A2(_01992_),
    .B1(_02008_),
    .X(_02009_));
 sky130_fd_sc_hd__o2bb2a_1 _07228_ (.A1_N(\genblk1[10].osc.clkdiv_C.cnt[7] ),
    .A2_N(_01235_),
    .B1(_01227_),
    .B2(\genblk1[10].osc.clkdiv_C.cnt[9] ),
    .X(_02010_));
 sky130_fd_sc_hd__nand2_4 _07229_ (.A(_01229_),
    .B(_01230_),
    .Y(_02011_));
 sky130_fd_sc_hd__xnor2_1 _07230_ (.A(\genblk1[10].osc.clkdiv_C.cnt[6] ),
    .B(_01432_),
    .Y(_02012_));
 sky130_fd_sc_hd__nor2_2 _07231_ (.A(_01225_),
    .B(_01354_),
    .Y(_02013_));
 sky130_fd_sc_hd__o2bb2a_1 _07232_ (.A1_N(\genblk1[10].osc.clkdiv_C.cnt[0] ),
    .A2_N(_01321_),
    .B1(_02013_),
    .B2(\genblk1[10].osc.clkdiv_C.cnt[3] ),
    .X(_02014_));
 sky130_fd_sc_hd__o21ba_1 _07233_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[16] ),
    .A2(_01363_),
    .B1_N(\genblk1[10].osc.clkdiv_C.cnt[15] ),
    .X(_02015_));
 sky130_fd_sc_hd__nor2_1 _07234_ (.A(\genblk1[10].osc.clkdiv_C.cnt[15] ),
    .B(_01359_),
    .Y(_02016_));
 sky130_fd_sc_hd__nor2_1 _07235_ (.A(\genblk1[10].osc.clkdiv_C.cnt[16] ),
    .B(_02016_),
    .Y(_02017_));
 sky130_fd_sc_hd__o2bb2a_1 _07236_ (.A1_N(\genblk1[10].osc.clkdiv_C.cnt[1] ),
    .A2_N(_02001_),
    .B1(_02002_),
    .B2(_02003_),
    .X(_02018_));
 sky130_fd_sc_hd__o221a_1 _07237_ (.A1(_01242_),
    .A2(_02015_),
    .B1(_02017_),
    .B2(_01197_),
    .C1(_02018_),
    .X(_02019_));
 sky130_fd_sc_hd__o2111a_1 _07238_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[12] ),
    .A2(_02011_),
    .B1(_02012_),
    .C1(_02014_),
    .D1(_02019_),
    .X(_02020_));
 sky130_fd_sc_hd__xnor2_1 _07239_ (.A(\genblk1[10].osc.clkdiv_C.cnt[10] ),
    .B(_01215_),
    .Y(_02021_));
 sky130_fd_sc_hd__a21oi_1 _07240_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[3] ),
    .A2(_02013_),
    .B1(_02021_),
    .Y(_02022_));
 sky130_fd_sc_hd__inv_2 _07241_ (.A(\genblk1[10].osc.clkdiv_C.cnt[12] ),
    .Y(_02023_));
 sky130_fd_sc_hd__o22a_1 _07242_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[0] ),
    .A2(_01321_),
    .B1(_01183_),
    .B2(_02023_),
    .X(_02024_));
 sky130_fd_sc_hd__o2111a_1 _07243_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[7] ),
    .A2(_01235_),
    .B1(_02020_),
    .C1(_02022_),
    .D1(_02024_),
    .X(_02025_));
 sky130_fd_sc_hd__o2111a_1 _07244_ (.A1(_01990_),
    .A2(_01991_),
    .B1(_02009_),
    .C1(_02010_),
    .D1(_02025_),
    .X(_02026_));
 sky130_fd_sc_hd__clkbuf_4 _07245_ (.A(_02026_),
    .X(_02027_));
 sky130_fd_sc_hd__nor2_1 _07246_ (.A(net1080),
    .B(_02027_),
    .Y(\genblk1[10].osc.clkdiv_C.next_cnt[0] ));
 sky130_fd_sc_hd__inv_2 _07247_ (.A(_02026_),
    .Y(_02028_));
 sky130_fd_sc_hd__or2_1 _07248_ (.A(\genblk1[10].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[10].osc.clkdiv_C.cnt[0] ),
    .X(_02029_));
 sky130_fd_sc_hd__nand2_1 _07249_ (.A(\genblk1[10].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[10].osc.clkdiv_C.cnt[0] ),
    .Y(_02030_));
 sky130_fd_sc_hd__and3_1 _07250_ (.A(_02028_),
    .B(_02029_),
    .C(_02030_),
    .X(_02031_));
 sky130_fd_sc_hd__clkbuf_1 _07251_ (.A(_02031_),
    .X(\genblk1[10].osc.clkdiv_C.next_cnt[1] ));
 sky130_fd_sc_hd__and3_1 _07252_ (.A(\genblk1[10].osc.clkdiv_C.cnt[2] ),
    .B(\genblk1[10].osc.clkdiv_C.cnt[1] ),
    .C(\genblk1[10].osc.clkdiv_C.cnt[0] ),
    .X(_02032_));
 sky130_fd_sc_hd__a21oi_1 _07253_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[1] ),
    .A2(\genblk1[10].osc.clkdiv_C.cnt[0] ),
    .B1(\genblk1[10].osc.clkdiv_C.cnt[2] ),
    .Y(_02033_));
 sky130_fd_sc_hd__nor3_1 _07254_ (.A(_02027_),
    .B(_02032_),
    .C(_02033_),
    .Y(\genblk1[10].osc.clkdiv_C.next_cnt[2] ));
 sky130_fd_sc_hd__and2_1 _07255_ (.A(\genblk1[10].osc.clkdiv_C.cnt[3] ),
    .B(_02032_),
    .X(_02034_));
 sky130_fd_sc_hd__nor2_1 _07256_ (.A(\genblk1[10].osc.clkdiv_C.cnt[3] ),
    .B(_02032_),
    .Y(_02035_));
 sky130_fd_sc_hd__nor3_1 _07257_ (.A(_02027_),
    .B(_02034_),
    .C(_02035_),
    .Y(\genblk1[10].osc.clkdiv_C.next_cnt[3] ));
 sky130_fd_sc_hd__nand2_1 _07258_ (.A(\genblk1[10].osc.clkdiv_C.cnt[4] ),
    .B(_02034_),
    .Y(_02036_));
 sky130_fd_sc_hd__or2_1 _07259_ (.A(\genblk1[10].osc.clkdiv_C.cnt[4] ),
    .B(_02034_),
    .X(_02037_));
 sky130_fd_sc_hd__and3_1 _07260_ (.A(_02028_),
    .B(_02036_),
    .C(_02037_),
    .X(_02038_));
 sky130_fd_sc_hd__clkbuf_1 _07261_ (.A(_02038_),
    .X(\genblk1[10].osc.clkdiv_C.next_cnt[4] ));
 sky130_fd_sc_hd__and3_1 _07262_ (.A(\genblk1[10].osc.clkdiv_C.cnt[5] ),
    .B(\genblk1[10].osc.clkdiv_C.cnt[4] ),
    .C(_02034_),
    .X(_02039_));
 sky130_fd_sc_hd__a21oi_1 _07263_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[4] ),
    .A2(_02034_),
    .B1(\genblk1[10].osc.clkdiv_C.cnt[5] ),
    .Y(_02040_));
 sky130_fd_sc_hd__nor3_1 _07264_ (.A(_02027_),
    .B(_02039_),
    .C(_02040_),
    .Y(\genblk1[10].osc.clkdiv_C.next_cnt[5] ));
 sky130_fd_sc_hd__and2_1 _07265_ (.A(\genblk1[10].osc.clkdiv_C.cnt[6] ),
    .B(_02039_),
    .X(_02041_));
 sky130_fd_sc_hd__nor2_1 _07266_ (.A(\genblk1[10].osc.clkdiv_C.cnt[6] ),
    .B(_02039_),
    .Y(_02042_));
 sky130_fd_sc_hd__nor3_1 _07267_ (.A(_02027_),
    .B(_02041_),
    .C(_02042_),
    .Y(\genblk1[10].osc.clkdiv_C.next_cnt[6] ));
 sky130_fd_sc_hd__nand2_1 _07268_ (.A(\genblk1[10].osc.clkdiv_C.cnt[7] ),
    .B(_02041_),
    .Y(_02043_));
 sky130_fd_sc_hd__or2_1 _07269_ (.A(\genblk1[10].osc.clkdiv_C.cnt[7] ),
    .B(_02041_),
    .X(_02044_));
 sky130_fd_sc_hd__and3_1 _07270_ (.A(_02028_),
    .B(_02043_),
    .C(_02044_),
    .X(_02045_));
 sky130_fd_sc_hd__clkbuf_1 _07271_ (.A(_02045_),
    .X(\genblk1[10].osc.clkdiv_C.next_cnt[7] ));
 sky130_fd_sc_hd__and3_1 _07272_ (.A(\genblk1[10].osc.clkdiv_C.cnt[8] ),
    .B(\genblk1[10].osc.clkdiv_C.cnt[7] ),
    .C(_02041_),
    .X(_02046_));
 sky130_fd_sc_hd__a21oi_1 _07273_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[7] ),
    .A2(_02041_),
    .B1(net1183),
    .Y(_02047_));
 sky130_fd_sc_hd__nor3_1 _07274_ (.A(_02027_),
    .B(_02046_),
    .C(_02047_),
    .Y(\genblk1[10].osc.clkdiv_C.next_cnt[8] ));
 sky130_fd_sc_hd__and2_1 _07275_ (.A(\genblk1[10].osc.clkdiv_C.cnt[9] ),
    .B(_02046_),
    .X(_02048_));
 sky130_fd_sc_hd__nor2_1 _07276_ (.A(\genblk1[10].osc.clkdiv_C.cnt[9] ),
    .B(_02046_),
    .Y(_02049_));
 sky130_fd_sc_hd__nor3_1 _07277_ (.A(_02027_),
    .B(_02048_),
    .C(_02049_),
    .Y(\genblk1[10].osc.clkdiv_C.next_cnt[9] ));
 sky130_fd_sc_hd__nand2_1 _07278_ (.A(\genblk1[10].osc.clkdiv_C.cnt[10] ),
    .B(_02048_),
    .Y(_02050_));
 sky130_fd_sc_hd__o211a_1 _07279_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[10] ),
    .A2(_02048_),
    .B1(_02050_),
    .C1(_02028_),
    .X(\genblk1[10].osc.clkdiv_C.next_cnt[10] ));
 sky130_fd_sc_hd__a21oi_1 _07280_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[10] ),
    .A2(_02048_),
    .B1(\genblk1[10].osc.clkdiv_C.cnt[11] ),
    .Y(_02051_));
 sky130_fd_sc_hd__and3_1 _07281_ (.A(\genblk1[10].osc.clkdiv_C.cnt[11] ),
    .B(\genblk1[10].osc.clkdiv_C.cnt[10] ),
    .C(_02048_),
    .X(_02052_));
 sky130_fd_sc_hd__nor3_1 _07282_ (.A(_02027_),
    .B(_02051_),
    .C(_02052_),
    .Y(\genblk1[10].osc.clkdiv_C.next_cnt[11] ));
 sky130_fd_sc_hd__and2_1 _07283_ (.A(\genblk1[10].osc.clkdiv_C.cnt[12] ),
    .B(_02052_),
    .X(_02053_));
 sky130_fd_sc_hd__nor2_1 _07284_ (.A(_02026_),
    .B(_02053_),
    .Y(_02054_));
 sky130_fd_sc_hd__o21a_1 _07285_ (.A1(net1119),
    .A2(_02052_),
    .B1(_02054_),
    .X(\genblk1[10].osc.clkdiv_C.next_cnt[12] ));
 sky130_fd_sc_hd__a21oi_1 _07286_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[13] ),
    .A2(_02053_),
    .B1(_02027_),
    .Y(_02055_));
 sky130_fd_sc_hd__o21a_1 _07287_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[13] ),
    .A2(_02053_),
    .B1(_02055_),
    .X(\genblk1[10].osc.clkdiv_C.next_cnt[13] ));
 sky130_fd_sc_hd__a21oi_1 _07288_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[13] ),
    .A2(_02053_),
    .B1(\genblk1[10].osc.clkdiv_C.cnt[14] ),
    .Y(_02056_));
 sky130_fd_sc_hd__and3_1 _07289_ (.A(\genblk1[10].osc.clkdiv_C.cnt[14] ),
    .B(\genblk1[10].osc.clkdiv_C.cnt[13] ),
    .C(_02053_),
    .X(_02057_));
 sky130_fd_sc_hd__nor3_1 _07290_ (.A(_02027_),
    .B(_02056_),
    .C(_02057_),
    .Y(\genblk1[10].osc.clkdiv_C.next_cnt[14] ));
 sky130_fd_sc_hd__and2_1 _07291_ (.A(\genblk1[10].osc.clkdiv_C.cnt[15] ),
    .B(_02057_),
    .X(_02058_));
 sky130_fd_sc_hd__nor2_1 _07292_ (.A(_02026_),
    .B(_02058_),
    .Y(_02059_));
 sky130_fd_sc_hd__o21a_1 _07293_ (.A1(net1143),
    .A2(_02057_),
    .B1(_02059_),
    .X(\genblk1[10].osc.clkdiv_C.next_cnt[15] ));
 sky130_fd_sc_hd__or2_1 _07294_ (.A(\genblk1[10].osc.clkdiv_C.cnt[16] ),
    .B(_02058_),
    .X(_02060_));
 sky130_fd_sc_hd__nand2_1 _07295_ (.A(\genblk1[10].osc.clkdiv_C.cnt[16] ),
    .B(_02058_),
    .Y(_02061_));
 sky130_fd_sc_hd__and3_1 _07296_ (.A(_02028_),
    .B(_02060_),
    .C(_02061_),
    .X(_02062_));
 sky130_fd_sc_hd__clkbuf_1 _07297_ (.A(_02062_),
    .X(\genblk1[10].osc.clkdiv_C.next_cnt[16] ));
 sky130_fd_sc_hd__xnor2_1 _07298_ (.A(net695),
    .B(_02061_),
    .Y(\genblk1[10].osc.clkdiv_C.next_cnt[17] ));
 sky130_fd_sc_hd__xnor2_1 _07299_ (.A(\genblk1[11].osc.clkdiv_C.cnt[9] ),
    .B(_01235_),
    .Y(_02063_));
 sky130_fd_sc_hd__nor2_4 _07300_ (.A(_01182_),
    .B(_01226_),
    .Y(_02064_));
 sky130_fd_sc_hd__nor2_1 _07301_ (.A(\genblk1[11].osc.clkdiv_C.cnt[6] ),
    .B(_01595_),
    .Y(_02065_));
 sky130_fd_sc_hd__a221o_1 _07302_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[13] ),
    .A2(_01256_),
    .B1(_02064_),
    .B2(\genblk1[11].osc.clkdiv_C.cnt[5] ),
    .C1(_02065_),
    .X(_02066_));
 sky130_fd_sc_hd__a2bb2o_1 _07303_ (.A1_N(\genblk1[11].osc.clkdiv_C.cnt[13] ),
    .A2_N(_01256_),
    .B1(_01595_),
    .B2(\genblk1[11].osc.clkdiv_C.cnt[6] ),
    .X(_02067_));
 sky130_fd_sc_hd__a2bb2o_1 _07304_ (.A1_N(\genblk1[11].osc.clkdiv_C.cnt[5] ),
    .A2_N(_02064_),
    .B1(_01925_),
    .B2(\genblk1[11].osc.clkdiv_C.cnt[2] ),
    .X(_02068_));
 sky130_fd_sc_hd__or4_1 _07305_ (.A(_02063_),
    .B(_02066_),
    .C(_02067_),
    .D(_02068_),
    .X(_02069_));
 sky130_fd_sc_hd__o21ai_1 _07306_ (.A1(_01223_),
    .A2(_01678_),
    .B1(\genblk1[11].osc.clkdiv_C.cnt[0] ),
    .Y(_02070_));
 sky130_fd_sc_hd__or3_1 _07307_ (.A(\genblk1[11].osc.clkdiv_C.cnt[0] ),
    .B(_01223_),
    .C(_01678_),
    .X(_02071_));
 sky130_fd_sc_hd__a22o_1 _07308_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[4] ),
    .A2(_01513_),
    .B1(_02070_),
    .B2(_02071_),
    .X(_02072_));
 sky130_fd_sc_hd__xnor2_1 _07309_ (.A(\genblk1[11].osc.clkdiv_C.cnt[7] ),
    .B(_01430_),
    .Y(_02073_));
 sky130_fd_sc_hd__xnor2_1 _07310_ (.A(\genblk1[11].osc.clkdiv_C.cnt[10] ),
    .B(_02002_),
    .Y(_02074_));
 sky130_fd_sc_hd__o2bb2a_1 _07311_ (.A1_N(\genblk1[11].osc.clkdiv_C.cnt[8] ),
    .A2_N(_01211_),
    .B1(_01262_),
    .B2(\genblk1[11].osc.clkdiv_C.cnt[11] ),
    .X(_02075_));
 sky130_fd_sc_hd__o221a_1 _07312_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[14] ),
    .A2(_01210_),
    .B1(_01578_),
    .B2(\genblk1[11].osc.clkdiv_C.cnt[16] ),
    .C1(_02075_),
    .X(_02076_));
 sky130_fd_sc_hd__nand2_2 _07313_ (.A(_01308_),
    .B(_01439_),
    .Y(_02077_));
 sky130_fd_sc_hd__a21oi_1 _07314_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[12] ),
    .A2(_02077_),
    .B1(\genblk1[11].osc.clkdiv_C.cnt[17] ),
    .Y(_02078_));
 sky130_fd_sc_hd__o221a_1 _07315_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[8] ),
    .A2(_01211_),
    .B1(_02077_),
    .B2(\genblk1[11].osc.clkdiv_C.cnt[12] ),
    .C1(_02078_),
    .X(_02079_));
 sky130_fd_sc_hd__inv_2 _07316_ (.A(\genblk1[11].osc.clkdiv_C.cnt[15] ),
    .Y(_02080_));
 sky130_fd_sc_hd__inv_2 _07317_ (.A(\genblk1[11].osc.clkdiv_C.cnt[14] ),
    .Y(_02081_));
 sky130_fd_sc_hd__nand2_1 _07318_ (.A(\genblk1[11].osc.clkdiv_C.cnt[11] ),
    .B(_01262_),
    .Y(_02082_));
 sky130_fd_sc_hd__o221a_1 _07319_ (.A1(_02080_),
    .A2(_01242_),
    .B1(_01423_),
    .B2(_02081_),
    .C1(_02082_),
    .X(_02083_));
 sky130_fd_sc_hd__o2111a_1 _07320_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[4] ),
    .A2(_01513_),
    .B1(_02076_),
    .C1(_02079_),
    .D1(_02083_),
    .X(_02084_));
 sky130_fd_sc_hd__nor2_1 _07321_ (.A(\genblk1[11].osc.clkdiv_C.cnt[15] ),
    .B(_01359_),
    .Y(_02085_));
 sky130_fd_sc_hd__nor2_1 _07322_ (.A(\genblk1[11].osc.clkdiv_C.cnt[16] ),
    .B(_02085_),
    .Y(_02086_));
 sky130_fd_sc_hd__o2bb2a_1 _07323_ (.A1_N(\genblk1[11].osc.clkdiv_C.cnt[3] ),
    .A2_N(_01334_),
    .B1(_01321_),
    .B2(\genblk1[11].osc.clkdiv_C.cnt[1] ),
    .X(_02087_));
 sky130_fd_sc_hd__o221a_1 _07324_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[3] ),
    .A2(_01334_),
    .B1(_02086_),
    .B2(_01197_),
    .C1(_02087_),
    .X(_02088_));
 sky130_fd_sc_hd__o2bb2a_1 _07325_ (.A1_N(\genblk1[11].osc.clkdiv_C.cnt[1] ),
    .A2_N(_01321_),
    .B1(_01925_),
    .B2(\genblk1[11].osc.clkdiv_C.cnt[2] ),
    .X(_02089_));
 sky130_fd_sc_hd__nand4_1 _07326_ (.A(_02074_),
    .B(_02084_),
    .C(_02088_),
    .D(_02089_),
    .Y(_02090_));
 sky130_fd_sc_hd__or4_4 _07327_ (.A(_02069_),
    .B(_02072_),
    .C(_02073_),
    .D(_02090_),
    .X(_02091_));
 sky130_fd_sc_hd__buf_2 _07328_ (.A(_02091_),
    .X(_02092_));
 sky130_fd_sc_hd__and2b_1 _07329_ (.A_N(\genblk1[11].osc.clkdiv_C.cnt[0] ),
    .B(_02092_),
    .X(_02093_));
 sky130_fd_sc_hd__clkbuf_1 _07330_ (.A(_02093_),
    .X(\genblk1[11].osc.clkdiv_C.next_cnt[0] ));
 sky130_fd_sc_hd__or2_1 _07331_ (.A(\genblk1[11].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[11].osc.clkdiv_C.cnt[0] ),
    .X(_02094_));
 sky130_fd_sc_hd__nand2_1 _07332_ (.A(\genblk1[11].osc.clkdiv_C.cnt[1] ),
    .B(\genblk1[11].osc.clkdiv_C.cnt[0] ),
    .Y(_02095_));
 sky130_fd_sc_hd__and3_1 _07333_ (.A(_02092_),
    .B(_02094_),
    .C(_02095_),
    .X(_02096_));
 sky130_fd_sc_hd__clkbuf_1 _07334_ (.A(_02096_),
    .X(\genblk1[11].osc.clkdiv_C.next_cnt[1] ));
 sky130_fd_sc_hd__and3_1 _07335_ (.A(\genblk1[11].osc.clkdiv_C.cnt[2] ),
    .B(\genblk1[11].osc.clkdiv_C.cnt[1] ),
    .C(\genblk1[11].osc.clkdiv_C.cnt[0] ),
    .X(_02097_));
 sky130_fd_sc_hd__inv_2 _07336_ (.A(_02097_),
    .Y(_02098_));
 sky130_fd_sc_hd__a21o_1 _07337_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[1] ),
    .A2(\genblk1[11].osc.clkdiv_C.cnt[0] ),
    .B1(\genblk1[11].osc.clkdiv_C.cnt[2] ),
    .X(_02099_));
 sky130_fd_sc_hd__and3_1 _07338_ (.A(_02092_),
    .B(_02098_),
    .C(_02099_),
    .X(_02100_));
 sky130_fd_sc_hd__clkbuf_1 _07339_ (.A(_02100_),
    .X(\genblk1[11].osc.clkdiv_C.next_cnt[2] ));
 sky130_fd_sc_hd__and2_1 _07340_ (.A(\genblk1[11].osc.clkdiv_C.cnt[3] ),
    .B(_02097_),
    .X(_02101_));
 sky130_fd_sc_hd__inv_2 _07341_ (.A(_02101_),
    .Y(_02102_));
 sky130_fd_sc_hd__or2_1 _07342_ (.A(\genblk1[11].osc.clkdiv_C.cnt[3] ),
    .B(_02097_),
    .X(_02103_));
 sky130_fd_sc_hd__and3_1 _07343_ (.A(_02092_),
    .B(_02102_),
    .C(_02103_),
    .X(_02104_));
 sky130_fd_sc_hd__clkbuf_1 _07344_ (.A(_02104_),
    .X(\genblk1[11].osc.clkdiv_C.next_cnt[3] ));
 sky130_fd_sc_hd__nand2_1 _07345_ (.A(\genblk1[11].osc.clkdiv_C.cnt[4] ),
    .B(_02101_),
    .Y(_02105_));
 sky130_fd_sc_hd__or2_1 _07346_ (.A(\genblk1[11].osc.clkdiv_C.cnt[4] ),
    .B(_02101_),
    .X(_02106_));
 sky130_fd_sc_hd__and3_1 _07347_ (.A(_02092_),
    .B(_02105_),
    .C(_02106_),
    .X(_02107_));
 sky130_fd_sc_hd__clkbuf_1 _07348_ (.A(_02107_),
    .X(\genblk1[11].osc.clkdiv_C.next_cnt[4] ));
 sky130_fd_sc_hd__and3_1 _07349_ (.A(\genblk1[11].osc.clkdiv_C.cnt[5] ),
    .B(\genblk1[11].osc.clkdiv_C.cnt[4] ),
    .C(_02101_),
    .X(_02108_));
 sky130_fd_sc_hd__inv_2 _07350_ (.A(_02108_),
    .Y(_02109_));
 sky130_fd_sc_hd__a31o_1 _07351_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[4] ),
    .A2(\genblk1[11].osc.clkdiv_C.cnt[3] ),
    .A3(_02097_),
    .B1(\genblk1[11].osc.clkdiv_C.cnt[5] ),
    .X(_02110_));
 sky130_fd_sc_hd__and3_1 _07352_ (.A(_02092_),
    .B(_02109_),
    .C(_02110_),
    .X(_02111_));
 sky130_fd_sc_hd__clkbuf_1 _07353_ (.A(_02111_),
    .X(\genblk1[11].osc.clkdiv_C.next_cnt[5] ));
 sky130_fd_sc_hd__and2_1 _07354_ (.A(\genblk1[11].osc.clkdiv_C.cnt[6] ),
    .B(_02108_),
    .X(_02112_));
 sky130_fd_sc_hd__inv_2 _07355_ (.A(_02112_),
    .Y(_02113_));
 sky130_fd_sc_hd__or2_1 _07356_ (.A(\genblk1[11].osc.clkdiv_C.cnt[6] ),
    .B(_02108_),
    .X(_02114_));
 sky130_fd_sc_hd__and3_1 _07357_ (.A(_02092_),
    .B(_02113_),
    .C(_02114_),
    .X(_02115_));
 sky130_fd_sc_hd__clkbuf_1 _07358_ (.A(_02115_),
    .X(\genblk1[11].osc.clkdiv_C.next_cnt[6] ));
 sky130_fd_sc_hd__nand2_1 _07359_ (.A(\genblk1[11].osc.clkdiv_C.cnt[7] ),
    .B(_02112_),
    .Y(_02116_));
 sky130_fd_sc_hd__or2_1 _07360_ (.A(\genblk1[11].osc.clkdiv_C.cnt[7] ),
    .B(_02112_),
    .X(_02117_));
 sky130_fd_sc_hd__and3_1 _07361_ (.A(_02091_),
    .B(_02116_),
    .C(_02117_),
    .X(_02118_));
 sky130_fd_sc_hd__clkbuf_1 _07362_ (.A(_02118_),
    .X(\genblk1[11].osc.clkdiv_C.next_cnt[7] ));
 sky130_fd_sc_hd__and3_1 _07363_ (.A(\genblk1[11].osc.clkdiv_C.cnt[8] ),
    .B(\genblk1[11].osc.clkdiv_C.cnt[7] ),
    .C(_02112_),
    .X(_02119_));
 sky130_fd_sc_hd__inv_2 _07364_ (.A(_02119_),
    .Y(_02120_));
 sky130_fd_sc_hd__a31o_1 _07365_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[7] ),
    .A2(\genblk1[11].osc.clkdiv_C.cnt[6] ),
    .A3(_02108_),
    .B1(\genblk1[11].osc.clkdiv_C.cnt[8] ),
    .X(_02121_));
 sky130_fd_sc_hd__and3_1 _07366_ (.A(_02091_),
    .B(_02120_),
    .C(_02121_),
    .X(_02122_));
 sky130_fd_sc_hd__clkbuf_1 _07367_ (.A(_02122_),
    .X(\genblk1[11].osc.clkdiv_C.next_cnt[8] ));
 sky130_fd_sc_hd__and2_1 _07368_ (.A(\genblk1[11].osc.clkdiv_C.cnt[9] ),
    .B(_02119_),
    .X(_02123_));
 sky130_fd_sc_hd__inv_2 _07369_ (.A(_02123_),
    .Y(_02124_));
 sky130_fd_sc_hd__or2_1 _07370_ (.A(\genblk1[11].osc.clkdiv_C.cnt[9] ),
    .B(_02119_),
    .X(_02125_));
 sky130_fd_sc_hd__and3_1 _07371_ (.A(_02091_),
    .B(_02124_),
    .C(_02125_),
    .X(_02126_));
 sky130_fd_sc_hd__clkbuf_1 _07372_ (.A(_02126_),
    .X(\genblk1[11].osc.clkdiv_C.next_cnt[9] ));
 sky130_fd_sc_hd__nand2_1 _07373_ (.A(\genblk1[11].osc.clkdiv_C.cnt[10] ),
    .B(_02123_),
    .Y(_02127_));
 sky130_fd_sc_hd__o211a_1 _07374_ (.A1(net1269),
    .A2(_02123_),
    .B1(_02127_),
    .C1(_02092_),
    .X(\genblk1[11].osc.clkdiv_C.next_cnt[10] ));
 sky130_fd_sc_hd__inv_2 _07375_ (.A(\genblk1[11].osc.clkdiv_C.cnt[11] ),
    .Y(_02128_));
 sky130_fd_sc_hd__nand2_1 _07376_ (.A(_02128_),
    .B(_02127_),
    .Y(_02129_));
 sky130_fd_sc_hd__o211a_1 _07377_ (.A1(_02128_),
    .A2(_02127_),
    .B1(_02129_),
    .C1(_02092_),
    .X(\genblk1[11].osc.clkdiv_C.next_cnt[11] ));
 sky130_fd_sc_hd__nor2_1 _07378_ (.A(_02128_),
    .B(_02127_),
    .Y(_02130_));
 sky130_fd_sc_hd__or2_1 _07379_ (.A(\genblk1[11].osc.clkdiv_C.cnt[12] ),
    .B(_02130_),
    .X(_02131_));
 sky130_fd_sc_hd__and2_1 _07380_ (.A(\genblk1[11].osc.clkdiv_C.cnt[12] ),
    .B(_02130_),
    .X(_02132_));
 sky130_fd_sc_hd__inv_2 _07381_ (.A(_02132_),
    .Y(_02133_));
 sky130_fd_sc_hd__and3_1 _07382_ (.A(_02091_),
    .B(_02131_),
    .C(_02133_),
    .X(_02134_));
 sky130_fd_sc_hd__clkbuf_1 _07383_ (.A(_02134_),
    .X(\genblk1[11].osc.clkdiv_C.next_cnt[12] ));
 sky130_fd_sc_hd__or2_1 _07384_ (.A(\genblk1[11].osc.clkdiv_C.cnt[13] ),
    .B(_02132_),
    .X(_02135_));
 sky130_fd_sc_hd__nand2_1 _07385_ (.A(\genblk1[11].osc.clkdiv_C.cnt[13] ),
    .B(_02132_),
    .Y(_02136_));
 sky130_fd_sc_hd__and3_1 _07386_ (.A(_02091_),
    .B(_02135_),
    .C(_02136_),
    .X(_02137_));
 sky130_fd_sc_hd__clkbuf_1 _07387_ (.A(_02137_),
    .X(\genblk1[11].osc.clkdiv_C.next_cnt[13] ));
 sky130_fd_sc_hd__nand2_1 _07388_ (.A(_02081_),
    .B(_02136_),
    .Y(_02138_));
 sky130_fd_sc_hd__nor2_1 _07389_ (.A(_02081_),
    .B(_02136_),
    .Y(_02139_));
 sky130_fd_sc_hd__inv_2 _07390_ (.A(_02139_),
    .Y(_02140_));
 sky130_fd_sc_hd__and3_1 _07391_ (.A(_02091_),
    .B(_02138_),
    .C(_02140_),
    .X(_02141_));
 sky130_fd_sc_hd__clkbuf_1 _07392_ (.A(_02141_),
    .X(\genblk1[11].osc.clkdiv_C.next_cnt[14] ));
 sky130_fd_sc_hd__or2_1 _07393_ (.A(\genblk1[11].osc.clkdiv_C.cnt[15] ),
    .B(_02139_),
    .X(_02142_));
 sky130_fd_sc_hd__o211a_1 _07394_ (.A1(_02080_),
    .A2(_02140_),
    .B1(_02142_),
    .C1(_02092_),
    .X(\genblk1[11].osc.clkdiv_C.next_cnt[15] ));
 sky130_fd_sc_hd__nor2_1 _07395_ (.A(_02080_),
    .B(_02140_),
    .Y(_02143_));
 sky130_fd_sc_hd__or2_1 _07396_ (.A(\genblk1[11].osc.clkdiv_C.cnt[16] ),
    .B(_02143_),
    .X(_02144_));
 sky130_fd_sc_hd__nand2_1 _07397_ (.A(\genblk1[11].osc.clkdiv_C.cnt[16] ),
    .B(_02143_),
    .Y(_02145_));
 sky130_fd_sc_hd__and3_1 _07398_ (.A(_02091_),
    .B(_02144_),
    .C(_02145_),
    .X(_02146_));
 sky130_fd_sc_hd__clkbuf_1 _07399_ (.A(_02146_),
    .X(\genblk1[11].osc.clkdiv_C.next_cnt[16] ));
 sky130_fd_sc_hd__xnor2_1 _07400_ (.A(net1220),
    .B(_02145_),
    .Y(\genblk1[11].osc.clkdiv_C.next_cnt[17] ));
 sky130_fd_sc_hd__buf_8 _07401_ (.A(\genblk2[0].wave_shpr.div.start ),
    .X(_02147_));
 sky130_fd_sc_hd__nand3b_1 _07402_ (.A_N(\genblk2[0].wave_shpr.div.i[2] ),
    .B(\genblk2[0].wave_shpr.div.i[3] ),
    .C(\genblk2[0].wave_shpr.div.i[0] ),
    .Y(_02148_));
 sky130_fd_sc_hd__or3b_1 _07403_ (.A(\genblk2[0].wave_shpr.div.i[1] ),
    .B(_02148_),
    .C_N(\genblk2[0].wave_shpr.div.i[4] ),
    .X(_02149_));
 sky130_fd_sc_hd__and2_1 _07404_ (.A(\genblk2[0].wave_shpr.div.busy ),
    .B(_02149_),
    .X(_02150_));
 sky130_fd_sc_hd__nor2_1 _07405_ (.A(_02147_),
    .B(_02150_),
    .Y(_02151_));
 sky130_fd_sc_hd__inv_2 _07406_ (.A(_02151_),
    .Y(_00000_));
 sky130_fd_sc_hd__inv_6 _07407_ (.A(\genblk2[0].wave_shpr.div.start ),
    .Y(_02152_));
 sky130_fd_sc_hd__buf_6 _07408_ (.A(_02152_),
    .X(_02153_));
 sky130_fd_sc_hd__and3b_1 _07409_ (.A_N(_02149_),
    .B(_02153_),
    .C(\genblk2[0].wave_shpr.div.busy ),
    .X(_02154_));
 sky130_fd_sc_hd__clkbuf_4 _07410_ (.A(_02154_),
    .X(_00001_));
 sky130_fd_sc_hd__buf_8 _07411_ (.A(\genblk2[0].wave_shpr.div.start ),
    .X(_02155_));
 sky130_fd_sc_hd__nand3b_1 _07412_ (.A_N(\genblk2[1].wave_shpr.div.i[2] ),
    .B(\genblk2[1].wave_shpr.div.i[3] ),
    .C(\genblk2[1].wave_shpr.div.i[0] ),
    .Y(_02156_));
 sky130_fd_sc_hd__or3b_1 _07413_ (.A(\genblk2[1].wave_shpr.div.i[1] ),
    .B(_02156_),
    .C_N(\genblk2[1].wave_shpr.div.i[4] ),
    .X(_02157_));
 sky130_fd_sc_hd__and2_1 _07414_ (.A(\genblk2[1].wave_shpr.div.busy ),
    .B(_02157_),
    .X(_02158_));
 sky130_fd_sc_hd__nor2_1 _07415_ (.A(_02155_),
    .B(_02158_),
    .Y(_02159_));
 sky130_fd_sc_hd__inv_2 _07416_ (.A(_02159_),
    .Y(_00006_));
 sky130_fd_sc_hd__and3b_2 _07417_ (.A_N(_02157_),
    .B(_02153_),
    .C(\genblk2[1].wave_shpr.div.busy ),
    .X(_02160_));
 sky130_fd_sc_hd__clkbuf_4 _07418_ (.A(_02160_),
    .X(_00007_));
 sky130_fd_sc_hd__nand3b_1 _07419_ (.A_N(\genblk2[2].wave_shpr.div.i[2] ),
    .B(\genblk2[2].wave_shpr.div.i[3] ),
    .C(\genblk2[2].wave_shpr.div.i[0] ),
    .Y(_02161_));
 sky130_fd_sc_hd__or3b_1 _07420_ (.A(\genblk2[2].wave_shpr.div.i[1] ),
    .B(_02161_),
    .C_N(\genblk2[2].wave_shpr.div.i[4] ),
    .X(_02162_));
 sky130_fd_sc_hd__and2_1 _07421_ (.A(\genblk2[2].wave_shpr.div.busy ),
    .B(_02162_),
    .X(_02163_));
 sky130_fd_sc_hd__nor2_1 _07422_ (.A(_02147_),
    .B(_02163_),
    .Y(_02164_));
 sky130_fd_sc_hd__inv_2 _07423_ (.A(_02164_),
    .Y(_00008_));
 sky130_fd_sc_hd__and3b_1 _07424_ (.A_N(_02162_),
    .B(_02153_),
    .C(\genblk2[2].wave_shpr.div.busy ),
    .X(_02165_));
 sky130_fd_sc_hd__buf_4 _07425_ (.A(_02165_),
    .X(_00009_));
 sky130_fd_sc_hd__nand3b_1 _07426_ (.A_N(\genblk2[3].wave_shpr.div.i[2] ),
    .B(\genblk2[3].wave_shpr.div.i[3] ),
    .C(\genblk2[3].wave_shpr.div.i[0] ),
    .Y(_02166_));
 sky130_fd_sc_hd__or3b_1 _07427_ (.A(\genblk2[3].wave_shpr.div.i[1] ),
    .B(_02166_),
    .C_N(\genblk2[3].wave_shpr.div.i[4] ),
    .X(_02167_));
 sky130_fd_sc_hd__and2_1 _07428_ (.A(\genblk2[3].wave_shpr.div.busy ),
    .B(_02167_),
    .X(_02168_));
 sky130_fd_sc_hd__nor2_1 _07429_ (.A(_02155_),
    .B(_02168_),
    .Y(_02169_));
 sky130_fd_sc_hd__inv_2 _07430_ (.A(_02169_),
    .Y(_00010_));
 sky130_fd_sc_hd__buf_6 _07431_ (.A(_02152_),
    .X(_02170_));
 sky130_fd_sc_hd__buf_8 _07432_ (.A(_02170_),
    .X(_02171_));
 sky130_fd_sc_hd__nor3b_1 _07433_ (.A(\genblk2[3].wave_shpr.div.i[1] ),
    .B(_02166_),
    .C_N(\genblk2[3].wave_shpr.div.i[4] ),
    .Y(_02172_));
 sky130_fd_sc_hd__and3_1 _07434_ (.A(_02171_),
    .B(\genblk2[3].wave_shpr.div.busy ),
    .C(_02172_),
    .X(_02173_));
 sky130_fd_sc_hd__buf_1 _07435_ (.A(_02173_),
    .X(_00011_));
 sky130_fd_sc_hd__nand3b_1 _07436_ (.A_N(\genblk2[4].wave_shpr.div.i[2] ),
    .B(\genblk2[4].wave_shpr.div.i[3] ),
    .C(\genblk2[4].wave_shpr.div.i[0] ),
    .Y(_02174_));
 sky130_fd_sc_hd__or3b_1 _07437_ (.A(\genblk2[4].wave_shpr.div.i[1] ),
    .B(_02174_),
    .C_N(\genblk2[4].wave_shpr.div.i[4] ),
    .X(_02175_));
 sky130_fd_sc_hd__and2_1 _07438_ (.A(\genblk2[4].wave_shpr.div.busy ),
    .B(_02175_),
    .X(_02176_));
 sky130_fd_sc_hd__nor2_1 _07439_ (.A(_02147_),
    .B(_02176_),
    .Y(_02177_));
 sky130_fd_sc_hd__inv_2 _07440_ (.A(_02177_),
    .Y(_00012_));
 sky130_fd_sc_hd__and3b_1 _07441_ (.A_N(_02175_),
    .B(_02153_),
    .C(\genblk2[4].wave_shpr.div.busy ),
    .X(_02178_));
 sky130_fd_sc_hd__clkbuf_4 _07442_ (.A(_02178_),
    .X(_00013_));
 sky130_fd_sc_hd__nand3b_1 _07443_ (.A_N(\genblk2[5].wave_shpr.div.i[2] ),
    .B(\genblk2[5].wave_shpr.div.i[3] ),
    .C(\genblk2[5].wave_shpr.div.i[0] ),
    .Y(_02179_));
 sky130_fd_sc_hd__or3b_1 _07444_ (.A(\genblk2[5].wave_shpr.div.i[1] ),
    .B(_02179_),
    .C_N(\genblk2[5].wave_shpr.div.i[4] ),
    .X(_02180_));
 sky130_fd_sc_hd__and2_1 _07445_ (.A(\genblk2[5].wave_shpr.div.busy ),
    .B(_02180_),
    .X(_02181_));
 sky130_fd_sc_hd__nor2_1 _07446_ (.A(_02147_),
    .B(_02181_),
    .Y(_02182_));
 sky130_fd_sc_hd__clkbuf_4 _07447_ (.A(_02182_),
    .X(_02183_));
 sky130_fd_sc_hd__inv_2 _07448_ (.A(_02183_),
    .Y(_00014_));
 sky130_fd_sc_hd__and3b_1 _07449_ (.A_N(_02180_),
    .B(_02153_),
    .C(\genblk2[5].wave_shpr.div.busy ),
    .X(_02184_));
 sky130_fd_sc_hd__clkbuf_4 _07450_ (.A(_02184_),
    .X(_00015_));
 sky130_fd_sc_hd__nand3b_1 _07451_ (.A_N(\genblk2[6].wave_shpr.div.i[2] ),
    .B(\genblk2[6].wave_shpr.div.i[3] ),
    .C(\genblk2[6].wave_shpr.div.i[0] ),
    .Y(_02185_));
 sky130_fd_sc_hd__or3b_1 _07452_ (.A(\genblk2[6].wave_shpr.div.i[1] ),
    .B(_02185_),
    .C_N(\genblk2[6].wave_shpr.div.i[4] ),
    .X(_02186_));
 sky130_fd_sc_hd__and2_1 _07453_ (.A(\genblk2[6].wave_shpr.div.busy ),
    .B(_02186_),
    .X(_02187_));
 sky130_fd_sc_hd__nor2_1 _07454_ (.A(_02147_),
    .B(_02187_),
    .Y(_02188_));
 sky130_fd_sc_hd__inv_2 _07455_ (.A(_02188_),
    .Y(_00016_));
 sky130_fd_sc_hd__and3b_1 _07456_ (.A_N(_02186_),
    .B(_02153_),
    .C(\genblk2[6].wave_shpr.div.busy ),
    .X(_02189_));
 sky130_fd_sc_hd__clkbuf_4 _07457_ (.A(_02189_),
    .X(_00017_));
 sky130_fd_sc_hd__nand3b_1 _07458_ (.A_N(\genblk2[7].wave_shpr.div.i[2] ),
    .B(\genblk2[7].wave_shpr.div.i[3] ),
    .C(\genblk2[7].wave_shpr.div.i[4] ),
    .Y(_02190_));
 sky130_fd_sc_hd__or3b_1 _07459_ (.A(_02190_),
    .B(\genblk2[7].wave_shpr.div.i[1] ),
    .C_N(\genblk2[7].wave_shpr.div.i[0] ),
    .X(_02191_));
 sky130_fd_sc_hd__and2_1 _07460_ (.A(\genblk2[7].wave_shpr.div.busy ),
    .B(_02191_),
    .X(_02192_));
 sky130_fd_sc_hd__nor2_1 _07461_ (.A(_02155_),
    .B(_02192_),
    .Y(_02193_));
 sky130_fd_sc_hd__inv_2 _07462_ (.A(_02193_),
    .Y(_00018_));
 sky130_fd_sc_hd__and3b_1 _07463_ (.A_N(_02191_),
    .B(_02153_),
    .C(\genblk2[7].wave_shpr.div.busy ),
    .X(_02194_));
 sky130_fd_sc_hd__clkbuf_4 _07464_ (.A(_02194_),
    .X(_00019_));
 sky130_fd_sc_hd__nand3b_1 _07465_ (.A_N(\genblk2[8].wave_shpr.div.i[2] ),
    .B(\genblk2[8].wave_shpr.div.i[3] ),
    .C(\genblk2[8].wave_shpr.div.i[4] ),
    .Y(_02195_));
 sky130_fd_sc_hd__or3b_1 _07466_ (.A(_02195_),
    .B(\genblk2[8].wave_shpr.div.i[1] ),
    .C_N(\genblk2[8].wave_shpr.div.i[0] ),
    .X(_02196_));
 sky130_fd_sc_hd__and2_1 _07467_ (.A(\genblk2[8].wave_shpr.div.busy ),
    .B(_02196_),
    .X(_02197_));
 sky130_fd_sc_hd__nor2_1 _07468_ (.A(_02147_),
    .B(_02197_),
    .Y(_02198_));
 sky130_fd_sc_hd__inv_2 _07469_ (.A(_02198_),
    .Y(_00020_));
 sky130_fd_sc_hd__and3b_1 _07470_ (.A_N(_02196_),
    .B(_02153_),
    .C(\genblk2[8].wave_shpr.div.busy ),
    .X(_02199_));
 sky130_fd_sc_hd__clkbuf_4 _07471_ (.A(_02199_),
    .X(_00021_));
 sky130_fd_sc_hd__nand3b_1 _07472_ (.A_N(\genblk2[9].wave_shpr.div.i[2] ),
    .B(\genblk2[9].wave_shpr.div.i[3] ),
    .C(\genblk2[9].wave_shpr.div.i[0] ),
    .Y(_02200_));
 sky130_fd_sc_hd__or3b_1 _07473_ (.A(\genblk2[9].wave_shpr.div.i[1] ),
    .B(_02200_),
    .C_N(\genblk2[9].wave_shpr.div.i[4] ),
    .X(_02201_));
 sky130_fd_sc_hd__and2_2 _07474_ (.A(\genblk2[9].wave_shpr.div.busy ),
    .B(_02201_),
    .X(_02202_));
 sky130_fd_sc_hd__nor2_4 _07475_ (.A(_02155_),
    .B(_02202_),
    .Y(_02203_));
 sky130_fd_sc_hd__inv_2 _07476_ (.A(_02203_),
    .Y(_00022_));
 sky130_fd_sc_hd__and3b_1 _07477_ (.A_N(_02201_),
    .B(_02153_),
    .C(\genblk2[9].wave_shpr.div.busy ),
    .X(_02204_));
 sky130_fd_sc_hd__clkbuf_4 _07478_ (.A(_02204_),
    .X(_00023_));
 sky130_fd_sc_hd__nand3b_1 _07479_ (.A_N(\genblk2[10].wave_shpr.div.i[2] ),
    .B(\genblk2[10].wave_shpr.div.i[3] ),
    .C(\genblk2[10].wave_shpr.div.i[0] ),
    .Y(_02205_));
 sky130_fd_sc_hd__or3b_1 _07480_ (.A(\genblk2[10].wave_shpr.div.i[1] ),
    .B(_02205_),
    .C_N(\genblk2[10].wave_shpr.div.i[4] ),
    .X(_02206_));
 sky130_fd_sc_hd__and2_1 _07481_ (.A(\genblk2[10].wave_shpr.div.busy ),
    .B(_02206_),
    .X(_02207_));
 sky130_fd_sc_hd__nor2_1 _07482_ (.A(_02147_),
    .B(_02207_),
    .Y(_02208_));
 sky130_fd_sc_hd__inv_2 _07483_ (.A(_02208_),
    .Y(_00002_));
 sky130_fd_sc_hd__and3b_2 _07484_ (.A_N(_02206_),
    .B(_02153_),
    .C(\genblk2[10].wave_shpr.div.busy ),
    .X(_02209_));
 sky130_fd_sc_hd__clkbuf_4 _07485_ (.A(_02209_),
    .X(_00003_));
 sky130_fd_sc_hd__nand3b_1 _07486_ (.A_N(\genblk2[11].wave_shpr.div.i[2] ),
    .B(\genblk2[11].wave_shpr.div.i[3] ),
    .C(\genblk2[11].wave_shpr.div.i[0] ),
    .Y(_02210_));
 sky130_fd_sc_hd__or3b_1 _07487_ (.A(\genblk2[11].wave_shpr.div.i[1] ),
    .B(_02210_),
    .C_N(\genblk2[11].wave_shpr.div.i[4] ),
    .X(_02211_));
 sky130_fd_sc_hd__and2_1 _07488_ (.A(\genblk2[11].wave_shpr.div.busy ),
    .B(_02211_),
    .X(_02212_));
 sky130_fd_sc_hd__nor2_1 _07489_ (.A(_02147_),
    .B(_02212_),
    .Y(_02213_));
 sky130_fd_sc_hd__inv_2 _07490_ (.A(_02213_),
    .Y(_00004_));
 sky130_fd_sc_hd__and3b_1 _07491_ (.A_N(_02211_),
    .B(_02152_),
    .C(\genblk2[11].wave_shpr.div.busy ),
    .X(_02214_));
 sky130_fd_sc_hd__clkbuf_4 _07492_ (.A(_02214_),
    .X(_00005_));
 sky130_fd_sc_hd__inv_2 _07493_ (.A(\modein.delay_in[0] ),
    .Y(_02215_));
 sky130_fd_sc_hd__buf_2 _07494_ (.A(net17),
    .X(_02216_));
 sky130_fd_sc_hd__buf_2 _07495_ (.A(_02216_),
    .X(_02217_));
 sky130_fd_sc_hd__o21ai_1 _07496_ (.A1(_02215_),
    .A2(net760),
    .B1(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__or3_1 _07497_ (.A(_02217_),
    .B(_02215_),
    .C(net760),
    .X(_02219_));
 sky130_fd_sc_hd__nand2_1 _07498_ (.A(_02218_),
    .B(_02219_),
    .Y(\FSM.next_mode[0] ));
 sky130_fd_sc_hd__or2b_1 _07499_ (.A(net18),
    .B_N(net17),
    .X(_02220_));
 sky130_fd_sc_hd__buf_4 _07500_ (.A(_02220_),
    .X(_02221_));
 sky130_fd_sc_hd__nand2b_4 _07501_ (.A_N(net17),
    .B(net18),
    .Y(_02222_));
 sky130_fd_sc_hd__buf_4 _07502_ (.A(_02222_),
    .X(_02223_));
 sky130_fd_sc_hd__clkbuf_4 _07503_ (.A(_02223_),
    .X(_02224_));
 sky130_fd_sc_hd__nor2b_2 _07504_ (.A(net18),
    .B_N(net17),
    .Y(_02225_));
 sky130_fd_sc_hd__o21a_1 _07505_ (.A1(_02215_),
    .A2(net760),
    .B1(_02225_),
    .X(_02226_));
 sky130_fd_sc_hd__a31oi_1 _07506_ (.A1(_02218_),
    .A2(_02221_),
    .A3(_02224_),
    .B1(_02226_),
    .Y(\FSM.next_mode[1] ));
 sky130_fd_sc_hd__inv_2 _07507_ (.A(\PWM.counter[7] ),
    .Y(_02227_));
 sky130_fd_sc_hd__inv_2 _07508_ (.A(\PWM.counter[6] ),
    .Y(_02228_));
 sky130_fd_sc_hd__and2_1 _07509_ (.A(_02228_),
    .B(\PWM.final_sample_in[6] ),
    .X(_02229_));
 sky130_fd_sc_hd__inv_2 _07510_ (.A(\PWM.counter[5] ),
    .Y(_02230_));
 sky130_fd_sc_hd__and2_1 _07511_ (.A(_02230_),
    .B(\PWM.final_sample_in[5] ),
    .X(_02231_));
 sky130_fd_sc_hd__inv_2 _07512_ (.A(\PWM.counter[3] ),
    .Y(_02232_));
 sky130_fd_sc_hd__or2_1 _07513_ (.A(_02232_),
    .B(\PWM.final_sample_in[3] ),
    .X(_02233_));
 sky130_fd_sc_hd__inv_2 _07514_ (.A(\PWM.counter[2] ),
    .Y(_02234_));
 sky130_fd_sc_hd__and2_1 _07515_ (.A(\PWM.next_counter[0] ),
    .B(\PWM.final_sample_in[0] ),
    .X(_02235_));
 sky130_fd_sc_hd__a21bo_1 _07516_ (.A1(\PWM.final_sample_in[1] ),
    .A2(_02235_),
    .B1_N(\PWM.counter[1] ),
    .X(_02236_));
 sky130_fd_sc_hd__o221a_1 _07517_ (.A1(_02234_),
    .A2(\PWM.final_sample_in[2] ),
    .B1(\PWM.final_sample_in[1] ),
    .B2(_02235_),
    .C1(_02236_),
    .X(_02237_));
 sky130_fd_sc_hd__a221o_1 _07518_ (.A1(_02232_),
    .A2(\PWM.final_sample_in[3] ),
    .B1(\PWM.final_sample_in[2] ),
    .B2(_02234_),
    .C1(_02237_),
    .X(_02238_));
 sky130_fd_sc_hd__a22o_1 _07519_ (.A1(_01163_),
    .A2(\PWM.final_sample_in[4] ),
    .B1(_02233_),
    .B2(_02238_),
    .X(_02239_));
 sky130_fd_sc_hd__o221a_1 _07520_ (.A1(_02230_),
    .A2(\PWM.final_sample_in[5] ),
    .B1(\PWM.final_sample_in[4] ),
    .B2(_01163_),
    .C1(_02239_),
    .X(_02240_));
 sky130_fd_sc_hd__o22a_1 _07521_ (.A1(_02228_),
    .A2(\PWM.final_sample_in[6] ),
    .B1(_02231_),
    .B2(_02240_),
    .X(_02241_));
 sky130_fd_sc_hd__o22a_1 _07522_ (.A1(_02227_),
    .A2(net286),
    .B1(_02229_),
    .B2(_02241_),
    .X(_02242_));
 sky130_fd_sc_hd__a21o_1 _07523_ (.A1(_02227_),
    .A2(net286),
    .B1(_02242_),
    .X(\PWM.next_pwm_out ));
 sky130_fd_sc_hd__and3b_1 _07524_ (.A_N(_01152_),
    .B(\sig_norm.i[0] ),
    .C(\sig_norm.busy ),
    .X(_02243_));
 sky130_fd_sc_hd__inv_2 _07525_ (.A(_02243_),
    .Y(_02244_));
 sky130_fd_sc_hd__o211a_1 _07526_ (.A1(\sig_norm.busy ),
    .A2(net939),
    .B1(_01099_),
    .C1(_02244_),
    .X(_00026_));
 sky130_fd_sc_hd__nand2_1 _07527_ (.A(\sig_norm.i[1] ),
    .B(_02243_),
    .Y(_02245_));
 sky130_fd_sc_hd__a21o_1 _07528_ (.A1(\sig_norm.busy ),
    .A2(\sig_norm.i[0] ),
    .B1(\sig_norm.i[1] ),
    .X(_02246_));
 sky130_fd_sc_hd__and3_1 _07529_ (.A(_01099_),
    .B(_02245_),
    .C(_02246_),
    .X(_02247_));
 sky130_fd_sc_hd__clkbuf_1 _07530_ (.A(_02247_),
    .X(_00027_));
 sky130_fd_sc_hd__buf_4 _07531_ (.A(_01155_),
    .X(_02248_));
 sky130_fd_sc_hd__nor2_1 _07532_ (.A(_01151_),
    .B(_02245_),
    .Y(_02249_));
 sky130_fd_sc_hd__or2_1 _07533_ (.A(_02248_),
    .B(_02249_),
    .X(_02250_));
 sky130_fd_sc_hd__a21oi_1 _07534_ (.A1(_01151_),
    .A2(_02245_),
    .B1(_02250_),
    .Y(_00028_));
 sky130_fd_sc_hd__o21ai_1 _07535_ (.A1(net279),
    .A2(_02249_),
    .B1(_01099_),
    .Y(_02251_));
 sky130_fd_sc_hd__a21oi_1 _07536_ (.A1(net279),
    .A2(_02249_),
    .B1(_02251_),
    .Y(_00029_));
 sky130_fd_sc_hd__mux2_1 _07537_ (.A0(net1111),
    .A1(\PWM.final_in[0] ),
    .S(\PWM.start ),
    .X(_02252_));
 sky130_fd_sc_hd__clkbuf_1 _07538_ (.A(net1112),
    .X(_00030_));
 sky130_fd_sc_hd__mux2_1 _07539_ (.A0(\PWM.final_sample_in[1] ),
    .A1(net1103),
    .S(\PWM.start ),
    .X(_02253_));
 sky130_fd_sc_hd__clkbuf_1 _07540_ (.A(_02253_),
    .X(_00031_));
 sky130_fd_sc_hd__mux2_1 _07541_ (.A0(\PWM.final_sample_in[2] ),
    .A1(net1102),
    .S(\PWM.start ),
    .X(_02254_));
 sky130_fd_sc_hd__clkbuf_1 _07542_ (.A(_02254_),
    .X(_00032_));
 sky130_fd_sc_hd__mux2_1 _07543_ (.A0(\PWM.final_sample_in[3] ),
    .A1(net1172),
    .S(\PWM.start ),
    .X(_02255_));
 sky130_fd_sc_hd__clkbuf_1 _07544_ (.A(_02255_),
    .X(_00033_));
 sky130_fd_sc_hd__mux2_1 _07545_ (.A0(\PWM.final_sample_in[4] ),
    .A1(net1150),
    .S(\PWM.start ),
    .X(_02256_));
 sky130_fd_sc_hd__clkbuf_1 _07546_ (.A(_02256_),
    .X(_00034_));
 sky130_fd_sc_hd__mux2_1 _07547_ (.A0(\PWM.final_sample_in[5] ),
    .A1(net1168),
    .S(\PWM.start ),
    .X(_02257_));
 sky130_fd_sc_hd__clkbuf_1 _07548_ (.A(net1169),
    .X(_00035_));
 sky130_fd_sc_hd__mux2_1 _07549_ (.A0(net1157),
    .A1(net1132),
    .S(\PWM.start ),
    .X(_02258_));
 sky130_fd_sc_hd__clkbuf_1 _07550_ (.A(_02258_),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_1 _07551_ (.A0(net1142),
    .A1(net1128),
    .S(\PWM.start ),
    .X(_02259_));
 sky130_fd_sc_hd__clkbuf_1 _07552_ (.A(_02259_),
    .X(_00037_));
 sky130_fd_sc_hd__clkbuf_4 _07553_ (.A(_01157_),
    .X(_02260_));
 sky130_fd_sc_hd__buf_4 _07554_ (.A(_02223_),
    .X(_02261_));
 sky130_fd_sc_hd__or2_1 _07555_ (.A(\genblk2[9].wave_shpr.div.fin_quo[0] ),
    .B(\genblk2[9].wave_shpr.div.fin_quo[1] ),
    .X(_02262_));
 sky130_fd_sc_hd__or2_1 _07556_ (.A(\genblk2[9].wave_shpr.div.fin_quo[2] ),
    .B(_02262_),
    .X(_02263_));
 sky130_fd_sc_hd__or2_1 _07557_ (.A(\genblk2[9].wave_shpr.div.fin_quo[3] ),
    .B(_02263_),
    .X(_02264_));
 sky130_fd_sc_hd__or2_1 _07558_ (.A(\genblk2[9].wave_shpr.div.fin_quo[4] ),
    .B(_02264_),
    .X(_02265_));
 sky130_fd_sc_hd__a211o_1 _07559_ (.A1(_01200_),
    .A2(\genblk1[9].osc.clkdiv_C.cnt[14] ),
    .B1(_01361_),
    .C1(\genblk1[9].osc.clkdiv_C.cnt[15] ),
    .X(_02266_));
 sky130_fd_sc_hd__o22a_1 _07560_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[13] ),
    .A2(_01245_),
    .B1(_01328_),
    .B2(\genblk1[9].osc.clkdiv_C.cnt[12] ),
    .X(_02267_));
 sky130_fd_sc_hd__inv_2 _07561_ (.A(\genblk1[9].osc.clkdiv_C.cnt[10] ),
    .Y(_02268_));
 sky130_fd_sc_hd__a2bb2o_1 _07562_ (.A1_N(\genblk1[9].osc.clkdiv_C.cnt[11] ),
    .A2_N(_01799_),
    .B1(_01731_),
    .B2(_02268_),
    .X(_02269_));
 sky130_fd_sc_hd__a32o_1 _07563_ (.A1(_01930_),
    .A2(_01556_),
    .A3(_01564_),
    .B1(_01801_),
    .B2(_01928_),
    .X(_02270_));
 sky130_fd_sc_hd__o221a_1 _07564_ (.A1(_01930_),
    .A2(_01227_),
    .B1(_01732_),
    .B2(_02268_),
    .C1(_02270_),
    .X(_02271_));
 sky130_fd_sc_hd__a22oi_1 _07565_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[12] ),
    .A2(_01328_),
    .B1(_01799_),
    .B2(\genblk1[9].osc.clkdiv_C.cnt[11] ),
    .Y(_02272_));
 sky130_fd_sc_hd__o21ai_1 _07566_ (.A1(_02269_),
    .A2(_02271_),
    .B1(_02272_),
    .Y(_02273_));
 sky130_fd_sc_hd__o21a_1 _07567_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[14] ),
    .A2(_01936_),
    .B1(_01349_),
    .X(_02274_));
 sky130_fd_sc_hd__a2bb2o_1 _07568_ (.A1_N(\genblk1[9].osc.clkdiv_C.cnt[14] ),
    .A2_N(_01349_),
    .B1(_01246_),
    .B2(\genblk1[9].osc.clkdiv_C.cnt[13] ),
    .X(_02275_));
 sky130_fd_sc_hd__a211o_1 _07569_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[15] ),
    .A2(_01577_),
    .B1(_02274_),
    .C1(_02275_),
    .X(_02276_));
 sky130_fd_sc_hd__a21o_1 _07570_ (.A1(_02267_),
    .A2(_02273_),
    .B1(_02276_),
    .X(_02277_));
 sky130_fd_sc_hd__or3_1 _07571_ (.A(\genblk1[9].osc.clkdiv_C.cnt[4] ),
    .B(_01186_),
    .C(_01355_),
    .X(_02278_));
 sky130_fd_sc_hd__or4_1 _07572_ (.A(\genblk1[9].osc.clkdiv_C.cnt[5] ),
    .B(_01186_),
    .C(_01437_),
    .D(_01225_),
    .X(_02279_));
 sky130_fd_sc_hd__nand2_1 _07573_ (.A(_02278_),
    .B(_02279_),
    .Y(_02280_));
 sky130_fd_sc_hd__o31a_1 _07574_ (.A1(_01336_),
    .A2(_01437_),
    .A3(_01226_),
    .B1(\genblk1[9].osc.clkdiv_C.cnt[5] ),
    .X(_02281_));
 sky130_fd_sc_hd__a211o_1 _07575_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[4] ),
    .A2(_01925_),
    .B1(_02280_),
    .C1(_02281_),
    .X(_02282_));
 sky130_fd_sc_hd__a2bb2o_1 _07576_ (.A1_N(\genblk1[9].osc.clkdiv_C.cnt[6] ),
    .A2_N(_01512_),
    .B1(_01234_),
    .B2(\genblk1[9].osc.clkdiv_C.cnt[7] ),
    .X(_02283_));
 sky130_fd_sc_hd__and2_1 _07577_ (.A(\genblk1[9].osc.clkdiv_C.cnt[6] ),
    .B(_01512_),
    .X(_02284_));
 sky130_fd_sc_hd__or2_1 _07578_ (.A(\genblk1[9].osc.clkdiv_C.cnt[7] ),
    .B(_01234_),
    .X(_02285_));
 sky130_fd_sc_hd__or3b_1 _07579_ (.A(_02283_),
    .B(_02284_),
    .C_N(_02285_),
    .X(_02286_));
 sky130_fd_sc_hd__a21o_1 _07580_ (.A1(_01432_),
    .A2(_01221_),
    .B1(\genblk1[9].osc.clkdiv_C.cnt[1] ),
    .X(_02287_));
 sky130_fd_sc_hd__o311a_1 _07581_ (.A1(_01186_),
    .A2(_01437_),
    .A3(_01226_),
    .B1(_01171_),
    .C1(\genblk1[9].osc.clkdiv_C.cnt[0] ),
    .X(_02288_));
 sky130_fd_sc_hd__and3_1 _07582_ (.A(\genblk1[9].osc.clkdiv_C.cnt[1] ),
    .B(_01230_),
    .C(_01221_),
    .X(_02289_));
 sky130_fd_sc_hd__a221o_1 _07583_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[2] ),
    .A2(_01234_),
    .B1(_02287_),
    .B2(_02288_),
    .C1(_02289_),
    .X(_02290_));
 sky130_fd_sc_hd__o22a_1 _07584_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[2] ),
    .A2(_01234_),
    .B1(_01310_),
    .B2(\genblk1[9].osc.clkdiv_C.cnt[3] ),
    .X(_02291_));
 sky130_fd_sc_hd__a22o_1 _07585_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[3] ),
    .A2(_01311_),
    .B1(_02290_),
    .B2(_02291_),
    .X(_02292_));
 sky130_fd_sc_hd__a21o_1 _07586_ (.A1(_02278_),
    .A2(_02279_),
    .B1(_02281_),
    .X(_02293_));
 sky130_fd_sc_hd__a211o_1 _07587_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[7] ),
    .A2(_01234_),
    .B1(_01513_),
    .C1(\genblk1[9].osc.clkdiv_C.cnt[6] ),
    .X(_02294_));
 sky130_fd_sc_hd__o311a_1 _07588_ (.A1(_02284_),
    .A2(_02283_),
    .A3(_02293_),
    .B1(_02294_),
    .C1(_02285_),
    .X(_02295_));
 sky130_fd_sc_hd__o31a_1 _07589_ (.A1(_02282_),
    .A2(_02286_),
    .A3(_02292_),
    .B1(_02295_),
    .X(_02296_));
 sky130_fd_sc_hd__a22o_1 _07590_ (.A1(\genblk1[9].osc.clkdiv_C.cnt[9] ),
    .A2(_01991_),
    .B1(_01923_),
    .B2(\genblk1[9].osc.clkdiv_C.cnt[10] ),
    .X(_02297_));
 sky130_fd_sc_hd__nor2_1 _07591_ (.A(_01928_),
    .B(_01801_),
    .Y(_02298_));
 sky130_fd_sc_hd__and4bb_1 _07592_ (.A_N(_02298_),
    .B_N(_02269_),
    .C(_02272_),
    .D(_02267_),
    .X(_02299_));
 sky130_fd_sc_hd__or3b_1 _07593_ (.A(_02270_),
    .B(_02297_),
    .C_N(_02299_),
    .X(_02300_));
 sky130_fd_sc_hd__or3_1 _07594_ (.A(_02276_),
    .B(_02296_),
    .C(_02300_),
    .X(_02301_));
 sky130_fd_sc_hd__a311oi_4 _07595_ (.A1(_02266_),
    .A2(_02277_),
    .A3(_02301_),
    .B1(\genblk1[9].osc.clkdiv_C.cnt[17] ),
    .C1(\genblk1[9].osc.clkdiv_C.cnt[16] ),
    .Y(_02302_));
 sky130_fd_sc_hd__buf_2 _07596_ (.A(net32),
    .X(_02303_));
 sky130_fd_sc_hd__or3b_1 _07597_ (.A(_02265_),
    .B(\genblk2[9].wave_shpr.div.fin_quo[5] ),
    .C_N(_02303_),
    .X(_02304_));
 sky130_fd_sc_hd__xor2_1 _07598_ (.A(\genblk2[9].wave_shpr.div.fin_quo[6] ),
    .B(_02304_),
    .X(_02305_));
 sky130_fd_sc_hd__nor2_1 _07599_ (.A(_02261_),
    .B(_02305_),
    .Y(_02306_));
 sky130_fd_sc_hd__and2_2 _07600_ (.A(net17),
    .B(net18),
    .X(_02307_));
 sky130_fd_sc_hd__buf_4 _07601_ (.A(_02307_),
    .X(_02308_));
 sky130_fd_sc_hd__buf_4 _07602_ (.A(_02308_),
    .X(_02309_));
 sky130_fd_sc_hd__nor2_2 _07603_ (.A(_02221_),
    .B(net32),
    .Y(_02310_));
 sky130_fd_sc_hd__a21o_1 _07604_ (.A1(\genblk2[9].wave_shpr.div.fin_quo[7] ),
    .A2(_02309_),
    .B1(_02310_),
    .X(_02311_));
 sky130_fd_sc_hd__or2_2 _07605_ (.A(net17),
    .B(net18),
    .X(_02312_));
 sky130_fd_sc_hd__and3_1 _07606_ (.A(net15),
    .B(net163),
    .C(_02312_),
    .X(_02313_));
 sky130_fd_sc_hd__buf_2 _07607_ (.A(_02313_),
    .X(_02314_));
 sky130_fd_sc_hd__o21a_1 _07608_ (.A1(_02306_),
    .A2(_02311_),
    .B1(_02314_),
    .X(_02315_));
 sky130_fd_sc_hd__clkbuf_4 _07609_ (.A(_02222_),
    .X(_02316_));
 sky130_fd_sc_hd__nand2_1 _07610_ (.A(\genblk1[11].osc.clkdiv_C.cnt[7] ),
    .B(_01211_),
    .Y(_02317_));
 sky130_fd_sc_hd__o31a_1 _07611_ (.A1(_01186_),
    .A2(_01437_),
    .A3(_01225_),
    .B1(\genblk1[11].osc.clkdiv_C.cnt[2] ),
    .X(_02318_));
 sky130_fd_sc_hd__o21a_1 _07612_ (.A1(_01186_),
    .A2(_01354_),
    .B1(\genblk1[11].osc.clkdiv_C.cnt[1] ),
    .X(_02319_));
 sky130_fd_sc_hd__o311a_1 _07613_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[1] ),
    .A2(_01186_),
    .A3(_01354_),
    .B1(_01321_),
    .C1(\genblk1[11].osc.clkdiv_C.cnt[0] ),
    .X(_02320_));
 sky130_fd_sc_hd__a31o_1 _07614_ (.A1(_01171_),
    .A2(_01192_),
    .A3(_01208_),
    .B1(\genblk1[11].osc.clkdiv_C.cnt[3] ),
    .X(_02321_));
 sky130_fd_sc_hd__or4_1 _07615_ (.A(\genblk1[11].osc.clkdiv_C.cnt[2] ),
    .B(_01186_),
    .C(_01437_),
    .D(_01225_),
    .X(_02322_));
 sky130_fd_sc_hd__o311a_1 _07616_ (.A1(_02318_),
    .A2(_02319_),
    .A3(_02320_),
    .B1(_02321_),
    .C1(_02322_),
    .X(_02323_));
 sky130_fd_sc_hd__a22o_1 _07617_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[3] ),
    .A2(_01513_),
    .B1(_02064_),
    .B2(\genblk1[11].osc.clkdiv_C.cnt[4] ),
    .X(_02324_));
 sky130_fd_sc_hd__or2_1 _07618_ (.A(\genblk1[11].osc.clkdiv_C.cnt[4] ),
    .B(_02064_),
    .X(_02325_));
 sky130_fd_sc_hd__o221a_1 _07619_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[5] ),
    .A2(_01595_),
    .B1(_02323_),
    .B2(_02324_),
    .C1(_02325_),
    .X(_02326_));
 sky130_fd_sc_hd__a22o_1 _07620_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[6] ),
    .A2(_01430_),
    .B1(_01595_),
    .B2(\genblk1[11].osc.clkdiv_C.cnt[5] ),
    .X(_02327_));
 sky130_fd_sc_hd__o22ai_1 _07621_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[6] ),
    .A2(_01430_),
    .B1(_02326_),
    .B2(_02327_),
    .Y(_02328_));
 sky130_fd_sc_hd__nor2_1 _07622_ (.A(\genblk1[11].osc.clkdiv_C.cnt[7] ),
    .B(_01211_),
    .Y(_02329_));
 sky130_fd_sc_hd__a21oi_2 _07623_ (.A1(_02317_),
    .A2(_02328_),
    .B1(_02329_),
    .Y(_02330_));
 sky130_fd_sc_hd__o21a_1 _07624_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[14] ),
    .A2(_02085_),
    .B1(_01172_),
    .X(_02331_));
 sky130_fd_sc_hd__a22o_1 _07625_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[13] ),
    .A2(_01208_),
    .B1(_01576_),
    .B2(\genblk1[11].osc.clkdiv_C.cnt[15] ),
    .X(_02332_));
 sky130_fd_sc_hd__a211o_1 _07626_ (.A1(_02081_),
    .A2(_01241_),
    .B1(_02331_),
    .C1(_02332_),
    .X(_02333_));
 sky130_fd_sc_hd__o22ai_1 _07627_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[13] ),
    .A2(_01209_),
    .B1(_01256_),
    .B2(\genblk1[11].osc.clkdiv_C.cnt[12] ),
    .Y(_02334_));
 sky130_fd_sc_hd__a211o_1 _07628_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[12] ),
    .A2(_01256_),
    .B1(_02333_),
    .C1(_02334_),
    .X(_02335_));
 sky130_fd_sc_hd__nand2_4 _07629_ (.A(_01174_),
    .B(_01177_),
    .Y(_02336_));
 sky130_fd_sc_hd__and3_1 _07630_ (.A(\genblk1[11].osc.clkdiv_C.cnt[8] ),
    .B(_02336_),
    .C(net34),
    .X(_02337_));
 sky130_fd_sc_hd__or3_1 _07631_ (.A(_02128_),
    .B(_01179_),
    .C(_01249_),
    .X(_02338_));
 sky130_fd_sc_hd__a21bo_1 _07632_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[10] ),
    .A2(_01262_),
    .B1_N(_02338_),
    .X(_02339_));
 sky130_fd_sc_hd__a2bb2o_1 _07633_ (.A1_N(\genblk1[11].osc.clkdiv_C.cnt[10] ),
    .A2_N(_01262_),
    .B1(_01494_),
    .B2(_02128_),
    .X(_02340_));
 sky130_fd_sc_hd__a211o_1 _07634_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[9] ),
    .A2(_01190_),
    .B1(_02339_),
    .C1(_02340_),
    .X(_02341_));
 sky130_fd_sc_hd__o22a_1 _07635_ (.A1(\genblk1[11].osc.clkdiv_C.cnt[9] ),
    .A2(_01190_),
    .B1(_01235_),
    .B2(\genblk1[11].osc.clkdiv_C.cnt[8] ),
    .X(_02342_));
 sky130_fd_sc_hd__or3b_1 _07636_ (.A(_02337_),
    .B(_02341_),
    .C_N(_02342_),
    .X(_02343_));
 sky130_fd_sc_hd__o2bb2a_1 _07637_ (.A1_N(_02338_),
    .A2_N(_02340_),
    .B1(_02341_),
    .B2(_02342_),
    .X(_02344_));
 sky130_fd_sc_hd__o21ai_1 _07638_ (.A1(_01229_),
    .A2(_02081_),
    .B1(_02085_),
    .Y(_02345_));
 sky130_fd_sc_hd__or2b_1 _07639_ (.A(_02333_),
    .B_N(_02334_),
    .X(_02346_));
 sky130_fd_sc_hd__o211a_1 _07640_ (.A1(_02335_),
    .A2(_02344_),
    .B1(_02345_),
    .C1(_02346_),
    .X(_02347_));
 sky130_fd_sc_hd__o31ai_4 _07641_ (.A1(_02330_),
    .A2(_02335_),
    .A3(_02343_),
    .B1(_02347_),
    .Y(_02348_));
 sky130_fd_sc_hd__clkbuf_4 _07642_ (.A(net33),
    .X(_02349_));
 sky130_fd_sc_hd__nor2_4 _07643_ (.A(\genblk1[11].osc.clkdiv_C.cnt[16] ),
    .B(\genblk1[11].osc.clkdiv_C.cnt[17] ),
    .Y(_02350_));
 sky130_fd_sc_hd__buf_2 _07644_ (.A(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__or2_1 _07645_ (.A(\genblk2[11].wave_shpr.div.fin_quo[0] ),
    .B(\genblk2[11].wave_shpr.div.fin_quo[1] ),
    .X(_02352_));
 sky130_fd_sc_hd__or2_1 _07646_ (.A(\genblk2[11].wave_shpr.div.fin_quo[2] ),
    .B(_02352_),
    .X(_02353_));
 sky130_fd_sc_hd__or2_1 _07647_ (.A(\genblk2[11].wave_shpr.div.fin_quo[3] ),
    .B(_02353_),
    .X(_02354_));
 sky130_fd_sc_hd__or2_1 _07648_ (.A(\genblk2[11].wave_shpr.div.fin_quo[4] ),
    .B(_02354_),
    .X(_02355_));
 sky130_fd_sc_hd__nor2_1 _07649_ (.A(\genblk2[11].wave_shpr.div.fin_quo[5] ),
    .B(_02355_),
    .Y(_02356_));
 sky130_fd_sc_hd__and4_1 _07650_ (.A(\genblk2[11].wave_shpr.div.fin_quo[6] ),
    .B(_02349_),
    .C(_02351_),
    .D(_02356_),
    .X(_02357_));
 sky130_fd_sc_hd__a31o_1 _07651_ (.A1(_02349_),
    .A2(_02351_),
    .A3(_02356_),
    .B1(\genblk2[11].wave_shpr.div.fin_quo[6] ),
    .X(_02358_));
 sky130_fd_sc_hd__or3b_1 _07652_ (.A(_02316_),
    .B(_02357_),
    .C_N(_02358_),
    .X(_02359_));
 sky130_fd_sc_hd__a21o_1 _07653_ (.A1(_02349_),
    .A2(_02351_),
    .B1(_02221_),
    .X(_02360_));
 sky130_fd_sc_hd__buf_4 _07654_ (.A(_02307_),
    .X(_02361_));
 sky130_fd_sc_hd__clkbuf_4 _07655_ (.A(_02361_),
    .X(_02362_));
 sky130_fd_sc_hd__nand2_1 _07656_ (.A(\genblk2[11].wave_shpr.div.fin_quo[7] ),
    .B(_02362_),
    .Y(_02363_));
 sky130_fd_sc_hd__clkbuf_4 _07657_ (.A(net136),
    .X(_02364_));
 sky130_fd_sc_hd__clkbuf_4 _07658_ (.A(_02312_),
    .X(_02365_));
 sky130_fd_sc_hd__nand3_2 _07659_ (.A(net3),
    .B(_02364_),
    .C(_02365_),
    .Y(_02366_));
 sky130_fd_sc_hd__a31o_1 _07660_ (.A1(_02359_),
    .A2(_02360_),
    .A3(_02363_),
    .B1(_02366_),
    .X(_02367_));
 sky130_fd_sc_hd__o22ai_1 _07661_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[7] ),
    .A2(_01190_),
    .B1(_01235_),
    .B2(\genblk1[10].osc.clkdiv_C.cnt[6] ),
    .Y(_02368_));
 sky130_fd_sc_hd__or2_1 _07662_ (.A(\genblk1[10].osc.clkdiv_C.cnt[5] ),
    .B(_01182_),
    .X(_02369_));
 sky130_fd_sc_hd__a211o_1 _07663_ (.A1(_01360_),
    .A2(_01224_),
    .B1(_01241_),
    .C1(\genblk1[10].osc.clkdiv_C.cnt[4] ),
    .X(_02370_));
 sky130_fd_sc_hd__a32o_1 _07664_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[6] ),
    .A2(_02336_),
    .A3(_01794_),
    .B1(\genblk1[10].osc.clkdiv_C.cnt[5] ),
    .B2(_01182_),
    .X(_02371_));
 sky130_fd_sc_hd__a21oi_1 _07665_ (.A1(_02369_),
    .A2(_02370_),
    .B1(_02371_),
    .Y(_02372_));
 sky130_fd_sc_hd__a2bb2o_1 _07666_ (.A1_N(_02368_),
    .A2_N(_02372_),
    .B1(\genblk1[10].osc.clkdiv_C.cnt[7] ),
    .B2(_01190_),
    .X(_02373_));
 sky130_fd_sc_hd__nor2_4 _07667_ (.A(_01308_),
    .B(_01187_),
    .Y(_02374_));
 sky130_fd_sc_hd__o22a_1 _07668_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[3] ),
    .A2(_02374_),
    .B1(_02013_),
    .B2(\genblk1[10].osc.clkdiv_C.cnt[2] ),
    .X(_02375_));
 sky130_fd_sc_hd__and3_1 _07669_ (.A(_01188_),
    .B(_01440_),
    .C(\genblk1[10].osc.clkdiv_C.cnt[3] ),
    .X(_02376_));
 sky130_fd_sc_hd__or2_1 _07670_ (.A(_02375_),
    .B(_02376_),
    .X(_02377_));
 sky130_fd_sc_hd__and2_1 _07671_ (.A(_01308_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[1] ),
    .X(_02378_));
 sky130_fd_sc_hd__or2_1 _07672_ (.A(_01308_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[1] ),
    .X(_02379_));
 sky130_fd_sc_hd__a32o_1 _07673_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[0] ),
    .A2(_02001_),
    .A3(_02379_),
    .B1(_02013_),
    .B2(\genblk1[10].osc.clkdiv_C.cnt[2] ),
    .X(_02380_));
 sky130_fd_sc_hd__or4b_1 _07674_ (.A(_02378_),
    .B(_02376_),
    .C(_02380_),
    .D_N(_02375_),
    .X(_02381_));
 sky130_fd_sc_hd__nand2_1 _07675_ (.A(_02369_),
    .B(_02370_),
    .Y(_02382_));
 sky130_fd_sc_hd__a221o_1 _07676_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[7] ),
    .A2(_01190_),
    .B1(_01992_),
    .B2(\genblk1[10].osc.clkdiv_C.cnt[4] ),
    .C1(_02371_),
    .X(_02383_));
 sky130_fd_sc_hd__a2111o_1 _07677_ (.A1(_02377_),
    .A2(_02381_),
    .B1(_02368_),
    .C1(_02382_),
    .D1(_02383_),
    .X(_02384_));
 sky130_fd_sc_hd__a2bb2o_1 _07678_ (.A1_N(\genblk1[10].osc.clkdiv_C.cnt[9] ),
    .A2_N(_01215_),
    .B1(_01991_),
    .B2(_02003_),
    .X(_02385_));
 sky130_fd_sc_hd__nor2_1 _07679_ (.A(_01489_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[13] ),
    .Y(_02386_));
 sky130_fd_sc_hd__nand2_1 _07680_ (.A(_01181_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[12] ),
    .Y(_02387_));
 sky130_fd_sc_hd__inv_2 _07681_ (.A(_02387_),
    .Y(_02388_));
 sky130_fd_sc_hd__a21oi_1 _07682_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[13] ),
    .A2(_01246_),
    .B1(_02386_),
    .Y(_02389_));
 sky130_fd_sc_hd__nand2_1 _07683_ (.A(_01174_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[14] ),
    .Y(_02390_));
 sky130_fd_sc_hd__mux2_1 _07684_ (.A0(_01179_),
    .A1(_01575_),
    .S(\genblk1[10].osc.clkdiv_C.cnt[15] ),
    .X(_02391_));
 sky130_fd_sc_hd__o2bb2a_1 _07685_ (.A1_N(_02390_),
    .A2_N(_02391_),
    .B1(_01995_),
    .B2(_02016_),
    .X(_02392_));
 sky130_fd_sc_hd__o221a_1 _07686_ (.A1(_02023_),
    .A2(_02386_),
    .B1(_02388_),
    .B2(_02389_),
    .C1(_02392_),
    .X(_02393_));
 sky130_fd_sc_hd__o22ai_2 _07687_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[11] ),
    .A2(_02011_),
    .B1(_02005_),
    .B2(\genblk1[10].osc.clkdiv_C.cnt[10] ),
    .Y(_02394_));
 sky130_fd_sc_hd__a22o_1 _07688_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[9] ),
    .A2(_01215_),
    .B1(_02011_),
    .B2(\genblk1[10].osc.clkdiv_C.cnt[11] ),
    .X(_02395_));
 sky130_fd_sc_hd__a211oi_1 _07689_ (.A1(\genblk1[10].osc.clkdiv_C.cnt[10] ),
    .A2(_02005_),
    .B1(_02394_),
    .C1(_02395_),
    .Y(_02396_));
 sky130_fd_sc_hd__o211ai_1 _07690_ (.A1(_02003_),
    .A2(_01991_),
    .B1(_02393_),
    .C1(_02396_),
    .Y(_02397_));
 sky130_fd_sc_hd__a211o_1 _07691_ (.A1(_02373_),
    .A2(_02384_),
    .B1(_02385_),
    .C1(_02397_),
    .X(_02398_));
 sky130_fd_sc_hd__nand2_1 _07692_ (.A(\genblk1[10].osc.clkdiv_C.cnt[11] ),
    .B(_02011_),
    .Y(_02399_));
 sky130_fd_sc_hd__a22o_1 _07693_ (.A1(_02399_),
    .A2(_02394_),
    .B1(_02385_),
    .B2(_02396_),
    .X(_02400_));
 sky130_fd_sc_hd__and3_1 _07694_ (.A(_02386_),
    .B(_02392_),
    .C(_02387_),
    .X(_02401_));
 sky130_fd_sc_hd__a221oi_2 _07695_ (.A1(_02016_),
    .A2(_02390_),
    .B1(_02393_),
    .B2(_02400_),
    .C1(_02401_),
    .Y(_02402_));
 sky130_fd_sc_hd__a211o_4 _07696_ (.A1(_02398_),
    .A2(_02402_),
    .B1(\genblk1[10].osc.clkdiv_C.cnt[16] ),
    .C1(\genblk1[10].osc.clkdiv_C.cnt[17] ),
    .X(_02403_));
 sky130_fd_sc_hd__buf_2 _07697_ (.A(_02403_),
    .X(_02404_));
 sky130_fd_sc_hd__inv_2 _07698_ (.A(\genblk2[10].wave_shpr.div.fin_quo[5] ),
    .Y(_02405_));
 sky130_fd_sc_hd__inv_2 _07699_ (.A(\genblk2[10].wave_shpr.div.fin_quo[3] ),
    .Y(_02406_));
 sky130_fd_sc_hd__nor2_1 _07700_ (.A(\genblk2[10].wave_shpr.div.fin_quo[0] ),
    .B(\genblk2[10].wave_shpr.div.fin_quo[1] ),
    .Y(_02407_));
 sky130_fd_sc_hd__and2b_1 _07701_ (.A_N(\genblk2[10].wave_shpr.div.fin_quo[2] ),
    .B(_02407_),
    .X(_02408_));
 sky130_fd_sc_hd__nand2_1 _07702_ (.A(_02406_),
    .B(_02408_),
    .Y(_02409_));
 sky130_fd_sc_hd__nor2_1 _07703_ (.A(\genblk2[10].wave_shpr.div.fin_quo[4] ),
    .B(_02409_),
    .Y(_02410_));
 sky130_fd_sc_hd__and4b_1 _07704_ (.A_N(_02404_),
    .B(_02405_),
    .C(\genblk2[10].wave_shpr.div.fin_quo[6] ),
    .D(_02410_),
    .X(_02411_));
 sky130_fd_sc_hd__inv_2 _07705_ (.A(\genblk2[10].wave_shpr.div.fin_quo[6] ),
    .Y(_02412_));
 sky130_fd_sc_hd__o41a_1 _07706_ (.A1(\genblk2[10].wave_shpr.div.fin_quo[4] ),
    .A2(\genblk2[10].wave_shpr.div.fin_quo[5] ),
    .A3(_02404_),
    .A4(_02409_),
    .B1(_02412_),
    .X(_02413_));
 sky130_fd_sc_hd__or3_1 _07707_ (.A(_02316_),
    .B(_02411_),
    .C(_02413_),
    .X(_02414_));
 sky130_fd_sc_hd__and2_1 _07708_ (.A(_02225_),
    .B(_02403_),
    .X(_02415_));
 sky130_fd_sc_hd__buf_2 _07709_ (.A(_02415_),
    .X(_02416_));
 sky130_fd_sc_hd__a21oi_1 _07710_ (.A1(\genblk2[10].wave_shpr.div.fin_quo[7] ),
    .A2(_02362_),
    .B1(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__and3_1 _07711_ (.A(net2),
    .B(net163),
    .C(_02312_),
    .X(_02418_));
 sky130_fd_sc_hd__buf_2 _07712_ (.A(_02418_),
    .X(_02419_));
 sky130_fd_sc_hd__a21bo_1 _07713_ (.A1(_02414_),
    .A2(_02417_),
    .B1_N(_02419_),
    .X(_02420_));
 sky130_fd_sc_hd__xor2_1 _07714_ (.A(_02367_),
    .B(_02420_),
    .X(_02421_));
 sky130_fd_sc_hd__nor2_1 _07715_ (.A(_02367_),
    .B(_02420_),
    .Y(_02422_));
 sky130_fd_sc_hd__a21o_1 _07716_ (.A1(_02315_),
    .A2(_02421_),
    .B1(_02422_),
    .X(_02423_));
 sky130_fd_sc_hd__nand3_2 _07717_ (.A(net7),
    .B(_02364_),
    .C(_02365_),
    .Y(_02424_));
 sky130_fd_sc_hd__nand2_4 _07718_ (.A(_01360_),
    .B(_01302_),
    .Y(_02425_));
 sky130_fd_sc_hd__o22ai_2 _07719_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[15] ),
    .A2(_01309_),
    .B1(_01209_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[14] ),
    .Y(_02426_));
 sky130_fd_sc_hd__a22o_1 _07720_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[15] ),
    .A2(_01309_),
    .B1(_01208_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[14] ),
    .X(_02427_));
 sky130_fd_sc_hd__a211oi_2 _07721_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[13] ),
    .A2(_02425_),
    .B1(_02426_),
    .C1(_02427_),
    .Y(_02428_));
 sky130_fd_sc_hd__o211ai_1 _07722_ (.A1(_01330_),
    .A2(_01262_),
    .B1(_01591_),
    .C1(_01172_),
    .Y(_02429_));
 sky130_fd_sc_hd__a22o_1 _07723_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[2] ),
    .A2(_01323_),
    .B1(_02429_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[1] ),
    .X(_02430_));
 sky130_fd_sc_hd__o22a_1 _07724_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[2] ),
    .A2(_01323_),
    .B1(_01313_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[3] ),
    .X(_02431_));
 sky130_fd_sc_hd__a22o_1 _07725_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[4] ),
    .A2(_01305_),
    .B1(_01313_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[3] ),
    .X(_02432_));
 sky130_fd_sc_hd__nor2_4 _07726_ (.A(_01342_),
    .B(_01241_),
    .Y(_02433_));
 sky130_fd_sc_hd__o22ai_1 _07727_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[5] ),
    .A2(_02433_),
    .B1(_01305_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[4] ),
    .Y(_02434_));
 sky130_fd_sc_hd__nor2_1 _07728_ (.A(_01342_),
    .B(\genblk1[1].osc.clkdiv_C.cnt[7] ),
    .Y(_02435_));
 sky130_fd_sc_hd__a21oi_1 _07729_ (.A1(_01360_),
    .A2(net37),
    .B1(\genblk1[1].osc.clkdiv_C.cnt[6] ),
    .Y(_02436_));
 sky130_fd_sc_hd__and2_1 _07730_ (.A(_01188_),
    .B(\genblk1[1].osc.clkdiv_C.cnt[7] ),
    .X(_02437_));
 sky130_fd_sc_hd__a31o_1 _07731_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[6] ),
    .A2(_01360_),
    .A3(net37),
    .B1(_02437_),
    .X(_02438_));
 sky130_fd_sc_hd__a2111o_1 _07732_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[5] ),
    .A2(_02433_),
    .B1(_02435_),
    .C1(_02436_),
    .D1(_02438_),
    .X(_02439_));
 sky130_fd_sc_hd__a2111o_1 _07733_ (.A1(_02430_),
    .A2(_02431_),
    .B1(_02432_),
    .C1(_02434_),
    .D1(_02439_),
    .X(_02440_));
 sky130_fd_sc_hd__nor2_1 _07734_ (.A(_02435_),
    .B(_02436_),
    .Y(_02441_));
 sky130_fd_sc_hd__o22a_1 _07735_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[5] ),
    .A2(_02433_),
    .B1(_01305_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[4] ),
    .X(_02442_));
 sky130_fd_sc_hd__o22a_1 _07736_ (.A1(_02441_),
    .A2(_02437_),
    .B1(_02439_),
    .B2(_02442_),
    .X(_02443_));
 sky130_fd_sc_hd__inv_2 _07737_ (.A(\genblk1[1].osc.clkdiv_C.cnt[8] ),
    .Y(_02444_));
 sky130_fd_sc_hd__nor2_1 _07738_ (.A(_02444_),
    .B(_02013_),
    .Y(_02445_));
 sky130_fd_sc_hd__a22o_1 _07739_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[9] ),
    .A2(_01334_),
    .B1(_01312_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[10] ),
    .X(_02446_));
 sky130_fd_sc_hd__o22a_1 _07740_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[9] ),
    .A2(_01334_),
    .B1(_01356_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[8] ),
    .X(_02447_));
 sky130_fd_sc_hd__o22a_1 _07741_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[11] ),
    .A2(_01337_),
    .B1(_01312_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[10] ),
    .X(_02448_));
 sky130_fd_sc_hd__or4bb_1 _07742_ (.A(_02445_),
    .B(_02446_),
    .C_N(_02447_),
    .D_N(_02448_),
    .X(_02449_));
 sky130_fd_sc_hd__a21oi_1 _07743_ (.A1(_02440_),
    .A2(_02443_),
    .B1(_02449_),
    .Y(_02450_));
 sky130_fd_sc_hd__o22ai_2 _07744_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[13] ),
    .A2(_02425_),
    .B1(_01344_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[12] ),
    .Y(_02451_));
 sky130_fd_sc_hd__a221oi_2 _07745_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[12] ),
    .A2(_01344_),
    .B1(_01337_),
    .B2(\genblk1[1].osc.clkdiv_C.cnt[11] ),
    .C1(_02451_),
    .Y(_02452_));
 sky130_fd_sc_hd__o21ai_1 _07746_ (.A1(_02447_),
    .A2(_02446_),
    .B1(_02448_),
    .Y(_02453_));
 sky130_fd_sc_hd__nand2_1 _07747_ (.A(\genblk1[1].osc.clkdiv_C.cnt[15] ),
    .B(_01172_),
    .Y(_02454_));
 sky130_fd_sc_hd__nor2_1 _07748_ (.A(\genblk1[1].osc.clkdiv_C.cnt[16] ),
    .B(_01576_),
    .Y(_02455_));
 sky130_fd_sc_hd__a221o_1 _07749_ (.A1(_02426_),
    .A2(_02454_),
    .B1(_02428_),
    .B2(_02451_),
    .C1(_02455_),
    .X(_02456_));
 sky130_fd_sc_hd__a31o_1 _07750_ (.A1(_02428_),
    .A2(_02453_),
    .A3(_02452_),
    .B1(_02456_),
    .X(_02457_));
 sky130_fd_sc_hd__a31o_4 _07751_ (.A1(_02428_),
    .A2(_02450_),
    .A3(_02452_),
    .B1(_02457_),
    .X(_02458_));
 sky130_fd_sc_hd__a21oi_4 _07752_ (.A1(\genblk1[1].osc.clkdiv_C.cnt[16] ),
    .A2(_01577_),
    .B1(\genblk1[1].osc.clkdiv_C.cnt[17] ),
    .Y(_02459_));
 sky130_fd_sc_hd__and2_1 _07753_ (.A(_02458_),
    .B(_02459_),
    .X(_02460_));
 sky130_fd_sc_hd__clkbuf_2 _07754_ (.A(_02460_),
    .X(_02461_));
 sky130_fd_sc_hd__or2_1 _07755_ (.A(\genblk2[1].wave_shpr.div.fin_quo[0] ),
    .B(\genblk2[1].wave_shpr.div.fin_quo[1] ),
    .X(_02462_));
 sky130_fd_sc_hd__or3_1 _07756_ (.A(\genblk2[1].wave_shpr.div.fin_quo[2] ),
    .B(\genblk2[1].wave_shpr.div.fin_quo[3] ),
    .C(_02462_),
    .X(_02463_));
 sky130_fd_sc_hd__or2_1 _07757_ (.A(\genblk2[1].wave_shpr.div.fin_quo[4] ),
    .B(_02463_),
    .X(_02464_));
 sky130_fd_sc_hd__a21oi_1 _07758_ (.A1(_02461_),
    .A2(_02464_),
    .B1(\genblk2[1].wave_shpr.div.fin_quo[5] ),
    .Y(_02465_));
 sky130_fd_sc_hd__a31o_1 _07759_ (.A1(\genblk2[1].wave_shpr.div.fin_quo[5] ),
    .A2(_02461_),
    .A3(_02464_),
    .B1(_02224_),
    .X(_02466_));
 sky130_fd_sc_hd__clkbuf_4 _07760_ (.A(_02362_),
    .X(_02467_));
 sky130_fd_sc_hd__clkbuf_4 _07761_ (.A(_02467_),
    .X(_02468_));
 sky130_fd_sc_hd__a21oi_4 _07762_ (.A1(_02458_),
    .A2(_02459_),
    .B1(_02220_),
    .Y(_02469_));
 sky130_fd_sc_hd__a21oi_1 _07763_ (.A1(\genblk2[1].wave_shpr.div.fin_quo[6] ),
    .A2(_02468_),
    .B1(_02469_),
    .Y(_02470_));
 sky130_fd_sc_hd__o21a_1 _07764_ (.A1(_02465_),
    .A2(_02466_),
    .B1(_02470_),
    .X(_02471_));
 sky130_fd_sc_hd__a22o_1 _07765_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[15] ),
    .A2(_01309_),
    .B1(_01208_),
    .B2(\genblk1[0].osc.clkdiv_C.cnt[14] ),
    .X(_02472_));
 sky130_fd_sc_hd__and2_1 _07766_ (.A(\genblk1[0].osc.clkdiv_C.cnt[13] ),
    .B(_01255_),
    .X(_02473_));
 sky130_fd_sc_hd__o22a_1 _07767_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[15] ),
    .A2(_01309_),
    .B1(_01208_),
    .B2(\genblk1[0].osc.clkdiv_C.cnt[14] ),
    .X(_02474_));
 sky130_fd_sc_hd__or3b_1 _07768_ (.A(_02472_),
    .B(_02473_),
    .C_N(_02474_),
    .X(_02475_));
 sky130_fd_sc_hd__o22a_1 _07769_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[13] ),
    .A2(_01256_),
    .B1(_01240_),
    .B2(\genblk1[0].osc.clkdiv_C.cnt[12] ),
    .X(_02476_));
 sky130_fd_sc_hd__a21bo_1 _07770_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[12] ),
    .A2(_01240_),
    .B1_N(_02476_),
    .X(_02477_));
 sky130_fd_sc_hd__or2_1 _07771_ (.A(_02475_),
    .B(_02477_),
    .X(_02478_));
 sky130_fd_sc_hd__o2111a_1 _07772_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[1] ),
    .A2(_01190_),
    .B1(net34),
    .C1(\genblk1[0].osc.clkdiv_C.cnt[0] ),
    .D1(_02336_),
    .X(_02479_));
 sky130_fd_sc_hd__a32o_1 _07773_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[2] ),
    .A2(_01556_),
    .A3(_01564_),
    .B1(_01190_),
    .B2(\genblk1[0].osc.clkdiv_C.cnt[1] ),
    .X(_02480_));
 sky130_fd_sc_hd__or2_1 _07774_ (.A(\genblk1[0].osc.clkdiv_C.cnt[3] ),
    .B(_01215_),
    .X(_02481_));
 sky130_fd_sc_hd__o221a_1 _07775_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[2] ),
    .A2(_01227_),
    .B1(_02479_),
    .B2(_02480_),
    .C1(_02481_),
    .X(_02482_));
 sky130_fd_sc_hd__nand2_1 _07776_ (.A(_01229_),
    .B(_01359_),
    .Y(_02483_));
 sky130_fd_sc_hd__xnor2_1 _07777_ (.A(\genblk1[0].osc.clkdiv_C.cnt[4] ),
    .B(_01258_),
    .Y(_02484_));
 sky130_fd_sc_hd__a21oi_1 _07778_ (.A1(_01181_),
    .A2(\genblk1[0].osc.clkdiv_C.cnt[7] ),
    .B1(_01198_),
    .Y(_02485_));
 sky130_fd_sc_hd__o21ai_1 _07779_ (.A1(_01181_),
    .A2(\genblk1[0].osc.clkdiv_C.cnt[7] ),
    .B1(_02485_),
    .Y(_02486_));
 sky130_fd_sc_hd__a2bb2o_1 _07780_ (.A1_N(\genblk1[0].osc.clkdiv_C.cnt[5] ),
    .A2_N(_02483_),
    .B1(_01215_),
    .B2(\genblk1[0].osc.clkdiv_C.cnt[3] ),
    .X(_02487_));
 sky130_fd_sc_hd__a2111o_1 _07781_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[5] ),
    .A2(_02483_),
    .B1(_02484_),
    .C1(_02486_),
    .D1(_02487_),
    .X(_02488_));
 sky130_fd_sc_hd__o21a_1 _07782_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[4] ),
    .A2(_01241_),
    .B1(_02483_),
    .X(_02489_));
 sky130_fd_sc_hd__a21o_1 _07783_ (.A1(_01200_),
    .A2(\genblk1[0].osc.clkdiv_C.cnt[6] ),
    .B1(\genblk1[0].osc.clkdiv_C.cnt[7] ),
    .X(_02490_));
 sky130_fd_sc_hd__o31ai_1 _07784_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[5] ),
    .A2(_02486_),
    .A3(_02489_),
    .B1(_02490_),
    .Y(_02491_));
 sky130_fd_sc_hd__o21ba_1 _07785_ (.A1(_02482_),
    .A2(_02488_),
    .B1_N(_02491_),
    .X(_02492_));
 sky130_fd_sc_hd__o22ai_1 _07786_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[8] ),
    .A2(_01193_),
    .B1(_01184_),
    .B2(\genblk1[0].osc.clkdiv_C.cnt[9] ),
    .Y(_02493_));
 sky130_fd_sc_hd__a22o_1 _07787_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[8] ),
    .A2(_01193_),
    .B1(_01184_),
    .B2(\genblk1[0].osc.clkdiv_C.cnt[9] ),
    .X(_02494_));
 sky130_fd_sc_hd__or2_1 _07788_ (.A(_02493_),
    .B(_02494_),
    .X(_02495_));
 sky130_fd_sc_hd__or2_1 _07789_ (.A(\genblk1[0].osc.clkdiv_C.cnt[11] ),
    .B(_01263_),
    .X(_02496_));
 sky130_fd_sc_hd__or3_1 _07790_ (.A(\genblk1[0].osc.clkdiv_C.cnt[10] ),
    .B(_01996_),
    .C(_01801_),
    .X(_02497_));
 sky130_fd_sc_hd__nand2_1 _07791_ (.A(\genblk1[0].osc.clkdiv_C.cnt[11] ),
    .B(_01263_),
    .Y(_02498_));
 sky130_fd_sc_hd__a31o_1 _07792_ (.A1(_01246_),
    .A2(_01439_),
    .A3(_01344_),
    .B1(_01169_),
    .X(_02499_));
 sky130_fd_sc_hd__and4_1 _07793_ (.A(_02496_),
    .B(_02497_),
    .C(_02498_),
    .D(_02499_),
    .X(_02500_));
 sky130_fd_sc_hd__or4b_1 _07794_ (.A(_02478_),
    .B(_02492_),
    .C(_02495_),
    .D_N(_02500_),
    .X(_02501_));
 sky130_fd_sc_hd__nand2_1 _07795_ (.A(\genblk1[0].osc.clkdiv_C.cnt[9] ),
    .B(_01184_),
    .Y(_02502_));
 sky130_fd_sc_hd__nand2_1 _07796_ (.A(_02496_),
    .B(_02497_),
    .Y(_02503_));
 sky130_fd_sc_hd__a32oi_1 _07797_ (.A1(_02493_),
    .A2(_02500_),
    .A3(_02502_),
    .B1(_02498_),
    .B2(_02503_),
    .Y(_02504_));
 sky130_fd_sc_hd__or3_1 _07798_ (.A(\genblk1[0].osc.clkdiv_C.cnt[15] ),
    .B(\genblk1[0].osc.clkdiv_C.cnt[14] ),
    .C(_01209_),
    .X(_02505_));
 sky130_fd_sc_hd__o221a_1 _07799_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[15] ),
    .A2(_01349_),
    .B1(_01577_),
    .B2(\genblk1[0].osc.clkdiv_C.cnt[16] ),
    .C1(_02505_),
    .X(_02506_));
 sky130_fd_sc_hd__o221a_1 _07800_ (.A1(_02475_),
    .A2(_02476_),
    .B1(_02478_),
    .B2(_02504_),
    .C1(_02506_),
    .X(_02507_));
 sky130_fd_sc_hd__a221oi_2 _07801_ (.A1(\genblk1[0].osc.clkdiv_C.cnt[16] ),
    .A2(_01577_),
    .B1(_02501_),
    .B2(_02507_),
    .C1(\genblk1[0].osc.clkdiv_C.cnt[17] ),
    .Y(_02508_));
 sky130_fd_sc_hd__nor2_2 _07802_ (.A(_02221_),
    .B(net31),
    .Y(_02509_));
 sky130_fd_sc_hd__buf_2 _07803_ (.A(net31),
    .X(_02510_));
 sky130_fd_sc_hd__or3_1 _07804_ (.A(\genblk2[0].wave_shpr.div.fin_quo[0] ),
    .B(\genblk2[0].wave_shpr.div.fin_quo[1] ),
    .C(\genblk2[0].wave_shpr.div.fin_quo[2] ),
    .X(_02511_));
 sky130_fd_sc_hd__or2_1 _07805_ (.A(\genblk2[0].wave_shpr.div.fin_quo[3] ),
    .B(_02511_),
    .X(_02512_));
 sky130_fd_sc_hd__or2_1 _07806_ (.A(\genblk2[0].wave_shpr.div.fin_quo[4] ),
    .B(_02512_),
    .X(_02513_));
 sky130_fd_sc_hd__a21oi_1 _07807_ (.A1(_02510_),
    .A2(_02513_),
    .B1(\genblk2[0].wave_shpr.div.fin_quo[5] ),
    .Y(_02514_));
 sky130_fd_sc_hd__a31o_1 _07808_ (.A1(\genblk2[0].wave_shpr.div.fin_quo[5] ),
    .A2(_02510_),
    .A3(_02513_),
    .B1(_02224_),
    .X(_02515_));
 sky130_fd_sc_hd__a2bb2o_1 _07809_ (.A1_N(_02514_),
    .A2_N(_02515_),
    .B1(\genblk2[0].wave_shpr.div.fin_quo[6] ),
    .B2(_02468_),
    .X(_02516_));
 sky130_fd_sc_hd__and3_1 _07810_ (.A(net1),
    .B(net150),
    .C(_02312_),
    .X(_02517_));
 sky130_fd_sc_hd__buf_2 _07811_ (.A(_02517_),
    .X(_02518_));
 sky130_fd_sc_hd__o21ai_1 _07812_ (.A1(_02509_),
    .A2(_02516_),
    .B1(_02518_),
    .Y(_02519_));
 sky130_fd_sc_hd__nor3_2 _07813_ (.A(_02424_),
    .B(_02471_),
    .C(_02519_),
    .Y(_02520_));
 sky130_fd_sc_hd__buf_4 _07814_ (.A(_02308_),
    .X(_02521_));
 sky130_fd_sc_hd__o21a_1 _07815_ (.A1(\genblk2[1].wave_shpr.div.fin_quo[2] ),
    .A2(_02462_),
    .B1(_02461_),
    .X(_02522_));
 sky130_fd_sc_hd__xor2_1 _07816_ (.A(\genblk2[1].wave_shpr.div.fin_quo[3] ),
    .B(_02522_),
    .X(_02523_));
 sky130_fd_sc_hd__and2b_2 _07817_ (.A_N(net17),
    .B(net18),
    .X(_02524_));
 sky130_fd_sc_hd__clkbuf_4 _07818_ (.A(_02524_),
    .X(_02525_));
 sky130_fd_sc_hd__clkbuf_4 _07819_ (.A(_02525_),
    .X(_02526_));
 sky130_fd_sc_hd__clkbuf_4 _07820_ (.A(_02526_),
    .X(_02527_));
 sky130_fd_sc_hd__a22o_1 _07821_ (.A1(\genblk2[1].wave_shpr.div.fin_quo[4] ),
    .A2(_02521_),
    .B1(_02523_),
    .B2(_02527_),
    .X(_02528_));
 sky130_fd_sc_hd__and3_2 _07822_ (.A(net7),
    .B(net150),
    .C(_02312_),
    .X(_02529_));
 sky130_fd_sc_hd__o21ai_1 _07823_ (.A1(_02469_),
    .A2(_02528_),
    .B1(_02529_),
    .Y(_02530_));
 sky130_fd_sc_hd__a21oi_1 _07824_ (.A1(_02510_),
    .A2(_02511_),
    .B1(\genblk2[0].wave_shpr.div.fin_quo[3] ),
    .Y(_02531_));
 sky130_fd_sc_hd__a31o_1 _07825_ (.A1(\genblk2[0].wave_shpr.div.fin_quo[3] ),
    .A2(_02510_),
    .A3(_02511_),
    .B1(_02223_),
    .X(_02532_));
 sky130_fd_sc_hd__nor2_1 _07826_ (.A(_02531_),
    .B(_02532_),
    .Y(_02533_));
 sky130_fd_sc_hd__a21o_1 _07827_ (.A1(\genblk2[0].wave_shpr.div.fin_quo[4] ),
    .A2(_02309_),
    .B1(_02509_),
    .X(_02534_));
 sky130_fd_sc_hd__o21ai_1 _07828_ (.A1(_02533_),
    .A2(_02534_),
    .B1(_02518_),
    .Y(_02535_));
 sky130_fd_sc_hd__nor2_1 _07829_ (.A(_02530_),
    .B(_02535_),
    .Y(_02536_));
 sky130_fd_sc_hd__a21oi_1 _07830_ (.A1(_02461_),
    .A2(_02463_),
    .B1(\genblk2[1].wave_shpr.div.fin_quo[4] ),
    .Y(_02537_));
 sky130_fd_sc_hd__a31o_1 _07831_ (.A1(\genblk2[1].wave_shpr.div.fin_quo[4] ),
    .A2(_02461_),
    .A3(_02463_),
    .B1(_02224_),
    .X(_02538_));
 sky130_fd_sc_hd__clkbuf_4 _07832_ (.A(_02309_),
    .X(_02539_));
 sky130_fd_sc_hd__a21oi_1 _07833_ (.A1(\genblk2[1].wave_shpr.div.fin_quo[5] ),
    .A2(_02539_),
    .B1(_02469_),
    .Y(_02540_));
 sky130_fd_sc_hd__o21a_1 _07834_ (.A1(_02537_),
    .A2(_02538_),
    .B1(_02540_),
    .X(_02541_));
 sky130_fd_sc_hd__a21oi_1 _07835_ (.A1(_02510_),
    .A2(_02512_),
    .B1(\genblk2[0].wave_shpr.div.fin_quo[4] ),
    .Y(_02542_));
 sky130_fd_sc_hd__a31o_1 _07836_ (.A1(\genblk2[0].wave_shpr.div.fin_quo[4] ),
    .A2(_02510_),
    .A3(_02512_),
    .B1(_02261_),
    .X(_02543_));
 sky130_fd_sc_hd__nor2_1 _07837_ (.A(_02542_),
    .B(_02543_),
    .Y(_02544_));
 sky130_fd_sc_hd__a211o_1 _07838_ (.A1(\genblk2[0].wave_shpr.div.fin_quo[5] ),
    .A2(_02539_),
    .B1(_02509_),
    .C1(_02544_),
    .X(_02545_));
 sky130_fd_sc_hd__and4b_1 _07839_ (.A_N(_02541_),
    .B(_02545_),
    .C(_02529_),
    .D(_02518_),
    .X(_02546_));
 sky130_fd_sc_hd__nor2_1 _07840_ (.A(_02536_),
    .B(_02546_),
    .Y(_02547_));
 sky130_fd_sc_hd__xnor2_1 _07841_ (.A(_02530_),
    .B(_02535_),
    .Y(_02548_));
 sky130_fd_sc_hd__o21a_1 _07842_ (.A1(\genblk2[0].wave_shpr.div.fin_quo[0] ),
    .A2(\genblk2[0].wave_shpr.div.fin_quo[1] ),
    .B1(_02510_),
    .X(_02549_));
 sky130_fd_sc_hd__o21ai_1 _07843_ (.A1(\genblk2[0].wave_shpr.div.fin_quo[2] ),
    .A2(_02549_),
    .B1(_02527_),
    .Y(_02550_));
 sky130_fd_sc_hd__a21oi_1 _07844_ (.A1(\genblk2[0].wave_shpr.div.fin_quo[2] ),
    .A2(_02549_),
    .B1(_02550_),
    .Y(_02551_));
 sky130_fd_sc_hd__buf_2 _07845_ (.A(net18),
    .X(_02552_));
 sky130_fd_sc_hd__clkbuf_2 _07846_ (.A(_02552_),
    .X(_02553_));
 sky130_fd_sc_hd__and3_1 _07847_ (.A(_02217_),
    .B(_02553_),
    .C(\genblk2[0].wave_shpr.div.fin_quo[3] ),
    .X(_02554_));
 sky130_fd_sc_hd__or3_1 _07848_ (.A(_02509_),
    .B(_02551_),
    .C(_02554_),
    .X(_02555_));
 sky130_fd_sc_hd__a21oi_1 _07849_ (.A1(_02461_),
    .A2(_02462_),
    .B1(\genblk2[1].wave_shpr.div.fin_quo[2] ),
    .Y(_02556_));
 sky130_fd_sc_hd__a31o_1 _07850_ (.A1(\genblk2[1].wave_shpr.div.fin_quo[2] ),
    .A2(_02461_),
    .A3(_02462_),
    .B1(_02316_),
    .X(_02557_));
 sky130_fd_sc_hd__or2_1 _07851_ (.A(_02556_),
    .B(_02557_),
    .X(_02558_));
 sky130_fd_sc_hd__a21oi_1 _07852_ (.A1(\genblk2[1].wave_shpr.div.fin_quo[3] ),
    .A2(_02309_),
    .B1(_02469_),
    .Y(_02559_));
 sky130_fd_sc_hd__a21oi_1 _07853_ (.A1(_02558_),
    .A2(_02559_),
    .B1(_02424_),
    .Y(_02560_));
 sky130_fd_sc_hd__a21oi_1 _07854_ (.A1(_02518_),
    .A2(_02555_),
    .B1(_02560_),
    .Y(_02561_));
 sky130_fd_sc_hd__o311a_1 _07855_ (.A1(_02509_),
    .A2(_02551_),
    .A3(_02554_),
    .B1(_02560_),
    .C1(_02518_),
    .X(_02562_));
 sky130_fd_sc_hd__a21o_1 _07856_ (.A1(\genblk2[0].wave_shpr.div.fin_quo[0] ),
    .A2(net31),
    .B1(\genblk2[0].wave_shpr.div.fin_quo[1] ),
    .X(_02563_));
 sky130_fd_sc_hd__a31oi_1 _07857_ (.A1(\genblk2[0].wave_shpr.div.fin_quo[0] ),
    .A2(\genblk2[0].wave_shpr.div.fin_quo[1] ),
    .A3(_02510_),
    .B1(_02316_),
    .Y(_02564_));
 sky130_fd_sc_hd__and3_1 _07858_ (.A(_02216_),
    .B(_02552_),
    .C(\genblk2[0].wave_shpr.div.fin_quo[2] ),
    .X(_02565_));
 sky130_fd_sc_hd__a211o_1 _07859_ (.A1(_02563_),
    .A2(_02564_),
    .B1(_02565_),
    .C1(_02509_),
    .X(_02566_));
 sky130_fd_sc_hd__nand4_1 _07860_ (.A(\genblk2[1].wave_shpr.div.fin_quo[0] ),
    .B(\genblk2[1].wave_shpr.div.fin_quo[1] ),
    .C(_02458_),
    .D(_02459_),
    .Y(_02567_));
 sky130_fd_sc_hd__a31o_1 _07861_ (.A1(\genblk2[1].wave_shpr.div.fin_quo[0] ),
    .A2(_02458_),
    .A3(_02459_),
    .B1(\genblk2[1].wave_shpr.div.fin_quo[1] ),
    .X(_02568_));
 sky130_fd_sc_hd__a32o_1 _07862_ (.A1(_02525_),
    .A2(_02567_),
    .A3(_02568_),
    .B1(_02361_),
    .B2(\genblk2[1].wave_shpr.div.fin_quo[2] ),
    .X(_02569_));
 sky130_fd_sc_hd__o21a_1 _07863_ (.A1(_02469_),
    .A2(_02569_),
    .B1(_02529_),
    .X(_02570_));
 sky130_fd_sc_hd__a21o_1 _07864_ (.A1(_02517_),
    .A2(_02566_),
    .B1(_02570_),
    .X(_02571_));
 sky130_fd_sc_hd__and3_1 _07865_ (.A(_02216_),
    .B(_02552_),
    .C(\genblk2[0].wave_shpr.div.fin_quo[0] ),
    .X(_02572_));
 sky130_fd_sc_hd__and3_1 _07866_ (.A(net17),
    .B(_02552_),
    .C(\genblk2[1].wave_shpr.div.fin_quo[0] ),
    .X(_02573_));
 sky130_fd_sc_hd__o21a_1 _07867_ (.A1(_02469_),
    .A2(_02573_),
    .B1(_02529_),
    .X(_02574_));
 sky130_fd_sc_hd__o211a_1 _07868_ (.A1(_02509_),
    .A2(_02572_),
    .B1(_02574_),
    .C1(_02517_),
    .X(_02575_));
 sky130_fd_sc_hd__a22o_1 _07869_ (.A1(\genblk2[0].wave_shpr.div.fin_quo[0] ),
    .A2(_02524_),
    .B1(_02307_),
    .B2(\genblk2[0].wave_shpr.div.fin_quo[1] ),
    .X(_02576_));
 sky130_fd_sc_hd__o21bai_1 _07870_ (.A1(_02221_),
    .A2(_02510_),
    .B1_N(_02576_),
    .Y(_02577_));
 sky130_fd_sc_hd__a22o_1 _07871_ (.A1(\genblk2[1].wave_shpr.div.fin_quo[0] ),
    .A2(_02524_),
    .B1(_02307_),
    .B2(\genblk2[1].wave_shpr.div.fin_quo[1] ),
    .X(_02578_));
 sky130_fd_sc_hd__o21a_1 _07872_ (.A1(_02469_),
    .A2(_02578_),
    .B1(_02529_),
    .X(_02579_));
 sky130_fd_sc_hd__a21o_1 _07873_ (.A1(_02517_),
    .A2(_02577_),
    .B1(_02579_),
    .X(_02580_));
 sky130_fd_sc_hd__and3_1 _07874_ (.A(_02517_),
    .B(_02579_),
    .C(_02577_),
    .X(_02581_));
 sky130_fd_sc_hd__a21o_1 _07875_ (.A1(_02575_),
    .A2(_02580_),
    .B1(_02581_),
    .X(_02582_));
 sky130_fd_sc_hd__and3_1 _07876_ (.A(_02517_),
    .B(_02570_),
    .C(_02566_),
    .X(_02583_));
 sky130_fd_sc_hd__a21o_1 _07877_ (.A1(_02571_),
    .A2(_02582_),
    .B1(_02583_),
    .X(_02584_));
 sky130_fd_sc_hd__nor2_1 _07878_ (.A(_02562_),
    .B(_02584_),
    .Y(_02585_));
 sky130_fd_sc_hd__or3_2 _07879_ (.A(_02548_),
    .B(_02561_),
    .C(_02585_),
    .X(_02586_));
 sky130_fd_sc_hd__o21a_1 _07880_ (.A1(_02424_),
    .A2(_02471_),
    .B1(_02519_),
    .X(_02587_));
 sky130_fd_sc_hd__o2bb2a_1 _07881_ (.A1_N(_02545_),
    .A2_N(_02518_),
    .B1(_02424_),
    .B2(_02541_),
    .X(_02588_));
 sky130_fd_sc_hd__a2111oi_1 _07882_ (.A1(_02547_),
    .A2(_02586_),
    .B1(_02520_),
    .C1(_02587_),
    .D1(_02588_),
    .Y(_02589_));
 sky130_fd_sc_hd__or3b_1 _07883_ (.A(_02464_),
    .B(\genblk2[1].wave_shpr.div.fin_quo[5] ),
    .C_N(_02461_),
    .X(_02590_));
 sky130_fd_sc_hd__xnor2_1 _07884_ (.A(\genblk2[1].wave_shpr.div.fin_quo[6] ),
    .B(_02590_),
    .Y(_02591_));
 sky130_fd_sc_hd__clkbuf_4 _07885_ (.A(_02526_),
    .X(_02592_));
 sky130_fd_sc_hd__a22o_1 _07886_ (.A1(\genblk2[1].wave_shpr.div.fin_quo[7] ),
    .A2(_02539_),
    .B1(_02591_),
    .B2(_02592_),
    .X(_02593_));
 sky130_fd_sc_hd__or2_1 _07887_ (.A(_02469_),
    .B(_02593_),
    .X(_02594_));
 sky130_fd_sc_hd__or3b_1 _07888_ (.A(_02513_),
    .B(\genblk2[0].wave_shpr.div.fin_quo[5] ),
    .C_N(_02510_),
    .X(_02595_));
 sky130_fd_sc_hd__xnor2_1 _07889_ (.A(\genblk2[0].wave_shpr.div.fin_quo[6] ),
    .B(_02595_),
    .Y(_02596_));
 sky130_fd_sc_hd__a22o_1 _07890_ (.A1(\genblk2[0].wave_shpr.div.fin_quo[7] ),
    .A2(_02539_),
    .B1(_02596_),
    .B2(_02592_),
    .X(_02597_));
 sky130_fd_sc_hd__or2_1 _07891_ (.A(_02509_),
    .B(_02597_),
    .X(_02598_));
 sky130_fd_sc_hd__and4_1 _07892_ (.A(_02529_),
    .B(_02594_),
    .C(_02518_),
    .D(_02598_),
    .X(_02599_));
 sky130_fd_sc_hd__a22o_1 _07893_ (.A1(_02529_),
    .A2(_02594_),
    .B1(_02518_),
    .B2(_02598_),
    .X(_02600_));
 sky130_fd_sc_hd__o31a_1 _07894_ (.A1(_02520_),
    .A2(net24),
    .A3(_02599_),
    .B1(_02600_),
    .X(_02601_));
 sky130_fd_sc_hd__nand2_1 _07895_ (.A(_02423_),
    .B(_02601_),
    .Y(_02602_));
 sky130_fd_sc_hd__and3_1 _07896_ (.A(net14),
    .B(net136),
    .C(_02365_),
    .X(_02603_));
 sky130_fd_sc_hd__buf_2 _07897_ (.A(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__a2bb2o_1 _07898_ (.A1_N(\genblk1[8].osc.clkdiv_C.cnt[14] ),
    .A2_N(_01309_),
    .B1(_01576_),
    .B2(\genblk1[8].osc.clkdiv_C.cnt[15] ),
    .X(_02605_));
 sky130_fd_sc_hd__a2bb2o_1 _07899_ (.A1_N(_01181_),
    .A2_N(_01852_),
    .B1(_01245_),
    .B2(\genblk1[8].osc.clkdiv_C.cnt[13] ),
    .X(_02606_));
 sky130_fd_sc_hd__a211o_1 _07900_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[14] ),
    .A2(_01172_),
    .B1(_02605_),
    .C1(_02606_),
    .X(_02607_));
 sky130_fd_sc_hd__o22ai_1 _07901_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[13] ),
    .A2(_01246_),
    .B1(_01328_),
    .B2(\genblk1[8].osc.clkdiv_C.cnt[12] ),
    .Y(_02608_));
 sky130_fd_sc_hd__a211o_1 _07902_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[12] ),
    .A2(_01328_),
    .B1(_02607_),
    .C1(_02608_),
    .X(_02609_));
 sky130_fd_sc_hd__and3_1 _07903_ (.A(\genblk1[8].osc.clkdiv_C.cnt[11] ),
    .B(_01360_),
    .C(_02011_),
    .X(_02610_));
 sky130_fd_sc_hd__nor2_1 _07904_ (.A(\genblk1[8].osc.clkdiv_C.cnt[11] ),
    .B(_01869_),
    .Y(_02611_));
 sky130_fd_sc_hd__xnor2_1 _07905_ (.A(\genblk1[8].osc.clkdiv_C.cnt[10] ),
    .B(_01870_),
    .Y(_02612_));
 sky130_fd_sc_hd__a2111o_1 _07906_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[9] ),
    .A2(_01859_),
    .B1(_02610_),
    .C1(_02611_),
    .D1(_02612_),
    .X(_02613_));
 sky130_fd_sc_hd__o22a_1 _07907_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[8] ),
    .A2(_01865_),
    .B1(_01859_),
    .B2(\genblk1[8].osc.clkdiv_C.cnt[9] ),
    .X(_02614_));
 sky130_fd_sc_hd__or3_1 _07908_ (.A(\genblk1[8].osc.clkdiv_C.cnt[10] ),
    .B(_01870_),
    .C(_02610_),
    .X(_02615_));
 sky130_fd_sc_hd__o221a_1 _07909_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[11] ),
    .A2(_01869_),
    .B1(_02613_),
    .B2(_02614_),
    .C1(_02615_),
    .X(_02616_));
 sky130_fd_sc_hd__a211oi_1 _07910_ (.A1(_01230_),
    .A2(_01564_),
    .B1(_01889_),
    .C1(_01238_),
    .Y(_02617_));
 sky130_fd_sc_hd__o41a_1 _07911_ (.A1(_01228_),
    .A2(_01308_),
    .A3(_01440_),
    .A4(_01889_),
    .B1(_01879_),
    .X(_02618_));
 sky130_fd_sc_hd__o21ba_1 _07912_ (.A1(_01233_),
    .A2(_02617_),
    .B1_N(_02618_),
    .X(_02619_));
 sky130_fd_sc_hd__a311o_1 _07913_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[0] ),
    .A2(_01309_),
    .A3(_01855_),
    .B1(\genblk1[8].osc.clkdiv_C.cnt[1] ),
    .C1(\genblk1[8].osc.clkdiv_C.cnt[2] ),
    .X(_02620_));
 sky130_fd_sc_hd__o221a_1 _07914_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[3] ),
    .A2(_01866_),
    .B1(_02619_),
    .B2(_01489_),
    .C1(_02620_),
    .X(_02621_));
 sky130_fd_sc_hd__a22o_1 _07915_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[3] ),
    .A2(_01866_),
    .B1(_01487_),
    .B2(\genblk1[8].osc.clkdiv_C.cnt[4] ),
    .X(_02622_));
 sky130_fd_sc_hd__or2_1 _07916_ (.A(\genblk1[8].osc.clkdiv_C.cnt[4] ),
    .B(_01487_),
    .X(_02623_));
 sky130_fd_sc_hd__o221a_1 _07917_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[5] ),
    .A2(_01858_),
    .B1(_02621_),
    .B2(_02622_),
    .C1(_02623_),
    .X(_02624_));
 sky130_fd_sc_hd__xor2_1 _07918_ (.A(_01489_),
    .B(\genblk1[8].osc.clkdiv_C.cnt[6] ),
    .X(_02625_));
 sky130_fd_sc_hd__a221o_1 _07919_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[7] ),
    .A2(_01430_),
    .B1(_01858_),
    .B2(\genblk1[8].osc.clkdiv_C.cnt[5] ),
    .C1(_02625_),
    .X(_02626_));
 sky130_fd_sc_hd__a211o_1 _07920_ (.A1(\genblk1[8].osc.clkdiv_C.cnt[7] ),
    .A2(_01430_),
    .B1(\genblk1[8].osc.clkdiv_C.cnt[6] ),
    .C1(_01441_),
    .X(_02627_));
 sky130_fd_sc_hd__or2_1 _07921_ (.A(\genblk1[8].osc.clkdiv_C.cnt[7] ),
    .B(_01430_),
    .X(_02628_));
 sky130_fd_sc_hd__o211a_1 _07922_ (.A1(_02624_),
    .A2(_02626_),
    .B1(_02627_),
    .C1(_02628_),
    .X(_02629_));
 sky130_fd_sc_hd__and2_1 _07923_ (.A(\genblk1[8].osc.clkdiv_C.cnt[8] ),
    .B(_01865_),
    .X(_02630_));
 sky130_fd_sc_hd__or4b_1 _07924_ (.A(_02609_),
    .B(_02613_),
    .C(_02630_),
    .D_N(_02614_),
    .X(_02631_));
 sky130_fd_sc_hd__o22a_1 _07925_ (.A1(_02609_),
    .A2(_02616_),
    .B1(_02629_),
    .B2(_02631_),
    .X(_02632_));
 sky130_fd_sc_hd__or2b_1 _07926_ (.A(_02607_),
    .B_N(_02608_),
    .X(_02633_));
 sky130_fd_sc_hd__a211o_1 _07927_ (.A1(_01200_),
    .A2(\genblk1[8].osc.clkdiv_C.cnt[14] ),
    .B1(_01362_),
    .C1(\genblk1[8].osc.clkdiv_C.cnt[15] ),
    .X(_02634_));
 sky130_fd_sc_hd__a311oi_2 _07928_ (.A1(_02632_),
    .A2(_02633_),
    .A3(_02634_),
    .B1(\genblk1[8].osc.clkdiv_C.cnt[17] ),
    .C1(\genblk1[8].osc.clkdiv_C.cnt[16] ),
    .Y(_02635_));
 sky130_fd_sc_hd__nor2_2 _07929_ (.A(_02221_),
    .B(net30),
    .Y(_02636_));
 sky130_fd_sc_hd__inv_2 _07930_ (.A(\genblk2[8].wave_shpr.div.fin_quo[5] ),
    .Y(_02637_));
 sky130_fd_sc_hd__buf_2 _07931_ (.A(net30),
    .X(_02638_));
 sky130_fd_sc_hd__or3_1 _07932_ (.A(\genblk2[8].wave_shpr.div.fin_quo[0] ),
    .B(\genblk2[8].wave_shpr.div.fin_quo[1] ),
    .C(\genblk2[8].wave_shpr.div.fin_quo[2] ),
    .X(_02639_));
 sky130_fd_sc_hd__or2_1 _07933_ (.A(\genblk2[8].wave_shpr.div.fin_quo[3] ),
    .B(_02639_),
    .X(_02640_));
 sky130_fd_sc_hd__nor2_1 _07934_ (.A(\genblk2[8].wave_shpr.div.fin_quo[4] ),
    .B(_02640_),
    .Y(_02641_));
 sky130_fd_sc_hd__a41o_1 _07935_ (.A1(_02637_),
    .A2(\genblk2[8].wave_shpr.div.fin_quo[6] ),
    .A3(_02638_),
    .A4(_02641_),
    .B1(_02223_),
    .X(_02642_));
 sky130_fd_sc_hd__a31o_1 _07936_ (.A1(_02637_),
    .A2(_02638_),
    .A3(_02641_),
    .B1(\genblk2[8].wave_shpr.div.fin_quo[6] ),
    .X(_02643_));
 sky130_fd_sc_hd__and2b_1 _07937_ (.A_N(_02642_),
    .B(_02643_),
    .X(_02644_));
 sky130_fd_sc_hd__a211o_1 _07938_ (.A1(\genblk2[8].wave_shpr.div.fin_quo[7] ),
    .A2(_02539_),
    .B1(_02636_),
    .C1(_02644_),
    .X(_02645_));
 sky130_fd_sc_hd__nor2_1 _07939_ (.A(_02217_),
    .B(_02553_),
    .Y(_02646_));
 sky130_fd_sc_hd__nand2_1 _07940_ (.A(net13),
    .B(_02364_),
    .Y(_02647_));
 sky130_fd_sc_hd__nor2_2 _07941_ (.A(_02646_),
    .B(_02647_),
    .Y(_02648_));
 sky130_fd_sc_hd__o22a_1 _07942_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[10] ),
    .A2(_01311_),
    .B1(_01925_),
    .B2(\genblk1[7].osc.clkdiv_C.cnt[11] ),
    .X(_02649_));
 sky130_fd_sc_hd__a21o_1 _07943_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[11] ),
    .A2(_01925_),
    .B1(_02649_),
    .X(_02650_));
 sky130_fd_sc_hd__o22a_1 _07944_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[8] ),
    .A2(_01920_),
    .B1(_01514_),
    .B2(\genblk1[7].osc.clkdiv_C.cnt[9] ),
    .X(_02651_));
 sky130_fd_sc_hd__o22a_1 _07945_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[5] ),
    .A2(_01802_),
    .B1(_01805_),
    .B2(\genblk1[7].osc.clkdiv_C.cnt[4] ),
    .X(_02652_));
 sky130_fd_sc_hd__a22o_1 _07946_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[6] ),
    .A2(_01574_),
    .B1(_01802_),
    .B2(\genblk1[7].osc.clkdiv_C.cnt[5] ),
    .X(_02653_));
 sky130_fd_sc_hd__or2_1 _07947_ (.A(\genblk1[7].osc.clkdiv_C.cnt[6] ),
    .B(_01574_),
    .X(_02654_));
 sky130_fd_sc_hd__o221a_1 _07948_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[7] ),
    .A2(_01947_),
    .B1(_02652_),
    .B2(_02653_),
    .C1(_02654_),
    .X(_02655_));
 sky130_fd_sc_hd__nand2_2 _07949_ (.A(_01172_),
    .B(_02011_),
    .Y(_02656_));
 sky130_fd_sc_hd__a21o_1 _07950_ (.A1(_01556_),
    .A2(_01564_),
    .B1(\genblk1[7].osc.clkdiv_C.cnt[1] ),
    .X(_02657_));
 sky130_fd_sc_hd__a32o_1 _07951_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[1] ),
    .A2(_01556_),
    .A3(_01564_),
    .B1(_01732_),
    .B2(\genblk1[7].osc.clkdiv_C.cnt[2] ),
    .X(_02658_));
 sky130_fd_sc_hd__a31o_1 _07952_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[0] ),
    .A2(_01801_),
    .A3(_02657_),
    .B1(_02658_),
    .X(_02659_));
 sky130_fd_sc_hd__o22a_1 _07953_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[2] ),
    .A2(_01732_),
    .B1(_02656_),
    .B2(\genblk1[7].osc.clkdiv_C.cnt[3] ),
    .X(_02660_));
 sky130_fd_sc_hd__and2_1 _07954_ (.A(\genblk1[7].osc.clkdiv_C.cnt[4] ),
    .B(_01805_),
    .X(_02661_));
 sky130_fd_sc_hd__or3b_1 _07955_ (.A(_02661_),
    .B(_02653_),
    .C_N(_02652_),
    .X(_02662_));
 sky130_fd_sc_hd__a221o_1 _07956_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[3] ),
    .A2(_02656_),
    .B1(_02659_),
    .B2(_02660_),
    .C1(_02662_),
    .X(_02663_));
 sky130_fd_sc_hd__a22o_1 _07957_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[8] ),
    .A2(_01920_),
    .B1(_01947_),
    .B2(\genblk1[7].osc.clkdiv_C.cnt[7] ),
    .X(_02664_));
 sky130_fd_sc_hd__a21o_1 _07958_ (.A1(_02655_),
    .A2(_02663_),
    .B1(_02664_),
    .X(_02665_));
 sky130_fd_sc_hd__a22o_1 _07959_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[10] ),
    .A2(_01311_),
    .B1(_01925_),
    .B2(\genblk1[7].osc.clkdiv_C.cnt[11] ),
    .X(_02666_));
 sky130_fd_sc_hd__a221o_1 _07960_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[9] ),
    .A2(_01514_),
    .B1(_02651_),
    .B2(_02665_),
    .C1(_02666_),
    .X(_02667_));
 sky130_fd_sc_hd__or2_1 _07961_ (.A(\genblk1[7].osc.clkdiv_C.cnt[14] ),
    .B(_01360_),
    .X(_02668_));
 sky130_fd_sc_hd__nand2_1 _07962_ (.A(\genblk1[7].osc.clkdiv_C.cnt[14] ),
    .B(_01361_),
    .Y(_02669_));
 sky130_fd_sc_hd__o311a_1 _07963_ (.A1(_01200_),
    .A2(\genblk1[7].osc.clkdiv_C.cnt[15] ),
    .A3(_01361_),
    .B1(_02668_),
    .C1(_02669_),
    .X(_02670_));
 sky130_fd_sc_hd__inv_2 _07964_ (.A(_02670_),
    .Y(_02671_));
 sky130_fd_sc_hd__a221o_1 _07965_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[15] ),
    .A2(_01577_),
    .B1(_01675_),
    .B2(\genblk1[7].osc.clkdiv_C.cnt[13] ),
    .C1(_02671_),
    .X(_02672_));
 sky130_fd_sc_hd__o22a_1 _07966_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[12] ),
    .A2(_01214_),
    .B1(_01675_),
    .B2(\genblk1[7].osc.clkdiv_C.cnt[13] ),
    .X(_02673_));
 sky130_fd_sc_hd__a21bo_1 _07967_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[12] ),
    .A2(_01214_),
    .B1_N(_02673_),
    .X(_02674_));
 sky130_fd_sc_hd__or2_1 _07968_ (.A(_02672_),
    .B(_02674_),
    .X(_02675_));
 sky130_fd_sc_hd__a21oi_2 _07969_ (.A1(_02650_),
    .A2(_02667_),
    .B1(_02675_),
    .Y(_02676_));
 sky130_fd_sc_hd__a21o_1 _07970_ (.A1(\genblk1[7].osc.clkdiv_C.cnt[15] ),
    .A2(_01577_),
    .B1(_02668_),
    .X(_02677_));
 sky130_fd_sc_hd__o31a_1 _07971_ (.A1(_01201_),
    .A2(\genblk1[7].osc.clkdiv_C.cnt[15] ),
    .A3(_01362_),
    .B1(_02677_),
    .X(_02678_));
 sky130_fd_sc_hd__o21ai_2 _07972_ (.A1(_02672_),
    .A2(_02673_),
    .B1(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__nor2_1 _07973_ (.A(\genblk1[7].osc.clkdiv_C.cnt[16] ),
    .B(\genblk1[7].osc.clkdiv_C.cnt[17] ),
    .Y(_02680_));
 sky130_fd_sc_hd__o21ai_2 _07974_ (.A1(_02676_),
    .A2(_02679_),
    .B1(_02680_),
    .Y(_02681_));
 sky130_fd_sc_hd__buf_2 _07975_ (.A(_02681_),
    .X(_02682_));
 sky130_fd_sc_hd__inv_2 _07976_ (.A(\genblk2[7].wave_shpr.div.fin_quo[5] ),
    .Y(_02683_));
 sky130_fd_sc_hd__inv_2 _07977_ (.A(\genblk2[7].wave_shpr.div.fin_quo[3] ),
    .Y(_02684_));
 sky130_fd_sc_hd__inv_2 _07978_ (.A(\genblk2[7].wave_shpr.div.fin_quo[2] ),
    .Y(_02685_));
 sky130_fd_sc_hd__nor2_1 _07979_ (.A(\genblk2[7].wave_shpr.div.fin_quo[0] ),
    .B(\genblk2[7].wave_shpr.div.fin_quo[1] ),
    .Y(_02686_));
 sky130_fd_sc_hd__and2_1 _07980_ (.A(_02685_),
    .B(_02686_),
    .X(_02687_));
 sky130_fd_sc_hd__nand2_1 _07981_ (.A(_02684_),
    .B(_02687_),
    .Y(_02688_));
 sky130_fd_sc_hd__nor2_1 _07982_ (.A(\genblk2[7].wave_shpr.div.fin_quo[4] ),
    .B(_02688_),
    .Y(_02689_));
 sky130_fd_sc_hd__nand2_1 _07983_ (.A(_02683_),
    .B(_02689_),
    .Y(_02690_));
 sky130_fd_sc_hd__inv_2 _07984_ (.A(\genblk2[7].wave_shpr.div.fin_quo[6] ),
    .Y(_02691_));
 sky130_fd_sc_hd__o21ai_1 _07985_ (.A1(_02682_),
    .A2(_02690_),
    .B1(_02691_),
    .Y(_02692_));
 sky130_fd_sc_hd__o31a_1 _07986_ (.A1(_02691_),
    .A2(_02682_),
    .A3(_02690_),
    .B1(_02527_),
    .X(_02693_));
 sky130_fd_sc_hd__and2_1 _07987_ (.A(_02225_),
    .B(_02681_),
    .X(_02694_));
 sky130_fd_sc_hd__and3_1 _07988_ (.A(_02217_),
    .B(_02553_),
    .C(\genblk2[7].wave_shpr.div.fin_quo[7] ),
    .X(_02695_));
 sky130_fd_sc_hd__a211o_1 _07989_ (.A1(_02692_),
    .A2(_02693_),
    .B1(_02694_),
    .C1(_02695_),
    .X(_02696_));
 sky130_fd_sc_hd__nand4_2 _07990_ (.A(_02604_),
    .B(_02645_),
    .C(_02648_),
    .D(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hd__a22o_1 _07991_ (.A1(_02604_),
    .A2(_02645_),
    .B1(_02648_),
    .B2(_02696_),
    .X(_02698_));
 sky130_fd_sc_hd__inv_2 _07992_ (.A(\genblk2[6].wave_shpr.div.fin_quo[5] ),
    .Y(_02699_));
 sky130_fd_sc_hd__o22a_1 _07993_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[10] ),
    .A2(_01484_),
    .B1(_01519_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[11] ),
    .X(_02700_));
 sky130_fd_sc_hd__o22a_1 _07994_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[8] ),
    .A2(_01732_),
    .B1(_01742_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[9] ),
    .X(_02701_));
 sky130_fd_sc_hd__a22oi_1 _07995_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[10] ),
    .A2(_01484_),
    .B1(_01742_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[9] ),
    .Y(_02702_));
 sky130_fd_sc_hd__or2b_1 _07996_ (.A(_02701_),
    .B_N(_02702_),
    .X(_02703_));
 sky130_fd_sc_hd__or2_1 _07997_ (.A(\genblk1[6].osc.clkdiv_C.cnt[14] ),
    .B(_01360_),
    .X(_02704_));
 sky130_fd_sc_hd__nand2_1 _07998_ (.A(\genblk1[6].osc.clkdiv_C.cnt[14] ),
    .B(_01361_),
    .Y(_02705_));
 sky130_fd_sc_hd__o311a_1 _07999_ (.A1(_01200_),
    .A2(\genblk1[6].osc.clkdiv_C.cnt[15] ),
    .A3(_01361_),
    .B1(_02704_),
    .C1(_02705_),
    .X(_02706_));
 sky130_fd_sc_hd__inv_2 _08000_ (.A(_02706_),
    .Y(_02707_));
 sky130_fd_sc_hd__a221o_1 _08001_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[15] ),
    .A2(_01577_),
    .B1(_01675_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[13] ),
    .C1(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__o22a_1 _08002_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[13] ),
    .A2(_01675_),
    .B1(_01666_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[12] ),
    .X(_02709_));
 sky130_fd_sc_hd__a21bo_1 _08003_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[12] ),
    .A2(_01666_),
    .B1_N(_02709_),
    .X(_02710_));
 sky130_fd_sc_hd__a211oi_1 _08004_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[11] ),
    .A2(_01519_),
    .B1(_02708_),
    .C1(_02710_),
    .Y(_02711_));
 sky130_fd_sc_hd__a21boi_1 _08005_ (.A1(_02700_),
    .A2(_02703_),
    .B1_N(_02711_),
    .Y(_02712_));
 sky130_fd_sc_hd__o211a_1 _08006_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[1] ),
    .A2(_01735_),
    .B1(_01738_),
    .C1(\genblk1[6].osc.clkdiv_C.cnt[0] ),
    .X(_02713_));
 sky130_fd_sc_hd__a2bb2o_1 _08007_ (.A1_N(_01729_),
    .A2_N(_01758_),
    .B1(_01735_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[1] ),
    .X(_02714_));
 sky130_fd_sc_hd__a2bb2o_1 _08008_ (.A1_N(\genblk1[6].osc.clkdiv_C.cnt[3] ),
    .A2_N(_01730_),
    .B1(_01758_),
    .B2(_01729_),
    .X(_02715_));
 sky130_fd_sc_hd__o21ba_1 _08009_ (.A1(_02713_),
    .A2(_02714_),
    .B1_N(_02715_),
    .X(_02716_));
 sky130_fd_sc_hd__o21a_1 _08010_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[5] ),
    .A2(_01365_),
    .B1(\genblk1[6].osc.clkdiv_C.cnt[3] ),
    .X(_02717_));
 sky130_fd_sc_hd__a221o_1 _08011_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[5] ),
    .A2(_01367_),
    .B1(_01747_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[4] ),
    .C1(_02717_),
    .X(_02718_));
 sky130_fd_sc_hd__or2_1 _08012_ (.A(\genblk1[6].osc.clkdiv_C.cnt[4] ),
    .B(_01747_),
    .X(_02719_));
 sky130_fd_sc_hd__o221a_1 _08013_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[5] ),
    .A2(_01367_),
    .B1(_02716_),
    .B2(_02718_),
    .C1(_02719_),
    .X(_02720_));
 sky130_fd_sc_hd__nand2_1 _08014_ (.A(\genblk1[6].osc.clkdiv_C.cnt[5] ),
    .B(_01367_),
    .Y(_02721_));
 sky130_fd_sc_hd__a2bb2o_1 _08015_ (.A1_N(_02721_),
    .A2_N(_02719_),
    .B1(\genblk1[6].osc.clkdiv_C.cnt[6] ),
    .B2(_01750_),
    .X(_02722_));
 sky130_fd_sc_hd__o22a_1 _08016_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[6] ),
    .A2(_01750_),
    .B1(_01739_),
    .B2(\genblk1[6].osc.clkdiv_C.cnt[7] ),
    .X(_02723_));
 sky130_fd_sc_hd__o21ai_1 _08017_ (.A1(_02720_),
    .A2(_02722_),
    .B1(_02723_),
    .Y(_02724_));
 sky130_fd_sc_hd__inv_2 _08018_ (.A(_01739_),
    .Y(_02725_));
 sky130_fd_sc_hd__o2bb2a_1 _08019_ (.A1_N(\genblk1[6].osc.clkdiv_C.cnt[8] ),
    .A2_N(_01732_),
    .B1(_02725_),
    .B2(_01753_),
    .X(_02726_));
 sky130_fd_sc_hd__and4_1 _08020_ (.A(_02700_),
    .B(_02702_),
    .C(_02701_),
    .D(_02726_),
    .X(_02727_));
 sky130_fd_sc_hd__a21o_1 _08021_ (.A1(\genblk1[6].osc.clkdiv_C.cnt[15] ),
    .A2(_01577_),
    .B1(_02704_),
    .X(_02728_));
 sky130_fd_sc_hd__o21ai_1 _08022_ (.A1(_02709_),
    .A2(_02708_),
    .B1(_02728_),
    .Y(_02729_));
 sky130_fd_sc_hd__a21o_1 _08023_ (.A1(_01229_),
    .A2(_01749_),
    .B1(_02729_),
    .X(_02730_));
 sky130_fd_sc_hd__a31o_1 _08024_ (.A1(_02711_),
    .A2(_02724_),
    .A3(_02727_),
    .B1(_02730_),
    .X(_02731_));
 sky130_fd_sc_hd__nor2_1 _08025_ (.A(\genblk1[6].osc.clkdiv_C.cnt[16] ),
    .B(\genblk1[6].osc.clkdiv_C.cnt[17] ),
    .Y(_02732_));
 sky130_fd_sc_hd__o21a_4 _08026_ (.A1(_02712_),
    .A2(_02731_),
    .B1(_02732_),
    .X(_02733_));
 sky130_fd_sc_hd__buf_2 _08027_ (.A(_02733_),
    .X(_02734_));
 sky130_fd_sc_hd__or2_1 _08028_ (.A(\genblk2[6].wave_shpr.div.fin_quo[0] ),
    .B(\genblk2[6].wave_shpr.div.fin_quo[1] ),
    .X(_02735_));
 sky130_fd_sc_hd__or2_1 _08029_ (.A(\genblk2[6].wave_shpr.div.fin_quo[2] ),
    .B(_02735_),
    .X(_02736_));
 sky130_fd_sc_hd__or2_1 _08030_ (.A(\genblk2[6].wave_shpr.div.fin_quo[3] ),
    .B(_02736_),
    .X(_02737_));
 sky130_fd_sc_hd__nor2_1 _08031_ (.A(\genblk2[6].wave_shpr.div.fin_quo[4] ),
    .B(_02737_),
    .Y(_02738_));
 sky130_fd_sc_hd__a41o_1 _08032_ (.A1(_02699_),
    .A2(\genblk2[6].wave_shpr.div.fin_quo[6] ),
    .A3(_02734_),
    .A4(_02738_),
    .B1(_02261_),
    .X(_02739_));
 sky130_fd_sc_hd__a31o_1 _08033_ (.A1(_02699_),
    .A2(_02734_),
    .A3(_02738_),
    .B1(\genblk2[6].wave_shpr.div.fin_quo[6] ),
    .X(_02740_));
 sky130_fd_sc_hd__and2b_1 _08034_ (.A_N(_02739_),
    .B(_02740_),
    .X(_02741_));
 sky130_fd_sc_hd__nor2_2 _08035_ (.A(_02221_),
    .B(_02733_),
    .Y(_02742_));
 sky130_fd_sc_hd__a21o_1 _08036_ (.A1(\genblk2[6].wave_shpr.div.fin_quo[7] ),
    .A2(_02539_),
    .B1(_02742_),
    .X(_02743_));
 sky130_fd_sc_hd__buf_2 _08037_ (.A(_02364_),
    .X(_02744_));
 sky130_fd_sc_hd__and3_2 _08038_ (.A(net12),
    .B(_02744_),
    .C(_02365_),
    .X(_02745_));
 sky130_fd_sc_hd__o21a_1 _08039_ (.A1(_02741_),
    .A2(_02743_),
    .B1(_02745_),
    .X(_02746_));
 sky130_fd_sc_hd__nand3_1 _08040_ (.A(_02697_),
    .B(_02698_),
    .C(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__and2_1 _08041_ (.A(\genblk1[5].osc.clkdiv_C.cnt[15] ),
    .B(_01576_),
    .X(_02748_));
 sky130_fd_sc_hd__or2_1 _08042_ (.A(\genblk1[5].osc.clkdiv_C.cnt[14] ),
    .B(_01359_),
    .X(_02749_));
 sky130_fd_sc_hd__nand2_1 _08043_ (.A(\genblk1[5].osc.clkdiv_C.cnt[14] ),
    .B(_01360_),
    .Y(_02750_));
 sky130_fd_sc_hd__o211ai_1 _08044_ (.A1(_01181_),
    .A2(_01680_),
    .B1(_02749_),
    .C1(_02750_),
    .Y(_02751_));
 sky130_fd_sc_hd__a211o_1 _08045_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[13] ),
    .A2(_01675_),
    .B1(_02748_),
    .C1(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__o22a_1 _08046_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[13] ),
    .A2(_01674_),
    .B1(_01666_),
    .B2(\genblk1[5].osc.clkdiv_C.cnt[12] ),
    .X(_02753_));
 sky130_fd_sc_hd__a21bo_1 _08047_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[12] ),
    .A2(_01666_),
    .B1_N(_02753_),
    .X(_02754_));
 sky130_fd_sc_hd__or2_1 _08048_ (.A(_02752_),
    .B(_02754_),
    .X(_02755_));
 sky130_fd_sc_hd__nor2_1 _08049_ (.A(\genblk1[5].osc.clkdiv_C.cnt[11] ),
    .B(_01355_),
    .Y(_02756_));
 sky130_fd_sc_hd__and2_1 _08050_ (.A(\genblk1[5].osc.clkdiv_C.cnt[11] ),
    .B(_01355_),
    .X(_02757_));
 sky130_fd_sc_hd__nor2_1 _08051_ (.A(\genblk1[5].osc.clkdiv_C.cnt[10] ),
    .B(_01667_),
    .Y(_02758_));
 sky130_fd_sc_hd__a32o_1 _08052_ (.A1(_01489_),
    .A2(\genblk1[5].osc.clkdiv_C.cnt[9] ),
    .A3(net37),
    .B1(_01667_),
    .B2(\genblk1[5].osc.clkdiv_C.cnt[10] ),
    .X(_02759_));
 sky130_fd_sc_hd__or4_1 _08053_ (.A(_02756_),
    .B(_02757_),
    .C(_02758_),
    .D(_02759_),
    .X(_02760_));
 sky130_fd_sc_hd__or2_1 _08054_ (.A(\genblk1[5].osc.clkdiv_C.cnt[7] ),
    .B(_01223_),
    .X(_02761_));
 sky130_fd_sc_hd__a21o_1 _08055_ (.A1(_01309_),
    .A2(_01180_),
    .B1(\genblk1[5].osc.clkdiv_C.cnt[6] ),
    .X(_02762_));
 sky130_fd_sc_hd__nand2_1 _08056_ (.A(_02761_),
    .B(_02762_),
    .Y(_02763_));
 sky130_fd_sc_hd__and2_1 _08057_ (.A(\genblk1[5].osc.clkdiv_C.cnt[7] ),
    .B(_01223_),
    .X(_02764_));
 sky130_fd_sc_hd__a31o_1 _08058_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[6] ),
    .A2(_01172_),
    .A3(_01180_),
    .B1(_02764_),
    .X(_02765_));
 sky130_fd_sc_hd__o22a_1 _08059_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[5] ),
    .A2(_01238_),
    .B1(net36),
    .B2(\genblk1[5].osc.clkdiv_C.cnt[4] ),
    .X(_02766_));
 sky130_fd_sc_hd__and2_1 _08060_ (.A(\genblk1[5].osc.clkdiv_C.cnt[5] ),
    .B(_01238_),
    .X(_02767_));
 sky130_fd_sc_hd__a21oi_1 _08061_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[4] ),
    .A2(net36),
    .B1(_02767_),
    .Y(_02768_));
 sky130_fd_sc_hd__nand2_1 _08062_ (.A(_02766_),
    .B(_02768_),
    .Y(_02769_));
 sky130_fd_sc_hd__or3_1 _08063_ (.A(\genblk1[5].osc.clkdiv_C.cnt[2] ),
    .B(_01238_),
    .C(net35),
    .X(_02770_));
 sky130_fd_sc_hd__or3_1 _08064_ (.A(\genblk1[5].osc.clkdiv_C.cnt[3] ),
    .B(_01195_),
    .C(_01254_),
    .X(_02771_));
 sky130_fd_sc_hd__nand2_1 _08065_ (.A(_02770_),
    .B(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__o311a_1 _08066_ (.A1(_01179_),
    .A2(_01222_),
    .A3(_01254_),
    .B1(_01171_),
    .C1(\genblk1[5].osc.clkdiv_C.cnt[0] ),
    .X(_02773_));
 sky130_fd_sc_hd__o21a_1 _08067_ (.A1(_01660_),
    .A2(_02773_),
    .B1(\genblk1[5].osc.clkdiv_C.cnt[1] ),
    .X(_02774_));
 sky130_fd_sc_hd__o21a_1 _08068_ (.A1(_01196_),
    .A2(_01254_),
    .B1(\genblk1[5].osc.clkdiv_C.cnt[3] ),
    .X(_02775_));
 sky130_fd_sc_hd__a21o_1 _08069_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[2] ),
    .A2(_01592_),
    .B1(_02775_),
    .X(_02776_));
 sky130_fd_sc_hd__a21o_1 _08070_ (.A1(_02770_),
    .A2(_02771_),
    .B1(_02775_),
    .X(_02777_));
 sky130_fd_sc_hd__o31a_1 _08071_ (.A1(_02772_),
    .A2(_02774_),
    .A3(_02776_),
    .B1(_02777_),
    .X(_02778_));
 sky130_fd_sc_hd__a311o_1 _08072_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[6] ),
    .A2(_01309_),
    .A3(_01180_),
    .B1(_02767_),
    .C1(_02766_),
    .X(_02779_));
 sky130_fd_sc_hd__a31o_1 _08073_ (.A1(_02761_),
    .A2(_02762_),
    .A3(_02779_),
    .B1(_02764_),
    .X(_02780_));
 sky130_fd_sc_hd__o41a_1 _08074_ (.A1(_02763_),
    .A2(_02765_),
    .A3(_02769_),
    .A4(_02778_),
    .B1(_02780_),
    .X(_02781_));
 sky130_fd_sc_hd__o22a_1 _08075_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[8] ),
    .A2(_01678_),
    .B1(_01726_),
    .B2(\genblk1[5].osc.clkdiv_C.cnt[9] ),
    .X(_02782_));
 sky130_fd_sc_hd__a21bo_1 _08076_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[8] ),
    .A2(_01678_),
    .B1_N(_02782_),
    .X(_02783_));
 sky130_fd_sc_hd__or4_1 _08077_ (.A(_02755_),
    .B(_02760_),
    .C(_02781_),
    .D(_02783_),
    .X(_02784_));
 sky130_fd_sc_hd__or3_1 _08078_ (.A(\genblk1[5].osc.clkdiv_C.cnt[10] ),
    .B(_01667_),
    .C(_02757_),
    .X(_02785_));
 sky130_fd_sc_hd__o221a_1 _08079_ (.A1(\genblk1[5].osc.clkdiv_C.cnt[11] ),
    .A2(_01355_),
    .B1(_02760_),
    .B2(_02782_),
    .C1(_02785_),
    .X(_02786_));
 sky130_fd_sc_hd__o22a_1 _08080_ (.A1(_01200_),
    .A2(_01680_),
    .B1(_02748_),
    .B2(_02749_),
    .X(_02787_));
 sky130_fd_sc_hd__o221a_1 _08081_ (.A1(_02752_),
    .A2(_02753_),
    .B1(_02755_),
    .B2(_02786_),
    .C1(_02787_),
    .X(_02788_));
 sky130_fd_sc_hd__a211o_4 _08082_ (.A1(_02784_),
    .A2(_02788_),
    .B1(\genblk1[5].osc.clkdiv_C.cnt[16] ),
    .C1(\genblk1[5].osc.clkdiv_C.cnt[17] ),
    .X(_02789_));
 sky130_fd_sc_hd__and2_1 _08083_ (.A(_02225_),
    .B(_02789_),
    .X(_02790_));
 sky130_fd_sc_hd__buf_2 _08084_ (.A(_02790_),
    .X(_02791_));
 sky130_fd_sc_hd__or4_1 _08085_ (.A(\genblk2[5].wave_shpr.div.fin_quo[0] ),
    .B(\genblk2[5].wave_shpr.div.fin_quo[1] ),
    .C(\genblk2[5].wave_shpr.div.fin_quo[2] ),
    .D(\genblk2[5].wave_shpr.div.fin_quo[3] ),
    .X(_02792_));
 sky130_fd_sc_hd__nor2_1 _08086_ (.A(\genblk2[5].wave_shpr.div.fin_quo[4] ),
    .B(_02792_),
    .Y(_02793_));
 sky130_fd_sc_hd__or3b_1 _08087_ (.A(\genblk2[5].wave_shpr.div.fin_quo[5] ),
    .B(_02789_),
    .C_N(_02793_),
    .X(_02794_));
 sky130_fd_sc_hd__xnor2_1 _08088_ (.A(\genblk2[5].wave_shpr.div.fin_quo[6] ),
    .B(_02794_),
    .Y(_02795_));
 sky130_fd_sc_hd__a22o_1 _08089_ (.A1(\genblk2[5].wave_shpr.div.fin_quo[7] ),
    .A2(_02309_),
    .B1(_02795_),
    .B2(_02527_),
    .X(_02796_));
 sky130_fd_sc_hd__and3_1 _08090_ (.A(net11),
    .B(_02364_),
    .C(_02365_),
    .X(_02797_));
 sky130_fd_sc_hd__buf_2 _08091_ (.A(_02797_),
    .X(_02798_));
 sky130_fd_sc_hd__o21ai_2 _08092_ (.A1(_02791_),
    .A2(_02796_),
    .B1(_02798_),
    .Y(_02799_));
 sky130_fd_sc_hd__nor2_1 _08093_ (.A(\genblk1[4].osc.clkdiv_C.cnt[14] ),
    .B(_01360_),
    .Y(_02800_));
 sky130_fd_sc_hd__a22o_1 _08094_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[14] ),
    .A2(_01359_),
    .B1(_01498_),
    .B2(\genblk1[4].osc.clkdiv_C.cnt[13] ),
    .X(_02801_));
 sky130_fd_sc_hd__nor2_1 _08095_ (.A(_01650_),
    .B(_01196_),
    .Y(_02802_));
 sky130_fd_sc_hd__or3_1 _08096_ (.A(_01174_),
    .B(\genblk1[4].osc.clkdiv_C.cnt[15] ),
    .C(_01359_),
    .X(_02803_));
 sky130_fd_sc_hd__or4b_1 _08097_ (.A(_02800_),
    .B(_02801_),
    .C(_02802_),
    .D_N(_02803_),
    .X(_02804_));
 sky130_fd_sc_hd__nand2_2 _08098_ (.A(_01440_),
    .B(_01576_),
    .Y(_02805_));
 sky130_fd_sc_hd__o22a_1 _08099_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[13] ),
    .A2(_01498_),
    .B1(_02805_),
    .B2(\genblk1[4].osc.clkdiv_C.cnt[12] ),
    .X(_02806_));
 sky130_fd_sc_hd__a21bo_1 _08100_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[12] ),
    .A2(_02805_),
    .B1_N(_02806_),
    .X(_02807_));
 sky130_fd_sc_hd__or2_1 _08101_ (.A(_02804_),
    .B(_02807_),
    .X(_02808_));
 sky130_fd_sc_hd__and2_1 _08102_ (.A(\genblk1[4].osc.clkdiv_C.cnt[11] ),
    .B(_01574_),
    .X(_02809_));
 sky130_fd_sc_hd__or2_1 _08103_ (.A(\genblk1[4].osc.clkdiv_C.cnt[11] ),
    .B(_01574_),
    .X(_02810_));
 sky130_fd_sc_hd__o22a_1 _08104_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[9] ),
    .A2(_01323_),
    .B1(_01592_),
    .B2(\genblk1[4].osc.clkdiv_C.cnt[8] ),
    .X(_02811_));
 sky130_fd_sc_hd__and3_1 _08105_ (.A(_01588_),
    .B(_01192_),
    .C(_01208_),
    .X(_02812_));
 sky130_fd_sc_hd__nor2_1 _08106_ (.A(\genblk1[4].osc.clkdiv_C.cnt[11] ),
    .B(_01574_),
    .Y(_02813_));
 sky130_fd_sc_hd__a21oi_1 _08107_ (.A1(_01192_),
    .A2(_01208_),
    .B1(_01588_),
    .Y(_02814_));
 sky130_fd_sc_hd__or4_1 _08108_ (.A(_02812_),
    .B(_02809_),
    .C(_02813_),
    .D(_02814_),
    .X(_02815_));
 sky130_fd_sc_hd__a211o_1 _08109_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[9] ),
    .A2(_01323_),
    .B1(_02811_),
    .C1(_02815_),
    .X(_02816_));
 sky130_fd_sc_hd__o311a_1 _08110_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[10] ),
    .A2(_01313_),
    .A3(_02809_),
    .B1(_02810_),
    .C1(_02816_),
    .X(_02817_));
 sky130_fd_sc_hd__o31a_1 _08111_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[14] ),
    .A2(_01361_),
    .A3(_02802_),
    .B1(_02803_),
    .X(_02818_));
 sky130_fd_sc_hd__o221a_1 _08112_ (.A1(_02804_),
    .A2(_02806_),
    .B1(_02808_),
    .B2(_02817_),
    .C1(_02818_),
    .X(_02819_));
 sky130_fd_sc_hd__a22oi_1 _08113_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[9] ),
    .A2(_01323_),
    .B1(_01592_),
    .B2(\genblk1[4].osc.clkdiv_C.cnt[8] ),
    .Y(_02820_));
 sky130_fd_sc_hd__nand2_1 _08114_ (.A(_02811_),
    .B(_02820_),
    .Y(_02821_));
 sky130_fd_sc_hd__a21oi_1 _08115_ (.A1(_01172_),
    .A2(_01180_),
    .B1(_01568_),
    .Y(_02822_));
 sky130_fd_sc_hd__o21a_1 _08116_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[1] ),
    .A2(_01866_),
    .B1(\genblk1[4].osc.clkdiv_C.cnt[0] ),
    .X(_02823_));
 sky130_fd_sc_hd__and2_1 _08117_ (.A(\genblk1[4].osc.clkdiv_C.cnt[2] ),
    .B(_01326_),
    .X(_02824_));
 sky130_fd_sc_hd__o22a_1 _08118_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[2] ),
    .A2(_01326_),
    .B1(_01213_),
    .B2(\genblk1[4].osc.clkdiv_C.cnt[3] ),
    .X(_02825_));
 sky130_fd_sc_hd__o31a_1 _08119_ (.A1(_02822_),
    .A2(_02823_),
    .A3(_02824_),
    .B1(_02825_),
    .X(_02826_));
 sky130_fd_sc_hd__o21a_1 _08120_ (.A1(_01224_),
    .A2(_01249_),
    .B1(\genblk1[4].osc.clkdiv_C.cnt[5] ),
    .X(_02827_));
 sky130_fd_sc_hd__a21o_1 _08121_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[3] ),
    .A2(_01439_),
    .B1(_02827_),
    .X(_02828_));
 sky130_fd_sc_hd__o22a_1 _08122_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[7] ),
    .A2(_01340_),
    .B1(_01304_),
    .B2(\genblk1[4].osc.clkdiv_C.cnt[6] ),
    .X(_02829_));
 sky130_fd_sc_hd__o32a_1 _08123_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[5] ),
    .A2(_01224_),
    .A3(_01249_),
    .B1(_01565_),
    .B2(\genblk1[4].osc.clkdiv_C.cnt[4] ),
    .X(_02830_));
 sky130_fd_sc_hd__a22oi_1 _08124_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[7] ),
    .A2(_01340_),
    .B1(_01304_),
    .B2(\genblk1[4].osc.clkdiv_C.cnt[6] ),
    .Y(_02831_));
 sky130_fd_sc_hd__o2111ai_1 _08125_ (.A1(_01570_),
    .A2(_01870_),
    .B1(_02829_),
    .C1(_02830_),
    .D1(_02831_),
    .Y(_02832_));
 sky130_fd_sc_hd__a21o_1 _08126_ (.A1(\genblk1[4].osc.clkdiv_C.cnt[7] ),
    .A2(_01340_),
    .B1(_02829_),
    .X(_02833_));
 sky130_fd_sc_hd__or4bb_1 _08127_ (.A(_02830_),
    .B(_02827_),
    .C_N(_02831_),
    .D_N(_02829_),
    .X(_02834_));
 sky130_fd_sc_hd__o311a_1 _08128_ (.A1(_02826_),
    .A2(_02828_),
    .A3(_02832_),
    .B1(_02833_),
    .C1(_02834_),
    .X(_02835_));
 sky130_fd_sc_hd__or4_2 _08129_ (.A(_02808_),
    .B(_02815_),
    .C(_02821_),
    .D(_02835_),
    .X(_02836_));
 sky130_fd_sc_hd__a211oi_4 _08130_ (.A1(_02819_),
    .A2(_02836_),
    .B1(\genblk1[4].osc.clkdiv_C.cnt[16] ),
    .C1(\genblk1[4].osc.clkdiv_C.cnt[17] ),
    .Y(_02837_));
 sky130_fd_sc_hd__nor2_2 _08131_ (.A(_02221_),
    .B(_02837_),
    .Y(_02838_));
 sky130_fd_sc_hd__or2_1 _08132_ (.A(\genblk2[4].wave_shpr.div.fin_quo[0] ),
    .B(\genblk2[4].wave_shpr.div.fin_quo[1] ),
    .X(_02839_));
 sky130_fd_sc_hd__or2_1 _08133_ (.A(\genblk2[4].wave_shpr.div.fin_quo[2] ),
    .B(_02839_),
    .X(_02840_));
 sky130_fd_sc_hd__or2_1 _08134_ (.A(\genblk2[4].wave_shpr.div.fin_quo[3] ),
    .B(_02840_),
    .X(_02841_));
 sky130_fd_sc_hd__or2_1 _08135_ (.A(\genblk2[4].wave_shpr.div.fin_quo[4] ),
    .B(_02841_),
    .X(_02842_));
 sky130_fd_sc_hd__or3b_1 _08136_ (.A(_02842_),
    .B(\genblk2[4].wave_shpr.div.fin_quo[5] ),
    .C_N(_02837_),
    .X(_02843_));
 sky130_fd_sc_hd__xnor2_1 _08137_ (.A(\genblk2[4].wave_shpr.div.fin_quo[6] ),
    .B(_02843_),
    .Y(_02844_));
 sky130_fd_sc_hd__a22o_1 _08138_ (.A1(\genblk2[4].wave_shpr.div.fin_quo[7] ),
    .A2(_02309_),
    .B1(_02844_),
    .B2(_02527_),
    .X(_02845_));
 sky130_fd_sc_hd__and3_2 _08139_ (.A(net10),
    .B(_02364_),
    .C(_02365_),
    .X(_02846_));
 sky130_fd_sc_hd__o21ai_2 _08140_ (.A1(_02838_),
    .A2(_02845_),
    .B1(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__xor2_2 _08141_ (.A(_02799_),
    .B(_02847_),
    .X(_02848_));
 sky130_fd_sc_hd__inv_2 _08142_ (.A(_02848_),
    .Y(_02849_));
 sky130_fd_sc_hd__inv_2 _08143_ (.A(\genblk2[3].wave_shpr.div.fin_quo[6] ),
    .Y(_02850_));
 sky130_fd_sc_hd__nor2_1 _08144_ (.A(\genblk1[3].osc.clkdiv_C.cnt[15] ),
    .B(_01576_),
    .Y(_02851_));
 sky130_fd_sc_hd__a211oi_1 _08145_ (.A1(_01201_),
    .A2(\genblk1[3].osc.clkdiv_C.cnt[15] ),
    .B1(\genblk1[3].osc.clkdiv_C.cnt[14] ),
    .C1(_01362_),
    .Y(_02852_));
 sky130_fd_sc_hd__nor2_1 _08146_ (.A(_02851_),
    .B(_02852_),
    .Y(_02853_));
 sky130_fd_sc_hd__o211a_1 _08147_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[1] ),
    .A2(_01496_),
    .B1(_01519_),
    .C1(\genblk1[3].osc.clkdiv_C.cnt[0] ),
    .X(_02854_));
 sky130_fd_sc_hd__a22o_1 _08148_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[1] ),
    .A2(_01496_),
    .B1(_01513_),
    .B2(\genblk1[3].osc.clkdiv_C.cnt[2] ),
    .X(_02855_));
 sky130_fd_sc_hd__or2_1 _08149_ (.A(\genblk1[3].osc.clkdiv_C.cnt[2] ),
    .B(_01513_),
    .X(_02856_));
 sky130_fd_sc_hd__o221a_1 _08150_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[3] ),
    .A2(_01234_),
    .B1(_02854_),
    .B2(_02855_),
    .C1(_02856_),
    .X(_02857_));
 sky130_fd_sc_hd__a221o_1 _08151_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[4] ),
    .A2(_01250_),
    .B1(_01514_),
    .B2(\genblk1[3].osc.clkdiv_C.cnt[3] ),
    .C1(_02857_),
    .X(_02858_));
 sky130_fd_sc_hd__o22a_1 _08152_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[5] ),
    .A2(_01500_),
    .B1(_01250_),
    .B2(\genblk1[3].osc.clkdiv_C.cnt[4] ),
    .X(_02859_));
 sky130_fd_sc_hd__a22o_1 _08153_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[5] ),
    .A2(_01500_),
    .B1(_01494_),
    .B2(\genblk1[3].osc.clkdiv_C.cnt[6] ),
    .X(_02860_));
 sky130_fd_sc_hd__a21o_1 _08154_ (.A1(_02858_),
    .A2(_02859_),
    .B1(_02860_),
    .X(_02861_));
 sky130_fd_sc_hd__o22a_1 _08155_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[7] ),
    .A2(_01483_),
    .B1(_01494_),
    .B2(\genblk1[3].osc.clkdiv_C.cnt[6] ),
    .X(_02862_));
 sky130_fd_sc_hd__a2bb2o_1 _08156_ (.A1_N(\genblk1[3].osc.clkdiv_C.cnt[14] ),
    .A2_N(_01361_),
    .B1(_01576_),
    .B2(\genblk1[3].osc.clkdiv_C.cnt[15] ),
    .X(_02863_));
 sky130_fd_sc_hd__a211o_1 _08157_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[14] ),
    .A2(_01361_),
    .B1(_02851_),
    .C1(_02863_),
    .X(_02864_));
 sky130_fd_sc_hd__a221o_1 _08158_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[7] ),
    .A2(_01483_),
    .B1(_01858_),
    .B2(_01486_),
    .C1(_02864_),
    .X(_02865_));
 sky130_fd_sc_hd__nand2_1 _08159_ (.A(_01489_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[12] ),
    .Y(_02866_));
 sky130_fd_sc_hd__or2_1 _08160_ (.A(_01489_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[12] ),
    .X(_02867_));
 sky130_fd_sc_hd__or2_1 _08161_ (.A(\genblk1[3].osc.clkdiv_C.cnt[13] ),
    .B(_01498_),
    .X(_02868_));
 sky130_fd_sc_hd__and3_1 _08162_ (.A(_02866_),
    .B(_02867_),
    .C(_02868_),
    .X(_02869_));
 sky130_fd_sc_hd__a21bo_1 _08163_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[13] ),
    .A2(_01498_),
    .B1_N(_02869_),
    .X(_02870_));
 sky130_fd_sc_hd__and3_1 _08164_ (.A(_01181_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[9] ),
    .C(_01182_),
    .X(_02871_));
 sky130_fd_sc_hd__or2_1 _08165_ (.A(\genblk1[3].osc.clkdiv_C.cnt[10] ),
    .B(_01508_),
    .X(_02872_));
 sky130_fd_sc_hd__or2_1 _08166_ (.A(\genblk1[3].osc.clkdiv_C.cnt[8] ),
    .B(_01423_),
    .X(_02873_));
 sky130_fd_sc_hd__or2_1 _08167_ (.A(\genblk1[3].osc.clkdiv_C.cnt[9] ),
    .B(_01231_),
    .X(_02874_));
 sky130_fd_sc_hd__nand3_1 _08168_ (.A(_02872_),
    .B(_02873_),
    .C(_02874_),
    .Y(_02875_));
 sky130_fd_sc_hd__a2111o_1 _08169_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[8] ),
    .A2(_01423_),
    .B1(_02870_),
    .C1(_02871_),
    .D1(_02875_),
    .X(_02876_));
 sky130_fd_sc_hd__a22o_1 _08170_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[10] ),
    .A2(_01508_),
    .B1(_01507_),
    .B2(\genblk1[3].osc.clkdiv_C.cnt[11] ),
    .X(_02877_));
 sky130_fd_sc_hd__a2111o_1 _08171_ (.A1(_02861_),
    .A2(_02862_),
    .B1(_02865_),
    .C1(_02876_),
    .D1(_02877_),
    .X(_02878_));
 sky130_fd_sc_hd__a21o_1 _08172_ (.A1(\genblk1[3].osc.clkdiv_C.cnt[13] ),
    .A2(_01498_),
    .B1(_02867_),
    .X(_02879_));
 sky130_fd_sc_hd__nand2_1 _08173_ (.A(_01486_),
    .B(_01858_),
    .Y(_02880_));
 sky130_fd_sc_hd__a21o_1 _08174_ (.A1(_02873_),
    .A2(_02874_),
    .B1(_02871_),
    .X(_02881_));
 sky130_fd_sc_hd__a21o_1 _08175_ (.A1(_02872_),
    .A2(_02881_),
    .B1(_02877_),
    .X(_02882_));
 sky130_fd_sc_hd__a21o_1 _08176_ (.A1(_02880_),
    .A2(_02882_),
    .B1(_02870_),
    .X(_02883_));
 sky130_fd_sc_hd__a31o_1 _08177_ (.A1(_02868_),
    .A2(_02879_),
    .A3(_02883_),
    .B1(_02864_),
    .X(_02884_));
 sky130_fd_sc_hd__a311o_4 _08178_ (.A1(_02853_),
    .A2(_02878_),
    .A3(_02884_),
    .B1(\genblk1[3].osc.clkdiv_C.cnt[17] ),
    .C1(\genblk1[3].osc.clkdiv_C.cnt[16] ),
    .X(_02885_));
 sky130_fd_sc_hd__or4_1 _08179_ (.A(\genblk2[3].wave_shpr.div.fin_quo[0] ),
    .B(\genblk2[3].wave_shpr.div.fin_quo[1] ),
    .C(\genblk2[3].wave_shpr.div.fin_quo[2] ),
    .D(\genblk2[3].wave_shpr.div.fin_quo[3] ),
    .X(_02886_));
 sky130_fd_sc_hd__nor2_1 _08180_ (.A(\genblk2[3].wave_shpr.div.fin_quo[4] ),
    .B(_02886_),
    .Y(_02887_));
 sky130_fd_sc_hd__or3b_1 _08181_ (.A(\genblk2[3].wave_shpr.div.fin_quo[5] ),
    .B(_02885_),
    .C_N(_02887_),
    .X(_02888_));
 sky130_fd_sc_hd__a21oi_1 _08182_ (.A1(_02850_),
    .A2(_02888_),
    .B1(_02224_),
    .Y(_02889_));
 sky130_fd_sc_hd__o21ai_1 _08183_ (.A1(_02850_),
    .A2(_02888_),
    .B1(_02889_),
    .Y(_02890_));
 sky130_fd_sc_hd__nand2_1 _08184_ (.A(_02225_),
    .B(_02885_),
    .Y(_02891_));
 sky130_fd_sc_hd__nand2_1 _08185_ (.A(\genblk2[3].wave_shpr.div.fin_quo[7] ),
    .B(_02539_),
    .Y(_02892_));
 sky130_fd_sc_hd__nand3_1 _08186_ (.A(net9),
    .B(_02744_),
    .C(_02365_),
    .Y(_02893_));
 sky130_fd_sc_hd__a31o_1 _08187_ (.A1(_02890_),
    .A2(_02891_),
    .A3(_02892_),
    .B1(_02893_),
    .X(_02894_));
 sky130_fd_sc_hd__or2_1 _08188_ (.A(_02799_),
    .B(_02847_),
    .X(_02895_));
 sky130_fd_sc_hd__o21a_1 _08189_ (.A1(_02849_),
    .A2(_02894_),
    .B1(_02895_),
    .X(_02896_));
 sky130_fd_sc_hd__a21oi_1 _08190_ (.A1(_02697_),
    .A2(_02747_),
    .B1(_02896_),
    .Y(_02897_));
 sky130_fd_sc_hd__and3_1 _08191_ (.A(_02697_),
    .B(_02747_),
    .C(_02896_),
    .X(_02898_));
 sky130_fd_sc_hd__or2_1 _08192_ (.A(_02897_),
    .B(_02898_),
    .X(_02899_));
 sky130_fd_sc_hd__xnor2_1 _08193_ (.A(_02423_),
    .B(_02601_),
    .Y(_02900_));
 sky130_fd_sc_hd__and3_1 _08194_ (.A(net3),
    .B(net163),
    .C(_02312_),
    .X(_02901_));
 sky130_fd_sc_hd__a31oi_1 _08195_ (.A1(_02349_),
    .A2(_02351_),
    .A3(_02355_),
    .B1(\genblk2[11].wave_shpr.div.fin_quo[5] ),
    .Y(_02902_));
 sky130_fd_sc_hd__a41o_1 _08196_ (.A1(\genblk2[11].wave_shpr.div.fin_quo[5] ),
    .A2(net33),
    .A3(_02350_),
    .A4(_02355_),
    .B1(_02222_),
    .X(_02903_));
 sky130_fd_sc_hd__nand2_1 _08197_ (.A(\genblk2[11].wave_shpr.div.fin_quo[6] ),
    .B(_02361_),
    .Y(_02904_));
 sky130_fd_sc_hd__o211ai_2 _08198_ (.A1(_02902_),
    .A2(_02903_),
    .B1(_02904_),
    .C1(_02360_),
    .Y(_02905_));
 sky130_fd_sc_hd__o21ai_1 _08199_ (.A1(_02404_),
    .A2(_02410_),
    .B1(_02405_),
    .Y(_02906_));
 sky130_fd_sc_hd__o31a_1 _08200_ (.A1(_02405_),
    .A2(_02403_),
    .A3(_02410_),
    .B1(_02524_),
    .X(_02907_));
 sky130_fd_sc_hd__and3_1 _08201_ (.A(net17),
    .B(_02552_),
    .C(\genblk2[10].wave_shpr.div.fin_quo[6] ),
    .X(_02908_));
 sky130_fd_sc_hd__a211o_1 _08202_ (.A1(_02906_),
    .A2(_02907_),
    .B1(_02908_),
    .C1(_02416_),
    .X(_02909_));
 sky130_fd_sc_hd__a22o_1 _08203_ (.A1(_02901_),
    .A2(_02905_),
    .B1(_02909_),
    .B2(_02419_),
    .X(_02910_));
 sky130_fd_sc_hd__a21oi_1 _08204_ (.A1(_02303_),
    .A2(_02265_),
    .B1(\genblk2[9].wave_shpr.div.fin_quo[5] ),
    .Y(_02911_));
 sky130_fd_sc_hd__a31o_1 _08205_ (.A1(\genblk2[9].wave_shpr.div.fin_quo[5] ),
    .A2(_02303_),
    .A3(_02265_),
    .B1(_02316_),
    .X(_02912_));
 sky130_fd_sc_hd__a2bb2o_1 _08206_ (.A1_N(_02911_),
    .A2_N(_02912_),
    .B1(\genblk2[9].wave_shpr.div.fin_quo[6] ),
    .B2(_02362_),
    .X(_02913_));
 sky130_fd_sc_hd__o21a_1 _08207_ (.A1(_02310_),
    .A2(_02913_),
    .B1(_02314_),
    .X(_02914_));
 sky130_fd_sc_hd__and4_1 _08208_ (.A(_02901_),
    .B(_02419_),
    .C(_02905_),
    .D(_02909_),
    .X(_02915_));
 sky130_fd_sc_hd__a21oi_1 _08209_ (.A1(_02910_),
    .A2(_02914_),
    .B1(_02915_),
    .Y(_02916_));
 sky130_fd_sc_hd__xor2_1 _08210_ (.A(_02315_),
    .B(_02421_),
    .X(_02917_));
 sky130_fd_sc_hd__or2b_1 _08211_ (.A(_02916_),
    .B_N(_02917_),
    .X(_02918_));
 sky130_fd_sc_hd__a21o_1 _08212_ (.A1(_02697_),
    .A2(_02698_),
    .B1(_02746_),
    .X(_02919_));
 sky130_fd_sc_hd__xnor2_1 _08213_ (.A(_02917_),
    .B(_02916_),
    .Y(_02920_));
 sky130_fd_sc_hd__nand3_1 _08214_ (.A(_02747_),
    .B(_02919_),
    .C(_02920_),
    .Y(_02921_));
 sky130_fd_sc_hd__nand2_1 _08215_ (.A(_02918_),
    .B(_02921_),
    .Y(_02922_));
 sky130_fd_sc_hd__xnor2_1 _08216_ (.A(_02900_),
    .B(_02922_),
    .Y(_02923_));
 sky130_fd_sc_hd__or2b_1 _08217_ (.A(_02899_),
    .B_N(_02923_),
    .X(_02924_));
 sky130_fd_sc_hd__and2b_1 _08218_ (.A_N(_02900_),
    .B(_02922_),
    .X(_02925_));
 sky130_fd_sc_hd__xor2_1 _08219_ (.A(_02602_),
    .B(_02924_),
    .X(_02926_));
 sky130_fd_sc_hd__o21ai_1 _08220_ (.A1(_02925_),
    .A2(_02926_),
    .B1(_02897_),
    .Y(_02927_));
 sky130_fd_sc_hd__or3b_1 _08221_ (.A(_02793_),
    .B(_02789_),
    .C_N(\genblk2[5].wave_shpr.div.fin_quo[5] ),
    .X(_02928_));
 sky130_fd_sc_hd__o21bai_1 _08222_ (.A1(_02789_),
    .A2(_02793_),
    .B1_N(\genblk2[5].wave_shpr.div.fin_quo[5] ),
    .Y(_02929_));
 sky130_fd_sc_hd__a21o_1 _08223_ (.A1(\genblk2[5].wave_shpr.div.fin_quo[6] ),
    .A2(_02308_),
    .B1(_02791_),
    .X(_02930_));
 sky130_fd_sc_hd__a31o_1 _08224_ (.A1(_02527_),
    .A2(_02928_),
    .A3(_02929_),
    .B1(_02930_),
    .X(_02931_));
 sky130_fd_sc_hd__buf_2 _08225_ (.A(_02837_),
    .X(_02932_));
 sky130_fd_sc_hd__a21oi_1 _08226_ (.A1(_02932_),
    .A2(_02842_),
    .B1(\genblk2[4].wave_shpr.div.fin_quo[5] ),
    .Y(_02933_));
 sky130_fd_sc_hd__a31o_1 _08227_ (.A1(\genblk2[4].wave_shpr.div.fin_quo[5] ),
    .A2(_02932_),
    .A3(_02842_),
    .B1(_02316_),
    .X(_02934_));
 sky130_fd_sc_hd__a2bb2o_1 _08228_ (.A1_N(_02933_),
    .A2_N(_02934_),
    .B1(\genblk2[4].wave_shpr.div.fin_quo[6] ),
    .B2(_02362_),
    .X(_02935_));
 sky130_fd_sc_hd__o21a_1 _08229_ (.A1(_02838_),
    .A2(_02935_),
    .B1(_02846_),
    .X(_02936_));
 sky130_fd_sc_hd__nand2_1 _08230_ (.A(_02798_),
    .B(_02931_),
    .Y(_02937_));
 sky130_fd_sc_hd__xnor2_1 _08231_ (.A(_02937_),
    .B(_02936_),
    .Y(_02938_));
 sky130_fd_sc_hd__and2_2 _08232_ (.A(_02225_),
    .B(_02885_),
    .X(_02939_));
 sky130_fd_sc_hd__or3b_1 _08233_ (.A(_02887_),
    .B(_02885_),
    .C_N(\genblk2[3].wave_shpr.div.fin_quo[5] ),
    .X(_02940_));
 sky130_fd_sc_hd__o21bai_1 _08234_ (.A1(_02885_),
    .A2(_02887_),
    .B1_N(\genblk2[3].wave_shpr.div.fin_quo[5] ),
    .Y(_02941_));
 sky130_fd_sc_hd__a32o_1 _08235_ (.A1(_02592_),
    .A2(_02940_),
    .A3(_02941_),
    .B1(_02467_),
    .B2(\genblk2[3].wave_shpr.div.fin_quo[6] ),
    .X(_02942_));
 sky130_fd_sc_hd__and3_1 _08236_ (.A(net9),
    .B(_02744_),
    .C(_02365_),
    .X(_02943_));
 sky130_fd_sc_hd__o21a_1 _08237_ (.A1(_02939_),
    .A2(_02942_),
    .B1(_02943_),
    .X(_02944_));
 sky130_fd_sc_hd__a32o_1 _08238_ (.A1(_02798_),
    .A2(_02931_),
    .A3(_02936_),
    .B1(_02938_),
    .B2(_02944_),
    .X(_02945_));
 sky130_fd_sc_hd__or2_1 _08239_ (.A(_02646_),
    .B(_02647_),
    .X(_02946_));
 sky130_fd_sc_hd__o21a_1 _08240_ (.A1(_02682_),
    .A2(_02689_),
    .B1(_02683_),
    .X(_02947_));
 sky130_fd_sc_hd__o31ai_1 _08241_ (.A1(_02683_),
    .A2(_02682_),
    .A3(_02689_),
    .B1(_02527_),
    .Y(_02948_));
 sky130_fd_sc_hd__nand2_1 _08242_ (.A(\genblk2[7].wave_shpr.div.fin_quo[6] ),
    .B(_02309_),
    .Y(_02949_));
 sky130_fd_sc_hd__nand2_1 _08243_ (.A(_02225_),
    .B(_02682_),
    .Y(_02950_));
 sky130_fd_sc_hd__o211a_1 _08244_ (.A1(_02947_),
    .A2(_02948_),
    .B1(_02949_),
    .C1(_02950_),
    .X(_02951_));
 sky130_fd_sc_hd__inv_2 _08245_ (.A(_02641_),
    .Y(_02952_));
 sky130_fd_sc_hd__a21oi_1 _08246_ (.A1(_02638_),
    .A2(_02952_),
    .B1(\genblk2[8].wave_shpr.div.fin_quo[5] ),
    .Y(_02953_));
 sky130_fd_sc_hd__a31o_1 _08247_ (.A1(\genblk2[8].wave_shpr.div.fin_quo[5] ),
    .A2(_02638_),
    .A3(_02952_),
    .B1(_02223_),
    .X(_02954_));
 sky130_fd_sc_hd__nor2_1 _08248_ (.A(_02953_),
    .B(_02954_),
    .Y(_02955_));
 sky130_fd_sc_hd__a21o_1 _08249_ (.A1(\genblk2[8].wave_shpr.div.fin_quo[6] ),
    .A2(_02309_),
    .B1(_02636_),
    .X(_02956_));
 sky130_fd_sc_hd__o21ai_1 _08250_ (.A1(_02955_),
    .A2(_02956_),
    .B1(_02604_),
    .Y(_02957_));
 sky130_fd_sc_hd__o21ai_1 _08251_ (.A1(_02946_),
    .A2(_02951_),
    .B1(_02957_),
    .Y(_02958_));
 sky130_fd_sc_hd__inv_2 _08252_ (.A(_02738_),
    .Y(_02959_));
 sky130_fd_sc_hd__a21oi_1 _08253_ (.A1(_02734_),
    .A2(_02959_),
    .B1(\genblk2[6].wave_shpr.div.fin_quo[5] ),
    .Y(_02960_));
 sky130_fd_sc_hd__a31o_1 _08254_ (.A1(\genblk2[6].wave_shpr.div.fin_quo[5] ),
    .A2(_02733_),
    .A3(_02959_),
    .B1(_02261_),
    .X(_02961_));
 sky130_fd_sc_hd__a2bb2o_1 _08255_ (.A1_N(_02960_),
    .A2_N(_02961_),
    .B1(\genblk2[6].wave_shpr.div.fin_quo[6] ),
    .B2(_02539_),
    .X(_02962_));
 sky130_fd_sc_hd__o21a_1 _08256_ (.A1(_02742_),
    .A2(_02962_),
    .B1(_02745_),
    .X(_02963_));
 sky130_fd_sc_hd__or3_1 _08257_ (.A(_02946_),
    .B(_02957_),
    .C(_02951_),
    .X(_02964_));
 sky130_fd_sc_hd__a21bo_1 _08258_ (.A1(_02958_),
    .A2(_02963_),
    .B1_N(_02964_),
    .X(_02965_));
 sky130_fd_sc_hd__xor2_2 _08259_ (.A(_02848_),
    .B(_02894_),
    .X(_02966_));
 sky130_fd_sc_hd__xnor2_1 _08260_ (.A(_02965_),
    .B(_02966_),
    .Y(_02967_));
 sky130_fd_sc_hd__and2b_1 _08261_ (.A_N(_02966_),
    .B(_02965_),
    .X(_02968_));
 sky130_fd_sc_hd__a21o_1 _08262_ (.A1(_02945_),
    .A2(_02967_),
    .B1(_02968_),
    .X(_02969_));
 sky130_fd_sc_hd__xnor2_1 _08263_ (.A(_02899_),
    .B(_02923_),
    .Y(_02970_));
 sky130_fd_sc_hd__or2b_1 _08264_ (.A(_02915_),
    .B_N(_02910_),
    .X(_02971_));
 sky130_fd_sc_hd__xor2_1 _08265_ (.A(_02971_),
    .B(_02914_),
    .X(_02972_));
 sky130_fd_sc_hd__a31oi_1 _08266_ (.A1(_02349_),
    .A2(_02351_),
    .A3(_02354_),
    .B1(\genblk2[11].wave_shpr.div.fin_quo[4] ),
    .Y(_02973_));
 sky130_fd_sc_hd__a41o_1 _08267_ (.A1(\genblk2[11].wave_shpr.div.fin_quo[4] ),
    .A2(net33),
    .A3(_02350_),
    .A4(_02354_),
    .B1(_02222_),
    .X(_02974_));
 sky130_fd_sc_hd__nand2_1 _08268_ (.A(\genblk2[11].wave_shpr.div.fin_quo[5] ),
    .B(_02361_),
    .Y(_02975_));
 sky130_fd_sc_hd__o211a_1 _08269_ (.A1(_02973_),
    .A2(_02974_),
    .B1(_02975_),
    .C1(_02360_),
    .X(_02976_));
 sky130_fd_sc_hd__nor2_1 _08270_ (.A(_02366_),
    .B(_02976_),
    .Y(_02977_));
 sky130_fd_sc_hd__inv_2 _08271_ (.A(_02409_),
    .Y(_02978_));
 sky130_fd_sc_hd__inv_2 _08272_ (.A(\genblk2[10].wave_shpr.div.fin_quo[4] ),
    .Y(_02979_));
 sky130_fd_sc_hd__o21ai_1 _08273_ (.A1(_02404_),
    .A2(_02978_),
    .B1(_02979_),
    .Y(_02980_));
 sky130_fd_sc_hd__o31a_1 _08274_ (.A1(_02979_),
    .A2(_02404_),
    .A3(_02978_),
    .B1(_02525_),
    .X(_02981_));
 sky130_fd_sc_hd__a22o_1 _08275_ (.A1(\genblk2[10].wave_shpr.div.fin_quo[5] ),
    .A2(_02361_),
    .B1(_02980_),
    .B2(_02981_),
    .X(_02982_));
 sky130_fd_sc_hd__o21ai_2 _08276_ (.A1(_02416_),
    .A2(_02982_),
    .B1(_02419_),
    .Y(_02983_));
 sky130_fd_sc_hd__and2b_1 _08277_ (.A_N(_02977_),
    .B(_02983_),
    .X(_02984_));
 sky130_fd_sc_hd__a21oi_1 _08278_ (.A1(_02303_),
    .A2(_02264_),
    .B1(\genblk2[9].wave_shpr.div.fin_quo[4] ),
    .Y(_02985_));
 sky130_fd_sc_hd__a31o_1 _08279_ (.A1(\genblk2[9].wave_shpr.div.fin_quo[4] ),
    .A2(_02303_),
    .A3(_02264_),
    .B1(_02223_),
    .X(_02986_));
 sky130_fd_sc_hd__nor2_1 _08280_ (.A(_02985_),
    .B(_02986_),
    .Y(_02987_));
 sky130_fd_sc_hd__a21o_1 _08281_ (.A1(\genblk2[9].wave_shpr.div.fin_quo[5] ),
    .A2(_02521_),
    .B1(_02310_),
    .X(_02988_));
 sky130_fd_sc_hd__o21ai_1 _08282_ (.A1(_02987_),
    .A2(_02988_),
    .B1(_02314_),
    .Y(_02989_));
 sky130_fd_sc_hd__or3_1 _08283_ (.A(_02366_),
    .B(_02976_),
    .C(_02983_),
    .X(_02990_));
 sky130_fd_sc_hd__o21ai_1 _08284_ (.A1(_02984_),
    .A2(_02989_),
    .B1(_02990_),
    .Y(_02991_));
 sky130_fd_sc_hd__and2b_1 _08285_ (.A_N(_02972_),
    .B(_02991_),
    .X(_02992_));
 sky130_fd_sc_hd__nand3_1 _08286_ (.A(_02964_),
    .B(_02958_),
    .C(_02963_),
    .Y(_02993_));
 sky130_fd_sc_hd__a21o_1 _08287_ (.A1(_02964_),
    .A2(_02958_),
    .B1(_02963_),
    .X(_02994_));
 sky130_fd_sc_hd__xnor2_1 _08288_ (.A(_02972_),
    .B(_02991_),
    .Y(_02995_));
 sky130_fd_sc_hd__and3_1 _08289_ (.A(_02993_),
    .B(_02994_),
    .C(_02995_),
    .X(_02996_));
 sky130_fd_sc_hd__a21o_1 _08290_ (.A1(_02747_),
    .A2(_02919_),
    .B1(_02920_),
    .X(_02997_));
 sky130_fd_sc_hd__o211a_1 _08291_ (.A1(_02992_),
    .A2(_02996_),
    .B1(_02921_),
    .C1(_02997_),
    .X(_02998_));
 sky130_fd_sc_hd__xnor2_1 _08292_ (.A(_02945_),
    .B(_02967_),
    .Y(_02999_));
 sky130_fd_sc_hd__a211oi_1 _08293_ (.A1(_02921_),
    .A2(_02997_),
    .B1(_02992_),
    .C1(_02996_),
    .Y(_03000_));
 sky130_fd_sc_hd__nor3_1 _08294_ (.A(_02998_),
    .B(_02999_),
    .C(_03000_),
    .Y(_03001_));
 sky130_fd_sc_hd__nor2_1 _08295_ (.A(_02998_),
    .B(_03001_),
    .Y(_03002_));
 sky130_fd_sc_hd__xnor2_1 _08296_ (.A(_02970_),
    .B(_03002_),
    .Y(_03003_));
 sky130_fd_sc_hd__and2b_1 _08297_ (.A_N(_03002_),
    .B(_02970_),
    .X(_03004_));
 sky130_fd_sc_hd__a21oi_1 _08298_ (.A1(_02969_),
    .A2(_03003_),
    .B1(_03004_),
    .Y(_03005_));
 sky130_fd_sc_hd__or3_1 _08299_ (.A(_02897_),
    .B(_02925_),
    .C(_02926_),
    .X(_03006_));
 sky130_fd_sc_hd__and2_1 _08300_ (.A(_02927_),
    .B(_03006_),
    .X(_03007_));
 sky130_fd_sc_hd__or2b_1 _08301_ (.A(_03005_),
    .B_N(_03007_),
    .X(_03008_));
 sky130_fd_sc_hd__o211a_1 _08302_ (.A1(_02602_),
    .A2(_02924_),
    .B1(_02927_),
    .C1(_03008_),
    .X(_03009_));
 sky130_fd_sc_hd__xnor2_1 _08303_ (.A(_03007_),
    .B(_03005_),
    .Y(_03010_));
 sky130_fd_sc_hd__xnor2_1 _08304_ (.A(_02969_),
    .B(_03003_),
    .Y(_03011_));
 sky130_fd_sc_hd__xnor2_1 _08305_ (.A(_02977_),
    .B(_02983_),
    .Y(_03012_));
 sky130_fd_sc_hd__xnor2_1 _08306_ (.A(_03012_),
    .B(_02989_),
    .Y(_03013_));
 sky130_fd_sc_hd__a31oi_1 _08307_ (.A1(_02349_),
    .A2(_02351_),
    .A3(_02353_),
    .B1(\genblk2[11].wave_shpr.div.fin_quo[3] ),
    .Y(_03014_));
 sky130_fd_sc_hd__a41o_1 _08308_ (.A1(\genblk2[11].wave_shpr.div.fin_quo[3] ),
    .A2(_02349_),
    .A3(_02351_),
    .A4(_02353_),
    .B1(_02222_),
    .X(_03015_));
 sky130_fd_sc_hd__nand2_1 _08309_ (.A(\genblk2[11].wave_shpr.div.fin_quo[4] ),
    .B(_02361_),
    .Y(_03016_));
 sky130_fd_sc_hd__o211a_1 _08310_ (.A1(_03014_),
    .A2(_03015_),
    .B1(_03016_),
    .C1(_02360_),
    .X(_03017_));
 sky130_fd_sc_hd__nor2_1 _08311_ (.A(_02366_),
    .B(_03017_),
    .Y(_03018_));
 sky130_fd_sc_hd__o21ai_1 _08312_ (.A1(_02404_),
    .A2(_02408_),
    .B1(_02406_),
    .Y(_03019_));
 sky130_fd_sc_hd__o31a_1 _08313_ (.A1(_02406_),
    .A2(_02404_),
    .A3(_02408_),
    .B1(_02525_),
    .X(_03020_));
 sky130_fd_sc_hd__and3_1 _08314_ (.A(_02216_),
    .B(_02552_),
    .C(\genblk2[10].wave_shpr.div.fin_quo[4] ),
    .X(_03021_));
 sky130_fd_sc_hd__a211o_1 _08315_ (.A1(_03019_),
    .A2(_03020_),
    .B1(_03021_),
    .C1(_02416_),
    .X(_03022_));
 sky130_fd_sc_hd__nand2_1 _08316_ (.A(_02419_),
    .B(_03022_),
    .Y(_03023_));
 sky130_fd_sc_hd__xnor2_2 _08317_ (.A(_03018_),
    .B(_03023_),
    .Y(_03024_));
 sky130_fd_sc_hd__a21oi_1 _08318_ (.A1(_02303_),
    .A2(_02263_),
    .B1(\genblk2[9].wave_shpr.div.fin_quo[3] ),
    .Y(_03025_));
 sky130_fd_sc_hd__a31o_1 _08319_ (.A1(\genblk2[9].wave_shpr.div.fin_quo[3] ),
    .A2(_02303_),
    .A3(_02263_),
    .B1(_02316_),
    .X(_03026_));
 sky130_fd_sc_hd__a2bb2o_1 _08320_ (.A1_N(_03025_),
    .A2_N(_03026_),
    .B1(\genblk2[9].wave_shpr.div.fin_quo[4] ),
    .B2(_02362_),
    .X(_03027_));
 sky130_fd_sc_hd__o21a_1 _08321_ (.A1(_02310_),
    .A2(_03027_),
    .B1(_02314_),
    .X(_03028_));
 sky130_fd_sc_hd__a32o_1 _08322_ (.A1(_02419_),
    .A2(_03018_),
    .A3(_03022_),
    .B1(_03024_),
    .B2(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__and2_1 _08323_ (.A(_03013_),
    .B(_03029_),
    .X(_03030_));
 sky130_fd_sc_hd__a21oi_1 _08324_ (.A1(_02638_),
    .A2(_02640_),
    .B1(\genblk2[8].wave_shpr.div.fin_quo[4] ),
    .Y(_03031_));
 sky130_fd_sc_hd__a31o_1 _08325_ (.A1(\genblk2[8].wave_shpr.div.fin_quo[4] ),
    .A2(_02638_),
    .A3(_02640_),
    .B1(_02223_),
    .X(_03032_));
 sky130_fd_sc_hd__nor2_1 _08326_ (.A(_03031_),
    .B(_03032_),
    .Y(_03033_));
 sky130_fd_sc_hd__a211o_1 _08327_ (.A1(\genblk2[8].wave_shpr.div.fin_quo[5] ),
    .A2(_02467_),
    .B1(_03033_),
    .C1(_02636_),
    .X(_03034_));
 sky130_fd_sc_hd__inv_2 _08328_ (.A(_02688_),
    .Y(_03035_));
 sky130_fd_sc_hd__inv_2 _08329_ (.A(\genblk2[7].wave_shpr.div.fin_quo[4] ),
    .Y(_03036_));
 sky130_fd_sc_hd__o21ai_1 _08330_ (.A1(_02682_),
    .A2(_03035_),
    .B1(_03036_),
    .Y(_03037_));
 sky130_fd_sc_hd__o31a_1 _08331_ (.A1(_03036_),
    .A2(_02682_),
    .A3(_03035_),
    .B1(_02526_),
    .X(_03038_));
 sky130_fd_sc_hd__and3_1 _08332_ (.A(_02217_),
    .B(_02553_),
    .C(\genblk2[7].wave_shpr.div.fin_quo[5] ),
    .X(_03039_));
 sky130_fd_sc_hd__a211o_1 _08333_ (.A1(_03037_),
    .A2(_03038_),
    .B1(_03039_),
    .C1(_02694_),
    .X(_03040_));
 sky130_fd_sc_hd__nand4_2 _08334_ (.A(_02604_),
    .B(_02648_),
    .C(_03034_),
    .D(_03040_),
    .Y(_03041_));
 sky130_fd_sc_hd__a22o_1 _08335_ (.A1(_02604_),
    .A2(_03034_),
    .B1(_03040_),
    .B2(_02648_),
    .X(_03042_));
 sky130_fd_sc_hd__a21oi_1 _08336_ (.A1(_02734_),
    .A2(_02737_),
    .B1(\genblk2[6].wave_shpr.div.fin_quo[4] ),
    .Y(_03043_));
 sky130_fd_sc_hd__a31o_1 _08337_ (.A1(\genblk2[6].wave_shpr.div.fin_quo[4] ),
    .A2(_02734_),
    .A3(_02737_),
    .B1(_02261_),
    .X(_03044_));
 sky130_fd_sc_hd__nor2_1 _08338_ (.A(_03043_),
    .B(_03044_),
    .Y(_03045_));
 sky130_fd_sc_hd__a21o_1 _08339_ (.A1(\genblk2[6].wave_shpr.div.fin_quo[5] ),
    .A2(_02467_),
    .B1(_02742_),
    .X(_03046_));
 sky130_fd_sc_hd__o21a_1 _08340_ (.A1(_03045_),
    .A2(_03046_),
    .B1(_02745_),
    .X(_03047_));
 sky130_fd_sc_hd__nand3_1 _08341_ (.A(_03041_),
    .B(_03042_),
    .C(_03047_),
    .Y(_03048_));
 sky130_fd_sc_hd__a21o_1 _08342_ (.A1(_03041_),
    .A2(_03042_),
    .B1(_03047_),
    .X(_03049_));
 sky130_fd_sc_hd__xor2_1 _08343_ (.A(_03013_),
    .B(_03029_),
    .X(_03050_));
 sky130_fd_sc_hd__and3_2 _08344_ (.A(_03048_),
    .B(_03049_),
    .C(_03050_),
    .X(_03051_));
 sky130_fd_sc_hd__nand3_1 _08345_ (.A(_02993_),
    .B(_02994_),
    .C(_02995_),
    .Y(_03052_));
 sky130_fd_sc_hd__a21o_1 _08346_ (.A1(_02993_),
    .A2(_02994_),
    .B1(_02995_),
    .X(_03053_));
 sky130_fd_sc_hd__o211a_1 _08347_ (.A1(_03030_),
    .A2(_03051_),
    .B1(_03052_),
    .C1(_03053_),
    .X(_03054_));
 sky130_fd_sc_hd__inv_2 _08348_ (.A(_03054_),
    .Y(_03055_));
 sky130_fd_sc_hd__and2b_1 _08349_ (.A_N(_02789_),
    .B(_02792_),
    .X(_03056_));
 sky130_fd_sc_hd__o21ai_1 _08350_ (.A1(\genblk2[5].wave_shpr.div.fin_quo[4] ),
    .A2(_03056_),
    .B1(_02527_),
    .Y(_03057_));
 sky130_fd_sc_hd__a21oi_1 _08351_ (.A1(\genblk2[5].wave_shpr.div.fin_quo[4] ),
    .A2(_03056_),
    .B1(_03057_),
    .Y(_03058_));
 sky130_fd_sc_hd__a21o_1 _08352_ (.A1(\genblk2[5].wave_shpr.div.fin_quo[5] ),
    .A2(_02521_),
    .B1(_02791_),
    .X(_03059_));
 sky130_fd_sc_hd__o21a_1 _08353_ (.A1(_03058_),
    .A2(_03059_),
    .B1(_02798_),
    .X(_03060_));
 sky130_fd_sc_hd__a21oi_1 _08354_ (.A1(_02932_),
    .A2(_02841_),
    .B1(\genblk2[4].wave_shpr.div.fin_quo[4] ),
    .Y(_03061_));
 sky130_fd_sc_hd__a31o_1 _08355_ (.A1(\genblk2[4].wave_shpr.div.fin_quo[4] ),
    .A2(_02932_),
    .A3(_02841_),
    .B1(_02222_),
    .X(_03062_));
 sky130_fd_sc_hd__nor2_1 _08356_ (.A(_03061_),
    .B(_03062_),
    .Y(_03063_));
 sky130_fd_sc_hd__a211o_1 _08357_ (.A1(\genblk2[4].wave_shpr.div.fin_quo[5] ),
    .A2(_02521_),
    .B1(_02838_),
    .C1(_03063_),
    .X(_03064_));
 sky130_fd_sc_hd__and2_1 _08358_ (.A(_02846_),
    .B(_03064_),
    .X(_03065_));
 sky130_fd_sc_hd__xor2_1 _08359_ (.A(_03060_),
    .B(_03065_),
    .X(_03066_));
 sky130_fd_sc_hd__or2b_1 _08360_ (.A(_02885_),
    .B_N(_02886_),
    .X(_03067_));
 sky130_fd_sc_hd__xnor2_1 _08361_ (.A(\genblk2[3].wave_shpr.div.fin_quo[4] ),
    .B(_03067_),
    .Y(_03068_));
 sky130_fd_sc_hd__a22o_1 _08362_ (.A1(\genblk2[3].wave_shpr.div.fin_quo[5] ),
    .A2(_02539_),
    .B1(_03068_),
    .B2(_02592_),
    .X(_03069_));
 sky130_fd_sc_hd__o21a_1 _08363_ (.A1(_02939_),
    .A2(_03069_),
    .B1(_02943_),
    .X(_03070_));
 sky130_fd_sc_hd__a32o_1 _08364_ (.A1(_02846_),
    .A2(_03060_),
    .A3(_03064_),
    .B1(_03066_),
    .B2(_03070_),
    .X(_03071_));
 sky130_fd_sc_hd__a21bo_1 _08365_ (.A1(_03042_),
    .A2(_03047_),
    .B1_N(_03041_),
    .X(_03072_));
 sky130_fd_sc_hd__xnor2_1 _08366_ (.A(_02938_),
    .B(_02944_),
    .Y(_03073_));
 sky130_fd_sc_hd__xnor2_1 _08367_ (.A(_03072_),
    .B(_03073_),
    .Y(_03074_));
 sky130_fd_sc_hd__xnor2_1 _08368_ (.A(_03071_),
    .B(_03074_),
    .Y(_03075_));
 sky130_fd_sc_hd__a211oi_1 _08369_ (.A1(_03052_),
    .A2(_03053_),
    .B1(_03030_),
    .C1(_03051_),
    .Y(_03076_));
 sky130_fd_sc_hd__or3_2 _08370_ (.A(_03054_),
    .B(_03075_),
    .C(_03076_),
    .X(_03077_));
 sky130_fd_sc_hd__o21a_1 _08371_ (.A1(_02998_),
    .A2(_03000_),
    .B1(_02999_),
    .X(_03078_));
 sky130_fd_sc_hd__a211oi_1 _08372_ (.A1(_03055_),
    .A2(_03077_),
    .B1(_03001_),
    .C1(_03078_),
    .Y(_03079_));
 sky130_fd_sc_hd__inv_2 _08373_ (.A(_02599_),
    .Y(_03080_));
 sky130_fd_sc_hd__o211ai_1 _08374_ (.A1(_02520_),
    .A2(net1354),
    .B1(_03080_),
    .C1(_02600_),
    .Y(_03081_));
 sky130_fd_sc_hd__a211o_1 _08375_ (.A1(_02600_),
    .A2(_03080_),
    .B1(net24),
    .C1(_02520_),
    .X(_03082_));
 sky130_fd_sc_hd__nand2_1 _08376_ (.A(_03081_),
    .B(_03082_),
    .Y(_03083_));
 sky130_fd_sc_hd__and2b_1 _08377_ (.A_N(_03073_),
    .B(_03072_),
    .X(_03084_));
 sky130_fd_sc_hd__a21oi_1 _08378_ (.A1(_03071_),
    .A2(_03074_),
    .B1(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__nand2_1 _08379_ (.A(\genblk1[2].osc.clkdiv_C.cnt[6] ),
    .B(_01433_),
    .Y(_03086_));
 sky130_fd_sc_hd__o211a_1 _08380_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[1] ),
    .A2(_01209_),
    .B1(_02425_),
    .C1(\genblk1[2].osc.clkdiv_C.cnt[0] ),
    .X(_03087_));
 sky130_fd_sc_hd__a22o_1 _08381_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[1] ),
    .A2(_01209_),
    .B1(_02336_),
    .B2(\genblk1[2].osc.clkdiv_C.cnt[2] ),
    .X(_03088_));
 sky130_fd_sc_hd__o22a_1 _08382_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[2] ),
    .A2(_02336_),
    .B1(_01418_),
    .B2(\genblk1[2].osc.clkdiv_C.cnt[3] ),
    .X(_03089_));
 sky130_fd_sc_hd__o21a_1 _08383_ (.A1(_03087_),
    .A2(_03088_),
    .B1(_03089_),
    .X(_03090_));
 sky130_fd_sc_hd__and2b_1 _08384_ (.A_N(_01437_),
    .B(\genblk1[2].osc.clkdiv_C.cnt[5] ),
    .X(_03091_));
 sky130_fd_sc_hd__a221o_1 _08385_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[4] ),
    .A2(_01439_),
    .B1(_01418_),
    .B2(\genblk1[2].osc.clkdiv_C.cnt[3] ),
    .C1(_03091_),
    .X(_03092_));
 sky130_fd_sc_hd__a211o_1 _08386_ (.A1(_01200_),
    .A2(\genblk1[2].osc.clkdiv_C.cnt[4] ),
    .B1(\genblk1[2].osc.clkdiv_C.cnt[5] ),
    .C1(_01441_),
    .X(_03093_));
 sky130_fd_sc_hd__o21a_1 _08387_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[6] ),
    .A2(_01433_),
    .B1(_03093_),
    .X(_03094_));
 sky130_fd_sc_hd__o21ai_1 _08388_ (.A1(_03090_),
    .A2(_03092_),
    .B1(_03094_),
    .Y(_03095_));
 sky130_fd_sc_hd__o2bb2a_1 _08389_ (.A1_N(_03086_),
    .A2_N(_03095_),
    .B1(\genblk1[2].osc.clkdiv_C.cnt[7] ),
    .B2(_02011_),
    .X(_03096_));
 sky130_fd_sc_hd__a22o_1 _08390_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[8] ),
    .A2(_01442_),
    .B1(_02011_),
    .B2(\genblk1[2].osc.clkdiv_C.cnt[7] ),
    .X(_03097_));
 sky130_fd_sc_hd__nand2_1 _08391_ (.A(_01412_),
    .B(_01302_),
    .Y(_03098_));
 sky130_fd_sc_hd__o221a_1 _08392_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[9] ),
    .A2(_01431_),
    .B1(_03096_),
    .B2(_03097_),
    .C1(_03098_),
    .X(_03099_));
 sky130_fd_sc_hd__a22o_1 _08393_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[10] ),
    .A2(_01420_),
    .B1(_01431_),
    .B2(\genblk1[2].osc.clkdiv_C.cnt[9] ),
    .X(_03100_));
 sky130_fd_sc_hd__or2_1 _08394_ (.A(\genblk1[2].osc.clkdiv_C.cnt[11] ),
    .B(_01411_),
    .X(_03101_));
 sky130_fd_sc_hd__o221a_1 _08395_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[10] ),
    .A2(_01420_),
    .B1(_03099_),
    .B2(_03100_),
    .C1(_03101_),
    .X(_03102_));
 sky130_fd_sc_hd__o22ai_1 _08396_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[15] ),
    .A2(_01349_),
    .B1(_01209_),
    .B2(\genblk1[2].osc.clkdiv_C.cnt[14] ),
    .Y(_03103_));
 sky130_fd_sc_hd__a22o_1 _08397_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[14] ),
    .A2(_01209_),
    .B1(_02425_),
    .B2(\genblk1[2].osc.clkdiv_C.cnt[13] ),
    .X(_03104_));
 sky130_fd_sc_hd__nand2_1 _08398_ (.A(\genblk1[2].osc.clkdiv_C.cnt[15] ),
    .B(_01349_),
    .Y(_03105_));
 sky130_fd_sc_hd__or3b_1 _08399_ (.A(_03103_),
    .B(_03104_),
    .C_N(_03105_),
    .X(_03106_));
 sky130_fd_sc_hd__o22a_1 _08400_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[13] ),
    .A2(_02425_),
    .B1(_01591_),
    .B2(\genblk1[2].osc.clkdiv_C.cnt[12] ),
    .X(_03107_));
 sky130_fd_sc_hd__a21bo_1 _08401_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[12] ),
    .A2(_01591_),
    .B1_N(_03107_),
    .X(_03108_));
 sky130_fd_sc_hd__a2111o_1 _08402_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[11] ),
    .A2(_01411_),
    .B1(_03102_),
    .C1(_03106_),
    .D1(_03108_),
    .X(_03109_));
 sky130_fd_sc_hd__o2bb2a_1 _08403_ (.A1_N(_03103_),
    .A2_N(_03105_),
    .B1(_03106_),
    .B2(_03107_),
    .X(_03110_));
 sky130_fd_sc_hd__o311a_1 _08404_ (.A1(_01201_),
    .A2(\genblk1[2].osc.clkdiv_C.cnt[16] ),
    .A3(_01362_),
    .B1(_03109_),
    .C1(_03110_),
    .X(_03111_));
 sky130_fd_sc_hd__a211oi_1 _08405_ (.A1(\genblk1[2].osc.clkdiv_C.cnt[16] ),
    .A2(_01578_),
    .B1(_03111_),
    .C1(\genblk1[2].osc.clkdiv_C.cnt[17] ),
    .Y(_03112_));
 sky130_fd_sc_hd__buf_2 _08406_ (.A(net25),
    .X(_03113_));
 sky130_fd_sc_hd__nor2_2 _08407_ (.A(_02221_),
    .B(_03113_),
    .Y(_03114_));
 sky130_fd_sc_hd__or2_1 _08408_ (.A(\genblk2[2].wave_shpr.div.fin_quo[0] ),
    .B(\genblk2[2].wave_shpr.div.fin_quo[1] ),
    .X(_03115_));
 sky130_fd_sc_hd__or2_1 _08409_ (.A(\genblk2[2].wave_shpr.div.fin_quo[2] ),
    .B(_03115_),
    .X(_03116_));
 sky130_fd_sc_hd__or2_1 _08410_ (.A(\genblk2[2].wave_shpr.div.fin_quo[3] ),
    .B(_03116_),
    .X(_03117_));
 sky130_fd_sc_hd__or2_1 _08411_ (.A(\genblk2[2].wave_shpr.div.fin_quo[4] ),
    .B(_03117_),
    .X(_03118_));
 sky130_fd_sc_hd__or3b_1 _08412_ (.A(_03118_),
    .B(\genblk2[2].wave_shpr.div.fin_quo[5] ),
    .C_N(net25),
    .X(_03119_));
 sky130_fd_sc_hd__xnor2_1 _08413_ (.A(\genblk2[2].wave_shpr.div.fin_quo[6] ),
    .B(_03119_),
    .Y(_03120_));
 sky130_fd_sc_hd__a22o_1 _08414_ (.A1(\genblk2[2].wave_shpr.div.fin_quo[7] ),
    .A2(_02468_),
    .B1(_03120_),
    .B2(_02592_),
    .X(_03121_));
 sky130_fd_sc_hd__and3_2 _08415_ (.A(net8),
    .B(_02744_),
    .C(_02365_),
    .X(_03122_));
 sky130_fd_sc_hd__o21ai_1 _08416_ (.A1(_03114_),
    .A2(_03121_),
    .B1(_03122_),
    .Y(_03123_));
 sky130_fd_sc_hd__xnor2_1 _08417_ (.A(_03085_),
    .B(_03123_),
    .Y(_03124_));
 sky130_fd_sc_hd__xnor2_1 _08418_ (.A(_03083_),
    .B(_03124_),
    .Y(_03125_));
 sky130_fd_sc_hd__o211a_1 _08419_ (.A1(_03001_),
    .A2(_03078_),
    .B1(_03055_),
    .C1(_03077_),
    .X(_03126_));
 sky130_fd_sc_hd__or3_1 _08420_ (.A(_03079_),
    .B(_03125_),
    .C(_03126_),
    .X(_03127_));
 sky130_fd_sc_hd__or2b_1 _08421_ (.A(_03079_),
    .B_N(_03127_),
    .X(_03128_));
 sky130_fd_sc_hd__and2b_1 _08422_ (.A_N(_03011_),
    .B(_03128_),
    .X(_03129_));
 sky130_fd_sc_hd__or2_1 _08423_ (.A(_03085_),
    .B(_03123_),
    .X(_03130_));
 sky130_fd_sc_hd__o21a_1 _08424_ (.A1(_03083_),
    .A2(_03124_),
    .B1(_03130_),
    .X(_03131_));
 sky130_fd_sc_hd__xnor2_1 _08425_ (.A(_03011_),
    .B(_03128_),
    .Y(_03132_));
 sky130_fd_sc_hd__and2b_1 _08426_ (.A_N(_03131_),
    .B(_03132_),
    .X(_03133_));
 sky130_fd_sc_hd__nor3_1 _08427_ (.A(_03010_),
    .B(_03129_),
    .C(_03133_),
    .Y(_03134_));
 sky130_fd_sc_hd__o21a_1 _08428_ (.A1(_03129_),
    .A2(_03133_),
    .B1(_03010_),
    .X(_03135_));
 sky130_fd_sc_hd__xor2_1 _08429_ (.A(_03131_),
    .B(_03132_),
    .X(_03136_));
 sky130_fd_sc_hd__a21oi_1 _08430_ (.A1(_02303_),
    .A2(_02262_),
    .B1(\genblk2[9].wave_shpr.div.fin_quo[2] ),
    .Y(_03137_));
 sky130_fd_sc_hd__a31o_1 _08431_ (.A1(\genblk2[9].wave_shpr.div.fin_quo[2] ),
    .A2(net32),
    .A3(_02262_),
    .B1(_02222_),
    .X(_03138_));
 sky130_fd_sc_hd__a2bb2o_1 _08432_ (.A1_N(_03137_),
    .A2_N(_03138_),
    .B1(\genblk2[9].wave_shpr.div.fin_quo[3] ),
    .B2(_02308_),
    .X(_03139_));
 sky130_fd_sc_hd__o21a_1 _08433_ (.A1(_02310_),
    .A2(_03139_),
    .B1(_02314_),
    .X(_03140_));
 sky130_fd_sc_hd__a21oi_2 _08434_ (.A1(_02349_),
    .A2(_02351_),
    .B1(_02221_),
    .Y(_03141_));
 sky130_fd_sc_hd__a31o_1 _08435_ (.A1(net33),
    .A2(_02350_),
    .A3(_02352_),
    .B1(\genblk2[11].wave_shpr.div.fin_quo[2] ),
    .X(_03142_));
 sky130_fd_sc_hd__nand4_1 _08436_ (.A(\genblk2[11].wave_shpr.div.fin_quo[2] ),
    .B(_02349_),
    .C(_02351_),
    .D(_02352_),
    .Y(_03143_));
 sky130_fd_sc_hd__a32o_1 _08437_ (.A1(_02525_),
    .A2(_03142_),
    .A3(_03143_),
    .B1(_02361_),
    .B2(\genblk2[11].wave_shpr.div.fin_quo[3] ),
    .X(_03144_));
 sky130_fd_sc_hd__o21a_1 _08438_ (.A1(_03141_),
    .A2(_03144_),
    .B1(_02901_),
    .X(_03145_));
 sky130_fd_sc_hd__o21bai_1 _08439_ (.A1(_02404_),
    .A2(_02407_),
    .B1_N(\genblk2[10].wave_shpr.div.fin_quo[2] ),
    .Y(_03146_));
 sky130_fd_sc_hd__or3b_1 _08440_ (.A(_02407_),
    .B(_02403_),
    .C_N(\genblk2[10].wave_shpr.div.fin_quo[2] ),
    .X(_03147_));
 sky130_fd_sc_hd__a32o_1 _08441_ (.A1(_02525_),
    .A2(_03146_),
    .A3(_03147_),
    .B1(_02361_),
    .B2(\genblk2[10].wave_shpr.div.fin_quo[3] ),
    .X(_03148_));
 sky130_fd_sc_hd__o21a_1 _08442_ (.A1(_02416_),
    .A2(_03148_),
    .B1(_02419_),
    .X(_03149_));
 sky130_fd_sc_hd__xor2_2 _08443_ (.A(_03145_),
    .B(_03149_),
    .X(_03150_));
 sky130_fd_sc_hd__nand2_1 _08444_ (.A(_03145_),
    .B(_03149_),
    .Y(_03151_));
 sky130_fd_sc_hd__a21boi_2 _08445_ (.A1(_03140_),
    .A2(_03150_),
    .B1_N(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__xor2_2 _08446_ (.A(_03024_),
    .B(_03028_),
    .X(_03153_));
 sky130_fd_sc_hd__or2b_1 _08447_ (.A(_03152_),
    .B_N(_03153_),
    .X(_03154_));
 sky130_fd_sc_hd__a21oi_1 _08448_ (.A1(_02638_),
    .A2(_02639_),
    .B1(\genblk2[8].wave_shpr.div.fin_quo[3] ),
    .Y(_03155_));
 sky130_fd_sc_hd__a31o_1 _08449_ (.A1(\genblk2[8].wave_shpr.div.fin_quo[3] ),
    .A2(net30),
    .A3(_02639_),
    .B1(_02316_),
    .X(_03156_));
 sky130_fd_sc_hd__a2bb2o_1 _08450_ (.A1_N(_03155_),
    .A2_N(_03156_),
    .B1(\genblk2[8].wave_shpr.div.fin_quo[4] ),
    .B2(_02521_),
    .X(_03157_));
 sky130_fd_sc_hd__o21ai_1 _08451_ (.A1(_02636_),
    .A2(_03157_),
    .B1(_02604_),
    .Y(_03158_));
 sky130_fd_sc_hd__o21ai_1 _08452_ (.A1(_02682_),
    .A2(_02687_),
    .B1(_02684_),
    .Y(_03159_));
 sky130_fd_sc_hd__o31a_1 _08453_ (.A1(_02684_),
    .A2(_02681_),
    .A3(_02687_),
    .B1(_02526_),
    .X(_03160_));
 sky130_fd_sc_hd__and3_1 _08454_ (.A(_02216_),
    .B(_02553_),
    .C(\genblk2[7].wave_shpr.div.fin_quo[4] ),
    .X(_03161_));
 sky130_fd_sc_hd__a211o_1 _08455_ (.A1(_03159_),
    .A2(_03160_),
    .B1(_03161_),
    .C1(_02694_),
    .X(_03162_));
 sky130_fd_sc_hd__or3b_2 _08456_ (.A(_02946_),
    .B(_03158_),
    .C_N(_03162_),
    .X(_03163_));
 sky130_fd_sc_hd__a21bo_1 _08457_ (.A1(_02648_),
    .A2(_03162_),
    .B1_N(_03158_),
    .X(_03164_));
 sky130_fd_sc_hd__a21oi_1 _08458_ (.A1(_02734_),
    .A2(_02736_),
    .B1(\genblk2[6].wave_shpr.div.fin_quo[3] ),
    .Y(_03165_));
 sky130_fd_sc_hd__a31o_1 _08459_ (.A1(\genblk2[6].wave_shpr.div.fin_quo[3] ),
    .A2(_02734_),
    .A3(_02736_),
    .B1(_02261_),
    .X(_03166_));
 sky130_fd_sc_hd__nor2_1 _08460_ (.A(_03165_),
    .B(_03166_),
    .Y(_03167_));
 sky130_fd_sc_hd__and3_1 _08461_ (.A(_02217_),
    .B(_02553_),
    .C(\genblk2[6].wave_shpr.div.fin_quo[4] ),
    .X(_03168_));
 sky130_fd_sc_hd__o31a_1 _08462_ (.A1(_02742_),
    .A2(_03167_),
    .A3(_03168_),
    .B1(_02745_),
    .X(_03169_));
 sky130_fd_sc_hd__nand3_2 _08463_ (.A(_03163_),
    .B(_03164_),
    .C(_03169_),
    .Y(_03170_));
 sky130_fd_sc_hd__a21o_1 _08464_ (.A1(_03163_),
    .A2(_03164_),
    .B1(_03169_),
    .X(_03171_));
 sky130_fd_sc_hd__xnor2_2 _08465_ (.A(_03153_),
    .B(_03152_),
    .Y(_03172_));
 sky130_fd_sc_hd__nand3_4 _08466_ (.A(_03170_),
    .B(_03171_),
    .C(_03172_),
    .Y(_03173_));
 sky130_fd_sc_hd__a21oi_2 _08467_ (.A1(_03048_),
    .A2(_03049_),
    .B1(_03050_),
    .Y(_03174_));
 sky130_fd_sc_hd__a211oi_4 _08468_ (.A1(_03154_),
    .A2(_03173_),
    .B1(_03051_),
    .C1(_03174_),
    .Y(_03175_));
 sky130_fd_sc_hd__inv_2 _08469_ (.A(\genblk2[5].wave_shpr.div.fin_quo[2] ),
    .Y(_03176_));
 sky130_fd_sc_hd__nor2_1 _08470_ (.A(\genblk2[5].wave_shpr.div.fin_quo[0] ),
    .B(\genblk2[5].wave_shpr.div.fin_quo[1] ),
    .Y(_03177_));
 sky130_fd_sc_hd__a21oi_1 _08471_ (.A1(_03176_),
    .A2(_03177_),
    .B1(_02789_),
    .Y(_03178_));
 sky130_fd_sc_hd__o21ai_1 _08472_ (.A1(\genblk2[5].wave_shpr.div.fin_quo[3] ),
    .A2(_03178_),
    .B1(_02526_),
    .Y(_03179_));
 sky130_fd_sc_hd__a21oi_1 _08473_ (.A1(\genblk2[5].wave_shpr.div.fin_quo[3] ),
    .A2(_03178_),
    .B1(_03179_),
    .Y(_03180_));
 sky130_fd_sc_hd__a21o_1 _08474_ (.A1(\genblk2[5].wave_shpr.div.fin_quo[4] ),
    .A2(_02308_),
    .B1(_02791_),
    .X(_03181_));
 sky130_fd_sc_hd__o21a_1 _08475_ (.A1(_03180_),
    .A2(_03181_),
    .B1(_02797_),
    .X(_03182_));
 sky130_fd_sc_hd__a21oi_1 _08476_ (.A1(_02932_),
    .A2(_02840_),
    .B1(\genblk2[4].wave_shpr.div.fin_quo[3] ),
    .Y(_03183_));
 sky130_fd_sc_hd__a31o_1 _08477_ (.A1(\genblk2[4].wave_shpr.div.fin_quo[3] ),
    .A2(_02932_),
    .A3(_02840_),
    .B1(_02222_),
    .X(_03184_));
 sky130_fd_sc_hd__a2bb2o_1 _08478_ (.A1_N(_03183_),
    .A2_N(_03184_),
    .B1(\genblk2[4].wave_shpr.div.fin_quo[4] ),
    .B2(_02308_),
    .X(_03185_));
 sky130_fd_sc_hd__o21a_1 _08479_ (.A1(_02838_),
    .A2(_03185_),
    .B1(_02846_),
    .X(_03186_));
 sky130_fd_sc_hd__xor2_1 _08480_ (.A(_03182_),
    .B(_03186_),
    .X(_03187_));
 sky130_fd_sc_hd__inv_2 _08481_ (.A(\genblk2[3].wave_shpr.div.fin_quo[0] ),
    .Y(_03188_));
 sky130_fd_sc_hd__inv_2 _08482_ (.A(\genblk2[3].wave_shpr.div.fin_quo[1] ),
    .Y(_03189_));
 sky130_fd_sc_hd__inv_2 _08483_ (.A(\genblk2[3].wave_shpr.div.fin_quo[2] ),
    .Y(_03190_));
 sky130_fd_sc_hd__a31o_1 _08484_ (.A1(_03188_),
    .A2(_03189_),
    .A3(_03190_),
    .B1(_02885_),
    .X(_03191_));
 sky130_fd_sc_hd__xnor2_1 _08485_ (.A(\genblk2[3].wave_shpr.div.fin_quo[3] ),
    .B(_03191_),
    .Y(_03192_));
 sky130_fd_sc_hd__a22o_1 _08486_ (.A1(\genblk2[3].wave_shpr.div.fin_quo[4] ),
    .A2(_02467_),
    .B1(_03192_),
    .B2(_02592_),
    .X(_03193_));
 sky130_fd_sc_hd__o21a_1 _08487_ (.A1(_02939_),
    .A2(_03193_),
    .B1(_02943_),
    .X(_03194_));
 sky130_fd_sc_hd__nand2_1 _08488_ (.A(_03187_),
    .B(_03194_),
    .Y(_03195_));
 sky130_fd_sc_hd__a21bo_1 _08489_ (.A1(_03182_),
    .A2(_03186_),
    .B1_N(_03195_),
    .X(_03196_));
 sky130_fd_sc_hd__a21bo_1 _08490_ (.A1(_03164_),
    .A2(_03169_),
    .B1_N(_03163_),
    .X(_03197_));
 sky130_fd_sc_hd__xnor2_1 _08491_ (.A(_03066_),
    .B(_03070_),
    .Y(_03198_));
 sky130_fd_sc_hd__xnor2_1 _08492_ (.A(_03197_),
    .B(_03198_),
    .Y(_03199_));
 sky130_fd_sc_hd__xnor2_1 _08493_ (.A(_03196_),
    .B(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__o211a_1 _08494_ (.A1(_03051_),
    .A2(_03174_),
    .B1(_03154_),
    .C1(_03173_),
    .X(_03201_));
 sky130_fd_sc_hd__nor3_2 _08495_ (.A(_03175_),
    .B(_03200_),
    .C(_03201_),
    .Y(_03202_));
 sky130_fd_sc_hd__o21ai_1 _08496_ (.A1(_03054_),
    .A2(_03076_),
    .B1(_03075_),
    .Y(_03203_));
 sky130_fd_sc_hd__o211a_1 _08497_ (.A1(_03175_),
    .A2(_03202_),
    .B1(_03077_),
    .C1(_03203_),
    .X(_03204_));
 sky130_fd_sc_hd__a211oi_1 _08498_ (.A1(_03077_),
    .A2(_03203_),
    .B1(_03175_),
    .C1(_03202_),
    .Y(_03205_));
 sky130_fd_sc_hd__a21o_1 _08499_ (.A1(_02547_),
    .A2(_02586_),
    .B1(_02588_),
    .X(_03206_));
 sky130_fd_sc_hd__o21ai_1 _08500_ (.A1(_02520_),
    .A2(_02587_),
    .B1(_03206_),
    .Y(_03207_));
 sky130_fd_sc_hd__or2b_1 _08501_ (.A(net24),
    .B_N(_03207_),
    .X(_03208_));
 sky130_fd_sc_hd__and2b_1 _08502_ (.A_N(_03198_),
    .B(_03197_),
    .X(_03209_));
 sky130_fd_sc_hd__a21oi_1 _08503_ (.A1(_03196_),
    .A2(_03199_),
    .B1(_03209_),
    .Y(_03210_));
 sky130_fd_sc_hd__a21oi_1 _08504_ (.A1(_03113_),
    .A2(_03118_),
    .B1(\genblk2[2].wave_shpr.div.fin_quo[5] ),
    .Y(_03211_));
 sky130_fd_sc_hd__a31o_1 _08505_ (.A1(\genblk2[2].wave_shpr.div.fin_quo[5] ),
    .A2(_03113_),
    .A3(_03118_),
    .B1(_02224_),
    .X(_03212_));
 sky130_fd_sc_hd__a2bb2o_1 _08506_ (.A1_N(_03211_),
    .A2_N(_03212_),
    .B1(\genblk2[2].wave_shpr.div.fin_quo[6] ),
    .B2(_02468_),
    .X(_03213_));
 sky130_fd_sc_hd__o21a_1 _08507_ (.A1(_03114_),
    .A2(_03213_),
    .B1(_03122_),
    .X(_03214_));
 sky130_fd_sc_hd__xnor2_1 _08508_ (.A(_03210_),
    .B(_03214_),
    .Y(_03215_));
 sky130_fd_sc_hd__xnor2_1 _08509_ (.A(_03208_),
    .B(_03215_),
    .Y(_03216_));
 sky130_fd_sc_hd__nor3b_2 _08510_ (.A(_03204_),
    .B(_03205_),
    .C_N(_03216_),
    .Y(_03217_));
 sky130_fd_sc_hd__o21ai_1 _08511_ (.A1(_03079_),
    .A2(_03126_),
    .B1(_03125_),
    .Y(_03218_));
 sky130_fd_sc_hd__o211a_1 _08512_ (.A1(_03204_),
    .A2(_03217_),
    .B1(_03127_),
    .C1(_03218_),
    .X(_03219_));
 sky130_fd_sc_hd__or2b_1 _08513_ (.A(_03210_),
    .B_N(_03214_),
    .X(_03220_));
 sky130_fd_sc_hd__or2b_1 _08514_ (.A(_03208_),
    .B_N(_03215_),
    .X(_03221_));
 sky130_fd_sc_hd__a211oi_2 _08515_ (.A1(_03127_),
    .A2(_03218_),
    .B1(_03204_),
    .C1(_03217_),
    .Y(_03222_));
 sky130_fd_sc_hd__a211oi_2 _08516_ (.A1(_03220_),
    .A2(_03221_),
    .B1(_03219_),
    .C1(_03222_),
    .Y(_03223_));
 sky130_fd_sc_hd__nor2_1 _08517_ (.A(_03219_),
    .B(_03223_),
    .Y(_03224_));
 sky130_fd_sc_hd__nor2_1 _08518_ (.A(_03136_),
    .B(_03224_),
    .Y(_03225_));
 sky130_fd_sc_hd__and3_1 _08519_ (.A(_02216_),
    .B(_02552_),
    .C(\genblk2[11].wave_shpr.div.fin_quo[0] ),
    .X(_03226_));
 sky130_fd_sc_hd__o211ai_2 _08520_ (.A1(_03141_),
    .A2(_03226_),
    .B1(net3),
    .C1(_02364_),
    .Y(_03227_));
 sky130_fd_sc_hd__and3_1 _08521_ (.A(_02216_),
    .B(_02552_),
    .C(\genblk2[10].wave_shpr.div.fin_quo[0] ),
    .X(_03228_));
 sky130_fd_sc_hd__o211a_1 _08522_ (.A1(_02416_),
    .A2(_03228_),
    .B1(net2),
    .C1(_02364_),
    .X(_03229_));
 sky130_fd_sc_hd__and2b_1 _08523_ (.A_N(_03227_),
    .B(_03229_),
    .X(_03230_));
 sky130_fd_sc_hd__and3_1 _08524_ (.A(_02216_),
    .B(_02552_),
    .C(\genblk2[9].wave_shpr.div.fin_quo[0] ),
    .X(_03231_));
 sky130_fd_sc_hd__o21a_1 _08525_ (.A1(_02310_),
    .A2(_03231_),
    .B1(_02314_),
    .X(_03232_));
 sky130_fd_sc_hd__xnor2_1 _08526_ (.A(_03227_),
    .B(_03229_),
    .Y(_03233_));
 sky130_fd_sc_hd__and2_1 _08527_ (.A(_03232_),
    .B(_03233_),
    .X(_03234_));
 sky130_fd_sc_hd__nor2_1 _08528_ (.A(_03230_),
    .B(_03234_),
    .Y(_03235_));
 sky130_fd_sc_hd__a22o_1 _08529_ (.A1(\genblk2[11].wave_shpr.div.fin_quo[0] ),
    .A2(_02524_),
    .B1(_02307_),
    .B2(\genblk2[11].wave_shpr.div.fin_quo[1] ),
    .X(_03236_));
 sky130_fd_sc_hd__o211a_1 _08530_ (.A1(_03141_),
    .A2(_03236_),
    .B1(net3),
    .C1(net163),
    .X(_03237_));
 sky130_fd_sc_hd__a22o_1 _08531_ (.A1(\genblk2[10].wave_shpr.div.fin_quo[0] ),
    .A2(_02525_),
    .B1(_02307_),
    .B2(\genblk2[10].wave_shpr.div.fin_quo[1] ),
    .X(_03238_));
 sky130_fd_sc_hd__o211a_1 _08532_ (.A1(_02416_),
    .A2(_03238_),
    .B1(net2),
    .C1(_02364_),
    .X(_03239_));
 sky130_fd_sc_hd__xnor2_1 _08533_ (.A(_03237_),
    .B(_03239_),
    .Y(_03240_));
 sky130_fd_sc_hd__a221o_1 _08534_ (.A1(\genblk2[9].wave_shpr.div.fin_quo[0] ),
    .A2(_02526_),
    .B1(_02308_),
    .B2(\genblk2[9].wave_shpr.div.fin_quo[1] ),
    .C1(_02310_),
    .X(_03241_));
 sky130_fd_sc_hd__nand2_1 _08535_ (.A(_02314_),
    .B(_03241_),
    .Y(_03242_));
 sky130_fd_sc_hd__or2_1 _08536_ (.A(_03240_),
    .B(_03242_),
    .X(_03243_));
 sky130_fd_sc_hd__nand2_1 _08537_ (.A(_03240_),
    .B(_03242_),
    .Y(_03244_));
 sky130_fd_sc_hd__and2_1 _08538_ (.A(_03243_),
    .B(_03244_),
    .X(_03245_));
 sky130_fd_sc_hd__or2b_1 _08539_ (.A(_03235_),
    .B_N(_03245_),
    .X(_03246_));
 sky130_fd_sc_hd__inv_2 _08540_ (.A(_02647_),
    .Y(_03247_));
 sky130_fd_sc_hd__a221o_1 _08541_ (.A1(\genblk2[8].wave_shpr.div.fin_quo[0] ),
    .A2(_02526_),
    .B1(_02308_),
    .B2(\genblk2[8].wave_shpr.div.fin_quo[1] ),
    .C1(_02636_),
    .X(_03248_));
 sky130_fd_sc_hd__a22o_1 _08542_ (.A1(\genblk2[7].wave_shpr.div.fin_quo[0] ),
    .A2(_02526_),
    .B1(_02308_),
    .B2(\genblk2[7].wave_shpr.div.fin_quo[1] ),
    .X(_03249_));
 sky130_fd_sc_hd__a21o_1 _08543_ (.A1(_02225_),
    .A2(_02682_),
    .B1(_03249_),
    .X(_03250_));
 sky130_fd_sc_hd__and4_1 _08544_ (.A(_02603_),
    .B(_03247_),
    .C(_03248_),
    .D(_03250_),
    .X(_03251_));
 sky130_fd_sc_hd__a22o_1 _08545_ (.A1(_02604_),
    .A2(_03248_),
    .B1(_03250_),
    .B2(_03247_),
    .X(_03252_));
 sky130_fd_sc_hd__and2b_1 _08546_ (.A_N(_03251_),
    .B(_03252_),
    .X(_03253_));
 sky130_fd_sc_hd__a22o_1 _08547_ (.A1(\genblk2[6].wave_shpr.div.fin_quo[0] ),
    .A2(_02527_),
    .B1(_02309_),
    .B2(\genblk2[6].wave_shpr.div.fin_quo[1] ),
    .X(_03254_));
 sky130_fd_sc_hd__o21a_1 _08548_ (.A1(_02742_),
    .A2(_03254_),
    .B1(_02745_),
    .X(_03255_));
 sky130_fd_sc_hd__xnor2_1 _08549_ (.A(_03253_),
    .B(_03255_),
    .Y(_03256_));
 sky130_fd_sc_hd__xor2_1 _08550_ (.A(_03245_),
    .B(_03235_),
    .X(_03257_));
 sky130_fd_sc_hd__or2_2 _08551_ (.A(_03256_),
    .B(_03257_),
    .X(_03258_));
 sky130_fd_sc_hd__a21oi_1 _08552_ (.A1(\genblk2[6].wave_shpr.div.fin_quo[0] ),
    .A2(_02734_),
    .B1(\genblk2[6].wave_shpr.div.fin_quo[1] ),
    .Y(_03259_));
 sky130_fd_sc_hd__a31o_1 _08553_ (.A1(\genblk2[6].wave_shpr.div.fin_quo[0] ),
    .A2(\genblk2[6].wave_shpr.div.fin_quo[1] ),
    .A3(_02734_),
    .B1(_02261_),
    .X(_03260_));
 sky130_fd_sc_hd__nor2_1 _08554_ (.A(_03259_),
    .B(_03260_),
    .Y(_03261_));
 sky130_fd_sc_hd__and3_1 _08555_ (.A(_02217_),
    .B(_02553_),
    .C(\genblk2[6].wave_shpr.div.fin_quo[2] ),
    .X(_03262_));
 sky130_fd_sc_hd__o31a_1 _08556_ (.A1(_02742_),
    .A2(_03261_),
    .A3(_03262_),
    .B1(_02745_),
    .X(_03263_));
 sky130_fd_sc_hd__a21oi_1 _08557_ (.A1(\genblk2[8].wave_shpr.div.fin_quo[0] ),
    .A2(_02638_),
    .B1(\genblk2[8].wave_shpr.div.fin_quo[1] ),
    .Y(_03264_));
 sky130_fd_sc_hd__a31o_1 _08558_ (.A1(\genblk2[8].wave_shpr.div.fin_quo[0] ),
    .A2(\genblk2[8].wave_shpr.div.fin_quo[1] ),
    .A3(_02638_),
    .B1(_02223_),
    .X(_03265_));
 sky130_fd_sc_hd__nor2_1 _08559_ (.A(_03264_),
    .B(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__a21o_1 _08560_ (.A1(\genblk2[8].wave_shpr.div.fin_quo[2] ),
    .A2(_02362_),
    .B1(_02636_),
    .X(_03267_));
 sky130_fd_sc_hd__o21ai_1 _08561_ (.A1(_03266_),
    .A2(_03267_),
    .B1(_02604_),
    .Y(_03268_));
 sky130_fd_sc_hd__o211a_1 _08562_ (.A1(_02676_),
    .A2(_02679_),
    .B1(_02680_),
    .C1(\genblk2[7].wave_shpr.div.fin_quo[0] ),
    .X(_03269_));
 sky130_fd_sc_hd__xnor2_1 _08563_ (.A(\genblk2[7].wave_shpr.div.fin_quo[1] ),
    .B(_03269_),
    .Y(_03270_));
 sky130_fd_sc_hd__nand2_1 _08564_ (.A(\genblk2[7].wave_shpr.div.fin_quo[2] ),
    .B(_02521_),
    .Y(_03271_));
 sky130_fd_sc_hd__o211a_1 _08565_ (.A1(_02261_),
    .A2(_03270_),
    .B1(_03271_),
    .C1(_02950_),
    .X(_03272_));
 sky130_fd_sc_hd__or3_1 _08566_ (.A(_02946_),
    .B(_03268_),
    .C(_03272_),
    .X(_03273_));
 sky130_fd_sc_hd__o21ai_1 _08567_ (.A1(_02946_),
    .A2(_03272_),
    .B1(_03268_),
    .Y(_03274_));
 sky130_fd_sc_hd__nand3_1 _08568_ (.A(_03263_),
    .B(_03273_),
    .C(_03274_),
    .Y(_03275_));
 sky130_fd_sc_hd__a21o_1 _08569_ (.A1(_03273_),
    .A2(_03274_),
    .B1(_03263_),
    .X(_03276_));
 sky130_fd_sc_hd__a21oi_1 _08570_ (.A1(\genblk2[9].wave_shpr.div.fin_quo[0] ),
    .A2(_02303_),
    .B1(\genblk2[9].wave_shpr.div.fin_quo[1] ),
    .Y(_03277_));
 sky130_fd_sc_hd__a31o_1 _08571_ (.A1(\genblk2[9].wave_shpr.div.fin_quo[0] ),
    .A2(\genblk2[9].wave_shpr.div.fin_quo[1] ),
    .A3(_02303_),
    .B1(_02316_),
    .X(_03278_));
 sky130_fd_sc_hd__a2bb2o_1 _08572_ (.A1_N(_03277_),
    .A2_N(_03278_),
    .B1(\genblk2[9].wave_shpr.div.fin_quo[2] ),
    .B2(_02362_),
    .X(_03279_));
 sky130_fd_sc_hd__o21a_1 _08573_ (.A1(_02310_),
    .A2(_03279_),
    .B1(_02314_),
    .X(_03280_));
 sky130_fd_sc_hd__a31o_1 _08574_ (.A1(\genblk2[11].wave_shpr.div.fin_quo[0] ),
    .A2(net33),
    .A3(_02350_),
    .B1(\genblk2[11].wave_shpr.div.fin_quo[1] ),
    .X(_03281_));
 sky130_fd_sc_hd__nand4_1 _08575_ (.A(\genblk2[11].wave_shpr.div.fin_quo[0] ),
    .B(\genblk2[11].wave_shpr.div.fin_quo[1] ),
    .C(_02349_),
    .D(_02351_),
    .Y(_03282_));
 sky130_fd_sc_hd__a32o_1 _08576_ (.A1(_02525_),
    .A2(_03281_),
    .A3(_03282_),
    .B1(_02361_),
    .B2(\genblk2[11].wave_shpr.div.fin_quo[2] ),
    .X(_03283_));
 sky130_fd_sc_hd__o21a_1 _08577_ (.A1(_03141_),
    .A2(_03283_),
    .B1(_02901_),
    .X(_03284_));
 sky130_fd_sc_hd__inv_2 _08578_ (.A(\genblk2[10].wave_shpr.div.fin_quo[0] ),
    .Y(_03285_));
 sky130_fd_sc_hd__nor2_1 _08579_ (.A(_03285_),
    .B(_02404_),
    .Y(_03286_));
 sky130_fd_sc_hd__inv_2 _08580_ (.A(\genblk2[10].wave_shpr.div.fin_quo[1] ),
    .Y(_03287_));
 sky130_fd_sc_hd__o31a_1 _08581_ (.A1(_03285_),
    .A2(_03287_),
    .A3(_02404_),
    .B1(_02525_),
    .X(_03288_));
 sky130_fd_sc_hd__o21a_1 _08582_ (.A1(\genblk2[10].wave_shpr.div.fin_quo[1] ),
    .A2(_03286_),
    .B1(_03288_),
    .X(_03289_));
 sky130_fd_sc_hd__a21o_1 _08583_ (.A1(\genblk2[10].wave_shpr.div.fin_quo[2] ),
    .A2(_02308_),
    .B1(_02416_),
    .X(_03290_));
 sky130_fd_sc_hd__o21ai_1 _08584_ (.A1(_03289_),
    .A2(_03290_),
    .B1(_02419_),
    .Y(_03291_));
 sky130_fd_sc_hd__xnor2_2 _08585_ (.A(_03284_),
    .B(_03291_),
    .Y(_03292_));
 sky130_fd_sc_hd__xnor2_2 _08586_ (.A(_03280_),
    .B(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hd__a21bo_1 _08587_ (.A1(_03237_),
    .A2(_03239_),
    .B1_N(_03243_),
    .X(_03294_));
 sky130_fd_sc_hd__xnor2_2 _08588_ (.A(_03293_),
    .B(_03294_),
    .Y(_03295_));
 sky130_fd_sc_hd__and3_1 _08589_ (.A(_03275_),
    .B(_03276_),
    .C(_03295_),
    .X(_03296_));
 sky130_fd_sc_hd__a21oi_1 _08590_ (.A1(_03275_),
    .A2(_03276_),
    .B1(_03295_),
    .Y(_03297_));
 sky130_fd_sc_hd__a211o_2 _08591_ (.A1(_03246_),
    .A2(_03258_),
    .B1(_03296_),
    .C1(_03297_),
    .X(_03298_));
 sky130_fd_sc_hd__a221o_1 _08592_ (.A1(\genblk2[5].wave_shpr.div.fin_quo[0] ),
    .A2(_02527_),
    .B1(_02521_),
    .B2(\genblk2[5].wave_shpr.div.fin_quo[1] ),
    .C1(_02791_),
    .X(_03299_));
 sky130_fd_sc_hd__a221o_1 _08593_ (.A1(\genblk2[4].wave_shpr.div.fin_quo[0] ),
    .A2(_02526_),
    .B1(_02361_),
    .B2(\genblk2[4].wave_shpr.div.fin_quo[1] ),
    .C1(_02838_),
    .X(_03300_));
 sky130_fd_sc_hd__and3_1 _08594_ (.A(net10),
    .B(_02364_),
    .C(_03300_),
    .X(_03301_));
 sky130_fd_sc_hd__and3_1 _08595_ (.A(_02798_),
    .B(_03299_),
    .C(_03301_),
    .X(_03302_));
 sky130_fd_sc_hd__a21oi_1 _08596_ (.A1(_02798_),
    .A2(_03299_),
    .B1(_03301_),
    .Y(_03303_));
 sky130_fd_sc_hd__nor2_1 _08597_ (.A(_03302_),
    .B(_03303_),
    .Y(_03304_));
 sky130_fd_sc_hd__a221o_1 _08598_ (.A1(\genblk2[3].wave_shpr.div.fin_quo[0] ),
    .A2(_02592_),
    .B1(_02467_),
    .B2(\genblk2[3].wave_shpr.div.fin_quo[1] ),
    .C1(_02939_),
    .X(_03305_));
 sky130_fd_sc_hd__and3_1 _08599_ (.A(net9),
    .B(_02744_),
    .C(_03305_),
    .X(_03306_));
 sky130_fd_sc_hd__a21o_1 _08600_ (.A1(_03304_),
    .A2(_03306_),
    .B1(_03302_),
    .X(_03307_));
 sky130_fd_sc_hd__and3b_1 _08601_ (.A_N(_03251_),
    .B(_03252_),
    .C(_03255_),
    .X(_03308_));
 sky130_fd_sc_hd__nor3_1 _08602_ (.A(_03188_),
    .B(_03189_),
    .C(_02885_),
    .Y(_03309_));
 sky130_fd_sc_hd__o21ai_1 _08603_ (.A1(_03188_),
    .A2(_02885_),
    .B1(_03189_),
    .Y(_03310_));
 sky130_fd_sc_hd__or3b_1 _08604_ (.A(_02261_),
    .B(_03309_),
    .C_N(_03310_),
    .X(_03311_));
 sky130_fd_sc_hd__nand2_1 _08605_ (.A(\genblk2[3].wave_shpr.div.fin_quo[2] ),
    .B(_02467_),
    .Y(_03312_));
 sky130_fd_sc_hd__a31o_1 _08606_ (.A1(_02891_),
    .A2(_03311_),
    .A3(_03312_),
    .B1(_02893_),
    .X(_03313_));
 sky130_fd_sc_hd__inv_2 _08607_ (.A(\genblk2[5].wave_shpr.div.fin_quo[0] ),
    .Y(_03314_));
 sky130_fd_sc_hd__inv_2 _08608_ (.A(\genblk2[5].wave_shpr.div.fin_quo[1] ),
    .Y(_03315_));
 sky130_fd_sc_hd__o21a_1 _08609_ (.A1(_03314_),
    .A2(_02789_),
    .B1(_03315_),
    .X(_03316_));
 sky130_fd_sc_hd__or3_1 _08610_ (.A(_03314_),
    .B(_03315_),
    .C(_02789_),
    .X(_03317_));
 sky130_fd_sc_hd__or3b_1 _08611_ (.A(_03316_),
    .B(_02223_),
    .C_N(_03317_),
    .X(_03318_));
 sky130_fd_sc_hd__a21oi_1 _08612_ (.A1(\genblk2[5].wave_shpr.div.fin_quo[2] ),
    .A2(_02521_),
    .B1(_02791_),
    .Y(_03319_));
 sky130_fd_sc_hd__a21bo_1 _08613_ (.A1(_03318_),
    .A2(_03319_),
    .B1_N(_02797_),
    .X(_03320_));
 sky130_fd_sc_hd__a21oi_1 _08614_ (.A1(\genblk2[4].wave_shpr.div.fin_quo[0] ),
    .A2(_02932_),
    .B1(\genblk2[4].wave_shpr.div.fin_quo[1] ),
    .Y(_03321_));
 sky130_fd_sc_hd__a31o_1 _08615_ (.A1(\genblk2[4].wave_shpr.div.fin_quo[0] ),
    .A2(\genblk2[4].wave_shpr.div.fin_quo[1] ),
    .A3(_02932_),
    .B1(_02223_),
    .X(_03322_));
 sky130_fd_sc_hd__nor2_1 _08616_ (.A(_03321_),
    .B(_03322_),
    .Y(_03323_));
 sky130_fd_sc_hd__a21o_1 _08617_ (.A1(\genblk2[4].wave_shpr.div.fin_quo[2] ),
    .A2(_02362_),
    .B1(_02838_),
    .X(_03324_));
 sky130_fd_sc_hd__o21ai_2 _08618_ (.A1(_03323_),
    .A2(_03324_),
    .B1(_02846_),
    .Y(_03325_));
 sky130_fd_sc_hd__xor2_1 _08619_ (.A(_03320_),
    .B(_03325_),
    .X(_03326_));
 sky130_fd_sc_hd__xnor2_1 _08620_ (.A(_03313_),
    .B(_03326_),
    .Y(_03327_));
 sky130_fd_sc_hd__o21a_1 _08621_ (.A1(_03251_),
    .A2(_03308_),
    .B1(_03327_),
    .X(_03328_));
 sky130_fd_sc_hd__nor3_1 _08622_ (.A(_03251_),
    .B(_03308_),
    .C(_03327_),
    .Y(_03329_));
 sky130_fd_sc_hd__nor2_1 _08623_ (.A(_03328_),
    .B(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__xnor2_1 _08624_ (.A(_03307_),
    .B(_03330_),
    .Y(_03331_));
 sky130_fd_sc_hd__o211ai_2 _08625_ (.A1(_03296_),
    .A2(_03297_),
    .B1(_03246_),
    .C1(_03258_),
    .Y(_03332_));
 sky130_fd_sc_hd__nand3b_2 _08626_ (.A_N(_03331_),
    .B(_03332_),
    .C(_03298_),
    .Y(_03333_));
 sky130_fd_sc_hd__or2b_1 _08627_ (.A(_03293_),
    .B_N(_03294_),
    .X(_03334_));
 sky130_fd_sc_hd__nand3_2 _08628_ (.A(_03275_),
    .B(_03276_),
    .C(_03295_),
    .Y(_03335_));
 sky130_fd_sc_hd__a21oi_1 _08629_ (.A1(_02734_),
    .A2(_02735_),
    .B1(\genblk2[6].wave_shpr.div.fin_quo[2] ),
    .Y(_03336_));
 sky130_fd_sc_hd__a31o_1 _08630_ (.A1(\genblk2[6].wave_shpr.div.fin_quo[2] ),
    .A2(_02733_),
    .A3(_02735_),
    .B1(_02261_),
    .X(_03337_));
 sky130_fd_sc_hd__nor2_1 _08631_ (.A(_03336_),
    .B(_03337_),
    .Y(_03338_));
 sky130_fd_sc_hd__and3_1 _08632_ (.A(_02217_),
    .B(_02553_),
    .C(\genblk2[6].wave_shpr.div.fin_quo[3] ),
    .X(_03339_));
 sky130_fd_sc_hd__o31a_1 _08633_ (.A1(_02742_),
    .A2(_03338_),
    .A3(_03339_),
    .B1(_02745_),
    .X(_03340_));
 sky130_fd_sc_hd__o21ai_1 _08634_ (.A1(\genblk2[8].wave_shpr.div.fin_quo[0] ),
    .A2(\genblk2[8].wave_shpr.div.fin_quo[1] ),
    .B1(_02638_),
    .Y(_03341_));
 sky130_fd_sc_hd__xnor2_1 _08635_ (.A(\genblk2[8].wave_shpr.div.fin_quo[2] ),
    .B(_03341_),
    .Y(_03342_));
 sky130_fd_sc_hd__and3_1 _08636_ (.A(_02216_),
    .B(_02552_),
    .C(\genblk2[8].wave_shpr.div.fin_quo[3] ),
    .X(_03343_));
 sky130_fd_sc_hd__a211o_1 _08637_ (.A1(_02592_),
    .A2(_03342_),
    .B1(_03343_),
    .C1(_02636_),
    .X(_03344_));
 sky130_fd_sc_hd__o21ai_1 _08638_ (.A1(_02682_),
    .A2(_02686_),
    .B1(_02685_),
    .Y(_03345_));
 sky130_fd_sc_hd__o31a_1 _08639_ (.A1(_02685_),
    .A2(_02681_),
    .A3(_02686_),
    .B1(_02526_),
    .X(_03346_));
 sky130_fd_sc_hd__and3_1 _08640_ (.A(_02216_),
    .B(_02553_),
    .C(\genblk2[7].wave_shpr.div.fin_quo[3] ),
    .X(_03347_));
 sky130_fd_sc_hd__a211o_1 _08641_ (.A1(_03345_),
    .A2(_03346_),
    .B1(_03347_),
    .C1(_02694_),
    .X(_03348_));
 sky130_fd_sc_hd__nand4_1 _08642_ (.A(_02604_),
    .B(_02648_),
    .C(_03344_),
    .D(_03348_),
    .Y(_03349_));
 sky130_fd_sc_hd__a22o_1 _08643_ (.A1(_02604_),
    .A2(_03344_),
    .B1(_03348_),
    .B2(_02648_),
    .X(_03350_));
 sky130_fd_sc_hd__nand3_1 _08644_ (.A(_03340_),
    .B(_03349_),
    .C(_03350_),
    .Y(_03351_));
 sky130_fd_sc_hd__a21o_1 _08645_ (.A1(_03349_),
    .A2(_03350_),
    .B1(_03340_),
    .X(_03352_));
 sky130_fd_sc_hd__xor2_1 _08646_ (.A(_03140_),
    .B(_03150_),
    .X(_03353_));
 sky130_fd_sc_hd__o211a_1 _08647_ (.A1(_03289_),
    .A2(_03290_),
    .B1(_02419_),
    .C1(_03284_),
    .X(_03354_));
 sky130_fd_sc_hd__a21oi_1 _08648_ (.A1(_03280_),
    .A2(_03292_),
    .B1(_03354_),
    .Y(_03355_));
 sky130_fd_sc_hd__xnor2_1 _08649_ (.A(_03353_),
    .B(_03355_),
    .Y(_03356_));
 sky130_fd_sc_hd__and3_2 _08650_ (.A(_03351_),
    .B(_03352_),
    .C(_03356_),
    .X(_03357_));
 sky130_fd_sc_hd__a21oi_2 _08651_ (.A1(_03351_),
    .A2(_03352_),
    .B1(_03356_),
    .Y(_03358_));
 sky130_fd_sc_hd__a211oi_4 _08652_ (.A1(_03334_),
    .A2(_03335_),
    .B1(_03357_),
    .C1(_03358_),
    .Y(_03359_));
 sky130_fd_sc_hd__and2b_1 _08653_ (.A_N(_03313_),
    .B(_03326_),
    .X(_03360_));
 sky130_fd_sc_hd__o21bai_2 _08654_ (.A1(_03320_),
    .A2(_03325_),
    .B1_N(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__a21boi_1 _08655_ (.A1(_03263_),
    .A2(_03274_),
    .B1_N(_03273_),
    .Y(_03362_));
 sky130_fd_sc_hd__a21o_1 _08656_ (.A1(_03188_),
    .A2(_03189_),
    .B1(_02885_),
    .X(_03363_));
 sky130_fd_sc_hd__xnor2_1 _08657_ (.A(\genblk2[3].wave_shpr.div.fin_quo[2] ),
    .B(_03363_),
    .Y(_03364_));
 sky130_fd_sc_hd__a22o_1 _08658_ (.A1(\genblk2[3].wave_shpr.div.fin_quo[3] ),
    .A2(_02467_),
    .B1(_03364_),
    .B2(_02592_),
    .X(_03365_));
 sky130_fd_sc_hd__o21ai_1 _08659_ (.A1(_02939_),
    .A2(_03365_),
    .B1(_02943_),
    .Y(_03366_));
 sky130_fd_sc_hd__nor2_1 _08660_ (.A(_02789_),
    .B(_03177_),
    .Y(_03367_));
 sky130_fd_sc_hd__o31a_1 _08661_ (.A1(_03176_),
    .A2(_02789_),
    .A3(_03177_),
    .B1(_02525_),
    .X(_03368_));
 sky130_fd_sc_hd__o21a_1 _08662_ (.A1(\genblk2[5].wave_shpr.div.fin_quo[2] ),
    .A2(_03367_),
    .B1(_03368_),
    .X(_03369_));
 sky130_fd_sc_hd__a211o_1 _08663_ (.A1(\genblk2[5].wave_shpr.div.fin_quo[3] ),
    .A2(_02521_),
    .B1(_02791_),
    .C1(_03369_),
    .X(_03370_));
 sky130_fd_sc_hd__nand2_1 _08664_ (.A(_02798_),
    .B(_03370_),
    .Y(_03371_));
 sky130_fd_sc_hd__a21oi_1 _08665_ (.A1(_02932_),
    .A2(_02839_),
    .B1(\genblk2[4].wave_shpr.div.fin_quo[2] ),
    .Y(_03372_));
 sky130_fd_sc_hd__a31o_1 _08666_ (.A1(\genblk2[4].wave_shpr.div.fin_quo[2] ),
    .A2(_02932_),
    .A3(_02839_),
    .B1(_02316_),
    .X(_03373_));
 sky130_fd_sc_hd__a2bb2o_1 _08667_ (.A1_N(_03372_),
    .A2_N(_03373_),
    .B1(\genblk2[4].wave_shpr.div.fin_quo[3] ),
    .B2(_02362_),
    .X(_03374_));
 sky130_fd_sc_hd__o21a_1 _08668_ (.A1(_02838_),
    .A2(_03374_),
    .B1(_02846_),
    .X(_03375_));
 sky130_fd_sc_hd__xnor2_1 _08669_ (.A(_03371_),
    .B(_03375_),
    .Y(_03376_));
 sky130_fd_sc_hd__xnor2_1 _08670_ (.A(_03366_),
    .B(_03376_),
    .Y(_03377_));
 sky130_fd_sc_hd__xnor2_1 _08671_ (.A(_03362_),
    .B(_03377_),
    .Y(_03378_));
 sky130_fd_sc_hd__xnor2_1 _08672_ (.A(_03361_),
    .B(_03378_),
    .Y(_03379_));
 sky130_fd_sc_hd__o211a_1 _08673_ (.A1(_03357_),
    .A2(_03358_),
    .B1(_03334_),
    .C1(_03335_),
    .X(_03380_));
 sky130_fd_sc_hd__nor3_2 _08674_ (.A(_03359_),
    .B(_03379_),
    .C(_03380_),
    .Y(_03381_));
 sky130_fd_sc_hd__o21a_1 _08675_ (.A1(_03359_),
    .A2(_03380_),
    .B1(_03379_),
    .X(_03382_));
 sky130_fd_sc_hd__a211o_1 _08676_ (.A1(_03298_),
    .A2(_03333_),
    .B1(_03381_),
    .C1(_03382_),
    .X(_03383_));
 sky130_fd_sc_hd__a211oi_1 _08677_ (.A1(_03298_),
    .A2(_03333_),
    .B1(_03381_),
    .C1(_03382_),
    .Y(_03384_));
 sky130_fd_sc_hd__or2_1 _08678_ (.A(_02561_),
    .B(_02562_),
    .X(_03385_));
 sky130_fd_sc_hd__xnor2_2 _08679_ (.A(_02584_),
    .B(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__a21oi_1 _08680_ (.A1(_03307_),
    .A2(_03330_),
    .B1(_03328_),
    .Y(_03387_));
 sky130_fd_sc_hd__a21oi_1 _08681_ (.A1(_03113_),
    .A2(_03115_),
    .B1(\genblk2[2].wave_shpr.div.fin_quo[2] ),
    .Y(_03388_));
 sky130_fd_sc_hd__a31o_1 _08682_ (.A1(\genblk2[2].wave_shpr.div.fin_quo[2] ),
    .A2(_03113_),
    .A3(_03115_),
    .B1(_02224_),
    .X(_03389_));
 sky130_fd_sc_hd__a2bb2o_1 _08683_ (.A1_N(_03388_),
    .A2_N(_03389_),
    .B1(\genblk2[2].wave_shpr.div.fin_quo[3] ),
    .B2(_02468_),
    .X(_03390_));
 sky130_fd_sc_hd__o21a_1 _08684_ (.A1(_03114_),
    .A2(_03390_),
    .B1(_03122_),
    .X(_03391_));
 sky130_fd_sc_hd__xnor2_1 _08685_ (.A(_03387_),
    .B(_03391_),
    .Y(_03392_));
 sky130_fd_sc_hd__xnor2_1 _08686_ (.A(_03386_),
    .B(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__o211a_1 _08687_ (.A1(_03381_),
    .A2(_03382_),
    .B1(_03298_),
    .C1(_03333_),
    .X(_03394_));
 sky130_fd_sc_hd__or3_2 _08688_ (.A(_03384_),
    .B(_03393_),
    .C(_03394_),
    .X(_03395_));
 sky130_fd_sc_hd__and2b_1 _08689_ (.A_N(_03366_),
    .B(_03376_),
    .X(_03396_));
 sky130_fd_sc_hd__a31o_1 _08690_ (.A1(_02798_),
    .A2(_03370_),
    .A3(_03375_),
    .B1(_03396_),
    .X(_03397_));
 sky130_fd_sc_hd__a21bo_1 _08691_ (.A1(_03340_),
    .A2(_03350_),
    .B1_N(_03349_),
    .X(_03398_));
 sky130_fd_sc_hd__xnor2_1 _08692_ (.A(_03187_),
    .B(_03194_),
    .Y(_03399_));
 sky130_fd_sc_hd__xnor2_1 _08693_ (.A(_03398_),
    .B(_03399_),
    .Y(_03400_));
 sky130_fd_sc_hd__xnor2_1 _08694_ (.A(_03397_),
    .B(_03400_),
    .Y(_03401_));
 sky130_fd_sc_hd__a21o_1 _08695_ (.A1(_03170_),
    .A2(_03171_),
    .B1(_03172_),
    .X(_03402_));
 sky130_fd_sc_hd__and2b_1 _08696_ (.A_N(_03355_),
    .B(_03353_),
    .X(_03403_));
 sky130_fd_sc_hd__a211o_1 _08697_ (.A1(_03173_),
    .A2(_03402_),
    .B1(_03403_),
    .C1(_03357_),
    .X(_03404_));
 sky130_fd_sc_hd__o211ai_4 _08698_ (.A1(_03403_),
    .A2(_03357_),
    .B1(_03173_),
    .C1(_03402_),
    .Y(_03405_));
 sky130_fd_sc_hd__nand3b_2 _08699_ (.A_N(_03401_),
    .B(_03404_),
    .C(_03405_),
    .Y(_03406_));
 sky130_fd_sc_hd__a21bo_1 _08700_ (.A1(_03405_),
    .A2(_03404_),
    .B1_N(_03401_),
    .X(_03407_));
 sky130_fd_sc_hd__o211ai_2 _08701_ (.A1(_03359_),
    .A2(_03381_),
    .B1(_03406_),
    .C1(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__o21ai_1 _08702_ (.A1(_02561_),
    .A2(_02585_),
    .B1(_02548_),
    .Y(_03409_));
 sky130_fd_sc_hd__nand2_1 _08703_ (.A(_02586_),
    .B(_03409_),
    .Y(_03410_));
 sky130_fd_sc_hd__and2b_1 _08704_ (.A_N(_03362_),
    .B(_03377_),
    .X(_03411_));
 sky130_fd_sc_hd__a21o_1 _08705_ (.A1(_03361_),
    .A2(_03378_),
    .B1(_03411_),
    .X(_03412_));
 sky130_fd_sc_hd__a21oi_1 _08706_ (.A1(_03113_),
    .A2(_03116_),
    .B1(\genblk2[2].wave_shpr.div.fin_quo[3] ),
    .Y(_03413_));
 sky130_fd_sc_hd__a31o_1 _08707_ (.A1(\genblk2[2].wave_shpr.div.fin_quo[3] ),
    .A2(net25),
    .A3(_03116_),
    .B1(_02224_),
    .X(_03414_));
 sky130_fd_sc_hd__a2bb2o_1 _08708_ (.A1_N(_03413_),
    .A2_N(_03414_),
    .B1(\genblk2[2].wave_shpr.div.fin_quo[4] ),
    .B2(_02468_),
    .X(_03415_));
 sky130_fd_sc_hd__o21a_1 _08709_ (.A1(_03114_),
    .A2(_03415_),
    .B1(_03122_),
    .X(_03416_));
 sky130_fd_sc_hd__xnor2_1 _08710_ (.A(_03412_),
    .B(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__xor2_1 _08711_ (.A(_03410_),
    .B(_03417_),
    .X(_03418_));
 sky130_fd_sc_hd__a211o_1 _08712_ (.A1(_03406_),
    .A2(_03407_),
    .B1(_03359_),
    .C1(_03381_),
    .X(_03419_));
 sky130_fd_sc_hd__and3_2 _08713_ (.A(_03408_),
    .B(_03418_),
    .C(_03419_),
    .X(_03420_));
 sky130_fd_sc_hd__a21oi_2 _08714_ (.A1(_03408_),
    .A2(_03419_),
    .B1(_03418_),
    .Y(_03421_));
 sky130_fd_sc_hd__a211o_1 _08715_ (.A1(_03383_),
    .A2(_03395_),
    .B1(_03420_),
    .C1(_03421_),
    .X(_03422_));
 sky130_fd_sc_hd__or2b_1 _08716_ (.A(_03387_),
    .B_N(_03391_),
    .X(_03423_));
 sky130_fd_sc_hd__nand2_1 _08717_ (.A(_03386_),
    .B(_03392_),
    .Y(_03424_));
 sky130_fd_sc_hd__a211oi_2 _08718_ (.A1(_03383_),
    .A2(_03395_),
    .B1(_03420_),
    .C1(_03421_),
    .Y(_03425_));
 sky130_fd_sc_hd__o211a_1 _08719_ (.A1(_03420_),
    .A2(_03421_),
    .B1(_03383_),
    .C1(_03395_),
    .X(_03426_));
 sky130_fd_sc_hd__a211o_1 _08720_ (.A1(_03423_),
    .A2(_03424_),
    .B1(_03425_),
    .C1(_03426_),
    .X(_03427_));
 sky130_fd_sc_hd__inv_2 _08721_ (.A(_03408_),
    .Y(_03428_));
 sky130_fd_sc_hd__nor2_1 _08722_ (.A(_02588_),
    .B(_02546_),
    .Y(_03429_));
 sky130_fd_sc_hd__and2b_1 _08723_ (.A_N(_02536_),
    .B(_02586_),
    .X(_03430_));
 sky130_fd_sc_hd__xnor2_2 _08724_ (.A(_03429_),
    .B(_03430_),
    .Y(_03431_));
 sky130_fd_sc_hd__and2b_1 _08725_ (.A_N(_03399_),
    .B(_03398_),
    .X(_03432_));
 sky130_fd_sc_hd__a21oi_1 _08726_ (.A1(_03397_),
    .A2(_03400_),
    .B1(_03432_),
    .Y(_03433_));
 sky130_fd_sc_hd__a21oi_1 _08727_ (.A1(_03113_),
    .A2(_03117_),
    .B1(\genblk2[2].wave_shpr.div.fin_quo[4] ),
    .Y(_03434_));
 sky130_fd_sc_hd__a31o_1 _08728_ (.A1(\genblk2[2].wave_shpr.div.fin_quo[4] ),
    .A2(_03113_),
    .A3(_03117_),
    .B1(_02224_),
    .X(_03435_));
 sky130_fd_sc_hd__a2bb2o_1 _08729_ (.A1_N(_03434_),
    .A2_N(_03435_),
    .B1(\genblk2[2].wave_shpr.div.fin_quo[5] ),
    .B2(_02468_),
    .X(_03436_));
 sky130_fd_sc_hd__o21a_1 _08730_ (.A1(_03114_),
    .A2(_03436_),
    .B1(_03122_),
    .X(_03437_));
 sky130_fd_sc_hd__xnor2_1 _08731_ (.A(_03433_),
    .B(_03437_),
    .Y(_03438_));
 sky130_fd_sc_hd__xnor2_1 _08732_ (.A(_03431_),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__o21a_1 _08733_ (.A1(_03175_),
    .A2(_03201_),
    .B1(_03200_),
    .X(_03440_));
 sky130_fd_sc_hd__o211ai_2 _08734_ (.A1(_03202_),
    .A2(_03440_),
    .B1(_03405_),
    .C1(_03406_),
    .Y(_03441_));
 sky130_fd_sc_hd__a211o_1 _08735_ (.A1(_03405_),
    .A2(_03406_),
    .B1(_03202_),
    .C1(_03440_),
    .X(_03442_));
 sky130_fd_sc_hd__nand3b_2 _08736_ (.A_N(_03439_),
    .B(_03441_),
    .C(_03442_),
    .Y(_03443_));
 sky130_fd_sc_hd__a21bo_1 _08737_ (.A1(_03442_),
    .A2(_03441_),
    .B1_N(_03439_),
    .X(_03444_));
 sky130_fd_sc_hd__o211a_2 _08738_ (.A1(_03428_),
    .A2(_03420_),
    .B1(_03443_),
    .C1(_03444_),
    .X(_03445_));
 sky130_fd_sc_hd__a211oi_2 _08739_ (.A1(_03443_),
    .A2(_03444_),
    .B1(_03428_),
    .C1(_03420_),
    .Y(_03446_));
 sky130_fd_sc_hd__nand2_1 _08740_ (.A(_03412_),
    .B(_03416_),
    .Y(_03447_));
 sky130_fd_sc_hd__or2_2 _08741_ (.A(_03410_),
    .B(_03417_),
    .X(_03448_));
 sky130_fd_sc_hd__o211a_1 _08742_ (.A1(_03445_),
    .A2(_03446_),
    .B1(_03447_),
    .C1(_03448_),
    .X(_03449_));
 sky130_fd_sc_hd__a211oi_4 _08743_ (.A1(_03447_),
    .A2(_03448_),
    .B1(_03445_),
    .C1(_03446_),
    .Y(_03450_));
 sky130_fd_sc_hd__a211oi_2 _08744_ (.A1(_03422_),
    .A2(_03427_),
    .B1(_03449_),
    .C1(_03450_),
    .Y(_03451_));
 sky130_fd_sc_hd__nand2_1 _08745_ (.A(_03256_),
    .B(_03257_),
    .Y(_03452_));
 sky130_fd_sc_hd__and3_1 _08746_ (.A(_02217_),
    .B(_02553_),
    .C(\genblk2[6].wave_shpr.div.fin_quo[0] ),
    .X(_03453_));
 sky130_fd_sc_hd__o21ai_2 _08747_ (.A1(_02742_),
    .A2(_03453_),
    .B1(_02745_),
    .Y(_03454_));
 sky130_fd_sc_hd__nand3_1 _08748_ (.A(net14),
    .B(_02744_),
    .C(_02365_),
    .Y(_03455_));
 sky130_fd_sc_hd__a21oi_1 _08749_ (.A1(\genblk2[8].wave_shpr.div.fin_quo[0] ),
    .A2(_02309_),
    .B1(_02636_),
    .Y(_03456_));
 sky130_fd_sc_hd__or2_1 _08750_ (.A(_03455_),
    .B(_03456_),
    .X(_03457_));
 sky130_fd_sc_hd__nand2_1 _08751_ (.A(\genblk2[7].wave_shpr.div.fin_quo[0] ),
    .B(_02467_),
    .Y(_03458_));
 sky130_fd_sc_hd__a21oi_1 _08752_ (.A1(_02950_),
    .A2(_03458_),
    .B1(_02647_),
    .Y(_03459_));
 sky130_fd_sc_hd__xnor2_1 _08753_ (.A(_03457_),
    .B(_03459_),
    .Y(_03460_));
 sky130_fd_sc_hd__xnor2_1 _08754_ (.A(_03454_),
    .B(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__nor2_1 _08755_ (.A(_03232_),
    .B(_03233_),
    .Y(_03462_));
 sky130_fd_sc_hd__nor2_1 _08756_ (.A(_03234_),
    .B(_03462_),
    .Y(_03463_));
 sky130_fd_sc_hd__and2_1 _08757_ (.A(_03461_),
    .B(_03463_),
    .X(_03464_));
 sky130_fd_sc_hd__and3_1 _08758_ (.A(_03258_),
    .B(_03452_),
    .C(_03464_),
    .X(_03465_));
 sky130_fd_sc_hd__a21o_1 _08759_ (.A1(\genblk2[5].wave_shpr.div.fin_quo[0] ),
    .A2(_02467_),
    .B1(_02791_),
    .X(_03466_));
 sky130_fd_sc_hd__a21o_1 _08760_ (.A1(\genblk2[4].wave_shpr.div.fin_quo[0] ),
    .A2(_02521_),
    .B1(_02838_),
    .X(_03467_));
 sky130_fd_sc_hd__and3_1 _08761_ (.A(net10),
    .B(_02744_),
    .C(_03467_),
    .X(_03468_));
 sky130_fd_sc_hd__a21o_1 _08762_ (.A1(\genblk2[3].wave_shpr.div.fin_quo[0] ),
    .A2(_02539_),
    .B1(_02939_),
    .X(_03469_));
 sky130_fd_sc_hd__and3_1 _08763_ (.A(net9),
    .B(_02744_),
    .C(_03469_),
    .X(_03470_));
 sky130_fd_sc_hd__nand2_1 _08764_ (.A(_02798_),
    .B(_03466_),
    .Y(_03471_));
 sky130_fd_sc_hd__xnor2_1 _08765_ (.A(_03471_),
    .B(_03468_),
    .Y(_03472_));
 sky130_fd_sc_hd__and2_1 _08766_ (.A(_03470_),
    .B(_03472_),
    .X(_03473_));
 sky130_fd_sc_hd__a31o_1 _08767_ (.A1(_02798_),
    .A2(_03466_),
    .A3(_03468_),
    .B1(_03473_),
    .X(_03474_));
 sky130_fd_sc_hd__o21ba_1 _08768_ (.A1(_03455_),
    .A2(_03456_),
    .B1_N(_03459_),
    .X(_03475_));
 sky130_fd_sc_hd__or2b_1 _08769_ (.A(_03457_),
    .B_N(_03459_),
    .X(_03476_));
 sky130_fd_sc_hd__o21ai_2 _08770_ (.A1(_03454_),
    .A2(_03475_),
    .B1(_03476_),
    .Y(_03477_));
 sky130_fd_sc_hd__xnor2_1 _08771_ (.A(_03304_),
    .B(_03306_),
    .Y(_03478_));
 sky130_fd_sc_hd__xnor2_1 _08772_ (.A(_03477_),
    .B(_03478_),
    .Y(_03479_));
 sky130_fd_sc_hd__xnor2_1 _08773_ (.A(_03474_),
    .B(_03479_),
    .Y(_03480_));
 sky130_fd_sc_hd__a21oi_1 _08774_ (.A1(_03258_),
    .A2(_03452_),
    .B1(_03464_),
    .Y(_03481_));
 sky130_fd_sc_hd__nor3_2 _08775_ (.A(_03465_),
    .B(_03480_),
    .C(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__a21bo_1 _08776_ (.A1(_03298_),
    .A2(_03332_),
    .B1_N(_03331_),
    .X(_03483_));
 sky130_fd_sc_hd__o211a_1 _08777_ (.A1(_03465_),
    .A2(_03482_),
    .B1(_03333_),
    .C1(_03483_),
    .X(_03484_));
 sky130_fd_sc_hd__a211oi_2 _08778_ (.A1(_03333_),
    .A2(_03483_),
    .B1(_03465_),
    .C1(_03482_),
    .Y(_03485_));
 sky130_fd_sc_hd__a21oi_1 _08779_ (.A1(_02518_),
    .A2(_02566_),
    .B1(_02570_),
    .Y(_03486_));
 sky130_fd_sc_hd__or3b_1 _08780_ (.A(_02583_),
    .B(_03486_),
    .C_N(_02582_),
    .X(_03487_));
 sky130_fd_sc_hd__o21bai_1 _08781_ (.A1(_02583_),
    .A2(_03486_),
    .B1_N(_02582_),
    .Y(_03488_));
 sky130_fd_sc_hd__nand2_1 _08782_ (.A(_03487_),
    .B(_03488_),
    .Y(_03489_));
 sky130_fd_sc_hd__and2b_1 _08783_ (.A_N(_03478_),
    .B(_03477_),
    .X(_03490_));
 sky130_fd_sc_hd__a21o_1 _08784_ (.A1(_03474_),
    .A2(_03479_),
    .B1(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__a21oi_1 _08785_ (.A1(\genblk2[2].wave_shpr.div.fin_quo[0] ),
    .A2(_03113_),
    .B1(\genblk2[2].wave_shpr.div.fin_quo[1] ),
    .Y(_03492_));
 sky130_fd_sc_hd__a31o_1 _08786_ (.A1(\genblk2[2].wave_shpr.div.fin_quo[0] ),
    .A2(\genblk2[2].wave_shpr.div.fin_quo[1] ),
    .A3(_03113_),
    .B1(_02224_),
    .X(_03493_));
 sky130_fd_sc_hd__a2bb2o_1 _08787_ (.A1_N(_03492_),
    .A2_N(_03493_),
    .B1(\genblk2[2].wave_shpr.div.fin_quo[2] ),
    .B2(_02468_),
    .X(_03494_));
 sky130_fd_sc_hd__o21a_1 _08788_ (.A1(_03114_),
    .A2(_03494_),
    .B1(_03122_),
    .X(_03495_));
 sky130_fd_sc_hd__xnor2_1 _08789_ (.A(_03491_),
    .B(_03495_),
    .Y(_03496_));
 sky130_fd_sc_hd__xor2_1 _08790_ (.A(_03489_),
    .B(_03496_),
    .X(_03497_));
 sky130_fd_sc_hd__nor3b_2 _08791_ (.A(_03484_),
    .B(_03485_),
    .C_N(_03497_),
    .Y(_03498_));
 sky130_fd_sc_hd__o21ai_1 _08792_ (.A1(_03384_),
    .A2(_03394_),
    .B1(_03393_),
    .Y(_03499_));
 sky130_fd_sc_hd__o211a_1 _08793_ (.A1(_03484_),
    .A2(_03498_),
    .B1(_03395_),
    .C1(_03499_),
    .X(_03500_));
 sky130_fd_sc_hd__nand2_1 _08794_ (.A(_03491_),
    .B(_03495_),
    .Y(_03501_));
 sky130_fd_sc_hd__or2_1 _08795_ (.A(_03489_),
    .B(_03496_),
    .X(_03502_));
 sky130_fd_sc_hd__a211oi_2 _08796_ (.A1(_03395_),
    .A2(_03499_),
    .B1(_03484_),
    .C1(_03498_),
    .Y(_03503_));
 sky130_fd_sc_hd__a211oi_1 _08797_ (.A1(_03501_),
    .A2(_03502_),
    .B1(_03500_),
    .C1(_03503_),
    .Y(_03504_));
 sky130_fd_sc_hd__o211ai_2 _08798_ (.A1(_03425_),
    .A2(_03426_),
    .B1(_03423_),
    .C1(_03424_),
    .Y(_03505_));
 sky130_fd_sc_hd__o211a_1 _08799_ (.A1(_03500_),
    .A2(_03504_),
    .B1(_03427_),
    .C1(_03505_),
    .X(_03506_));
 sky130_fd_sc_hd__o211a_1 _08800_ (.A1(_03450_),
    .A2(_03449_),
    .B1(_03427_),
    .C1(_03422_),
    .X(_03507_));
 sky130_fd_sc_hd__o21bai_1 _08801_ (.A1(_03451_),
    .A2(_03506_),
    .B1_N(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__o211a_1 _08802_ (.A1(_03219_),
    .A2(_03222_),
    .B1(_03220_),
    .C1(_03221_),
    .X(_03509_));
 sky130_fd_sc_hd__o21ba_1 _08803_ (.A1(_03204_),
    .A2(_03205_),
    .B1_N(_03216_),
    .X(_03510_));
 sky130_fd_sc_hd__a211oi_2 _08804_ (.A1(_03442_),
    .A2(_03443_),
    .B1(_03217_),
    .C1(_03510_),
    .Y(_03511_));
 sky130_fd_sc_hd__inv_2 _08805_ (.A(_03511_),
    .Y(_03512_));
 sky130_fd_sc_hd__or2b_1 _08806_ (.A(_03433_),
    .B_N(_03437_),
    .X(_03513_));
 sky130_fd_sc_hd__nand2_1 _08807_ (.A(_03431_),
    .B(_03438_),
    .Y(_03514_));
 sky130_fd_sc_hd__o211a_1 _08808_ (.A1(_03217_),
    .A2(_03510_),
    .B1(_03442_),
    .C1(_03443_),
    .X(_03515_));
 sky130_fd_sc_hd__a211o_1 _08809_ (.A1(_03513_),
    .A2(_03514_),
    .B1(_03511_),
    .C1(_03515_),
    .X(_03516_));
 sky130_fd_sc_hd__o211a_1 _08810_ (.A1(_03223_),
    .A2(_03509_),
    .B1(_03512_),
    .C1(_03516_),
    .X(_03517_));
 sky130_fd_sc_hd__a211o_1 _08811_ (.A1(_03512_),
    .A2(_03516_),
    .B1(_03223_),
    .C1(_03509_),
    .X(_03518_));
 sky130_fd_sc_hd__or2b_1 _08812_ (.A(_03517_),
    .B_N(_03518_),
    .X(_03519_));
 sky130_fd_sc_hd__o211ai_2 _08813_ (.A1(_03511_),
    .A2(_03515_),
    .B1(_03513_),
    .C1(_03514_),
    .Y(_03520_));
 sky130_fd_sc_hd__o211ai_2 _08814_ (.A1(_03445_),
    .A2(_03450_),
    .B1(_03516_),
    .C1(_03520_),
    .Y(_03521_));
 sky130_fd_sc_hd__a211o_1 _08815_ (.A1(_03516_),
    .A2(_03520_),
    .B1(_03445_),
    .C1(_03450_),
    .X(_03522_));
 sky130_fd_sc_hd__nand2_1 _08816_ (.A(_03521_),
    .B(_03522_),
    .Y(_03523_));
 sky130_fd_sc_hd__a21o_1 _08817_ (.A1(_03518_),
    .A2(_03521_),
    .B1(_03517_),
    .X(_03524_));
 sky130_fd_sc_hd__o31a_1 _08818_ (.A1(_03508_),
    .A2(_03519_),
    .A3(_03523_),
    .B1(_03524_),
    .X(_03525_));
 sky130_fd_sc_hd__nor2_1 _08819_ (.A(_03461_),
    .B(_03463_),
    .Y(_03526_));
 sky130_fd_sc_hd__nor2_1 _08820_ (.A(_03470_),
    .B(_03472_),
    .Y(_03527_));
 sky130_fd_sc_hd__or2_1 _08821_ (.A(_03473_),
    .B(_03527_),
    .X(_03528_));
 sky130_fd_sc_hd__or3_1 _08822_ (.A(_03464_),
    .B(_03526_),
    .C(_03528_),
    .X(_03529_));
 sky130_fd_sc_hd__o21a_1 _08823_ (.A1(_03465_),
    .A2(_03481_),
    .B1(_03480_),
    .X(_03530_));
 sky130_fd_sc_hd__or3_1 _08824_ (.A(_03482_),
    .B(_03529_),
    .C(_03530_),
    .X(_03531_));
 sky130_fd_sc_hd__or2b_1 _08825_ (.A(_02581_),
    .B_N(_02580_),
    .X(_03532_));
 sky130_fd_sc_hd__xor2_2 _08826_ (.A(_02575_),
    .B(_03532_),
    .X(_03533_));
 sky130_fd_sc_hd__a221o_1 _08827_ (.A1(\genblk2[2].wave_shpr.div.fin_quo[0] ),
    .A2(_02592_),
    .B1(_02468_),
    .B2(\genblk2[2].wave_shpr.div.fin_quo[1] ),
    .C1(_03114_),
    .X(_03534_));
 sky130_fd_sc_hd__and3_1 _08828_ (.A(net8),
    .B(_02744_),
    .C(_03534_),
    .X(_03535_));
 sky130_fd_sc_hd__xnor2_1 _08829_ (.A(_03533_),
    .B(_03535_),
    .Y(_03536_));
 sky130_fd_sc_hd__o21ai_1 _08830_ (.A1(_03482_),
    .A2(_03530_),
    .B1(_03529_),
    .Y(_03537_));
 sky130_fd_sc_hd__and3_1 _08831_ (.A(_03531_),
    .B(_03536_),
    .C(_03537_),
    .X(_03538_));
 sky130_fd_sc_hd__a21oi_1 _08832_ (.A1(_03531_),
    .A2(_03537_),
    .B1(_03536_),
    .Y(_03539_));
 sky130_fd_sc_hd__nor2_1 _08833_ (.A(_03538_),
    .B(_03539_),
    .Y(_03540_));
 sky130_fd_sc_hd__a21o_1 _08834_ (.A1(\genblk2[2].wave_shpr.div.fin_quo[0] ),
    .A2(_02468_),
    .B1(_03114_),
    .X(_03541_));
 sky130_fd_sc_hd__and3_1 _08835_ (.A(net8),
    .B(_02744_),
    .C(_03541_),
    .X(_03542_));
 sky130_fd_sc_hd__o21ai_1 _08836_ (.A1(_02509_),
    .A2(_02572_),
    .B1(_02518_),
    .Y(_03543_));
 sky130_fd_sc_hd__xnor2_2 _08837_ (.A(_02574_),
    .B(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__and2_1 _08838_ (.A(_03542_),
    .B(_03544_),
    .X(_03545_));
 sky130_fd_sc_hd__nand2_1 _08839_ (.A(_03540_),
    .B(_03545_),
    .Y(_03546_));
 sky130_fd_sc_hd__o21ai_1 _08840_ (.A1(_03464_),
    .A2(_03526_),
    .B1(_03528_),
    .Y(_03547_));
 sky130_fd_sc_hd__or2_1 _08841_ (.A(_03542_),
    .B(_03544_),
    .X(_03548_));
 sky130_fd_sc_hd__and2b_1 _08842_ (.A_N(_03545_),
    .B(_03548_),
    .X(_03549_));
 sky130_fd_sc_hd__and3_1 _08843_ (.A(_03529_),
    .B(_03547_),
    .C(_03549_),
    .X(_03550_));
 sky130_fd_sc_hd__nand2_1 _08844_ (.A(_03540_),
    .B(_03550_),
    .Y(_03551_));
 sky130_fd_sc_hd__and2b_1 _08845_ (.A_N(_03533_),
    .B(_03535_),
    .X(_03552_));
 sky130_fd_sc_hd__o21ba_1 _08846_ (.A1(_03484_),
    .A2(_03485_),
    .B1_N(_03497_),
    .X(_03553_));
 sky130_fd_sc_hd__a21boi_1 _08847_ (.A1(_03536_),
    .A2(_03537_),
    .B1_N(_03531_),
    .Y(_03554_));
 sky130_fd_sc_hd__or3_1 _08848_ (.A(_03498_),
    .B(_03553_),
    .C(_03554_),
    .X(_03555_));
 sky130_fd_sc_hd__o21ai_1 _08849_ (.A1(_03498_),
    .A2(_03553_),
    .B1(_03554_),
    .Y(_03556_));
 sky130_fd_sc_hd__and3_1 _08850_ (.A(_03552_),
    .B(_03555_),
    .C(_03556_),
    .X(_03557_));
 sky130_fd_sc_hd__a21oi_1 _08851_ (.A1(_03555_),
    .A2(_03556_),
    .B1(_03552_),
    .Y(_03558_));
 sky130_fd_sc_hd__a211oi_2 _08852_ (.A1(_03546_),
    .A2(_03551_),
    .B1(_03557_),
    .C1(_03558_),
    .Y(_03559_));
 sky130_fd_sc_hd__a211o_1 _08853_ (.A1(_03501_),
    .A2(_03502_),
    .B1(_03500_),
    .C1(_03503_),
    .X(_03560_));
 sky130_fd_sc_hd__o211ai_1 _08854_ (.A1(_03500_),
    .A2(_03503_),
    .B1(_03501_),
    .C1(_03502_),
    .Y(_03561_));
 sky130_fd_sc_hd__nor3_1 _08855_ (.A(_03498_),
    .B(_03553_),
    .C(_03554_),
    .Y(_03562_));
 sky130_fd_sc_hd__a211o_1 _08856_ (.A1(_03560_),
    .A2(_03561_),
    .B1(_03562_),
    .C1(_03557_),
    .X(_03563_));
 sky130_fd_sc_hd__o211a_1 _08857_ (.A1(_03562_),
    .A2(_03557_),
    .B1(_03560_),
    .C1(_03561_),
    .X(_03564_));
 sky130_fd_sc_hd__a21oi_1 _08858_ (.A1(_03559_),
    .A2(_03563_),
    .B1(_03564_),
    .Y(_03565_));
 sky130_fd_sc_hd__a211oi_1 _08859_ (.A1(_03427_),
    .A2(_03505_),
    .B1(_03500_),
    .C1(_03504_),
    .Y(_03566_));
 sky130_fd_sc_hd__or4_1 _08860_ (.A(_03507_),
    .B(_03451_),
    .C(_03506_),
    .D(_03566_),
    .X(_03567_));
 sky130_fd_sc_hd__or4_1 _08861_ (.A(_03565_),
    .B(_03567_),
    .C(_03519_),
    .D(_03523_),
    .X(_03568_));
 sky130_fd_sc_hd__xnor2_1 _08862_ (.A(_03136_),
    .B(_03224_),
    .Y(_03569_));
 sky130_fd_sc_hd__a21oi_1 _08863_ (.A1(_03525_),
    .A2(_03568_),
    .B1(_03569_),
    .Y(_03570_));
 sky130_fd_sc_hd__nor3_1 _08864_ (.A(_03135_),
    .B(_03225_),
    .C(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hd__o31ai_2 _08865_ (.A1(_03009_),
    .A2(_03134_),
    .A3(_03571_),
    .B1(_02248_),
    .Y(_03572_));
 sky130_fd_sc_hd__o211a_1 _08866_ (.A1(net428),
    .A2(_02248_),
    .B1(_00024_),
    .C1(_03572_),
    .X(_03573_));
 sky130_fd_sc_hd__a21o_1 _08867_ (.A1(net1131),
    .A2(_02260_),
    .B1(_03573_),
    .X(_00038_));
 sky130_fd_sc_hd__clkbuf_4 _08868_ (.A(_01156_),
    .X(_03574_));
 sky130_fd_sc_hd__inv_2 _08869_ (.A(\sig_norm.b1[3] ),
    .Y(_03575_));
 sky130_fd_sc_hd__inv_2 _08870_ (.A(\sig_norm.b1[2] ),
    .Y(_03576_));
 sky130_fd_sc_hd__or2b_1 _08871_ (.A(\sig_norm.b1[1] ),
    .B_N(\sig_norm.acc[1] ),
    .X(_03577_));
 sky130_fd_sc_hd__inv_2 _08872_ (.A(\sig_norm.acc[0] ),
    .Y(_03578_));
 sky130_fd_sc_hd__or2b_1 _08873_ (.A(\sig_norm.acc[1] ),
    .B_N(\sig_norm.b1[1] ),
    .X(_03579_));
 sky130_fd_sc_hd__nand2_1 _08874_ (.A(_03577_),
    .B(_03579_),
    .Y(_03580_));
 sky130_fd_sc_hd__a21o_1 _08875_ (.A1(\sig_norm.b1[0] ),
    .A2(_03578_),
    .B1(_03580_),
    .X(_03581_));
 sky130_fd_sc_hd__xor2_1 _08876_ (.A(\sig_norm.b1[2] ),
    .B(\sig_norm.acc[2] ),
    .X(_03582_));
 sky130_fd_sc_hd__a21oi_1 _08877_ (.A1(_03577_),
    .A2(_03581_),
    .B1(_03582_),
    .Y(_03583_));
 sky130_fd_sc_hd__a21o_1 _08878_ (.A1(_03576_),
    .A2(\sig_norm.acc[2] ),
    .B1(_03583_),
    .X(_03584_));
 sky130_fd_sc_hd__o21a_1 _08879_ (.A1(_03575_),
    .A2(\sig_norm.acc[3] ),
    .B1(_03584_),
    .X(_03585_));
 sky130_fd_sc_hd__a21o_1 _08880_ (.A1(_03575_),
    .A2(\sig_norm.acc[3] ),
    .B1(_03585_),
    .X(_03586_));
 sky130_fd_sc_hd__or2_1 _08881_ (.A(\sig_norm.acc[4] ),
    .B(_03586_),
    .X(_03587_));
 sky130_fd_sc_hd__or4_1 _08882_ (.A(\sig_norm.acc[7] ),
    .B(\sig_norm.acc[6] ),
    .C(\sig_norm.acc[5] ),
    .D(_03587_),
    .X(_03588_));
 sky130_fd_sc_hd__or2_1 _08883_ (.A(\sig_norm.acc[8] ),
    .B(_03588_),
    .X(_03589_));
 sky130_fd_sc_hd__or2_1 _08884_ (.A(\sig_norm.acc[9] ),
    .B(_03589_),
    .X(_03590_));
 sky130_fd_sc_hd__or2_1 _08885_ (.A(\sig_norm.acc[10] ),
    .B(_03590_),
    .X(_03591_));
 sky130_fd_sc_hd__xnor2_1 _08886_ (.A(\sig_norm.b1[3] ),
    .B(\sig_norm.acc[3] ),
    .Y(_03592_));
 sky130_fd_sc_hd__o21ai_1 _08887_ (.A1(\sig_norm.b1[0] ),
    .A2(_03578_),
    .B1(_03592_),
    .Y(_03593_));
 sky130_fd_sc_hd__nor3_1 _08888_ (.A(_03582_),
    .B(_03581_),
    .C(_03593_),
    .Y(_03594_));
 sky130_fd_sc_hd__or4_1 _08889_ (.A(\sig_norm.acc[11] ),
    .B(\sig_norm.acc[12] ),
    .C(_03591_),
    .D(_03594_),
    .X(_03595_));
 sky130_fd_sc_hd__buf_2 _08890_ (.A(_03595_),
    .X(_03596_));
 sky130_fd_sc_hd__nand2_1 _08891_ (.A(\sig_norm.b1[0] ),
    .B(_03596_),
    .Y(_03597_));
 sky130_fd_sc_hd__xnor2_1 _08892_ (.A(\sig_norm.acc[0] ),
    .B(_03597_),
    .Y(_03598_));
 sky130_fd_sc_hd__and3_1 _08893_ (.A(_01099_),
    .B(_03574_),
    .C(_03598_),
    .X(_03599_));
 sky130_fd_sc_hd__a21o_1 _08894_ (.A1(net629),
    .A2(_02260_),
    .B1(_03599_),
    .X(_00039_));
 sky130_fd_sc_hd__or2_1 _08895_ (.A(net629),
    .B(_03596_),
    .X(_03600_));
 sky130_fd_sc_hd__nand3_1 _08896_ (.A(\sig_norm.b1[0] ),
    .B(_03578_),
    .C(_03580_),
    .Y(_03601_));
 sky130_fd_sc_hd__nor4_2 _08897_ (.A(\sig_norm.acc[11] ),
    .B(\sig_norm.acc[12] ),
    .C(_03591_),
    .D(_03594_),
    .Y(_03602_));
 sky130_fd_sc_hd__a21o_1 _08898_ (.A1(_03581_),
    .A2(_03601_),
    .B1(net26),
    .X(_03603_));
 sky130_fd_sc_hd__a32o_1 _08899_ (.A1(_03574_),
    .A2(_03600_),
    .A3(_03603_),
    .B1(_01157_),
    .B2(net1069),
    .X(_00040_));
 sky130_fd_sc_hd__or2_1 _08900_ (.A(\sig_norm.acc[2] ),
    .B(_03596_),
    .X(_03604_));
 sky130_fd_sc_hd__and3_1 _08901_ (.A(_03582_),
    .B(_03577_),
    .C(_03581_),
    .X(_03605_));
 sky130_fd_sc_hd__o21ai_1 _08902_ (.A1(_03583_),
    .A2(_03605_),
    .B1(_03596_),
    .Y(_03606_));
 sky130_fd_sc_hd__a32o_1 _08903_ (.A1(_03574_),
    .A2(_03604_),
    .A3(_03606_),
    .B1(_01157_),
    .B2(net1065),
    .X(_00041_));
 sky130_fd_sc_hd__xnor2_1 _08904_ (.A(_03584_),
    .B(_03592_),
    .Y(_03607_));
 sky130_fd_sc_hd__a21oi_1 _08905_ (.A1(_03596_),
    .A2(_03607_),
    .B1(_02248_),
    .Y(_03608_));
 sky130_fd_sc_hd__o21a_1 _08906_ (.A1(\sig_norm.acc[3] ),
    .A2(_03596_),
    .B1(_03608_),
    .X(_03609_));
 sky130_fd_sc_hd__mux2_1 _08907_ (.A0(_03609_),
    .A1(net1240),
    .S(_01157_),
    .X(_03610_));
 sky130_fd_sc_hd__clkbuf_1 _08908_ (.A(_03610_),
    .X(_00042_));
 sky130_fd_sc_hd__or2_1 _08909_ (.A(_03587_),
    .B(net26),
    .X(_03611_));
 sky130_fd_sc_hd__o21ai_1 _08910_ (.A1(_03586_),
    .A2(net26),
    .B1(\sig_norm.acc[4] ),
    .Y(_03612_));
 sky130_fd_sc_hd__nand2_1 _08911_ (.A(_03611_),
    .B(_03612_),
    .Y(_03613_));
 sky130_fd_sc_hd__a22o_1 _08912_ (.A1(net1027),
    .A2(_02260_),
    .B1(_03613_),
    .B2(_03574_),
    .X(_00043_));
 sky130_fd_sc_hd__or2_1 _08913_ (.A(\sig_norm.acc[5] ),
    .B(_03611_),
    .X(_03614_));
 sky130_fd_sc_hd__nand2_1 _08914_ (.A(\sig_norm.acc[5] ),
    .B(_03611_),
    .Y(_03615_));
 sky130_fd_sc_hd__nand2_1 _08915_ (.A(_03614_),
    .B(_03615_),
    .Y(_03616_));
 sky130_fd_sc_hd__a22o_1 _08916_ (.A1(net1155),
    .A2(_02260_),
    .B1(_03616_),
    .B2(_03574_),
    .X(_00044_));
 sky130_fd_sc_hd__xnor2_1 _08917_ (.A(\sig_norm.acc[6] ),
    .B(_03614_),
    .Y(_03617_));
 sky130_fd_sc_hd__a22o_1 _08918_ (.A1(net612),
    .A2(_02260_),
    .B1(_03617_),
    .B2(_03574_),
    .X(_00045_));
 sky130_fd_sc_hd__o21ai_1 _08919_ (.A1(\sig_norm.acc[6] ),
    .A2(_03614_),
    .B1(net612),
    .Y(_03618_));
 sky130_fd_sc_hd__o21ai_1 _08920_ (.A1(_03588_),
    .A2(_03602_),
    .B1(_03618_),
    .Y(_03619_));
 sky130_fd_sc_hd__a22o_1 _08921_ (.A1(net678),
    .A2(_02260_),
    .B1(_03619_),
    .B2(_03574_),
    .X(_00046_));
 sky130_fd_sc_hd__nand2_1 _08922_ (.A(net678),
    .B(_03588_),
    .Y(_03620_));
 sky130_fd_sc_hd__o21ai_1 _08923_ (.A1(_03589_),
    .A2(_03602_),
    .B1(_03620_),
    .Y(_03621_));
 sky130_fd_sc_hd__a22o_1 _08924_ (.A1(net717),
    .A2(_02260_),
    .B1(_03621_),
    .B2(_03574_),
    .X(_00047_));
 sky130_fd_sc_hd__nor2_1 _08925_ (.A(_03590_),
    .B(_03602_),
    .Y(_03622_));
 sky130_fd_sc_hd__a21o_1 _08926_ (.A1(\sig_norm.acc[9] ),
    .A2(_03589_),
    .B1(_03622_),
    .X(_03623_));
 sky130_fd_sc_hd__and3_1 _08927_ (.A(_01099_),
    .B(_01156_),
    .C(_03623_),
    .X(_03624_));
 sky130_fd_sc_hd__a21o_1 _08928_ (.A1(net663),
    .A2(_02260_),
    .B1(_03624_),
    .X(_00048_));
 sky130_fd_sc_hd__and2b_1 _08929_ (.A_N(\sig_norm.acc[10] ),
    .B(_03622_),
    .X(_03625_));
 sky130_fd_sc_hd__a21o_1 _08930_ (.A1(\sig_norm.acc[10] ),
    .A2(_03590_),
    .B1(_03625_),
    .X(_03626_));
 sky130_fd_sc_hd__a22o_1 _08931_ (.A1(net1141),
    .A2(_02260_),
    .B1(_03626_),
    .B2(_03574_),
    .X(_00049_));
 sky130_fd_sc_hd__mux2_1 _08932_ (.A0(_03625_),
    .A1(_03591_),
    .S(\sig_norm.acc[11] ),
    .X(_03627_));
 sky130_fd_sc_hd__and2_1 _08933_ (.A(\sig_norm.acc[12] ),
    .B(_01157_),
    .X(_03628_));
 sky130_fd_sc_hd__a31o_1 _08934_ (.A1(_01099_),
    .A2(_00024_),
    .A3(_03627_),
    .B1(_03628_),
    .X(_00050_));
 sky130_fd_sc_hd__a22o_1 _08935_ (.A1(net1083),
    .A2(_02260_),
    .B1(_03596_),
    .B2(_03574_),
    .X(_00051_));
 sky130_fd_sc_hd__a21o_1 _08936_ (.A1(_03529_),
    .A2(_03547_),
    .B1(_03549_),
    .X(_03629_));
 sky130_fd_sc_hd__nor2_1 _08937_ (.A(_01098_),
    .B(_03550_),
    .Y(_03630_));
 sky130_fd_sc_hd__a22o_1 _08938_ (.A1(\sig_norm.quo[0] ),
    .A2(_01098_),
    .B1(_03629_),
    .B2(_03630_),
    .X(_03631_));
 sky130_fd_sc_hd__mux2_1 _08939_ (.A0(\sig_norm.quo[1] ),
    .A1(_03631_),
    .S(_00024_),
    .X(_03632_));
 sky130_fd_sc_hd__clkbuf_1 _08940_ (.A(_03632_),
    .X(_00052_));
 sky130_fd_sc_hd__or2_1 _08941_ (.A(_03540_),
    .B(_03550_),
    .X(_03633_));
 sky130_fd_sc_hd__and2_1 _08942_ (.A(_03551_),
    .B(_03633_),
    .X(_03634_));
 sky130_fd_sc_hd__o211a_1 _08943_ (.A1(_03545_),
    .A2(_03634_),
    .B1(_03546_),
    .C1(_01155_),
    .X(_03635_));
 sky130_fd_sc_hd__a21o_1 _08944_ (.A1(\sig_norm.quo[1] ),
    .A2(_01098_),
    .B1(_03635_),
    .X(_03636_));
 sky130_fd_sc_hd__mux2_1 _08945_ (.A0(\sig_norm.quo[2] ),
    .A1(_03636_),
    .S(_00024_),
    .X(_03637_));
 sky130_fd_sc_hd__clkbuf_1 _08946_ (.A(_03637_),
    .X(_00053_));
 sky130_fd_sc_hd__o211a_1 _08947_ (.A1(_03557_),
    .A2(_03558_),
    .B1(_03546_),
    .C1(_03551_),
    .X(_03638_));
 sky130_fd_sc_hd__or2_1 _08948_ (.A(_01098_),
    .B(_03559_),
    .X(_03639_));
 sky130_fd_sc_hd__a2bb2o_1 _08949_ (.A1_N(_03638_),
    .A2_N(_03639_),
    .B1(\sig_norm.quo[2] ),
    .B2(_01098_),
    .X(_03640_));
 sky130_fd_sc_hd__mux2_1 _08950_ (.A0(\sig_norm.quo[3] ),
    .A1(_03640_),
    .S(_00024_),
    .X(_03641_));
 sky130_fd_sc_hd__clkbuf_1 _08951_ (.A(_03641_),
    .X(_00054_));
 sky130_fd_sc_hd__or2b_1 _08952_ (.A(_03564_),
    .B_N(_03563_),
    .X(_03642_));
 sky130_fd_sc_hd__xnor2_1 _08953_ (.A(_03559_),
    .B(_03642_),
    .Y(_03643_));
 sky130_fd_sc_hd__mux2_1 _08954_ (.A0(\sig_norm.quo[3] ),
    .A1(_03643_),
    .S(_02248_),
    .X(_03644_));
 sky130_fd_sc_hd__mux2_1 _08955_ (.A0(net1339),
    .A1(_03644_),
    .S(_00024_),
    .X(_03645_));
 sky130_fd_sc_hd__clkbuf_1 _08956_ (.A(_03645_),
    .X(_00055_));
 sky130_fd_sc_hd__nor2_1 _08957_ (.A(_03506_),
    .B(_03566_),
    .Y(_03646_));
 sky130_fd_sc_hd__xnor2_1 _08958_ (.A(_03565_),
    .B(_03646_),
    .Y(_03647_));
 sky130_fd_sc_hd__mux2_1 _08959_ (.A0(\sig_norm.quo[4] ),
    .A1(_03647_),
    .S(_02248_),
    .X(_03648_));
 sky130_fd_sc_hd__mux2_1 _08960_ (.A0(\sig_norm.quo[5] ),
    .A1(_03648_),
    .S(_00024_),
    .X(_03649_));
 sky130_fd_sc_hd__clkbuf_1 _08961_ (.A(_03649_),
    .X(_00056_));
 sky130_fd_sc_hd__nor2_1 _08962_ (.A(_03507_),
    .B(_03451_),
    .Y(_03650_));
 sky130_fd_sc_hd__a21o_1 _08963_ (.A1(_03559_),
    .A2(_03563_),
    .B1(_03564_),
    .X(_03651_));
 sky130_fd_sc_hd__a21oi_1 _08964_ (.A1(_03651_),
    .A2(_03646_),
    .B1(_03506_),
    .Y(_03652_));
 sky130_fd_sc_hd__xnor2_1 _08965_ (.A(_03650_),
    .B(_03652_),
    .Y(_03653_));
 sky130_fd_sc_hd__mux2_1 _08966_ (.A0(\sig_norm.quo[5] ),
    .A1(_03653_),
    .S(_01155_),
    .X(_03654_));
 sky130_fd_sc_hd__mux2_1 _08967_ (.A0(\sig_norm.quo[6] ),
    .A1(_03654_),
    .S(_00024_),
    .X(_03655_));
 sky130_fd_sc_hd__clkbuf_1 _08968_ (.A(_03655_),
    .X(_00057_));
 sky130_fd_sc_hd__o21a_1 _08969_ (.A1(_03565_),
    .A2(_03567_),
    .B1(_03508_),
    .X(_03656_));
 sky130_fd_sc_hd__nor2_1 _08970_ (.A(_03656_),
    .B(_03523_),
    .Y(_03657_));
 sky130_fd_sc_hd__a21o_1 _08971_ (.A1(_03656_),
    .A2(_03523_),
    .B1(_01098_),
    .X(_03658_));
 sky130_fd_sc_hd__a2bb2o_1 _08972_ (.A1_N(_03657_),
    .A2_N(_03658_),
    .B1(\sig_norm.quo[6] ),
    .B2(_01098_),
    .X(_03659_));
 sky130_fd_sc_hd__mux2_1 _08973_ (.A0(net1300),
    .A1(_03659_),
    .S(_01158_),
    .X(_03660_));
 sky130_fd_sc_hd__clkbuf_1 _08974_ (.A(_03660_),
    .X(_00058_));
 sky130_fd_sc_hd__inv_2 _08975_ (.A(\sig_norm.quo[7] ),
    .Y(_03661_));
 sky130_fd_sc_hd__o21a_1 _08976_ (.A1(_03656_),
    .A2(_03523_),
    .B1(_03521_),
    .X(_03662_));
 sky130_fd_sc_hd__xnor2_1 _08977_ (.A(_03519_),
    .B(_03662_),
    .Y(_03663_));
 sky130_fd_sc_hd__mux2_1 _08978_ (.A0(_03661_),
    .A1(_03663_),
    .S(_02248_),
    .X(_03664_));
 sky130_fd_sc_hd__nand2_1 _08979_ (.A(net372),
    .B(_01157_),
    .Y(_03665_));
 sky130_fd_sc_hd__o21ai_1 _08980_ (.A1(_01157_),
    .A2(_03664_),
    .B1(_03665_),
    .Y(_00059_));
 sky130_fd_sc_hd__and3_1 _08981_ (.A(_03525_),
    .B(_03568_),
    .C(_03569_),
    .X(_03666_));
 sky130_fd_sc_hd__or3_1 _08982_ (.A(_01097_),
    .B(_03570_),
    .C(_03666_),
    .X(_03667_));
 sky130_fd_sc_hd__a21bo_1 _08983_ (.A1(\sig_norm.quo[8] ),
    .A2(_01098_),
    .B1_N(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__mux2_1 _08984_ (.A0(net1156),
    .A1(_03668_),
    .S(_01158_),
    .X(_03669_));
 sky130_fd_sc_hd__clkbuf_1 _08985_ (.A(_03669_),
    .X(_00060_));
 sky130_fd_sc_hd__nor2_1 _08986_ (.A(_03225_),
    .B(_03570_),
    .Y(_03670_));
 sky130_fd_sc_hd__nor2_1 _08987_ (.A(_03134_),
    .B(_03135_),
    .Y(_03671_));
 sky130_fd_sc_hd__xnor2_1 _08988_ (.A(_03670_),
    .B(_03671_),
    .Y(_03672_));
 sky130_fd_sc_hd__mux2_1 _08989_ (.A0(\sig_norm.quo[9] ),
    .A1(_03672_),
    .S(_01155_),
    .X(_03673_));
 sky130_fd_sc_hd__mux2_1 _08990_ (.A0(net1261),
    .A1(_03673_),
    .S(_01158_),
    .X(_03674_));
 sky130_fd_sc_hd__clkbuf_1 _08991_ (.A(_03674_),
    .X(_00061_));
 sky130_fd_sc_hd__o21a_1 _08992_ (.A1(_03134_),
    .A2(_03571_),
    .B1(_03009_),
    .X(_03675_));
 sky130_fd_sc_hd__nor2_1 _08993_ (.A(_03572_),
    .B(_03675_),
    .Y(_03676_));
 sky130_fd_sc_hd__a21o_1 _08994_ (.A1(\sig_norm.quo[10] ),
    .A2(_01099_),
    .B1(_01157_),
    .X(_03677_));
 sky130_fd_sc_hd__o22a_1 _08995_ (.A1(net428),
    .A2(_00024_),
    .B1(_03676_),
    .B2(_03677_),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _08996_ (.A0(net1134),
    .A1(_03596_),
    .S(_01154_),
    .X(_03678_));
 sky130_fd_sc_hd__clkbuf_1 _08997_ (.A(_03678_),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _08998_ (.A0(net1103),
    .A1(\sig_norm.quo[0] ),
    .S(_01154_),
    .X(_03679_));
 sky130_fd_sc_hd__clkbuf_1 _08999_ (.A(_03679_),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _09000_ (.A0(net1102),
    .A1(net1126),
    .S(_01154_),
    .X(_03680_));
 sky130_fd_sc_hd__clkbuf_1 _09001_ (.A(_03680_),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _09002_ (.A0(net1172),
    .A1(net1176),
    .S(_01154_),
    .X(_03681_));
 sky130_fd_sc_hd__clkbuf_1 _09003_ (.A(_03681_),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _09004_ (.A0(net1150),
    .A1(\sig_norm.quo[3] ),
    .S(_01154_),
    .X(_03682_));
 sky130_fd_sc_hd__clkbuf_1 _09005_ (.A(net1151),
    .X(_00067_));
 sky130_fd_sc_hd__mux2_1 _09006_ (.A0(net1168),
    .A1(net1170),
    .S(_01154_),
    .X(_03683_));
 sky130_fd_sc_hd__clkbuf_1 _09007_ (.A(_03683_),
    .X(_00068_));
 sky130_fd_sc_hd__mux2_1 _09008_ (.A0(net1132),
    .A1(\sig_norm.quo[5] ),
    .S(_01154_),
    .X(_03684_));
 sky130_fd_sc_hd__clkbuf_1 _09009_ (.A(_03684_),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _09010_ (.A0(net1128),
    .A1(\sig_norm.quo[6] ),
    .S(_01154_),
    .X(_03685_));
 sky130_fd_sc_hd__clkbuf_1 _09011_ (.A(_03685_),
    .X(_00070_));
 sky130_fd_sc_hd__nand2_1 _09012_ (.A(\genblk2[9].wave_shpr.div.i[0] ),
    .B(_02202_),
    .Y(_03686_));
 sky130_fd_sc_hd__buf_6 _09013_ (.A(_02171_),
    .X(_03687_));
 sky130_fd_sc_hd__o211a_1 _09014_ (.A1(\genblk2[9].wave_shpr.div.busy ),
    .A2(\genblk2[9].wave_shpr.div.i[0] ),
    .B1(_03686_),
    .C1(_03687_),
    .X(_00071_));
 sky130_fd_sc_hd__a21oi_1 _09015_ (.A1(\genblk2[9].wave_shpr.div.i[0] ),
    .A2(_02202_),
    .B1(\genblk2[9].wave_shpr.div.i[1] ),
    .Y(_03688_));
 sky130_fd_sc_hd__buf_4 _09016_ (.A(_02155_),
    .X(_03689_));
 sky130_fd_sc_hd__buf_8 _09017_ (.A(_03689_),
    .X(_03690_));
 sky130_fd_sc_hd__a311oi_1 _09018_ (.A1(\genblk2[9].wave_shpr.div.busy ),
    .A2(net1039),
    .A3(\genblk2[9].wave_shpr.div.i[0] ),
    .B1(_03688_),
    .C1(_03690_),
    .Y(_00072_));
 sky130_fd_sc_hd__a21o_1 _09019_ (.A1(\genblk2[9].wave_shpr.div.i[1] ),
    .A2(\genblk2[9].wave_shpr.div.i[0] ),
    .B1(\genblk2[9].wave_shpr.div.i[2] ),
    .X(_03691_));
 sky130_fd_sc_hd__and3_1 _09020_ (.A(_02152_),
    .B(\genblk2[9].wave_shpr.div.busy ),
    .C(_02201_),
    .X(_03692_));
 sky130_fd_sc_hd__clkbuf_4 _09021_ (.A(_03692_),
    .X(_03693_));
 sky130_fd_sc_hd__clkbuf_4 _09022_ (.A(_03693_),
    .X(_03694_));
 sky130_fd_sc_hd__nand3_1 _09023_ (.A(\genblk2[9].wave_shpr.div.i[1] ),
    .B(\genblk2[9].wave_shpr.div.i[0] ),
    .C(\genblk2[9].wave_shpr.div.i[2] ),
    .Y(_03695_));
 sky130_fd_sc_hd__clkbuf_4 _09024_ (.A(_02203_),
    .X(_03696_));
 sky130_fd_sc_hd__a32o_1 _09025_ (.A1(_03691_),
    .A2(_03694_),
    .A3(_03695_),
    .B1(_03696_),
    .B2(net1149),
    .X(_00073_));
 sky130_fd_sc_hd__a31o_1 _09026_ (.A1(\genblk2[9].wave_shpr.div.i[1] ),
    .A2(\genblk2[9].wave_shpr.div.i[0] ),
    .A3(\genblk2[9].wave_shpr.div.i[2] ),
    .B1(\genblk2[9].wave_shpr.div.i[3] ),
    .X(_03697_));
 sky130_fd_sc_hd__and4_1 _09027_ (.A(\genblk2[9].wave_shpr.div.i[1] ),
    .B(\genblk2[9].wave_shpr.div.i[0] ),
    .C(\genblk2[9].wave_shpr.div.i[2] ),
    .D(\genblk2[9].wave_shpr.div.i[3] ),
    .X(_03698_));
 sky130_fd_sc_hd__inv_2 _09028_ (.A(_03698_),
    .Y(_03699_));
 sky130_fd_sc_hd__a32o_1 _09029_ (.A1(_03694_),
    .A2(_03697_),
    .A3(_03699_),
    .B1(_03696_),
    .B2(net789),
    .X(_00074_));
 sky130_fd_sc_hd__a21oi_1 _09030_ (.A1(\genblk2[9].wave_shpr.div.busy ),
    .A2(_03698_),
    .B1(net817),
    .Y(_03700_));
 sky130_fd_sc_hd__buf_8 _09031_ (.A(_02155_),
    .X(_03701_));
 sky130_fd_sc_hd__buf_8 _09032_ (.A(_03701_),
    .X(_03702_));
 sky130_fd_sc_hd__a31o_1 _09033_ (.A1(net817),
    .A2(_02202_),
    .A3(_03698_),
    .B1(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__nor2_1 _09034_ (.A(_03700_),
    .B(_03703_),
    .Y(_00075_));
 sky130_fd_sc_hd__buf_6 _09035_ (.A(_02171_),
    .X(_03704_));
 sky130_fd_sc_hd__nand2_8 _09036_ (.A(_03702_),
    .B(_01432_),
    .Y(_03705_));
 sky130_fd_sc_hd__a21bo_1 _09037_ (.A1(_03704_),
    .A2(net861),
    .B1_N(_03705_),
    .X(_00076_));
 sky130_fd_sc_hd__nand2_2 _09038_ (.A(_02336_),
    .B(net34),
    .Y(_03706_));
 sky130_fd_sc_hd__clkbuf_8 _09039_ (.A(_02147_),
    .X(_03707_));
 sky130_fd_sc_hd__buf_8 _09040_ (.A(_03707_),
    .X(_03708_));
 sky130_fd_sc_hd__mux2_1 _09041_ (.A0(net1243),
    .A1(_03706_),
    .S(_03708_),
    .X(_03709_));
 sky130_fd_sc_hd__clkbuf_1 _09042_ (.A(_03709_),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _09043_ (.A0(\genblk2[0].wave_shpr.div.b1[2] ),
    .A1(_02002_),
    .S(_03708_),
    .X(_03710_));
 sky130_fd_sc_hd__clkbuf_1 _09044_ (.A(_03710_),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _09045_ (.A0(net1238),
    .A1(_01991_),
    .S(_03708_),
    .X(_03711_));
 sky130_fd_sc_hd__clkbuf_1 _09046_ (.A(_03711_),
    .X(_00079_));
 sky130_fd_sc_hd__nor2_2 _09047_ (.A(_01248_),
    .B(_02374_),
    .Y(_03712_));
 sky130_fd_sc_hd__mux2_1 _09048_ (.A0(\genblk2[0].wave_shpr.div.b1[4] ),
    .A1(_03712_),
    .S(_03708_),
    .X(_03713_));
 sky130_fd_sc_hd__clkbuf_1 _09049_ (.A(_03713_),
    .X(_00080_));
 sky130_fd_sc_hd__buf_8 _09050_ (.A(_03708_),
    .X(_03714_));
 sky130_fd_sc_hd__nand2_1 _09051_ (.A(_03702_),
    .B(_01257_),
    .Y(_03715_));
 sky130_fd_sc_hd__nand2_2 _09052_ (.A(_03689_),
    .B(_01242_),
    .Y(_03716_));
 sky130_fd_sc_hd__buf_8 _09053_ (.A(_03716_),
    .X(_03717_));
 sky130_fd_sc_hd__o211a_1 _09054_ (.A1(_03714_),
    .A2(net727),
    .B1(_03715_),
    .C1(_03717_),
    .X(_00081_));
 sky130_fd_sc_hd__a21bo_1 _09055_ (.A1(_03704_),
    .A2(net394),
    .B1_N(_03715_),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _09056_ (.A0(net1289),
    .A1(_01201_),
    .S(_03708_),
    .X(_03718_));
 sky130_fd_sc_hd__clkbuf_1 _09057_ (.A(_03718_),
    .X(_00083_));
 sky130_fd_sc_hd__buf_6 _09058_ (.A(_02170_),
    .X(_03719_));
 sky130_fd_sc_hd__mux2_1 _09059_ (.A0(_01229_),
    .A1(\genblk2[0].wave_shpr.div.b1[8] ),
    .S(_03719_),
    .X(_03720_));
 sky130_fd_sc_hd__clkbuf_1 _09060_ (.A(_03720_),
    .X(_00084_));
 sky130_fd_sc_hd__inv_2 _09061_ (.A(_01193_),
    .Y(_03721_));
 sky130_fd_sc_hd__buf_4 _09062_ (.A(_03701_),
    .X(_03722_));
 sky130_fd_sc_hd__mux2_1 _09063_ (.A0(net1276),
    .A1(_03721_),
    .S(_03722_),
    .X(_03723_));
 sky130_fd_sc_hd__clkbuf_1 _09064_ (.A(_03723_),
    .X(_00085_));
 sky130_fd_sc_hd__mux2_1 _09065_ (.A0(net1184),
    .A1(_01185_),
    .S(_03722_),
    .X(_03724_));
 sky130_fd_sc_hd__clkbuf_1 _09066_ (.A(_03724_),
    .X(_00086_));
 sky130_fd_sc_hd__buf_2 _09067_ (.A(_02155_),
    .X(_03725_));
 sky130_fd_sc_hd__buf_8 _09068_ (.A(_03725_),
    .X(_03726_));
 sky130_fd_sc_hd__nand2_8 _09069_ (.A(_03701_),
    .B(_01221_),
    .Y(_03727_));
 sky130_fd_sc_hd__nand2_4 _09070_ (.A(_03702_),
    .B(_01996_),
    .Y(_03728_));
 sky130_fd_sc_hd__o221a_1 _09071_ (.A1(_03726_),
    .A2(net1084),
    .B1(_01302_),
    .B2(_03727_),
    .C1(_03728_),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _09072_ (.A0(\genblk2[0].wave_shpr.div.b1[12] ),
    .A1(_01340_),
    .S(_03722_),
    .X(_03729_));
 sky130_fd_sc_hd__clkbuf_1 _09073_ (.A(_03729_),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _09074_ (.A0(\genblk2[0].wave_shpr.div.b1[13] ),
    .A1(_01592_),
    .S(_03722_),
    .X(_03730_));
 sky130_fd_sc_hd__clkbuf_1 _09075_ (.A(_03730_),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _09076_ (.A0(net1291),
    .A1(_01483_),
    .S(_03722_),
    .X(_03731_));
 sky130_fd_sc_hd__clkbuf_1 _09077_ (.A(_03731_),
    .X(_00090_));
 sky130_fd_sc_hd__buf_8 _09078_ (.A(_03702_),
    .X(_03732_));
 sky130_fd_sc_hd__nand2_8 _09079_ (.A(_03708_),
    .B(_01210_),
    .Y(_03733_));
 sky130_fd_sc_hd__o21a_1 _09080_ (.A1(_03732_),
    .A2(net577),
    .B1(_03733_),
    .X(_00091_));
 sky130_fd_sc_hd__a21bo_1 _09081_ (.A1(_03704_),
    .A2(net396),
    .B1_N(_03717_),
    .X(_00092_));
 sky130_fd_sc_hd__inv_2 _09082_ (.A(net702),
    .Y(_03734_));
 sky130_fd_sc_hd__or3_4 _09083_ (.A(_02170_),
    .B(_01201_),
    .C(_01363_),
    .X(_03735_));
 sky130_fd_sc_hd__buf_8 _09084_ (.A(_03735_),
    .X(_03736_));
 sky130_fd_sc_hd__o21ai_1 _09085_ (.A1(_03714_),
    .A2(_03734_),
    .B1(_03736_),
    .Y(_00093_));
 sky130_fd_sc_hd__inv_2 _09086_ (.A(\modein.delay_octave_down_in[0] ),
    .Y(_03737_));
 sky130_fd_sc_hd__and2b_1 _09087_ (.A_N(\modein.delay_octave_up_in[1] ),
    .B(\modein.delay_octave_up_in[0] ),
    .X(_03738_));
 sky130_fd_sc_hd__o211a_1 _09088_ (.A1(_03737_),
    .A2(\modein.delay_octave_down_in[1] ),
    .B1(_01591_),
    .C1(_03738_),
    .X(_03739_));
 sky130_fd_sc_hd__or4_1 _09089_ (.A(_03737_),
    .B(\modein.delay_octave_down_in[1] ),
    .C(_01197_),
    .D(_03738_),
    .X(_03740_));
 sky130_fd_sc_hd__nor2b_1 _09090_ (.A(_03739_),
    .B_N(_03740_),
    .Y(_03741_));
 sky130_fd_sc_hd__xnor2_1 _09091_ (.A(_01201_),
    .B(_03741_),
    .Y(_00094_));
 sky130_fd_sc_hd__nor2_1 _09092_ (.A(_01367_),
    .B(_03740_),
    .Y(_03742_));
 sky130_fd_sc_hd__a221o_1 _09093_ (.A1(_01367_),
    .A2(_03739_),
    .B1(_03741_),
    .B2(_01342_),
    .C1(_03742_),
    .X(_00095_));
 sky130_fd_sc_hd__or2_1 _09094_ (.A(_01367_),
    .B(_03739_),
    .X(_03743_));
 sky130_fd_sc_hd__mux2_1 _09095_ (.A0(_01211_),
    .A1(_01556_),
    .S(_03743_),
    .X(_03744_));
 sky130_fd_sc_hd__mux2_1 _09096_ (.A0(_03744_),
    .A1(_01490_),
    .S(_03741_),
    .X(_03745_));
 sky130_fd_sc_hd__clkbuf_1 _09097_ (.A(_03745_),
    .X(_00096_));
 sky130_fd_sc_hd__or2_1 _09098_ (.A(_03734_),
    .B(\genblk2[0].wave_shpr.div.acc[17] ),
    .X(_03746_));
 sky130_fd_sc_hd__or2b_1 _09099_ (.A(\genblk2[0].wave_shpr.div.acc[16] ),
    .B_N(\genblk2[0].wave_shpr.div.b1[16] ),
    .X(_03747_));
 sky130_fd_sc_hd__or2b_1 _09100_ (.A(\genblk2[0].wave_shpr.div.acc[15] ),
    .B_N(\genblk2[0].wave_shpr.div.b1[15] ),
    .X(_03748_));
 sky130_fd_sc_hd__or2b_1 _09101_ (.A(\genblk2[0].wave_shpr.div.acc[14] ),
    .B_N(\genblk2[0].wave_shpr.div.b1[14] ),
    .X(_03749_));
 sky130_fd_sc_hd__or2b_1 _09102_ (.A(\genblk2[0].wave_shpr.div.acc[13] ),
    .B_N(\genblk2[0].wave_shpr.div.b1[13] ),
    .X(_03750_));
 sky130_fd_sc_hd__or2b_1 _09103_ (.A(\genblk2[0].wave_shpr.div.acc[12] ),
    .B_N(\genblk2[0].wave_shpr.div.b1[12] ),
    .X(_03751_));
 sky130_fd_sc_hd__or2b_1 _09104_ (.A(\genblk2[0].wave_shpr.div.acc[11] ),
    .B_N(\genblk2[0].wave_shpr.div.b1[11] ),
    .X(_03752_));
 sky130_fd_sc_hd__or2b_1 _09105_ (.A(\genblk2[0].wave_shpr.div.acc[10] ),
    .B_N(\genblk2[0].wave_shpr.div.b1[10] ),
    .X(_03753_));
 sky130_fd_sc_hd__or2b_1 _09106_ (.A(\genblk2[0].wave_shpr.div.acc[9] ),
    .B_N(\genblk2[0].wave_shpr.div.b1[9] ),
    .X(_03754_));
 sky130_fd_sc_hd__or2b_1 _09107_ (.A(\genblk2[0].wave_shpr.div.acc[8] ),
    .B_N(\genblk2[0].wave_shpr.div.b1[8] ),
    .X(_03755_));
 sky130_fd_sc_hd__or2b_1 _09108_ (.A(\genblk2[0].wave_shpr.div.acc[7] ),
    .B_N(\genblk2[0].wave_shpr.div.b1[7] ),
    .X(_03756_));
 sky130_fd_sc_hd__or2b_1 _09109_ (.A(\genblk2[0].wave_shpr.div.acc[6] ),
    .B_N(\genblk2[0].wave_shpr.div.b1[6] ),
    .X(_03757_));
 sky130_fd_sc_hd__or2b_1 _09110_ (.A(\genblk2[0].wave_shpr.div.acc[5] ),
    .B_N(\genblk2[0].wave_shpr.div.b1[5] ),
    .X(_03758_));
 sky130_fd_sc_hd__or2b_1 _09111_ (.A(\genblk2[0].wave_shpr.div.acc[4] ),
    .B_N(\genblk2[0].wave_shpr.div.b1[4] ),
    .X(_03759_));
 sky130_fd_sc_hd__or2b_1 _09112_ (.A(\genblk2[0].wave_shpr.div.acc[3] ),
    .B_N(\genblk2[0].wave_shpr.div.b1[3] ),
    .X(_03760_));
 sky130_fd_sc_hd__inv_2 _09113_ (.A(\genblk2[0].wave_shpr.div.b1[2] ),
    .Y(_03761_));
 sky130_fd_sc_hd__or2b_1 _09114_ (.A(\genblk2[0].wave_shpr.div.b1[1] ),
    .B_N(\genblk2[0].wave_shpr.div.acc[1] ),
    .X(_03762_));
 sky130_fd_sc_hd__or2b_1 _09115_ (.A(\genblk2[0].wave_shpr.div.acc[1] ),
    .B_N(\genblk2[0].wave_shpr.div.b1[1] ),
    .X(_03763_));
 sky130_fd_sc_hd__nand2_1 _09116_ (.A(_03762_),
    .B(_03763_),
    .Y(_03764_));
 sky130_fd_sc_hd__and2b_1 _09117_ (.A_N(\genblk2[0].wave_shpr.div.acc[0] ),
    .B(\genblk2[0].wave_shpr.div.b1[0] ),
    .X(_03765_));
 sky130_fd_sc_hd__o21ai_1 _09118_ (.A1(_03764_),
    .A2(_03765_),
    .B1(_03762_),
    .Y(_03766_));
 sky130_fd_sc_hd__o21a_1 _09119_ (.A1(_03761_),
    .A2(\genblk2[0].wave_shpr.div.acc[2] ),
    .B1(_03766_),
    .X(_03767_));
 sky130_fd_sc_hd__a21o_1 _09120_ (.A1(_03761_),
    .A2(\genblk2[0].wave_shpr.div.acc[2] ),
    .B1(_03767_),
    .X(_03768_));
 sky130_fd_sc_hd__and2b_1 _09121_ (.A_N(\genblk2[0].wave_shpr.div.b1[3] ),
    .B(\genblk2[0].wave_shpr.div.acc[3] ),
    .X(_03769_));
 sky130_fd_sc_hd__a21o_1 _09122_ (.A1(_03760_),
    .A2(_03768_),
    .B1(_03769_),
    .X(_03770_));
 sky130_fd_sc_hd__and2b_1 _09123_ (.A_N(\genblk2[0].wave_shpr.div.b1[4] ),
    .B(\genblk2[0].wave_shpr.div.acc[4] ),
    .X(_03771_));
 sky130_fd_sc_hd__a21o_1 _09124_ (.A1(_03759_),
    .A2(_03770_),
    .B1(_03771_),
    .X(_03772_));
 sky130_fd_sc_hd__and2b_1 _09125_ (.A_N(\genblk2[0].wave_shpr.div.b1[5] ),
    .B(\genblk2[0].wave_shpr.div.acc[5] ),
    .X(_03773_));
 sky130_fd_sc_hd__a21o_1 _09126_ (.A1(_03758_),
    .A2(_03772_),
    .B1(_03773_),
    .X(_03774_));
 sky130_fd_sc_hd__and2b_1 _09127_ (.A_N(\genblk2[0].wave_shpr.div.b1[6] ),
    .B(\genblk2[0].wave_shpr.div.acc[6] ),
    .X(_03775_));
 sky130_fd_sc_hd__a21o_1 _09128_ (.A1(_03757_),
    .A2(_03774_),
    .B1(_03775_),
    .X(_03776_));
 sky130_fd_sc_hd__and2b_1 _09129_ (.A_N(\genblk2[0].wave_shpr.div.b1[7] ),
    .B(\genblk2[0].wave_shpr.div.acc[7] ),
    .X(_03777_));
 sky130_fd_sc_hd__a21o_1 _09130_ (.A1(_03756_),
    .A2(_03776_),
    .B1(_03777_),
    .X(_03778_));
 sky130_fd_sc_hd__and2b_1 _09131_ (.A_N(\genblk2[0].wave_shpr.div.b1[8] ),
    .B(\genblk2[0].wave_shpr.div.acc[8] ),
    .X(_03779_));
 sky130_fd_sc_hd__a21o_1 _09132_ (.A1(_03755_),
    .A2(_03778_),
    .B1(_03779_),
    .X(_03780_));
 sky130_fd_sc_hd__and2b_1 _09133_ (.A_N(\genblk2[0].wave_shpr.div.b1[9] ),
    .B(\genblk2[0].wave_shpr.div.acc[9] ),
    .X(_03781_));
 sky130_fd_sc_hd__a21o_1 _09134_ (.A1(_03754_),
    .A2(_03780_),
    .B1(_03781_),
    .X(_03782_));
 sky130_fd_sc_hd__and2b_1 _09135_ (.A_N(\genblk2[0].wave_shpr.div.b1[10] ),
    .B(\genblk2[0].wave_shpr.div.acc[10] ),
    .X(_03783_));
 sky130_fd_sc_hd__a21o_1 _09136_ (.A1(_03753_),
    .A2(_03782_),
    .B1(_03783_),
    .X(_03784_));
 sky130_fd_sc_hd__and2b_1 _09137_ (.A_N(\genblk2[0].wave_shpr.div.b1[11] ),
    .B(\genblk2[0].wave_shpr.div.acc[11] ),
    .X(_03785_));
 sky130_fd_sc_hd__a21o_1 _09138_ (.A1(_03752_),
    .A2(_03784_),
    .B1(_03785_),
    .X(_03786_));
 sky130_fd_sc_hd__and2b_1 _09139_ (.A_N(\genblk2[0].wave_shpr.div.b1[12] ),
    .B(\genblk2[0].wave_shpr.div.acc[12] ),
    .X(_03787_));
 sky130_fd_sc_hd__a21o_1 _09140_ (.A1(_03751_),
    .A2(_03786_),
    .B1(_03787_),
    .X(_03788_));
 sky130_fd_sc_hd__and2b_1 _09141_ (.A_N(\genblk2[0].wave_shpr.div.b1[13] ),
    .B(\genblk2[0].wave_shpr.div.acc[13] ),
    .X(_03789_));
 sky130_fd_sc_hd__a21o_1 _09142_ (.A1(_03750_),
    .A2(_03788_),
    .B1(_03789_),
    .X(_03790_));
 sky130_fd_sc_hd__and2b_1 _09143_ (.A_N(\genblk2[0].wave_shpr.div.b1[14] ),
    .B(\genblk2[0].wave_shpr.div.acc[14] ),
    .X(_03791_));
 sky130_fd_sc_hd__a21o_1 _09144_ (.A1(_03749_),
    .A2(_03790_),
    .B1(_03791_),
    .X(_03792_));
 sky130_fd_sc_hd__and2b_1 _09145_ (.A_N(\genblk2[0].wave_shpr.div.b1[15] ),
    .B(\genblk2[0].wave_shpr.div.acc[15] ),
    .X(_03793_));
 sky130_fd_sc_hd__a21o_1 _09146_ (.A1(_03748_),
    .A2(_03792_),
    .B1(_03793_),
    .X(_03794_));
 sky130_fd_sc_hd__and2b_1 _09147_ (.A_N(\genblk2[0].wave_shpr.div.b1[16] ),
    .B(\genblk2[0].wave_shpr.div.acc[16] ),
    .X(_03795_));
 sky130_fd_sc_hd__a21o_1 _09148_ (.A1(_03747_),
    .A2(_03794_),
    .B1(_03795_),
    .X(_03796_));
 sky130_fd_sc_hd__and2_1 _09149_ (.A(_03734_),
    .B(\genblk2[0].wave_shpr.div.acc[17] ),
    .X(_03797_));
 sky130_fd_sc_hd__a21o_1 _09150_ (.A1(_03746_),
    .A2(_03796_),
    .B1(_03797_),
    .X(_03798_));
 sky130_fd_sc_hd__or2_1 _09151_ (.A(\genblk2[0].wave_shpr.div.acc[18] ),
    .B(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__or2_1 _09152_ (.A(\genblk2[0].wave_shpr.div.acc[19] ),
    .B(_03799_),
    .X(_03800_));
 sky130_fd_sc_hd__or4_1 _09153_ (.A(\genblk2[0].wave_shpr.div.acc[22] ),
    .B(\genblk2[0].wave_shpr.div.acc[21] ),
    .C(\genblk2[0].wave_shpr.div.acc[20] ),
    .D(_03800_),
    .X(_03801_));
 sky130_fd_sc_hd__or2_2 _09154_ (.A(\genblk2[0].wave_shpr.div.acc[23] ),
    .B(_03801_),
    .X(_03802_));
 sky130_fd_sc_hd__or4_2 _09155_ (.A(\genblk2[0].wave_shpr.div.acc[25] ),
    .B(\genblk2[0].wave_shpr.div.acc[24] ),
    .C(\genblk2[0].wave_shpr.div.acc[26] ),
    .D(_03802_),
    .X(_03803_));
 sky130_fd_sc_hd__buf_4 _09156_ (.A(_03803_),
    .X(_03804_));
 sky130_fd_sc_hd__mux2_1 _09157_ (.A0(\genblk2[0].wave_shpr.div.fin_quo[0] ),
    .A1(_03804_),
    .S(_00001_),
    .X(_03805_));
 sky130_fd_sc_hd__clkbuf_1 _09158_ (.A(_03805_),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _09159_ (.A0(\genblk2[0].wave_shpr.div.fin_quo[1] ),
    .A1(\genblk2[0].wave_shpr.div.quo[0] ),
    .S(_00001_),
    .X(_03806_));
 sky130_fd_sc_hd__clkbuf_1 _09160_ (.A(_03806_),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _09161_ (.A0(\genblk2[0].wave_shpr.div.fin_quo[2] ),
    .A1(net1322),
    .S(_00001_),
    .X(_03807_));
 sky130_fd_sc_hd__clkbuf_1 _09162_ (.A(_03807_),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _09163_ (.A0(\genblk2[0].wave_shpr.div.fin_quo[3] ),
    .A1(net1314),
    .S(_00001_),
    .X(_03808_));
 sky130_fd_sc_hd__clkbuf_1 _09164_ (.A(_03808_),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _09165_ (.A0(\genblk2[0].wave_shpr.div.fin_quo[4] ),
    .A1(\genblk2[0].wave_shpr.div.quo[3] ),
    .S(_00001_),
    .X(_03809_));
 sky130_fd_sc_hd__clkbuf_1 _09166_ (.A(_03809_),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _09167_ (.A0(\genblk2[0].wave_shpr.div.fin_quo[5] ),
    .A1(net1334),
    .S(_00001_),
    .X(_03810_));
 sky130_fd_sc_hd__clkbuf_1 _09168_ (.A(_03810_),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_1 _09169_ (.A0(\genblk2[0].wave_shpr.div.fin_quo[6] ),
    .A1(net652),
    .S(_00001_),
    .X(_03811_));
 sky130_fd_sc_hd__clkbuf_1 _09170_ (.A(_03811_),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _09171_ (.A0(net1218),
    .A1(\genblk2[0].wave_shpr.div.quo[6] ),
    .S(_00001_),
    .X(_03812_));
 sky130_fd_sc_hd__clkbuf_1 _09172_ (.A(net1219),
    .X(_00104_));
 sky130_fd_sc_hd__nor2_2 _09173_ (.A(_01342_),
    .B(_01441_),
    .Y(_03813_));
 sky130_fd_sc_hd__mux2_1 _09174_ (.A0(\genblk2[10].wave_shpr.div.b1[0] ),
    .A1(_03813_),
    .S(_03722_),
    .X(_03814_));
 sky130_fd_sc_hd__clkbuf_1 _09175_ (.A(_03814_),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_1 _09176_ (.A0(\genblk2[10].wave_shpr.div.b1[1] ),
    .A1(_01368_),
    .S(_03722_),
    .X(_03815_));
 sky130_fd_sc_hd__clkbuf_1 _09177_ (.A(_03815_),
    .X(_00106_));
 sky130_fd_sc_hd__mux2_1 _09178_ (.A0(net1171),
    .A1(_01342_),
    .S(_03722_),
    .X(_03816_));
 sky130_fd_sc_hd__clkbuf_1 _09179_ (.A(_03816_),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _09180_ (.A0(net1249),
    .A1(_01356_),
    .S(_03722_),
    .X(_03817_));
 sky130_fd_sc_hd__clkbuf_1 _09181_ (.A(_03817_),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _09182_ (.A0(net1273),
    .A1(_01214_),
    .S(_03722_),
    .X(_03818_));
 sky130_fd_sc_hd__clkbuf_1 _09183_ (.A(_03818_),
    .X(_00109_));
 sky130_fd_sc_hd__clkbuf_8 _09184_ (.A(_03719_),
    .X(_03819_));
 sky130_fd_sc_hd__a21oi_1 _09185_ (.A1(_01430_),
    .A2(_01344_),
    .B1(_03819_),
    .Y(_03820_));
 sky130_fd_sc_hd__a21o_1 _09186_ (.A1(_03704_),
    .A2(net651),
    .B1(_03820_),
    .X(_00110_));
 sky130_fd_sc_hd__inv_2 _09187_ (.A(net1173),
    .Y(_03821_));
 sky130_fd_sc_hd__o21ai_1 _09188_ (.A1(_03714_),
    .A2(_03821_),
    .B1(_03705_),
    .Y(_00111_));
 sky130_fd_sc_hd__clkbuf_8 _09189_ (.A(_03701_),
    .X(_03822_));
 sky130_fd_sc_hd__mux2_1 _09190_ (.A0(net1254),
    .A1(_03706_),
    .S(_03822_),
    .X(_03823_));
 sky130_fd_sc_hd__clkbuf_1 _09191_ (.A(_03823_),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _09192_ (.A0(net1244),
    .A1(_02002_),
    .S(_03822_),
    .X(_03824_));
 sky130_fd_sc_hd__clkbuf_1 _09193_ (.A(_03824_),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _09194_ (.A0(net1284),
    .A1(_01991_),
    .S(_03822_),
    .X(_03825_));
 sky130_fd_sc_hd__clkbuf_1 _09195_ (.A(_03825_),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _09196_ (.A0(net1224),
    .A1(_03712_),
    .S(_03822_),
    .X(_03826_));
 sky130_fd_sc_hd__clkbuf_1 _09197_ (.A(_03826_),
    .X(_00115_));
 sky130_fd_sc_hd__inv_2 _09198_ (.A(_02005_),
    .Y(_03827_));
 sky130_fd_sc_hd__mux2_1 _09199_ (.A0(net1292),
    .A1(_03827_),
    .S(_03822_),
    .X(_03828_));
 sky130_fd_sc_hd__clkbuf_1 _09200_ (.A(_03828_),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _09201_ (.A0(net1199),
    .A1(_01183_),
    .S(_03822_),
    .X(_03829_));
 sky130_fd_sc_hd__clkbuf_1 _09202_ (.A(_03829_),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_1 _09203_ (.A0(net1251),
    .A1(_01302_),
    .S(_03822_),
    .X(_03830_));
 sky130_fd_sc_hd__clkbuf_1 _09204_ (.A(_03830_),
    .X(_00118_));
 sky130_fd_sc_hd__a21bo_1 _09205_ (.A1(_03704_),
    .A2(net759),
    .B1_N(_03728_),
    .X(_00119_));
 sky130_fd_sc_hd__buf_8 _09206_ (.A(_02171_),
    .X(_03831_));
 sky130_fd_sc_hd__a21bo_1 _09207_ (.A1(_03831_),
    .A2(net674),
    .B1_N(_03717_),
    .X(_00120_));
 sky130_fd_sc_hd__inv_2 _09208_ (.A(net959),
    .Y(_03832_));
 sky130_fd_sc_hd__o21ai_1 _09209_ (.A1(_03714_),
    .A2(_03832_),
    .B1(_03736_),
    .Y(_00121_));
 sky130_fd_sc_hd__clkbuf_8 _09210_ (.A(_02170_),
    .X(_03833_));
 sky130_fd_sc_hd__and2_1 _09211_ (.A(_03833_),
    .B(net1302),
    .X(_03834_));
 sky130_fd_sc_hd__clkbuf_1 _09212_ (.A(_03834_),
    .X(_00122_));
 sky130_fd_sc_hd__buf_2 _09213_ (.A(_02151_),
    .X(_03835_));
 sky130_fd_sc_hd__clkbuf_4 _09214_ (.A(_03835_),
    .X(_03836_));
 sky130_fd_sc_hd__and3_1 _09215_ (.A(_02152_),
    .B(\genblk2[0].wave_shpr.div.busy ),
    .C(_02149_),
    .X(_03837_));
 sky130_fd_sc_hd__clkbuf_4 _09216_ (.A(_03837_),
    .X(_03838_));
 sky130_fd_sc_hd__clkbuf_4 _09217_ (.A(_03838_),
    .X(_03839_));
 sky130_fd_sc_hd__a22o_1 _09218_ (.A1(net804),
    .A2(_03836_),
    .B1(_03804_),
    .B2(_03839_),
    .X(_00123_));
 sky130_fd_sc_hd__clkbuf_4 _09219_ (.A(_03838_),
    .X(_03840_));
 sky130_fd_sc_hd__a22o_1 _09220_ (.A1(net655),
    .A2(_03836_),
    .B1(_03840_),
    .B2(net804),
    .X(_00124_));
 sky130_fd_sc_hd__a22o_1 _09221_ (.A1(net558),
    .A2(_03836_),
    .B1(_03840_),
    .B2(net655),
    .X(_00125_));
 sky130_fd_sc_hd__a22o_1 _09222_ (.A1(\genblk2[0].wave_shpr.div.quo[3] ),
    .A2(_03836_),
    .B1(_03840_),
    .B2(net558),
    .X(_00126_));
 sky130_fd_sc_hd__a22o_1 _09223_ (.A1(net600),
    .A2(_03836_),
    .B1(_03840_),
    .B2(net728),
    .X(_00127_));
 sky130_fd_sc_hd__a22o_1 _09224_ (.A1(\genblk2[0].wave_shpr.div.quo[5] ),
    .A2(_03836_),
    .B1(_03840_),
    .B2(net600),
    .X(_00128_));
 sky130_fd_sc_hd__a22o_1 _09225_ (.A1(net269),
    .A2(_03836_),
    .B1(_03840_),
    .B2(net652),
    .X(_00129_));
 sky130_fd_sc_hd__a22o_1 _09226_ (.A1(\genblk2[0].wave_shpr.div.quo[7] ),
    .A2(_03836_),
    .B1(_03840_),
    .B2(net269),
    .X(_00130_));
 sky130_fd_sc_hd__a22o_1 _09227_ (.A1(net277),
    .A2(_03836_),
    .B1(_03840_),
    .B2(net379),
    .X(_00131_));
 sky130_fd_sc_hd__clkbuf_4 _09228_ (.A(_03835_),
    .X(_03841_));
 sky130_fd_sc_hd__and2_1 _09229_ (.A(_03725_),
    .B(\genblk1[0].osc.clkdiv_C.cnt[0] ),
    .X(_03842_));
 sky130_fd_sc_hd__a221o_1 _09230_ (.A1(\genblk2[0].wave_shpr.div.quo[9] ),
    .A2(_03841_),
    .B1(_03839_),
    .B2(net277),
    .C1(_03842_),
    .X(_00132_));
 sky130_fd_sc_hd__and2_1 _09231_ (.A(_03725_),
    .B(\genblk1[0].osc.clkdiv_C.cnt[1] ),
    .X(_03843_));
 sky130_fd_sc_hd__a221o_1 _09232_ (.A1(net569),
    .A2(_03841_),
    .B1(_03839_),
    .B2(net598),
    .C1(_03843_),
    .X(_00133_));
 sky130_fd_sc_hd__and2_1 _09233_ (.A(_03725_),
    .B(\genblk1[0].osc.clkdiv_C.cnt[2] ),
    .X(_03844_));
 sky130_fd_sc_hd__a221o_1 _09234_ (.A1(\genblk2[0].wave_shpr.div.quo[11] ),
    .A2(_03841_),
    .B1(_03839_),
    .B2(net569),
    .C1(_03844_),
    .X(_00134_));
 sky130_fd_sc_hd__clkbuf_4 _09235_ (.A(_03835_),
    .X(_03845_));
 sky130_fd_sc_hd__and2_1 _09236_ (.A(_03725_),
    .B(\genblk1[0].osc.clkdiv_C.cnt[3] ),
    .X(_03846_));
 sky130_fd_sc_hd__a221o_1 _09237_ (.A1(net584),
    .A2(_03845_),
    .B1(_03839_),
    .B2(net599),
    .C1(_03846_),
    .X(_00135_));
 sky130_fd_sc_hd__buf_2 _09238_ (.A(_03838_),
    .X(_03847_));
 sky130_fd_sc_hd__and2_1 _09239_ (.A(_03725_),
    .B(\genblk1[0].osc.clkdiv_C.cnt[4] ),
    .X(_03848_));
 sky130_fd_sc_hd__a221o_1 _09240_ (.A1(net495),
    .A2(_03845_),
    .B1(_03847_),
    .B2(net584),
    .C1(_03848_),
    .X(_00136_));
 sky130_fd_sc_hd__and2_1 _09241_ (.A(_03725_),
    .B(\genblk1[0].osc.clkdiv_C.cnt[5] ),
    .X(_03849_));
 sky130_fd_sc_hd__a221o_1 _09242_ (.A1(\genblk2[0].wave_shpr.div.quo[14] ),
    .A2(_03845_),
    .B1(_03847_),
    .B2(net495),
    .C1(_03849_),
    .X(_00137_));
 sky130_fd_sc_hd__and2_1 _09243_ (.A(_03725_),
    .B(\genblk1[0].osc.clkdiv_C.cnt[6] ),
    .X(_03850_));
 sky130_fd_sc_hd__a221o_1 _09244_ (.A1(net543),
    .A2(_03845_),
    .B1(_03847_),
    .B2(\genblk2[0].wave_shpr.div.quo[14] ),
    .C1(_03850_),
    .X(_00138_));
 sky130_fd_sc_hd__and2_1 _09245_ (.A(_03725_),
    .B(\genblk1[0].osc.clkdiv_C.cnt[7] ),
    .X(_03851_));
 sky130_fd_sc_hd__a221o_1 _09246_ (.A1(net522),
    .A2(_03845_),
    .B1(_03847_),
    .B2(net543),
    .C1(_03851_),
    .X(_00139_));
 sky130_fd_sc_hd__and2_1 _09247_ (.A(_03725_),
    .B(\genblk1[0].osc.clkdiv_C.cnt[8] ),
    .X(_03852_));
 sky130_fd_sc_hd__a221o_1 _09248_ (.A1(net410),
    .A2(_03845_),
    .B1(_03847_),
    .B2(net522),
    .C1(_03852_),
    .X(_00140_));
 sky130_fd_sc_hd__clkbuf_4 _09249_ (.A(_03707_),
    .X(_03853_));
 sky130_fd_sc_hd__and2_1 _09250_ (.A(_03853_),
    .B(\genblk1[0].osc.clkdiv_C.cnt[9] ),
    .X(_03854_));
 sky130_fd_sc_hd__a221o_1 _09251_ (.A1(\genblk2[0].wave_shpr.div.quo[18] ),
    .A2(_03845_),
    .B1(_03847_),
    .B2(net410),
    .C1(_03854_),
    .X(_00141_));
 sky130_fd_sc_hd__buf_6 _09252_ (.A(_03719_),
    .X(_03855_));
 sky130_fd_sc_hd__nor2_1 _09253_ (.A(_03855_),
    .B(_01169_),
    .Y(_03856_));
 sky130_fd_sc_hd__a221o_1 _09254_ (.A1(net298),
    .A2(_03845_),
    .B1(_03847_),
    .B2(net466),
    .C1(_03856_),
    .X(_00142_));
 sky130_fd_sc_hd__and2_1 _09255_ (.A(_03853_),
    .B(\genblk1[0].osc.clkdiv_C.cnt[11] ),
    .X(_03857_));
 sky130_fd_sc_hd__a221o_1 _09256_ (.A1(\genblk2[0].wave_shpr.div.quo[20] ),
    .A2(_03845_),
    .B1(_03847_),
    .B2(net298),
    .C1(_03857_),
    .X(_00143_));
 sky130_fd_sc_hd__and2_1 _09257_ (.A(_03853_),
    .B(\genblk1[0].osc.clkdiv_C.cnt[12] ),
    .X(_03858_));
 sky130_fd_sc_hd__a221o_1 _09258_ (.A1(net265),
    .A2(_03845_),
    .B1(_03847_),
    .B2(net636),
    .C1(_03858_),
    .X(_00144_));
 sky130_fd_sc_hd__and2_1 _09259_ (.A(_03853_),
    .B(\genblk1[0].osc.clkdiv_C.cnt[13] ),
    .X(_03859_));
 sky130_fd_sc_hd__a221o_1 _09260_ (.A1(\genblk2[0].wave_shpr.div.quo[22] ),
    .A2(_03835_),
    .B1(_03847_),
    .B2(net265),
    .C1(_03859_),
    .X(_00145_));
 sky130_fd_sc_hd__and2_1 _09261_ (.A(_03853_),
    .B(\genblk1[0].osc.clkdiv_C.cnt[14] ),
    .X(_03860_));
 sky130_fd_sc_hd__a221o_1 _09262_ (.A1(net454),
    .A2(_03835_),
    .B1(_03838_),
    .B2(net476),
    .C1(_03860_),
    .X(_00146_));
 sky130_fd_sc_hd__and2_1 _09263_ (.A(_03853_),
    .B(\genblk1[0].osc.clkdiv_C.cnt[15] ),
    .X(_03861_));
 sky130_fd_sc_hd__a221o_1 _09264_ (.A1(\genblk2[0].wave_shpr.div.quo[24] ),
    .A2(_03835_),
    .B1(_03838_),
    .B2(net454),
    .C1(_03861_),
    .X(_00147_));
 sky130_fd_sc_hd__and2_1 _09265_ (.A(_03853_),
    .B(\genblk1[0].osc.clkdiv_C.cnt[16] ),
    .X(_03862_));
 sky130_fd_sc_hd__a221o_1 _09266_ (.A1(net578),
    .A2(_03835_),
    .B1(_03838_),
    .B2(\genblk2[0].wave_shpr.div.quo[24] ),
    .C1(_03862_),
    .X(_00148_));
 sky130_fd_sc_hd__inv_2 _09267_ (.A(_03838_),
    .Y(_03863_));
 sky130_fd_sc_hd__or2_1 _09268_ (.A(_02171_),
    .B(\genblk1[0].osc.clkdiv_C.cnt[17] ),
    .X(_03864_));
 sky130_fd_sc_hd__o221a_1 _09269_ (.A1(net715),
    .A2(_00000_),
    .B1(_03863_),
    .B2(net578),
    .C1(_03864_),
    .X(_00149_));
 sky130_fd_sc_hd__a21oi_1 _09270_ (.A1(\genblk2[0].wave_shpr.div.b1[0] ),
    .A2(_03804_),
    .B1(\genblk2[0].wave_shpr.div.acc[0] ),
    .Y(_03865_));
 sky130_fd_sc_hd__a31o_1 _09271_ (.A1(\genblk2[0].wave_shpr.div.b1[0] ),
    .A2(\genblk2[0].wave_shpr.div.acc[0] ),
    .A3(_03804_),
    .B1(_03863_),
    .X(_03866_));
 sky130_fd_sc_hd__a2bb2o_1 _09272_ (.A1_N(_03865_),
    .A2_N(_03866_),
    .B1(net1066),
    .B2(_03836_),
    .X(_00150_));
 sky130_fd_sc_hd__or2_1 _09273_ (.A(\genblk2[0].wave_shpr.div.acc[1] ),
    .B(_03803_),
    .X(_03867_));
 sky130_fd_sc_hd__xnor2_1 _09274_ (.A(_03764_),
    .B(_03765_),
    .Y(_03868_));
 sky130_fd_sc_hd__nand2_1 _09275_ (.A(_03804_),
    .B(_03868_),
    .Y(_03869_));
 sky130_fd_sc_hd__a32o_1 _09276_ (.A1(_03839_),
    .A2(_03867_),
    .A3(_03869_),
    .B1(_03841_),
    .B2(net1139),
    .X(_00151_));
 sky130_fd_sc_hd__clkbuf_4 _09277_ (.A(_03835_),
    .X(_03870_));
 sky130_fd_sc_hd__xor2_1 _09278_ (.A(\genblk2[0].wave_shpr.div.b1[2] ),
    .B(\genblk2[0].wave_shpr.div.acc[2] ),
    .X(_03871_));
 sky130_fd_sc_hd__xnor2_1 _09279_ (.A(_03766_),
    .B(_03871_),
    .Y(_03872_));
 sky130_fd_sc_hd__mux2_1 _09280_ (.A0(\genblk2[0].wave_shpr.div.acc[2] ),
    .A1(_03872_),
    .S(_03804_),
    .X(_03873_));
 sky130_fd_sc_hd__a22o_1 _09281_ (.A1(net854),
    .A2(_03870_),
    .B1(_03840_),
    .B2(_03873_),
    .X(_00152_));
 sky130_fd_sc_hd__or2b_1 _09282_ (.A(_03769_),
    .B_N(_03760_),
    .X(_03874_));
 sky130_fd_sc_hd__xnor2_1 _09283_ (.A(_03768_),
    .B(_03874_),
    .Y(_03875_));
 sky130_fd_sc_hd__mux2_1 _09284_ (.A0(\genblk2[0].wave_shpr.div.acc[3] ),
    .A1(_03875_),
    .S(_03804_),
    .X(_03876_));
 sky130_fd_sc_hd__a22o_1 _09285_ (.A1(net1033),
    .A2(_03870_),
    .B1(_03840_),
    .B2(_03876_),
    .X(_00153_));
 sky130_fd_sc_hd__clkbuf_4 _09286_ (.A(_03838_),
    .X(_03877_));
 sky130_fd_sc_hd__or2b_1 _09287_ (.A(_03771_),
    .B_N(_03759_),
    .X(_03878_));
 sky130_fd_sc_hd__xnor2_1 _09288_ (.A(_03878_),
    .B(_03770_),
    .Y(_03879_));
 sky130_fd_sc_hd__mux2_1 _09289_ (.A0(\genblk2[0].wave_shpr.div.acc[4] ),
    .A1(_03879_),
    .S(_03804_),
    .X(_03880_));
 sky130_fd_sc_hd__a22o_1 _09290_ (.A1(net823),
    .A2(_03870_),
    .B1(_03877_),
    .B2(_03880_),
    .X(_00154_));
 sky130_fd_sc_hd__or2b_1 _09291_ (.A(_03773_),
    .B_N(_03758_),
    .X(_03881_));
 sky130_fd_sc_hd__xnor2_1 _09292_ (.A(_03881_),
    .B(_03772_),
    .Y(_03882_));
 sky130_fd_sc_hd__mux2_1 _09293_ (.A0(\genblk2[0].wave_shpr.div.acc[5] ),
    .A1(_03882_),
    .S(_03804_),
    .X(_03883_));
 sky130_fd_sc_hd__a22o_1 _09294_ (.A1(net866),
    .A2(_03870_),
    .B1(_03877_),
    .B2(_03883_),
    .X(_00155_));
 sky130_fd_sc_hd__or2b_1 _09295_ (.A(_03775_),
    .B_N(_03757_),
    .X(_03884_));
 sky130_fd_sc_hd__xnor2_1 _09296_ (.A(_03774_),
    .B(_03884_),
    .Y(_03885_));
 sky130_fd_sc_hd__mux2_1 _09297_ (.A0(\genblk2[0].wave_shpr.div.acc[6] ),
    .A1(_03885_),
    .S(_03804_),
    .X(_03886_));
 sky130_fd_sc_hd__a22o_1 _09298_ (.A1(net964),
    .A2(_03870_),
    .B1(_03877_),
    .B2(_03886_),
    .X(_00156_));
 sky130_fd_sc_hd__or2b_1 _09299_ (.A(_03777_),
    .B_N(_03756_),
    .X(_03887_));
 sky130_fd_sc_hd__xnor2_1 _09300_ (.A(_03776_),
    .B(_03887_),
    .Y(_03888_));
 sky130_fd_sc_hd__buf_4 _09301_ (.A(_03803_),
    .X(_03889_));
 sky130_fd_sc_hd__mux2_1 _09302_ (.A0(\genblk2[0].wave_shpr.div.acc[7] ),
    .A1(_03888_),
    .S(_03889_),
    .X(_03890_));
 sky130_fd_sc_hd__a22o_1 _09303_ (.A1(net1049),
    .A2(_03870_),
    .B1(_03877_),
    .B2(_03890_),
    .X(_00157_));
 sky130_fd_sc_hd__or2b_1 _09304_ (.A(_03779_),
    .B_N(_03755_),
    .X(_03891_));
 sky130_fd_sc_hd__xnor2_1 _09305_ (.A(_03778_),
    .B(_03891_),
    .Y(_03892_));
 sky130_fd_sc_hd__mux2_1 _09306_ (.A0(\genblk2[0].wave_shpr.div.acc[8] ),
    .A1(_03892_),
    .S(_03889_),
    .X(_03893_));
 sky130_fd_sc_hd__a22o_1 _09307_ (.A1(net956),
    .A2(_03870_),
    .B1(_03877_),
    .B2(_03893_),
    .X(_00158_));
 sky130_fd_sc_hd__or2b_1 _09308_ (.A(_03781_),
    .B_N(_03754_),
    .X(_03894_));
 sky130_fd_sc_hd__xnor2_1 _09309_ (.A(_03780_),
    .B(_03894_),
    .Y(_03895_));
 sky130_fd_sc_hd__mux2_1 _09310_ (.A0(\genblk2[0].wave_shpr.div.acc[9] ),
    .A1(_03895_),
    .S(_03889_),
    .X(_03896_));
 sky130_fd_sc_hd__a22o_1 _09311_ (.A1(net934),
    .A2(_03870_),
    .B1(_03877_),
    .B2(_03896_),
    .X(_00159_));
 sky130_fd_sc_hd__or2b_1 _09312_ (.A(_03783_),
    .B_N(_03753_),
    .X(_03897_));
 sky130_fd_sc_hd__xnor2_1 _09313_ (.A(_03782_),
    .B(_03897_),
    .Y(_03898_));
 sky130_fd_sc_hd__mux2_1 _09314_ (.A0(\genblk2[0].wave_shpr.div.acc[10] ),
    .A1(_03898_),
    .S(_03889_),
    .X(_03899_));
 sky130_fd_sc_hd__a22o_1 _09315_ (.A1(net1004),
    .A2(_03870_),
    .B1(_03877_),
    .B2(_03899_),
    .X(_00160_));
 sky130_fd_sc_hd__or2b_1 _09316_ (.A(_03785_),
    .B_N(_03752_),
    .X(_03900_));
 sky130_fd_sc_hd__xnor2_1 _09317_ (.A(_03784_),
    .B(_03900_),
    .Y(_03901_));
 sky130_fd_sc_hd__mux2_1 _09318_ (.A0(\genblk2[0].wave_shpr.div.acc[11] ),
    .A1(_03901_),
    .S(_03889_),
    .X(_03902_));
 sky130_fd_sc_hd__a22o_1 _09319_ (.A1(net889),
    .A2(_03870_),
    .B1(_03877_),
    .B2(_03902_),
    .X(_00161_));
 sky130_fd_sc_hd__clkbuf_4 _09320_ (.A(_03835_),
    .X(_03903_));
 sky130_fd_sc_hd__or2b_1 _09321_ (.A(_03787_),
    .B_N(_03751_),
    .X(_03904_));
 sky130_fd_sc_hd__xnor2_1 _09322_ (.A(_03786_),
    .B(_03904_),
    .Y(_03905_));
 sky130_fd_sc_hd__mux2_1 _09323_ (.A0(\genblk2[0].wave_shpr.div.acc[12] ),
    .A1(_03905_),
    .S(_03889_),
    .X(_03906_));
 sky130_fd_sc_hd__a22o_1 _09324_ (.A1(net920),
    .A2(_03903_),
    .B1(_03877_),
    .B2(_03906_),
    .X(_00162_));
 sky130_fd_sc_hd__or2b_1 _09325_ (.A(_03789_),
    .B_N(_03750_),
    .X(_03907_));
 sky130_fd_sc_hd__xnor2_1 _09326_ (.A(_03788_),
    .B(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__mux2_1 _09327_ (.A0(\genblk2[0].wave_shpr.div.acc[13] ),
    .A1(_03908_),
    .S(_03889_),
    .X(_03909_));
 sky130_fd_sc_hd__a22o_1 _09328_ (.A1(net913),
    .A2(_03903_),
    .B1(_03877_),
    .B2(_03909_),
    .X(_00163_));
 sky130_fd_sc_hd__clkbuf_4 _09329_ (.A(_03838_),
    .X(_03910_));
 sky130_fd_sc_hd__or2b_1 _09330_ (.A(_03791_),
    .B_N(_03749_),
    .X(_03911_));
 sky130_fd_sc_hd__xnor2_1 _09331_ (.A(_03790_),
    .B(_03911_),
    .Y(_03912_));
 sky130_fd_sc_hd__mux2_1 _09332_ (.A0(\genblk2[0].wave_shpr.div.acc[14] ),
    .A1(_03912_),
    .S(_03889_),
    .X(_03913_));
 sky130_fd_sc_hd__a22o_1 _09333_ (.A1(net840),
    .A2(_03903_),
    .B1(_03910_),
    .B2(_03913_),
    .X(_00164_));
 sky130_fd_sc_hd__or2b_1 _09334_ (.A(_03793_),
    .B_N(_03748_),
    .X(_03914_));
 sky130_fd_sc_hd__xnor2_1 _09335_ (.A(_03792_),
    .B(_03914_),
    .Y(_03915_));
 sky130_fd_sc_hd__mux2_1 _09336_ (.A0(\genblk2[0].wave_shpr.div.acc[15] ),
    .A1(_03915_),
    .S(_03889_),
    .X(_03916_));
 sky130_fd_sc_hd__a22o_1 _09337_ (.A1(net1050),
    .A2(_03903_),
    .B1(_03910_),
    .B2(_03916_),
    .X(_00165_));
 sky130_fd_sc_hd__or2b_1 _09338_ (.A(_03795_),
    .B_N(_03747_),
    .X(_03917_));
 sky130_fd_sc_hd__xnor2_1 _09339_ (.A(_03917_),
    .B(_03794_),
    .Y(_03918_));
 sky130_fd_sc_hd__mux2_1 _09340_ (.A0(\genblk2[0].wave_shpr.div.acc[16] ),
    .A1(_03918_),
    .S(_03889_),
    .X(_03919_));
 sky130_fd_sc_hd__a22o_1 _09341_ (.A1(net786),
    .A2(_03903_),
    .B1(_03910_),
    .B2(_03919_),
    .X(_00166_));
 sky130_fd_sc_hd__or2b_1 _09342_ (.A(_03797_),
    .B_N(_03746_),
    .X(_03920_));
 sky130_fd_sc_hd__xnor2_1 _09343_ (.A(_03796_),
    .B(_03920_),
    .Y(_03921_));
 sky130_fd_sc_hd__mux2_1 _09344_ (.A0(\genblk2[0].wave_shpr.div.acc[17] ),
    .A1(_03921_),
    .S(_03803_),
    .X(_03922_));
 sky130_fd_sc_hd__a22o_1 _09345_ (.A1(net604),
    .A2(_03903_),
    .B1(_03910_),
    .B2(_03922_),
    .X(_00167_));
 sky130_fd_sc_hd__nor4_1 _09346_ (.A(\genblk2[0].wave_shpr.div.acc[25] ),
    .B(\genblk2[0].wave_shpr.div.acc[24] ),
    .C(\genblk2[0].wave_shpr.div.acc[26] ),
    .D(_03802_),
    .Y(_03923_));
 sky130_fd_sc_hd__or2_1 _09347_ (.A(_03799_),
    .B(net23),
    .X(_03924_));
 sky130_fd_sc_hd__o21ai_1 _09348_ (.A1(_03798_),
    .A2(net23),
    .B1(\genblk2[0].wave_shpr.div.acc[18] ),
    .Y(_03925_));
 sky130_fd_sc_hd__nand2_1 _09349_ (.A(_03924_),
    .B(_03925_),
    .Y(_03926_));
 sky130_fd_sc_hd__a22o_1 _09350_ (.A1(net688),
    .A2(_03903_),
    .B1(_03910_),
    .B2(_03926_),
    .X(_00168_));
 sky130_fd_sc_hd__nor2_1 _09351_ (.A(_03800_),
    .B(net23),
    .Y(_03927_));
 sky130_fd_sc_hd__a21o_1 _09352_ (.A1(\genblk2[0].wave_shpr.div.acc[19] ),
    .A2(_03924_),
    .B1(_03927_),
    .X(_03928_));
 sky130_fd_sc_hd__a22o_1 _09353_ (.A1(net1175),
    .A2(_03903_),
    .B1(_03910_),
    .B2(_03928_),
    .X(_00169_));
 sky130_fd_sc_hd__xor2_1 _09354_ (.A(\genblk2[0].wave_shpr.div.acc[20] ),
    .B(_03927_),
    .X(_03929_));
 sky130_fd_sc_hd__a22o_1 _09355_ (.A1(net1032),
    .A2(_03903_),
    .B1(_03910_),
    .B2(_03929_),
    .X(_00170_));
 sky130_fd_sc_hd__or3_1 _09356_ (.A(\genblk2[0].wave_shpr.div.acc[20] ),
    .B(_03800_),
    .C(net1352),
    .X(_03930_));
 sky130_fd_sc_hd__or4_1 _09357_ (.A(\genblk2[0].wave_shpr.div.acc[21] ),
    .B(\genblk2[0].wave_shpr.div.acc[20] ),
    .C(_03800_),
    .D(net1352),
    .X(_03931_));
 sky130_fd_sc_hd__a21bo_1 _09358_ (.A1(\genblk2[0].wave_shpr.div.acc[21] ),
    .A2(_03930_),
    .B1_N(_03931_),
    .X(_03932_));
 sky130_fd_sc_hd__a22o_1 _09359_ (.A1(net933),
    .A2(_03903_),
    .B1(_03910_),
    .B2(_03932_),
    .X(_00171_));
 sky130_fd_sc_hd__xnor2_1 _09360_ (.A(\genblk2[0].wave_shpr.div.acc[22] ),
    .B(_03931_),
    .Y(_03933_));
 sky130_fd_sc_hd__a22o_1 _09361_ (.A1(net653),
    .A2(_03841_),
    .B1(_03910_),
    .B2(_03933_),
    .X(_00172_));
 sky130_fd_sc_hd__nor2_1 _09362_ (.A(_03802_),
    .B(_03923_),
    .Y(_03934_));
 sky130_fd_sc_hd__a21o_1 _09363_ (.A1(\genblk2[0].wave_shpr.div.acc[23] ),
    .A2(_03801_),
    .B1(_03934_),
    .X(_03935_));
 sky130_fd_sc_hd__a22o_1 _09364_ (.A1(net1305),
    .A2(_03841_),
    .B1(_03910_),
    .B2(_03935_),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _09365_ (.A0(_03934_),
    .A1(_03802_),
    .S(\genblk2[0].wave_shpr.div.acc[24] ),
    .X(_03936_));
 sky130_fd_sc_hd__a22o_1 _09366_ (.A1(net1082),
    .A2(_03841_),
    .B1(_03839_),
    .B2(_03936_),
    .X(_00174_));
 sky130_fd_sc_hd__o21ai_1 _09367_ (.A1(\genblk2[0].wave_shpr.div.acc[24] ),
    .A2(_03802_),
    .B1(\genblk2[0].wave_shpr.div.acc[25] ),
    .Y(_03937_));
 sky130_fd_sc_hd__or4b_1 _09368_ (.A(\genblk2[0].wave_shpr.div.acc[25] ),
    .B(_03802_),
    .C(\genblk2[0].wave_shpr.div.acc[24] ),
    .D_N(\genblk2[0].wave_shpr.div.acc[26] ),
    .X(_03938_));
 sky130_fd_sc_hd__nand2_1 _09369_ (.A(_03937_),
    .B(_03938_),
    .Y(_03939_));
 sky130_fd_sc_hd__a22o_1 _09370_ (.A1(net821),
    .A2(_03841_),
    .B1(_03839_),
    .B2(_03939_),
    .X(_00175_));
 sky130_fd_sc_hd__and3_1 _09371_ (.A(_02170_),
    .B(\genblk2[11].wave_shpr.div.busy ),
    .C(_02211_),
    .X(_03940_));
 sky130_fd_sc_hd__buf_4 _09372_ (.A(_03940_),
    .X(_03941_));
 sky130_fd_sc_hd__buf_4 _09373_ (.A(_02213_),
    .X(_03942_));
 sky130_fd_sc_hd__mux2_1 _09374_ (.A0(_03941_),
    .A1(_03942_),
    .S(\genblk2[11].wave_shpr.div.i[0] ),
    .X(_03943_));
 sky130_fd_sc_hd__clkbuf_1 _09375_ (.A(_03943_),
    .X(_00176_));
 sky130_fd_sc_hd__clkbuf_4 _09376_ (.A(_03940_),
    .X(_03944_));
 sky130_fd_sc_hd__or2_1 _09377_ (.A(\genblk2[11].wave_shpr.div.i[1] ),
    .B(\genblk2[11].wave_shpr.div.i[0] ),
    .X(_03945_));
 sky130_fd_sc_hd__nand2_1 _09378_ (.A(\genblk2[11].wave_shpr.div.i[1] ),
    .B(\genblk2[11].wave_shpr.div.i[0] ),
    .Y(_03946_));
 sky130_fd_sc_hd__clkbuf_4 _09379_ (.A(_03942_),
    .X(_03947_));
 sky130_fd_sc_hd__a32o_1 _09380_ (.A1(_03944_),
    .A2(_03945_),
    .A3(_03946_),
    .B1(_03947_),
    .B2(net1124),
    .X(_00177_));
 sky130_fd_sc_hd__a21o_1 _09381_ (.A1(\genblk2[11].wave_shpr.div.i[1] ),
    .A2(\genblk2[11].wave_shpr.div.i[0] ),
    .B1(\genblk2[11].wave_shpr.div.i[2] ),
    .X(_03948_));
 sky130_fd_sc_hd__and3_1 _09382_ (.A(\genblk2[11].wave_shpr.div.i[1] ),
    .B(\genblk2[11].wave_shpr.div.i[0] ),
    .C(\genblk2[11].wave_shpr.div.i[2] ),
    .X(_03949_));
 sky130_fd_sc_hd__inv_2 _09383_ (.A(_03949_),
    .Y(_03950_));
 sky130_fd_sc_hd__a32o_1 _09384_ (.A1(_03944_),
    .A2(_03948_),
    .A3(_03950_),
    .B1(_03947_),
    .B2(net741),
    .X(_00178_));
 sky130_fd_sc_hd__a21oi_1 _09385_ (.A1(_00004_),
    .A2(_03949_),
    .B1(net1163),
    .Y(_03951_));
 sky130_fd_sc_hd__and3_1 _09386_ (.A(\genblk2[11].wave_shpr.div.i[3] ),
    .B(_02212_),
    .C(_03949_),
    .X(_03952_));
 sky130_fd_sc_hd__nor3_1 _09387_ (.A(_03726_),
    .B(_03951_),
    .C(_03952_),
    .Y(_00179_));
 sky130_fd_sc_hd__o21ai_1 _09388_ (.A1(net288),
    .A2(_03952_),
    .B1(_03819_),
    .Y(_03953_));
 sky130_fd_sc_hd__a21oi_1 _09389_ (.A1(net288),
    .A2(_03952_),
    .B1(_03953_),
    .Y(_00180_));
 sky130_fd_sc_hd__or2b_1 _09390_ (.A(\genblk2[1].wave_shpr.div.acc[17] ),
    .B_N(\genblk2[1].wave_shpr.div.b1[17] ),
    .X(_03954_));
 sky130_fd_sc_hd__and2b_1 _09391_ (.A_N(\genblk2[1].wave_shpr.div.acc[16] ),
    .B(\genblk2[1].wave_shpr.div.b1[16] ),
    .X(_03955_));
 sky130_fd_sc_hd__or2b_1 _09392_ (.A(\genblk2[1].wave_shpr.div.acc[15] ),
    .B_N(\genblk2[1].wave_shpr.div.b1[15] ),
    .X(_03956_));
 sky130_fd_sc_hd__or2b_1 _09393_ (.A(\genblk2[1].wave_shpr.div.acc[14] ),
    .B_N(\genblk2[1].wave_shpr.div.b1[14] ),
    .X(_03957_));
 sky130_fd_sc_hd__or2b_1 _09394_ (.A(\genblk2[1].wave_shpr.div.acc[13] ),
    .B_N(\genblk2[1].wave_shpr.div.b1[13] ),
    .X(_03958_));
 sky130_fd_sc_hd__or2b_1 _09395_ (.A(\genblk2[1].wave_shpr.div.acc[12] ),
    .B_N(\genblk2[1].wave_shpr.div.b1[12] ),
    .X(_03959_));
 sky130_fd_sc_hd__or2b_1 _09396_ (.A(\genblk2[1].wave_shpr.div.acc[11] ),
    .B_N(\genblk2[1].wave_shpr.div.b1[11] ),
    .X(_03960_));
 sky130_fd_sc_hd__or2b_1 _09397_ (.A(\genblk2[1].wave_shpr.div.acc[10] ),
    .B_N(\genblk2[1].wave_shpr.div.b1[10] ),
    .X(_03961_));
 sky130_fd_sc_hd__or2b_1 _09398_ (.A(\genblk2[1].wave_shpr.div.acc[9] ),
    .B_N(\genblk2[1].wave_shpr.div.b1[9] ),
    .X(_03962_));
 sky130_fd_sc_hd__or2b_1 _09399_ (.A(\genblk2[1].wave_shpr.div.acc[8] ),
    .B_N(\genblk2[1].wave_shpr.div.b1[8] ),
    .X(_03963_));
 sky130_fd_sc_hd__or2b_1 _09400_ (.A(\genblk2[1].wave_shpr.div.acc[7] ),
    .B_N(\genblk2[1].wave_shpr.div.b1[7] ),
    .X(_03964_));
 sky130_fd_sc_hd__inv_2 _09401_ (.A(\genblk2[1].wave_shpr.div.b1[6] ),
    .Y(_03965_));
 sky130_fd_sc_hd__and2b_1 _09402_ (.A_N(\genblk2[1].wave_shpr.div.acc[5] ),
    .B(\genblk2[1].wave_shpr.div.b1[5] ),
    .X(_03966_));
 sky130_fd_sc_hd__and2b_1 _09403_ (.A_N(\genblk2[1].wave_shpr.div.acc[4] ),
    .B(\genblk2[1].wave_shpr.div.b1[4] ),
    .X(_03967_));
 sky130_fd_sc_hd__or2b_1 _09404_ (.A(\genblk2[1].wave_shpr.div.acc[3] ),
    .B_N(\genblk2[1].wave_shpr.div.b1[3] ),
    .X(_03968_));
 sky130_fd_sc_hd__or2b_1 _09405_ (.A(\genblk2[1].wave_shpr.div.acc[2] ),
    .B_N(\genblk2[1].wave_shpr.div.b1[2] ),
    .X(_03969_));
 sky130_fd_sc_hd__xnor2_1 _09406_ (.A(\genblk2[1].wave_shpr.div.acc[1] ),
    .B(\genblk2[1].wave_shpr.div.b1[1] ),
    .Y(_03970_));
 sky130_fd_sc_hd__or2b_1 _09407_ (.A(\genblk2[1].wave_shpr.div.acc[0] ),
    .B_N(\genblk2[1].wave_shpr.div.b1[0] ),
    .X(_03971_));
 sky130_fd_sc_hd__and2b_1 _09408_ (.A_N(\genblk2[1].wave_shpr.div.b1[1] ),
    .B(\genblk2[1].wave_shpr.div.acc[1] ),
    .X(_03972_));
 sky130_fd_sc_hd__a21o_1 _09409_ (.A1(_03970_),
    .A2(_03971_),
    .B1(_03972_),
    .X(_03973_));
 sky130_fd_sc_hd__and2b_1 _09410_ (.A_N(\genblk2[1].wave_shpr.div.b1[2] ),
    .B(\genblk2[1].wave_shpr.div.acc[2] ),
    .X(_03974_));
 sky130_fd_sc_hd__a21o_1 _09411_ (.A1(_03969_),
    .A2(_03973_),
    .B1(_03974_),
    .X(_03975_));
 sky130_fd_sc_hd__and2b_1 _09412_ (.A_N(\genblk2[1].wave_shpr.div.b1[3] ),
    .B(\genblk2[1].wave_shpr.div.acc[3] ),
    .X(_03976_));
 sky130_fd_sc_hd__a21oi_1 _09413_ (.A1(_03968_),
    .A2(_03975_),
    .B1(_03976_),
    .Y(_03977_));
 sky130_fd_sc_hd__and2b_1 _09414_ (.A_N(\genblk2[1].wave_shpr.div.b1[4] ),
    .B(\genblk2[1].wave_shpr.div.acc[4] ),
    .X(_03978_));
 sky130_fd_sc_hd__o21ba_1 _09415_ (.A1(_03967_),
    .A2(_03977_),
    .B1_N(_03978_),
    .X(_03979_));
 sky130_fd_sc_hd__and2b_1 _09416_ (.A_N(\genblk2[1].wave_shpr.div.b1[5] ),
    .B(\genblk2[1].wave_shpr.div.acc[5] ),
    .X(_03980_));
 sky130_fd_sc_hd__o21bai_1 _09417_ (.A1(_03966_),
    .A2(_03979_),
    .B1_N(_03980_),
    .Y(_03981_));
 sky130_fd_sc_hd__o21a_1 _09418_ (.A1(_03965_),
    .A2(\genblk2[1].wave_shpr.div.acc[6] ),
    .B1(_03981_),
    .X(_03982_));
 sky130_fd_sc_hd__a21o_1 _09419_ (.A1(_03965_),
    .A2(\genblk2[1].wave_shpr.div.acc[6] ),
    .B1(_03982_),
    .X(_03983_));
 sky130_fd_sc_hd__and2b_1 _09420_ (.A_N(\genblk2[1].wave_shpr.div.b1[7] ),
    .B(\genblk2[1].wave_shpr.div.acc[7] ),
    .X(_03984_));
 sky130_fd_sc_hd__a21o_1 _09421_ (.A1(_03964_),
    .A2(_03983_),
    .B1(_03984_),
    .X(_03985_));
 sky130_fd_sc_hd__and2b_1 _09422_ (.A_N(\genblk2[1].wave_shpr.div.b1[8] ),
    .B(\genblk2[1].wave_shpr.div.acc[8] ),
    .X(_03986_));
 sky130_fd_sc_hd__a21o_1 _09423_ (.A1(_03963_),
    .A2(_03985_),
    .B1(_03986_),
    .X(_03987_));
 sky130_fd_sc_hd__and2b_1 _09424_ (.A_N(\genblk2[1].wave_shpr.div.b1[9] ),
    .B(\genblk2[1].wave_shpr.div.acc[9] ),
    .X(_03988_));
 sky130_fd_sc_hd__a21o_1 _09425_ (.A1(_03962_),
    .A2(_03987_),
    .B1(_03988_),
    .X(_03989_));
 sky130_fd_sc_hd__and2b_1 _09426_ (.A_N(\genblk2[1].wave_shpr.div.b1[10] ),
    .B(\genblk2[1].wave_shpr.div.acc[10] ),
    .X(_03990_));
 sky130_fd_sc_hd__a21o_1 _09427_ (.A1(_03961_),
    .A2(_03989_),
    .B1(_03990_),
    .X(_03991_));
 sky130_fd_sc_hd__and2b_1 _09428_ (.A_N(\genblk2[1].wave_shpr.div.b1[11] ),
    .B(\genblk2[1].wave_shpr.div.acc[11] ),
    .X(_03992_));
 sky130_fd_sc_hd__a21o_1 _09429_ (.A1(_03960_),
    .A2(_03991_),
    .B1(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__and2b_1 _09430_ (.A_N(\genblk2[1].wave_shpr.div.b1[12] ),
    .B(\genblk2[1].wave_shpr.div.acc[12] ),
    .X(_03994_));
 sky130_fd_sc_hd__a21o_1 _09431_ (.A1(_03959_),
    .A2(_03993_),
    .B1(_03994_),
    .X(_03995_));
 sky130_fd_sc_hd__and2b_1 _09432_ (.A_N(\genblk2[1].wave_shpr.div.b1[13] ),
    .B(\genblk2[1].wave_shpr.div.acc[13] ),
    .X(_03996_));
 sky130_fd_sc_hd__a21o_1 _09433_ (.A1(_03958_),
    .A2(_03995_),
    .B1(_03996_),
    .X(_03997_));
 sky130_fd_sc_hd__and2b_1 _09434_ (.A_N(\genblk2[1].wave_shpr.div.b1[14] ),
    .B(\genblk2[1].wave_shpr.div.acc[14] ),
    .X(_03998_));
 sky130_fd_sc_hd__a21o_1 _09435_ (.A1(_03957_),
    .A2(_03997_),
    .B1(_03998_),
    .X(_03999_));
 sky130_fd_sc_hd__and2b_1 _09436_ (.A_N(\genblk2[1].wave_shpr.div.b1[15] ),
    .B(\genblk2[1].wave_shpr.div.acc[15] ),
    .X(_04000_));
 sky130_fd_sc_hd__a21oi_1 _09437_ (.A1(_03956_),
    .A2(_03999_),
    .B1(_04000_),
    .Y(_04001_));
 sky130_fd_sc_hd__and2b_1 _09438_ (.A_N(\genblk2[1].wave_shpr.div.b1[16] ),
    .B(\genblk2[1].wave_shpr.div.acc[16] ),
    .X(_04002_));
 sky130_fd_sc_hd__o21bai_1 _09439_ (.A1(_03955_),
    .A2(_04001_),
    .B1_N(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__and2b_1 _09440_ (.A_N(\genblk2[1].wave_shpr.div.b1[17] ),
    .B(\genblk2[1].wave_shpr.div.acc[17] ),
    .X(_04004_));
 sky130_fd_sc_hd__a21o_1 _09441_ (.A1(_03954_),
    .A2(_04003_),
    .B1(_04004_),
    .X(_04005_));
 sky130_fd_sc_hd__or2_1 _09442_ (.A(\genblk2[1].wave_shpr.div.acc[18] ),
    .B(_04005_),
    .X(_04006_));
 sky130_fd_sc_hd__or3_1 _09443_ (.A(\genblk2[1].wave_shpr.div.acc[20] ),
    .B(\genblk2[1].wave_shpr.div.acc[19] ),
    .C(_04006_),
    .X(_04007_));
 sky130_fd_sc_hd__or4_1 _09444_ (.A(\genblk2[1].wave_shpr.div.acc[23] ),
    .B(\genblk2[1].wave_shpr.div.acc[22] ),
    .C(\genblk2[1].wave_shpr.div.acc[21] ),
    .D(_04007_),
    .X(_04008_));
 sky130_fd_sc_hd__or2_2 _09445_ (.A(\genblk2[1].wave_shpr.div.acc[24] ),
    .B(_04008_),
    .X(_04009_));
 sky130_fd_sc_hd__or3_2 _09446_ (.A(\genblk2[1].wave_shpr.div.acc[25] ),
    .B(\genblk2[1].wave_shpr.div.acc[26] ),
    .C(_04009_),
    .X(_04010_));
 sky130_fd_sc_hd__clkbuf_8 _09447_ (.A(_04010_),
    .X(_04011_));
 sky130_fd_sc_hd__mux2_1 _09448_ (.A0(\genblk2[1].wave_shpr.div.fin_quo[0] ),
    .A1(_04011_),
    .S(_00007_),
    .X(_04012_));
 sky130_fd_sc_hd__clkbuf_1 _09449_ (.A(_04012_),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _09450_ (.A0(\genblk2[1].wave_shpr.div.fin_quo[1] ),
    .A1(\genblk2[1].wave_shpr.div.quo[0] ),
    .S(_00007_),
    .X(_04013_));
 sky130_fd_sc_hd__clkbuf_1 _09451_ (.A(_04013_),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _09452_ (.A0(\genblk2[1].wave_shpr.div.fin_quo[2] ),
    .A1(net1312),
    .S(_00007_),
    .X(_04014_));
 sky130_fd_sc_hd__clkbuf_1 _09453_ (.A(_04014_),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _09454_ (.A0(\genblk2[1].wave_shpr.div.fin_quo[3] ),
    .A1(\genblk2[1].wave_shpr.div.quo[2] ),
    .S(_00007_),
    .X(_04015_));
 sky130_fd_sc_hd__clkbuf_1 _09455_ (.A(_04015_),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _09456_ (.A0(\genblk2[1].wave_shpr.div.fin_quo[4] ),
    .A1(net1316),
    .S(_00007_),
    .X(_04016_));
 sky130_fd_sc_hd__clkbuf_1 _09457_ (.A(_04016_),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _09458_ (.A0(\genblk2[1].wave_shpr.div.fin_quo[5] ),
    .A1(net414),
    .S(_00007_),
    .X(_04017_));
 sky130_fd_sc_hd__clkbuf_1 _09459_ (.A(_04017_),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _09460_ (.A0(\genblk2[1].wave_shpr.div.fin_quo[6] ),
    .A1(\genblk2[1].wave_shpr.div.quo[5] ),
    .S(_00007_),
    .X(_04018_));
 sky130_fd_sc_hd__clkbuf_1 _09461_ (.A(_04018_),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _09462_ (.A0(\genblk2[1].wave_shpr.div.fin_quo[7] ),
    .A1(\genblk2[1].wave_shpr.div.quo[6] ),
    .S(_00007_),
    .X(_04019_));
 sky130_fd_sc_hd__clkbuf_1 _09463_ (.A(_04019_),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _09464_ (.A0(\genblk2[2].wave_shpr.div.b1[0] ),
    .A1(net35),
    .S(_03822_),
    .X(_04020_));
 sky130_fd_sc_hd__clkbuf_1 _09465_ (.A(_04020_),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _09466_ (.A0(net1247),
    .A1(_01327_),
    .S(_03822_),
    .X(_04021_));
 sky130_fd_sc_hd__clkbuf_1 _09467_ (.A(_04021_),
    .X(_00190_));
 sky130_fd_sc_hd__o21a_1 _09468_ (.A1(_03732_),
    .A2(net1047),
    .B1(_03733_),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _09469_ (.A0(\genblk2[2].wave_shpr.div.b1[3] ),
    .A1(_01231_),
    .S(_03822_),
    .X(_04022_));
 sky130_fd_sc_hd__clkbuf_1 _09470_ (.A(_04022_),
    .X(_00192_));
 sky130_fd_sc_hd__inv_2 _09471_ (.A(_01418_),
    .Y(_04023_));
 sky130_fd_sc_hd__clkbuf_4 _09472_ (.A(_03701_),
    .X(_04024_));
 sky130_fd_sc_hd__mux2_1 _09473_ (.A0(\genblk2[2].wave_shpr.div.b1[4] ),
    .A1(_04023_),
    .S(_04024_),
    .X(_04025_));
 sky130_fd_sc_hd__clkbuf_1 _09474_ (.A(_04025_),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _09475_ (.A0(\genblk2[2].wave_shpr.div.b1[5] ),
    .A1(_01248_),
    .S(_04024_),
    .X(_04026_));
 sky130_fd_sc_hd__clkbuf_1 _09476_ (.A(_04026_),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _09477_ (.A0(\genblk2[2].wave_shpr.div.b1[6] ),
    .A1(_01437_),
    .S(_04024_),
    .X(_04027_));
 sky130_fd_sc_hd__clkbuf_1 _09478_ (.A(_04027_),
    .X(_00195_));
 sky130_fd_sc_hd__inv_2 _09479_ (.A(_01433_),
    .Y(_04028_));
 sky130_fd_sc_hd__mux2_1 _09480_ (.A0(\genblk2[2].wave_shpr.div.b1[7] ),
    .A1(_04028_),
    .S(_04024_),
    .X(_04029_));
 sky130_fd_sc_hd__clkbuf_1 _09481_ (.A(_04029_),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _09482_ (.A0(\genblk2[2].wave_shpr.div.b1[8] ),
    .A1(_01183_),
    .S(_04024_),
    .X(_04030_));
 sky130_fd_sc_hd__clkbuf_1 _09483_ (.A(_04030_),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _09484_ (.A0(\genblk2[2].wave_shpr.div.b1[9] ),
    .A1(_01302_),
    .S(_04024_),
    .X(_04031_));
 sky130_fd_sc_hd__clkbuf_1 _09485_ (.A(_04031_),
    .X(_00198_));
 sky130_fd_sc_hd__inv_2 _09486_ (.A(_01431_),
    .Y(_04032_));
 sky130_fd_sc_hd__mux2_1 _09487_ (.A0(net1304),
    .A1(_04032_),
    .S(_04024_),
    .X(_04033_));
 sky130_fd_sc_hd__clkbuf_1 _09488_ (.A(_04033_),
    .X(_00199_));
 sky130_fd_sc_hd__inv_2 _09489_ (.A(_01420_),
    .Y(_04034_));
 sky130_fd_sc_hd__mux2_1 _09490_ (.A0(\genblk2[2].wave_shpr.div.b1[11] ),
    .A1(_04034_),
    .S(_04024_),
    .X(_04035_));
 sky130_fd_sc_hd__clkbuf_1 _09491_ (.A(_04035_),
    .X(_00200_));
 sky130_fd_sc_hd__inv_2 _09492_ (.A(_01411_),
    .Y(_04036_));
 sky130_fd_sc_hd__mux2_1 _09493_ (.A0(net1277),
    .A1(_04036_),
    .S(_04024_),
    .X(_04037_));
 sky130_fd_sc_hd__clkbuf_1 _09494_ (.A(_04037_),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _09495_ (.A0(net1271),
    .A1(net35),
    .S(_04024_),
    .X(_04038_));
 sky130_fd_sc_hd__clkbuf_1 _09496_ (.A(_04038_),
    .X(_00202_));
 sky130_fd_sc_hd__clkbuf_4 _09497_ (.A(_03701_),
    .X(_04039_));
 sky130_fd_sc_hd__mux2_1 _09498_ (.A0(net1282),
    .A1(_01327_),
    .S(_04039_),
    .X(_04040_));
 sky130_fd_sc_hd__clkbuf_1 _09499_ (.A(_04040_),
    .X(_00203_));
 sky130_fd_sc_hd__o21a_1 _09500_ (.A1(_03732_),
    .A2(net369),
    .B1(_03733_),
    .X(_00204_));
 sky130_fd_sc_hd__a21bo_1 _09501_ (.A1(_03831_),
    .A2(net1025),
    .B1_N(_03717_),
    .X(_00205_));
 sky130_fd_sc_hd__inv_2 _09502_ (.A(net761),
    .Y(_04041_));
 sky130_fd_sc_hd__o21ai_1 _09503_ (.A1(_03714_),
    .A2(_04041_),
    .B1(_03736_),
    .Y(_00206_));
 sky130_fd_sc_hd__clkbuf_4 _09504_ (.A(_02159_),
    .X(_04042_));
 sky130_fd_sc_hd__buf_4 _09505_ (.A(_04042_),
    .X(_04043_));
 sky130_fd_sc_hd__and3_1 _09506_ (.A(_02170_),
    .B(\genblk2[1].wave_shpr.div.busy ),
    .C(_02157_),
    .X(_04044_));
 sky130_fd_sc_hd__clkbuf_4 _09507_ (.A(_04044_),
    .X(_04045_));
 sky130_fd_sc_hd__a22o_1 _09508_ (.A1(\genblk2[1].wave_shpr.div.quo[0] ),
    .A2(_04043_),
    .B1(_04011_),
    .B2(_04045_),
    .X(_00207_));
 sky130_fd_sc_hd__clkbuf_4 _09509_ (.A(_04044_),
    .X(_04046_));
 sky130_fd_sc_hd__buf_4 _09510_ (.A(_04046_),
    .X(_04047_));
 sky130_fd_sc_hd__a22o_1 _09511_ (.A1(net684),
    .A2(_04043_),
    .B1(_04047_),
    .B2(net764),
    .X(_00208_));
 sky130_fd_sc_hd__a22o_1 _09512_ (.A1(\genblk2[1].wave_shpr.div.quo[2] ),
    .A2(_04043_),
    .B1(_04047_),
    .B2(net684),
    .X(_00209_));
 sky130_fd_sc_hd__a22o_1 _09513_ (.A1(net701),
    .A2(_04043_),
    .B1(_04047_),
    .B2(net755),
    .X(_00210_));
 sky130_fd_sc_hd__a22o_1 _09514_ (.A1(net414),
    .A2(_04043_),
    .B1(_04047_),
    .B2(net701),
    .X(_00211_));
 sky130_fd_sc_hd__a22o_1 _09515_ (.A1(\genblk2[1].wave_shpr.div.quo[5] ),
    .A2(_04043_),
    .B1(_04047_),
    .B2(net414),
    .X(_00212_));
 sky130_fd_sc_hd__a22o_1 _09516_ (.A1(net292),
    .A2(_04043_),
    .B1(_04047_),
    .B2(net771),
    .X(_00213_));
 sky130_fd_sc_hd__a22o_1 _09517_ (.A1(\genblk2[1].wave_shpr.div.quo[7] ),
    .A2(_04043_),
    .B1(_04047_),
    .B2(net292),
    .X(_00214_));
 sky130_fd_sc_hd__a22o_1 _09518_ (.A1(net460),
    .A2(_04043_),
    .B1(_04047_),
    .B2(\genblk2[1].wave_shpr.div.quo[7] ),
    .X(_00215_));
 sky130_fd_sc_hd__clkbuf_4 _09519_ (.A(_04042_),
    .X(_04048_));
 sky130_fd_sc_hd__nor2_1 _09520_ (.A(_03855_),
    .B(_01330_),
    .Y(_04049_));
 sky130_fd_sc_hd__a221o_1 _09521_ (.A1(net517),
    .A2(_04048_),
    .B1(_04045_),
    .B2(net460),
    .C1(_04049_),
    .X(_00216_));
 sky130_fd_sc_hd__and2_1 _09522_ (.A(_03853_),
    .B(\genblk1[1].osc.clkdiv_C.cnt[1] ),
    .X(_04050_));
 sky130_fd_sc_hd__a221o_1 _09523_ (.A1(net610),
    .A2(_04048_),
    .B1(_04045_),
    .B2(net517),
    .C1(_04050_),
    .X(_00217_));
 sky130_fd_sc_hd__and2_1 _09524_ (.A(_03853_),
    .B(\genblk1[1].osc.clkdiv_C.cnt[2] ),
    .X(_04051_));
 sky130_fd_sc_hd__a221o_1 _09525_ (.A1(net645),
    .A2(_04048_),
    .B1(_04045_),
    .B2(net610),
    .C1(_04051_),
    .X(_00218_));
 sky130_fd_sc_hd__buf_2 _09526_ (.A(_04042_),
    .X(_04052_));
 sky130_fd_sc_hd__buf_2 _09527_ (.A(_04046_),
    .X(_04053_));
 sky130_fd_sc_hd__and2_1 _09528_ (.A(_03853_),
    .B(\genblk1[1].osc.clkdiv_C.cnt[3] ),
    .X(_04054_));
 sky130_fd_sc_hd__a221o_1 _09529_ (.A1(net537),
    .A2(_04052_),
    .B1(_04053_),
    .B2(net645),
    .C1(_04054_),
    .X(_00219_));
 sky130_fd_sc_hd__clkbuf_2 _09530_ (.A(_03707_),
    .X(_04055_));
 sky130_fd_sc_hd__and2_1 _09531_ (.A(_04055_),
    .B(\genblk1[1].osc.clkdiv_C.cnt[4] ),
    .X(_04056_));
 sky130_fd_sc_hd__a221o_1 _09532_ (.A1(net519),
    .A2(_04052_),
    .B1(_04053_),
    .B2(net537),
    .C1(_04056_),
    .X(_00220_));
 sky130_fd_sc_hd__and2_1 _09533_ (.A(_04055_),
    .B(\genblk1[1].osc.clkdiv_C.cnt[5] ),
    .X(_04057_));
 sky130_fd_sc_hd__a221o_1 _09534_ (.A1(net511),
    .A2(_04052_),
    .B1(_04053_),
    .B2(net519),
    .C1(_04057_),
    .X(_00221_));
 sky130_fd_sc_hd__buf_4 _09535_ (.A(_03719_),
    .X(_04058_));
 sky130_fd_sc_hd__nor2_1 _09536_ (.A(_04058_),
    .B(_01307_),
    .Y(_04059_));
 sky130_fd_sc_hd__a221o_1 _09537_ (.A1(\genblk2[1].wave_shpr.div.quo[15] ),
    .A2(_04052_),
    .B1(_04053_),
    .B2(net511),
    .C1(_04059_),
    .X(_00222_));
 sky130_fd_sc_hd__and2_1 _09538_ (.A(_04055_),
    .B(\genblk1[1].osc.clkdiv_C.cnt[7] ),
    .X(_04060_));
 sky130_fd_sc_hd__a221o_1 _09539_ (.A1(net462),
    .A2(_04052_),
    .B1(_04053_),
    .B2(\genblk2[1].wave_shpr.div.quo[15] ),
    .C1(_04060_),
    .X(_00223_));
 sky130_fd_sc_hd__nor2_1 _09540_ (.A(_04058_),
    .B(_02444_),
    .Y(_04061_));
 sky130_fd_sc_hd__a221o_1 _09541_ (.A1(net552),
    .A2(_04052_),
    .B1(_04053_),
    .B2(net462),
    .C1(_04061_),
    .X(_00224_));
 sky130_fd_sc_hd__and2_1 _09542_ (.A(_04055_),
    .B(\genblk1[1].osc.clkdiv_C.cnt[9] ),
    .X(_04062_));
 sky130_fd_sc_hd__a221o_1 _09543_ (.A1(net426),
    .A2(_04052_),
    .B1(_04053_),
    .B2(\genblk2[1].wave_shpr.div.quo[17] ),
    .C1(_04062_),
    .X(_00225_));
 sky130_fd_sc_hd__and2_1 _09544_ (.A(_04055_),
    .B(\genblk1[1].osc.clkdiv_C.cnt[10] ),
    .X(_04063_));
 sky130_fd_sc_hd__a221o_1 _09545_ (.A1(net417),
    .A2(_04052_),
    .B1(_04053_),
    .B2(net426),
    .C1(_04063_),
    .X(_00226_));
 sky130_fd_sc_hd__and2_1 _09546_ (.A(_04055_),
    .B(\genblk1[1].osc.clkdiv_C.cnt[11] ),
    .X(_04064_));
 sky130_fd_sc_hd__a221o_1 _09547_ (.A1(net257),
    .A2(_04052_),
    .B1(_04053_),
    .B2(net417),
    .C1(_04064_),
    .X(_00227_));
 sky130_fd_sc_hd__and2_1 _09548_ (.A(_04055_),
    .B(\genblk1[1].osc.clkdiv_C.cnt[12] ),
    .X(_04065_));
 sky130_fd_sc_hd__a221o_1 _09549_ (.A1(\genblk2[1].wave_shpr.div.quo[21] ),
    .A2(_04052_),
    .B1(_04053_),
    .B2(net257),
    .C1(_04065_),
    .X(_00228_));
 sky130_fd_sc_hd__and2_1 _09550_ (.A(_04055_),
    .B(\genblk1[1].osc.clkdiv_C.cnt[13] ),
    .X(_04066_));
 sky130_fd_sc_hd__a221o_1 _09551_ (.A1(net340),
    .A2(_04042_),
    .B1(_04046_),
    .B2(net608),
    .C1(_04066_),
    .X(_00229_));
 sky130_fd_sc_hd__and2_1 _09552_ (.A(_04055_),
    .B(\genblk1[1].osc.clkdiv_C.cnt[14] ),
    .X(_04067_));
 sky130_fd_sc_hd__a221o_1 _09553_ (.A1(\genblk2[1].wave_shpr.div.quo[23] ),
    .A2(_04042_),
    .B1(_04046_),
    .B2(net340),
    .C1(_04067_),
    .X(_00230_));
 sky130_fd_sc_hd__and2_1 _09554_ (.A(_04055_),
    .B(\genblk1[1].osc.clkdiv_C.cnt[15] ),
    .X(_04068_));
 sky130_fd_sc_hd__a221o_1 _09555_ (.A1(net632),
    .A2(_04042_),
    .B1(_04046_),
    .B2(\genblk2[1].wave_shpr.div.quo[23] ),
    .C1(_04068_),
    .X(_00231_));
 sky130_fd_sc_hd__clkbuf_4 _09556_ (.A(_03707_),
    .X(_04069_));
 sky130_fd_sc_hd__and2_1 _09557_ (.A(_04069_),
    .B(\genblk1[1].osc.clkdiv_C.cnt[16] ),
    .X(_04070_));
 sky130_fd_sc_hd__a221o_1 _09558_ (.A1(net588),
    .A2(_04042_),
    .B1(_04046_),
    .B2(\genblk2[1].wave_shpr.div.quo[24] ),
    .C1(_04070_),
    .X(_00232_));
 sky130_fd_sc_hd__or2b_1 _09559_ (.A(net588),
    .B_N(_04046_),
    .X(_04071_));
 sky130_fd_sc_hd__o221a_1 _09560_ (.A1(_03819_),
    .A2(\genblk1[1].osc.clkdiv_C.cnt[17] ),
    .B1(_00006_),
    .B2(net752),
    .C1(_04071_),
    .X(_00233_));
 sky130_fd_sc_hd__nand3_1 _09561_ (.A(\genblk2[1].wave_shpr.div.b1[0] ),
    .B(net752),
    .C(_04011_),
    .Y(_04072_));
 sky130_fd_sc_hd__a21o_1 _09562_ (.A1(\genblk2[1].wave_shpr.div.b1[0] ),
    .A2(_04011_),
    .B1(net752),
    .X(_04073_));
 sky130_fd_sc_hd__a32o_1 _09563_ (.A1(_04045_),
    .A2(_04072_),
    .A3(_04073_),
    .B1(_04048_),
    .B2(\genblk2[1].wave_shpr.div.acc[1] ),
    .X(_00234_));
 sky130_fd_sc_hd__xor2_1 _09564_ (.A(_03970_),
    .B(_03971_),
    .X(_04074_));
 sky130_fd_sc_hd__mux2_1 _09565_ (.A0(\genblk2[1].wave_shpr.div.acc[1] ),
    .A1(_04074_),
    .S(_04011_),
    .X(_04075_));
 sky130_fd_sc_hd__a22o_1 _09566_ (.A1(net990),
    .A2(_04043_),
    .B1(_04047_),
    .B2(_04075_),
    .X(_00235_));
 sky130_fd_sc_hd__clkbuf_4 _09567_ (.A(_04042_),
    .X(_04076_));
 sky130_fd_sc_hd__or2b_1 _09568_ (.A(_03974_),
    .B_N(_03969_),
    .X(_04077_));
 sky130_fd_sc_hd__xnor2_1 _09569_ (.A(_03973_),
    .B(_04077_),
    .Y(_04078_));
 sky130_fd_sc_hd__mux2_1 _09570_ (.A0(\genblk2[1].wave_shpr.div.acc[2] ),
    .A1(_04078_),
    .S(_04011_),
    .X(_04079_));
 sky130_fd_sc_hd__a22o_1 _09571_ (.A1(net965),
    .A2(_04076_),
    .B1(_04047_),
    .B2(_04079_),
    .X(_00236_));
 sky130_fd_sc_hd__clkbuf_4 _09572_ (.A(_04046_),
    .X(_04080_));
 sky130_fd_sc_hd__or2b_1 _09573_ (.A(_03976_),
    .B_N(_03968_),
    .X(_04081_));
 sky130_fd_sc_hd__xnor2_1 _09574_ (.A(_03975_),
    .B(_04081_),
    .Y(_04082_));
 sky130_fd_sc_hd__mux2_1 _09575_ (.A0(\genblk2[1].wave_shpr.div.acc[3] ),
    .A1(_04082_),
    .S(_04011_),
    .X(_04083_));
 sky130_fd_sc_hd__a22o_1 _09576_ (.A1(net829),
    .A2(_04076_),
    .B1(_04080_),
    .B2(_04083_),
    .X(_00237_));
 sky130_fd_sc_hd__nor2_1 _09577_ (.A(_03978_),
    .B(_03967_),
    .Y(_04084_));
 sky130_fd_sc_hd__xnor2_1 _09578_ (.A(_04084_),
    .B(_03977_),
    .Y(_04085_));
 sky130_fd_sc_hd__mux2_1 _09579_ (.A0(\genblk2[1].wave_shpr.div.acc[4] ),
    .A1(_04085_),
    .S(_04011_),
    .X(_04086_));
 sky130_fd_sc_hd__a22o_1 _09580_ (.A1(net825),
    .A2(_04076_),
    .B1(_04080_),
    .B2(_04086_),
    .X(_00238_));
 sky130_fd_sc_hd__nor2_1 _09581_ (.A(_03980_),
    .B(_03966_),
    .Y(_04087_));
 sky130_fd_sc_hd__xnor2_1 _09582_ (.A(_04087_),
    .B(_03979_),
    .Y(_04088_));
 sky130_fd_sc_hd__mux2_1 _09583_ (.A0(\genblk2[1].wave_shpr.div.acc[5] ),
    .A1(_04088_),
    .S(_04011_),
    .X(_04089_));
 sky130_fd_sc_hd__a22o_1 _09584_ (.A1(net1260),
    .A2(_04076_),
    .B1(_04080_),
    .B2(_04089_),
    .X(_00239_));
 sky130_fd_sc_hd__xor2_1 _09585_ (.A(\genblk2[1].wave_shpr.div.b1[6] ),
    .B(\genblk2[1].wave_shpr.div.acc[6] ),
    .X(_04090_));
 sky130_fd_sc_hd__xnor2_1 _09586_ (.A(_03981_),
    .B(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__mux2_1 _09587_ (.A0(\genblk2[1].wave_shpr.div.acc[6] ),
    .A1(_04091_),
    .S(_04011_),
    .X(_04092_));
 sky130_fd_sc_hd__a22o_1 _09588_ (.A1(net995),
    .A2(_04076_),
    .B1(_04080_),
    .B2(_04092_),
    .X(_00240_));
 sky130_fd_sc_hd__or2b_1 _09589_ (.A(_03984_),
    .B_N(_03964_),
    .X(_04093_));
 sky130_fd_sc_hd__xnor2_1 _09590_ (.A(_03983_),
    .B(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hd__buf_4 _09591_ (.A(_04010_),
    .X(_04095_));
 sky130_fd_sc_hd__mux2_1 _09592_ (.A0(\genblk2[1].wave_shpr.div.acc[7] ),
    .A1(_04094_),
    .S(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__a22o_1 _09593_ (.A1(net827),
    .A2(_04076_),
    .B1(_04080_),
    .B2(_04096_),
    .X(_00241_));
 sky130_fd_sc_hd__or2b_1 _09594_ (.A(_03986_),
    .B_N(_03963_),
    .X(_04097_));
 sky130_fd_sc_hd__xnor2_1 _09595_ (.A(_03985_),
    .B(_04097_),
    .Y(_04098_));
 sky130_fd_sc_hd__mux2_1 _09596_ (.A0(\genblk2[1].wave_shpr.div.acc[8] ),
    .A1(_04098_),
    .S(_04095_),
    .X(_04099_));
 sky130_fd_sc_hd__a22o_1 _09597_ (.A1(net847),
    .A2(_04076_),
    .B1(_04080_),
    .B2(_04099_),
    .X(_00242_));
 sky130_fd_sc_hd__or2b_1 _09598_ (.A(_03988_),
    .B_N(_03962_),
    .X(_04100_));
 sky130_fd_sc_hd__xnor2_1 _09599_ (.A(_03987_),
    .B(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__mux2_1 _09600_ (.A0(\genblk2[1].wave_shpr.div.acc[9] ),
    .A1(_04101_),
    .S(_04095_),
    .X(_04102_));
 sky130_fd_sc_hd__a22o_1 _09601_ (.A1(net813),
    .A2(_04076_),
    .B1(_04080_),
    .B2(_04102_),
    .X(_00243_));
 sky130_fd_sc_hd__or2b_1 _09602_ (.A(_03990_),
    .B_N(_03961_),
    .X(_04103_));
 sky130_fd_sc_hd__xnor2_1 _09603_ (.A(_03989_),
    .B(_04103_),
    .Y(_04104_));
 sky130_fd_sc_hd__mux2_1 _09604_ (.A0(\genblk2[1].wave_shpr.div.acc[10] ),
    .A1(_04104_),
    .S(_04095_),
    .X(_04105_));
 sky130_fd_sc_hd__a22o_1 _09605_ (.A1(net366),
    .A2(_04076_),
    .B1(_04080_),
    .B2(_04105_),
    .X(_00244_));
 sky130_fd_sc_hd__or2b_1 _09606_ (.A(_03992_),
    .B_N(_03960_),
    .X(_04106_));
 sky130_fd_sc_hd__xnor2_1 _09607_ (.A(_03991_),
    .B(_04106_),
    .Y(_04107_));
 sky130_fd_sc_hd__mux2_1 _09608_ (.A0(net366),
    .A1(_04107_),
    .S(_04095_),
    .X(_04108_));
 sky130_fd_sc_hd__a22o_1 _09609_ (.A1(\genblk2[1].wave_shpr.div.acc[12] ),
    .A2(_04076_),
    .B1(_04080_),
    .B2(_04108_),
    .X(_00245_));
 sky130_fd_sc_hd__buf_2 _09610_ (.A(_04042_),
    .X(_04109_));
 sky130_fd_sc_hd__or2b_1 _09611_ (.A(_03994_),
    .B_N(_03959_),
    .X(_04110_));
 sky130_fd_sc_hd__xnor2_1 _09612_ (.A(_03993_),
    .B(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__mux2_1 _09613_ (.A0(\genblk2[1].wave_shpr.div.acc[12] ),
    .A1(_04111_),
    .S(_04095_),
    .X(_04112_));
 sky130_fd_sc_hd__a22o_1 _09614_ (.A1(net865),
    .A2(_04109_),
    .B1(_04080_),
    .B2(_04112_),
    .X(_00246_));
 sky130_fd_sc_hd__buf_2 _09615_ (.A(_04046_),
    .X(_04113_));
 sky130_fd_sc_hd__or2b_1 _09616_ (.A(_03996_),
    .B_N(_03958_),
    .X(_04114_));
 sky130_fd_sc_hd__xnor2_1 _09617_ (.A(_03995_),
    .B(_04114_),
    .Y(_04115_));
 sky130_fd_sc_hd__mux2_1 _09618_ (.A0(\genblk2[1].wave_shpr.div.acc[13] ),
    .A1(_04115_),
    .S(_04095_),
    .X(_04116_));
 sky130_fd_sc_hd__a22o_1 _09619_ (.A1(net1019),
    .A2(_04109_),
    .B1(_04113_),
    .B2(_04116_),
    .X(_00247_));
 sky130_fd_sc_hd__or2b_1 _09620_ (.A(_03998_),
    .B_N(_03957_),
    .X(_04117_));
 sky130_fd_sc_hd__xnor2_1 _09621_ (.A(_03997_),
    .B(_04117_),
    .Y(_04118_));
 sky130_fd_sc_hd__mux2_1 _09622_ (.A0(\genblk2[1].wave_shpr.div.acc[14] ),
    .A1(_04118_),
    .S(_04095_),
    .X(_04119_));
 sky130_fd_sc_hd__a22o_1 _09623_ (.A1(net905),
    .A2(_04109_),
    .B1(_04113_),
    .B2(_04119_),
    .X(_00248_));
 sky130_fd_sc_hd__or2b_1 _09624_ (.A(_04000_),
    .B_N(_03956_),
    .X(_04120_));
 sky130_fd_sc_hd__xnor2_1 _09625_ (.A(_03999_),
    .B(_04120_),
    .Y(_04121_));
 sky130_fd_sc_hd__mux2_1 _09626_ (.A0(\genblk2[1].wave_shpr.div.acc[15] ),
    .A1(_04121_),
    .S(_04095_),
    .X(_04122_));
 sky130_fd_sc_hd__a22o_1 _09627_ (.A1(net774),
    .A2(_04109_),
    .B1(_04113_),
    .B2(_04122_),
    .X(_00249_));
 sky130_fd_sc_hd__nor2_1 _09628_ (.A(_04002_),
    .B(_03955_),
    .Y(_04123_));
 sky130_fd_sc_hd__xnor2_1 _09629_ (.A(_04123_),
    .B(_04001_),
    .Y(_04124_));
 sky130_fd_sc_hd__mux2_1 _09630_ (.A0(\genblk2[1].wave_shpr.div.acc[16] ),
    .A1(_04124_),
    .S(_04095_),
    .X(_04125_));
 sky130_fd_sc_hd__a22o_1 _09631_ (.A1(net973),
    .A2(_04109_),
    .B1(_04113_),
    .B2(_04125_),
    .X(_00250_));
 sky130_fd_sc_hd__or2b_1 _09632_ (.A(_04004_),
    .B_N(_03954_),
    .X(_04126_));
 sky130_fd_sc_hd__xnor2_1 _09633_ (.A(_04003_),
    .B(_04126_),
    .Y(_04127_));
 sky130_fd_sc_hd__mux2_1 _09634_ (.A0(\genblk2[1].wave_shpr.div.acc[17] ),
    .A1(_04127_),
    .S(_04010_),
    .X(_04128_));
 sky130_fd_sc_hd__a22o_1 _09635_ (.A1(net664),
    .A2(_04109_),
    .B1(_04113_),
    .B2(_04128_),
    .X(_00251_));
 sky130_fd_sc_hd__nor3_2 _09636_ (.A(\genblk2[1].wave_shpr.div.acc[25] ),
    .B(\genblk2[1].wave_shpr.div.acc[26] ),
    .C(_04009_),
    .Y(_04129_));
 sky130_fd_sc_hd__or2_1 _09637_ (.A(_04006_),
    .B(_04129_),
    .X(_04130_));
 sky130_fd_sc_hd__o21ai_1 _09638_ (.A1(_04005_),
    .A2(_04129_),
    .B1(\genblk2[1].wave_shpr.div.acc[18] ),
    .Y(_04131_));
 sky130_fd_sc_hd__nand2_1 _09639_ (.A(_04130_),
    .B(_04131_),
    .Y(_04132_));
 sky130_fd_sc_hd__a22o_1 _09640_ (.A1(net983),
    .A2(_04109_),
    .B1(_04113_),
    .B2(_04132_),
    .X(_00252_));
 sky130_fd_sc_hd__or2_1 _09641_ (.A(\genblk2[1].wave_shpr.div.acc[19] ),
    .B(_04130_),
    .X(_04133_));
 sky130_fd_sc_hd__nand2_1 _09642_ (.A(\genblk2[1].wave_shpr.div.acc[19] ),
    .B(_04130_),
    .Y(_04134_));
 sky130_fd_sc_hd__nand2_1 _09643_ (.A(_04133_),
    .B(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__a22o_1 _09644_ (.A1(net874),
    .A2(_04109_),
    .B1(_04113_),
    .B2(_04135_),
    .X(_00253_));
 sky130_fd_sc_hd__nor2_1 _09645_ (.A(_04007_),
    .B(_04129_),
    .Y(_04136_));
 sky130_fd_sc_hd__a21o_1 _09646_ (.A1(\genblk2[1].wave_shpr.div.acc[20] ),
    .A2(_04133_),
    .B1(_04136_),
    .X(_04137_));
 sky130_fd_sc_hd__a22o_1 _09647_ (.A1(net1109),
    .A2(_04109_),
    .B1(_04113_),
    .B2(_04137_),
    .X(_00254_));
 sky130_fd_sc_hd__xor2_1 _09648_ (.A(\genblk2[1].wave_shpr.div.acc[21] ),
    .B(_04136_),
    .X(_04138_));
 sky130_fd_sc_hd__a22o_1 _09649_ (.A1(\genblk2[1].wave_shpr.div.acc[22] ),
    .A2(_04109_),
    .B1(_04113_),
    .B2(_04138_),
    .X(_00255_));
 sky130_fd_sc_hd__or3_1 _09650_ (.A(\genblk2[1].wave_shpr.div.acc[21] ),
    .B(_04007_),
    .C(_04129_),
    .X(_04139_));
 sky130_fd_sc_hd__xnor2_1 _09651_ (.A(\genblk2[1].wave_shpr.div.acc[22] ),
    .B(_04139_),
    .Y(_04140_));
 sky130_fd_sc_hd__a22o_1 _09652_ (.A1(net803),
    .A2(_04048_),
    .B1(_04113_),
    .B2(_04140_),
    .X(_00256_));
 sky130_fd_sc_hd__or3b_1 _09653_ (.A(\genblk2[1].wave_shpr.div.acc[22] ),
    .B(_04139_),
    .C_N(\genblk2[1].wave_shpr.div.acc[23] ),
    .X(_04141_));
 sky130_fd_sc_hd__o21bai_1 _09654_ (.A1(\genblk2[1].wave_shpr.div.acc[22] ),
    .A2(_04139_),
    .B1_N(\genblk2[1].wave_shpr.div.acc[23] ),
    .Y(_04142_));
 sky130_fd_sc_hd__a32o_1 _09655_ (.A1(_04045_),
    .A2(_04141_),
    .A3(_04142_),
    .B1(_04048_),
    .B2(net448),
    .X(_00257_));
 sky130_fd_sc_hd__nand2_1 _09656_ (.A(\genblk2[1].wave_shpr.div.acc[24] ),
    .B(_04008_),
    .Y(_04143_));
 sky130_fd_sc_hd__o21ai_1 _09657_ (.A1(_04009_),
    .A2(_04129_),
    .B1(_04143_),
    .Y(_04144_));
 sky130_fd_sc_hd__a22o_1 _09658_ (.A1(net1228),
    .A2(_04048_),
    .B1(_04045_),
    .B2(_04144_),
    .X(_00258_));
 sky130_fd_sc_hd__or3b_1 _09659_ (.A(_04009_),
    .B(\genblk2[1].wave_shpr.div.acc[25] ),
    .C_N(\genblk2[1].wave_shpr.div.acc[26] ),
    .X(_04145_));
 sky130_fd_sc_hd__a21bo_1 _09660_ (.A1(\genblk2[1].wave_shpr.div.acc[25] ),
    .A2(_04009_),
    .B1_N(_04145_),
    .X(_04146_));
 sky130_fd_sc_hd__a22o_1 _09661_ (.A1(net1107),
    .A2(_04048_),
    .B1(_04045_),
    .B2(_04146_),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _09662_ (.A0(_04046_),
    .A1(_04042_),
    .S(\genblk2[1].wave_shpr.div.i[0] ),
    .X(_04147_));
 sky130_fd_sc_hd__clkbuf_1 _09663_ (.A(_04147_),
    .X(_00260_));
 sky130_fd_sc_hd__or2_1 _09664_ (.A(\genblk2[1].wave_shpr.div.i[1] ),
    .B(\genblk2[1].wave_shpr.div.i[0] ),
    .X(_04148_));
 sky130_fd_sc_hd__nand2_1 _09665_ (.A(\genblk2[1].wave_shpr.div.i[1] ),
    .B(\genblk2[1].wave_shpr.div.i[0] ),
    .Y(_04149_));
 sky130_fd_sc_hd__a32o_1 _09666_ (.A1(_04045_),
    .A2(_04148_),
    .A3(_04149_),
    .B1(_04048_),
    .B2(net1091),
    .X(_00261_));
 sky130_fd_sc_hd__a21o_1 _09667_ (.A1(\genblk2[1].wave_shpr.div.i[1] ),
    .A2(\genblk2[1].wave_shpr.div.i[0] ),
    .B1(\genblk2[1].wave_shpr.div.i[2] ),
    .X(_04150_));
 sky130_fd_sc_hd__and3_1 _09668_ (.A(\genblk2[1].wave_shpr.div.i[1] ),
    .B(\genblk2[1].wave_shpr.div.i[0] ),
    .C(\genblk2[1].wave_shpr.div.i[2] ),
    .X(_04151_));
 sky130_fd_sc_hd__inv_2 _09669_ (.A(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__a32o_1 _09670_ (.A1(_04045_),
    .A2(_04150_),
    .A3(_04152_),
    .B1(_04048_),
    .B2(net757),
    .X(_00262_));
 sky130_fd_sc_hd__a21oi_1 _09671_ (.A1(_00006_),
    .A2(_04151_),
    .B1(net1174),
    .Y(_04153_));
 sky130_fd_sc_hd__and3_1 _09672_ (.A(\genblk2[1].wave_shpr.div.i[3] ),
    .B(_02158_),
    .C(_04151_),
    .X(_04154_));
 sky130_fd_sc_hd__nor3_1 _09673_ (.A(_03690_),
    .B(_04153_),
    .C(_04154_),
    .Y(_00263_));
 sky130_fd_sc_hd__o21ai_1 _09674_ (.A1(net285),
    .A2(_04154_),
    .B1(_03819_),
    .Y(_04155_));
 sky130_fd_sc_hd__a21oi_1 _09675_ (.A1(net285),
    .A2(_04154_),
    .B1(_04155_),
    .Y(_00264_));
 sky130_fd_sc_hd__or2_1 _09676_ (.A(\genblk2[2].wave_shpr.div.acc[17] ),
    .B(_04041_),
    .X(_04156_));
 sky130_fd_sc_hd__or2b_1 _09677_ (.A(\genblk2[2].wave_shpr.div.acc[16] ),
    .B_N(\genblk2[2].wave_shpr.div.b1[16] ),
    .X(_04157_));
 sky130_fd_sc_hd__or2b_1 _09678_ (.A(\genblk2[2].wave_shpr.div.acc[15] ),
    .B_N(\genblk2[2].wave_shpr.div.b1[15] ),
    .X(_04158_));
 sky130_fd_sc_hd__or2b_1 _09679_ (.A(\genblk2[2].wave_shpr.div.acc[14] ),
    .B_N(\genblk2[2].wave_shpr.div.b1[14] ),
    .X(_04159_));
 sky130_fd_sc_hd__or2b_1 _09680_ (.A(\genblk2[2].wave_shpr.div.acc[13] ),
    .B_N(\genblk2[2].wave_shpr.div.b1[13] ),
    .X(_04160_));
 sky130_fd_sc_hd__or2b_1 _09681_ (.A(\genblk2[2].wave_shpr.div.acc[12] ),
    .B_N(\genblk2[2].wave_shpr.div.b1[12] ),
    .X(_04161_));
 sky130_fd_sc_hd__or2b_1 _09682_ (.A(\genblk2[2].wave_shpr.div.acc[11] ),
    .B_N(\genblk2[2].wave_shpr.div.b1[11] ),
    .X(_04162_));
 sky130_fd_sc_hd__or2b_1 _09683_ (.A(\genblk2[2].wave_shpr.div.acc[10] ),
    .B_N(\genblk2[2].wave_shpr.div.b1[10] ),
    .X(_04163_));
 sky130_fd_sc_hd__or2b_1 _09684_ (.A(\genblk2[2].wave_shpr.div.acc[9] ),
    .B_N(\genblk2[2].wave_shpr.div.b1[9] ),
    .X(_04164_));
 sky130_fd_sc_hd__or2b_1 _09685_ (.A(\genblk2[2].wave_shpr.div.acc[8] ),
    .B_N(\genblk2[2].wave_shpr.div.b1[8] ),
    .X(_04165_));
 sky130_fd_sc_hd__or2b_1 _09686_ (.A(\genblk2[2].wave_shpr.div.acc[7] ),
    .B_N(\genblk2[2].wave_shpr.div.b1[7] ),
    .X(_04166_));
 sky130_fd_sc_hd__or2b_1 _09687_ (.A(\genblk2[2].wave_shpr.div.acc[6] ),
    .B_N(\genblk2[2].wave_shpr.div.b1[6] ),
    .X(_04167_));
 sky130_fd_sc_hd__or2b_1 _09688_ (.A(\genblk2[2].wave_shpr.div.acc[5] ),
    .B_N(\genblk2[2].wave_shpr.div.b1[5] ),
    .X(_04168_));
 sky130_fd_sc_hd__or2b_1 _09689_ (.A(\genblk2[2].wave_shpr.div.acc[4] ),
    .B_N(\genblk2[2].wave_shpr.div.b1[4] ),
    .X(_04169_));
 sky130_fd_sc_hd__or2b_1 _09690_ (.A(\genblk2[2].wave_shpr.div.acc[3] ),
    .B_N(\genblk2[2].wave_shpr.div.b1[3] ),
    .X(_04170_));
 sky130_fd_sc_hd__inv_2 _09691_ (.A(\genblk2[2].wave_shpr.div.b1[2] ),
    .Y(_04171_));
 sky130_fd_sc_hd__or2b_1 _09692_ (.A(\genblk2[2].wave_shpr.div.b1[1] ),
    .B_N(\genblk2[2].wave_shpr.div.acc[1] ),
    .X(_04172_));
 sky130_fd_sc_hd__or2b_1 _09693_ (.A(\genblk2[2].wave_shpr.div.acc[1] ),
    .B_N(\genblk2[2].wave_shpr.div.b1[1] ),
    .X(_04173_));
 sky130_fd_sc_hd__nand2_1 _09694_ (.A(_04172_),
    .B(_04173_),
    .Y(_04174_));
 sky130_fd_sc_hd__and2b_1 _09695_ (.A_N(\genblk2[2].wave_shpr.div.acc[0] ),
    .B(\genblk2[2].wave_shpr.div.b1[0] ),
    .X(_04175_));
 sky130_fd_sc_hd__o21ai_1 _09696_ (.A1(_04174_),
    .A2(_04175_),
    .B1(_04172_),
    .Y(_04176_));
 sky130_fd_sc_hd__o21a_1 _09697_ (.A1(_04171_),
    .A2(\genblk2[2].wave_shpr.div.acc[2] ),
    .B1(_04176_),
    .X(_04177_));
 sky130_fd_sc_hd__a21o_1 _09698_ (.A1(_04171_),
    .A2(\genblk2[2].wave_shpr.div.acc[2] ),
    .B1(_04177_),
    .X(_04178_));
 sky130_fd_sc_hd__and2b_1 _09699_ (.A_N(\genblk2[2].wave_shpr.div.b1[3] ),
    .B(\genblk2[2].wave_shpr.div.acc[3] ),
    .X(_04179_));
 sky130_fd_sc_hd__a21o_1 _09700_ (.A1(_04170_),
    .A2(_04178_),
    .B1(_04179_),
    .X(_04180_));
 sky130_fd_sc_hd__and2b_1 _09701_ (.A_N(\genblk2[2].wave_shpr.div.b1[4] ),
    .B(\genblk2[2].wave_shpr.div.acc[4] ),
    .X(_04181_));
 sky130_fd_sc_hd__a21o_1 _09702_ (.A1(_04169_),
    .A2(_04180_),
    .B1(_04181_),
    .X(_04182_));
 sky130_fd_sc_hd__and2b_1 _09703_ (.A_N(\genblk2[2].wave_shpr.div.b1[5] ),
    .B(\genblk2[2].wave_shpr.div.acc[5] ),
    .X(_04183_));
 sky130_fd_sc_hd__a21o_1 _09704_ (.A1(_04168_),
    .A2(_04182_),
    .B1(_04183_),
    .X(_04184_));
 sky130_fd_sc_hd__and2b_1 _09705_ (.A_N(\genblk2[2].wave_shpr.div.b1[6] ),
    .B(\genblk2[2].wave_shpr.div.acc[6] ),
    .X(_04185_));
 sky130_fd_sc_hd__a21o_1 _09706_ (.A1(_04167_),
    .A2(_04184_),
    .B1(_04185_),
    .X(_04186_));
 sky130_fd_sc_hd__and2b_1 _09707_ (.A_N(\genblk2[2].wave_shpr.div.b1[7] ),
    .B(\genblk2[2].wave_shpr.div.acc[7] ),
    .X(_04187_));
 sky130_fd_sc_hd__a21o_1 _09708_ (.A1(_04166_),
    .A2(_04186_),
    .B1(_04187_),
    .X(_04188_));
 sky130_fd_sc_hd__and2b_1 _09709_ (.A_N(\genblk2[2].wave_shpr.div.b1[8] ),
    .B(\genblk2[2].wave_shpr.div.acc[8] ),
    .X(_04189_));
 sky130_fd_sc_hd__a21o_1 _09710_ (.A1(_04165_),
    .A2(_04188_),
    .B1(_04189_),
    .X(_04190_));
 sky130_fd_sc_hd__and2b_1 _09711_ (.A_N(\genblk2[2].wave_shpr.div.b1[9] ),
    .B(\genblk2[2].wave_shpr.div.acc[9] ),
    .X(_04191_));
 sky130_fd_sc_hd__a21o_1 _09712_ (.A1(_04164_),
    .A2(_04190_),
    .B1(_04191_),
    .X(_04192_));
 sky130_fd_sc_hd__and2b_1 _09713_ (.A_N(\genblk2[2].wave_shpr.div.b1[10] ),
    .B(\genblk2[2].wave_shpr.div.acc[10] ),
    .X(_04193_));
 sky130_fd_sc_hd__a21o_1 _09714_ (.A1(_04163_),
    .A2(_04192_),
    .B1(_04193_),
    .X(_04194_));
 sky130_fd_sc_hd__and2b_1 _09715_ (.A_N(\genblk2[2].wave_shpr.div.b1[11] ),
    .B(\genblk2[2].wave_shpr.div.acc[11] ),
    .X(_04195_));
 sky130_fd_sc_hd__a21o_1 _09716_ (.A1(_04162_),
    .A2(_04194_),
    .B1(_04195_),
    .X(_04196_));
 sky130_fd_sc_hd__and2b_1 _09717_ (.A_N(\genblk2[2].wave_shpr.div.b1[12] ),
    .B(\genblk2[2].wave_shpr.div.acc[12] ),
    .X(_04197_));
 sky130_fd_sc_hd__a21o_1 _09718_ (.A1(_04161_),
    .A2(_04196_),
    .B1(_04197_),
    .X(_04198_));
 sky130_fd_sc_hd__and2b_1 _09719_ (.A_N(\genblk2[2].wave_shpr.div.b1[13] ),
    .B(\genblk2[2].wave_shpr.div.acc[13] ),
    .X(_04199_));
 sky130_fd_sc_hd__a21o_1 _09720_ (.A1(_04160_),
    .A2(_04198_),
    .B1(_04199_),
    .X(_04200_));
 sky130_fd_sc_hd__and2b_1 _09721_ (.A_N(\genblk2[2].wave_shpr.div.b1[14] ),
    .B(\genblk2[2].wave_shpr.div.acc[14] ),
    .X(_04201_));
 sky130_fd_sc_hd__a21o_1 _09722_ (.A1(_04159_),
    .A2(_04200_),
    .B1(_04201_),
    .X(_04202_));
 sky130_fd_sc_hd__and2b_1 _09723_ (.A_N(\genblk2[2].wave_shpr.div.b1[15] ),
    .B(\genblk2[2].wave_shpr.div.acc[15] ),
    .X(_04203_));
 sky130_fd_sc_hd__a21o_1 _09724_ (.A1(_04158_),
    .A2(_04202_),
    .B1(_04203_),
    .X(_04204_));
 sky130_fd_sc_hd__and2b_1 _09725_ (.A_N(\genblk2[2].wave_shpr.div.b1[16] ),
    .B(\genblk2[2].wave_shpr.div.acc[16] ),
    .X(_04205_));
 sky130_fd_sc_hd__a21o_1 _09726_ (.A1(_04157_),
    .A2(_04204_),
    .B1(_04205_),
    .X(_04206_));
 sky130_fd_sc_hd__and2_1 _09727_ (.A(\genblk2[2].wave_shpr.div.acc[17] ),
    .B(_04041_),
    .X(_04207_));
 sky130_fd_sc_hd__a21o_1 _09728_ (.A1(_04156_),
    .A2(_04206_),
    .B1(_04207_),
    .X(_04208_));
 sky130_fd_sc_hd__or2_1 _09729_ (.A(\genblk2[2].wave_shpr.div.acc[18] ),
    .B(_04208_),
    .X(_04209_));
 sky130_fd_sc_hd__or2_1 _09730_ (.A(\genblk2[2].wave_shpr.div.acc[19] ),
    .B(_04209_),
    .X(_04210_));
 sky130_fd_sc_hd__or4_1 _09731_ (.A(\genblk2[2].wave_shpr.div.acc[22] ),
    .B(\genblk2[2].wave_shpr.div.acc[21] ),
    .C(\genblk2[2].wave_shpr.div.acc[20] ),
    .D(_04210_),
    .X(_04211_));
 sky130_fd_sc_hd__or2_2 _09732_ (.A(\genblk2[2].wave_shpr.div.acc[23] ),
    .B(_04211_),
    .X(_04212_));
 sky130_fd_sc_hd__or4_2 _09733_ (.A(\genblk2[2].wave_shpr.div.acc[25] ),
    .B(\genblk2[2].wave_shpr.div.acc[24] ),
    .C(\genblk2[2].wave_shpr.div.acc[26] ),
    .D(_04212_),
    .X(_04213_));
 sky130_fd_sc_hd__clkbuf_4 _09734_ (.A(_04213_),
    .X(_04214_));
 sky130_fd_sc_hd__mux2_1 _09735_ (.A0(\genblk2[2].wave_shpr.div.fin_quo[0] ),
    .A1(_04214_),
    .S(_00009_),
    .X(_04215_));
 sky130_fd_sc_hd__clkbuf_1 _09736_ (.A(_04215_),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _09737_ (.A0(\genblk2[2].wave_shpr.div.fin_quo[1] ),
    .A1(net1348),
    .S(_00009_),
    .X(_04216_));
 sky130_fd_sc_hd__clkbuf_1 _09738_ (.A(_04216_),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _09739_ (.A0(\genblk2[2].wave_shpr.div.fin_quo[2] ),
    .A1(net1343),
    .S(_00009_),
    .X(_04217_));
 sky130_fd_sc_hd__clkbuf_1 _09740_ (.A(_04217_),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _09741_ (.A0(\genblk2[2].wave_shpr.div.fin_quo[3] ),
    .A1(net1329),
    .S(_00009_),
    .X(_04218_));
 sky130_fd_sc_hd__clkbuf_1 _09742_ (.A(_04218_),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _09743_ (.A0(\genblk2[2].wave_shpr.div.fin_quo[4] ),
    .A1(net1327),
    .S(_00009_),
    .X(_04219_));
 sky130_fd_sc_hd__clkbuf_1 _09744_ (.A(_04219_),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _09745_ (.A0(\genblk2[2].wave_shpr.div.fin_quo[5] ),
    .A1(\genblk2[2].wave_shpr.div.quo[4] ),
    .S(_00009_),
    .X(_04220_));
 sky130_fd_sc_hd__clkbuf_1 _09746_ (.A(_04220_),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _09747_ (.A0(\genblk2[2].wave_shpr.div.fin_quo[6] ),
    .A1(\genblk2[2].wave_shpr.div.quo[5] ),
    .S(_00009_),
    .X(_04221_));
 sky130_fd_sc_hd__clkbuf_1 _09748_ (.A(_04221_),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _09749_ (.A0(\genblk2[2].wave_shpr.div.fin_quo[7] ),
    .A1(net1197),
    .S(_00009_),
    .X(_04222_));
 sky130_fd_sc_hd__clkbuf_1 _09750_ (.A(net1198),
    .X(_00272_));
 sky130_fd_sc_hd__nor2_2 _09751_ (.A(_01211_),
    .B(_01302_),
    .Y(_04223_));
 sky130_fd_sc_hd__mux2_1 _09752_ (.A0(\genblk2[3].wave_shpr.div.b1[0] ),
    .A1(_04223_),
    .S(_04039_),
    .X(_04224_));
 sky130_fd_sc_hd__clkbuf_1 _09753_ (.A(_04224_),
    .X(_00273_));
 sky130_fd_sc_hd__nand2_2 _09754_ (.A(_01436_),
    .B(_01925_),
    .Y(_04225_));
 sky130_fd_sc_hd__mux2_1 _09755_ (.A0(\genblk2[3].wave_shpr.div.b1[1] ),
    .A1(_04225_),
    .S(_04039_),
    .X(_04226_));
 sky130_fd_sc_hd__clkbuf_1 _09756_ (.A(_04226_),
    .X(_00274_));
 sky130_fd_sc_hd__inv_2 _09757_ (.A(_01496_),
    .Y(_04227_));
 sky130_fd_sc_hd__mux2_1 _09758_ (.A0(\genblk2[3].wave_shpr.div.b1[2] ),
    .A1(_04227_),
    .S(_04039_),
    .X(_04228_));
 sky130_fd_sc_hd__clkbuf_1 _09759_ (.A(_04228_),
    .X(_00275_));
 sky130_fd_sc_hd__nor2_4 _09760_ (.A(_01325_),
    .B(_01423_),
    .Y(_04229_));
 sky130_fd_sc_hd__nand2_4 _09761_ (.A(_01436_),
    .B(_04229_),
    .Y(_04230_));
 sky130_fd_sc_hd__mux2_1 _09762_ (.A0(net1290),
    .A1(_04230_),
    .S(_04039_),
    .X(_04231_));
 sky130_fd_sc_hd__clkbuf_1 _09763_ (.A(_04231_),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _09764_ (.A0(net1245),
    .A1(_01794_),
    .S(_04039_),
    .X(_04232_));
 sky130_fd_sc_hd__clkbuf_1 _09765_ (.A(_04232_),
    .X(_00277_));
 sky130_fd_sc_hd__nor2_4 _09766_ (.A(_01302_),
    .B(_03727_),
    .Y(_04233_));
 sky130_fd_sc_hd__a21o_1 _09767_ (.A1(_03704_),
    .A2(net1099),
    .B1(_04233_),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _09768_ (.A0(\genblk2[3].wave_shpr.div.b1[6] ),
    .A1(_01262_),
    .S(_04039_),
    .X(_04234_));
 sky130_fd_sc_hd__clkbuf_1 _09769_ (.A(_04234_),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _09770_ (.A0(\genblk2[3].wave_shpr.div.b1[7] ),
    .A1(_02077_),
    .S(_04039_),
    .X(_04235_));
 sky130_fd_sc_hd__clkbuf_1 _09771_ (.A(_04235_),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _09772_ (.A0(net1298),
    .A1(_01256_),
    .S(_04039_),
    .X(_04236_));
 sky130_fd_sc_hd__clkbuf_1 _09773_ (.A(_04236_),
    .X(_00281_));
 sky130_fd_sc_hd__a21bo_1 _09774_ (.A1(_03831_),
    .A2(net614),
    .B1_N(_03733_),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _09775_ (.A0(\genblk2[3].wave_shpr.div.b1[10] ),
    .A1(_02336_),
    .S(_04039_),
    .X(_04237_));
 sky130_fd_sc_hd__clkbuf_1 _09776_ (.A(_04237_),
    .X(_00283_));
 sky130_fd_sc_hd__buf_4 _09777_ (.A(_03701_),
    .X(_04238_));
 sky130_fd_sc_hd__mux2_1 _09778_ (.A0(net1297),
    .A1(_01487_),
    .S(_04238_),
    .X(_04239_));
 sky130_fd_sc_hd__clkbuf_1 _09779_ (.A(_04239_),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _09780_ (.A0(net1285),
    .A1(_01858_),
    .S(_04238_),
    .X(_04240_));
 sky130_fd_sc_hd__clkbuf_1 _09781_ (.A(_04240_),
    .X(_00285_));
 sky130_fd_sc_hd__nand2_4 _09782_ (.A(_03702_),
    .B(_01490_),
    .Y(_04241_));
 sky130_fd_sc_hd__o21a_1 _09783_ (.A1(_03732_),
    .A2(net1152),
    .B1(_04241_),
    .X(_00286_));
 sky130_fd_sc_hd__nor2_4 _09784_ (.A(_01490_),
    .B(_01233_),
    .Y(_04242_));
 sky130_fd_sc_hd__mux2_1 _09785_ (.A0(\genblk2[3].wave_shpr.div.b1[14] ),
    .A1(_04242_),
    .S(_04238_),
    .X(_04243_));
 sky130_fd_sc_hd__clkbuf_1 _09786_ (.A(_04243_),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _09787_ (.A0(\genblk2[3].wave_shpr.div.b1[15] ),
    .A1(_01365_),
    .S(_04238_),
    .X(_04244_));
 sky130_fd_sc_hd__clkbuf_1 _09788_ (.A(_04244_),
    .X(_00288_));
 sky130_fd_sc_hd__inv_2 _09789_ (.A(net730),
    .Y(_04245_));
 sky130_fd_sc_hd__o21ai_1 _09790_ (.A1(_03714_),
    .A2(_04245_),
    .B1(_03736_),
    .Y(_00289_));
 sky130_fd_sc_hd__and2_1 _09791_ (.A(_03833_),
    .B(net1190),
    .X(_04246_));
 sky130_fd_sc_hd__clkbuf_1 _09792_ (.A(_04246_),
    .X(_00290_));
 sky130_fd_sc_hd__clkbuf_4 _09793_ (.A(_02164_),
    .X(_04247_));
 sky130_fd_sc_hd__clkbuf_4 _09794_ (.A(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__and3_1 _09795_ (.A(_02152_),
    .B(\genblk2[2].wave_shpr.div.busy ),
    .C(_02162_),
    .X(_04249_));
 sky130_fd_sc_hd__buf_4 _09796_ (.A(_04249_),
    .X(_04250_));
 sky130_fd_sc_hd__clkbuf_4 _09797_ (.A(_04250_),
    .X(_04251_));
 sky130_fd_sc_hd__a22o_1 _09798_ (.A1(net1054),
    .A2(_04248_),
    .B1(_04214_),
    .B2(_04251_),
    .X(_00291_));
 sky130_fd_sc_hd__clkbuf_4 _09799_ (.A(_04250_),
    .X(_04252_));
 sky130_fd_sc_hd__a22o_1 _09800_ (.A1(net812),
    .A2(_04248_),
    .B1(_04252_),
    .B2(net1054),
    .X(_00292_));
 sky130_fd_sc_hd__a22o_1 _09801_ (.A1(net719),
    .A2(_04248_),
    .B1(_04252_),
    .B2(net812),
    .X(_00293_));
 sky130_fd_sc_hd__a22o_1 _09802_ (.A1(net336),
    .A2(_04248_),
    .B1(_04252_),
    .B2(net719),
    .X(_00294_));
 sky130_fd_sc_hd__a22o_1 _09803_ (.A1(\genblk2[2].wave_shpr.div.quo[4] ),
    .A2(_04248_),
    .B1(_04252_),
    .B2(net336),
    .X(_00295_));
 sky130_fd_sc_hd__a22o_1 _09804_ (.A1(\genblk2[2].wave_shpr.div.quo[5] ),
    .A2(_04248_),
    .B1(_04252_),
    .B2(net696),
    .X(_00296_));
 sky130_fd_sc_hd__a22o_1 _09805_ (.A1(net449),
    .A2(_04248_),
    .B1(_04252_),
    .B2(net716),
    .X(_00297_));
 sky130_fd_sc_hd__a22o_1 _09806_ (.A1(net275),
    .A2(_04248_),
    .B1(_04252_),
    .B2(net449),
    .X(_00298_));
 sky130_fd_sc_hd__a22o_1 _09807_ (.A1(\genblk2[2].wave_shpr.div.quo[8] ),
    .A2(_04248_),
    .B1(_04252_),
    .B2(net275),
    .X(_00299_));
 sky130_fd_sc_hd__clkbuf_4 _09808_ (.A(_04247_),
    .X(_04253_));
 sky130_fd_sc_hd__and2_1 _09809_ (.A(_04069_),
    .B(\genblk1[2].osc.clkdiv_C.cnt[0] ),
    .X(_04254_));
 sky130_fd_sc_hd__a221o_1 _09810_ (.A1(\genblk2[2].wave_shpr.div.quo[9] ),
    .A2(_04253_),
    .B1(_04251_),
    .B2(net300),
    .C1(_04254_),
    .X(_00300_));
 sky130_fd_sc_hd__and2_1 _09811_ (.A(_04069_),
    .B(\genblk1[2].osc.clkdiv_C.cnt[1] ),
    .X(_04255_));
 sky130_fd_sc_hd__a221o_1 _09812_ (.A1(net441),
    .A2(_04253_),
    .B1(_04251_),
    .B2(net574),
    .C1(_04255_),
    .X(_00301_));
 sky130_fd_sc_hd__nor2_1 _09813_ (.A(_04058_),
    .B(_01414_),
    .Y(_04256_));
 sky130_fd_sc_hd__a221o_1 _09814_ (.A1(\genblk2[2].wave_shpr.div.quo[11] ),
    .A2(_04253_),
    .B1(_04251_),
    .B2(net441),
    .C1(_04256_),
    .X(_00302_));
 sky130_fd_sc_hd__clkbuf_4 _09815_ (.A(_04247_),
    .X(_04257_));
 sky130_fd_sc_hd__nor2_1 _09816_ (.A(_04058_),
    .B(_01410_),
    .Y(_04258_));
 sky130_fd_sc_hd__a221o_1 _09817_ (.A1(net553),
    .A2(_04257_),
    .B1(_04251_),
    .B2(\genblk2[2].wave_shpr.div.quo[11] ),
    .C1(_04258_),
    .X(_00303_));
 sky130_fd_sc_hd__clkbuf_4 _09818_ (.A(_04250_),
    .X(_04259_));
 sky130_fd_sc_hd__and2_1 _09819_ (.A(_04069_),
    .B(\genblk1[2].osc.clkdiv_C.cnt[4] ),
    .X(_04260_));
 sky130_fd_sc_hd__a221o_1 _09820_ (.A1(net457),
    .A2(_04257_),
    .B1(_04259_),
    .B2(net553),
    .C1(_04260_),
    .X(_00304_));
 sky130_fd_sc_hd__and2_1 _09821_ (.A(_04069_),
    .B(\genblk1[2].osc.clkdiv_C.cnt[5] ),
    .X(_04261_));
 sky130_fd_sc_hd__a221o_1 _09822_ (.A1(\genblk2[2].wave_shpr.div.quo[14] ),
    .A2(_04257_),
    .B1(_04259_),
    .B2(net457),
    .C1(_04261_),
    .X(_00305_));
 sky130_fd_sc_hd__and2_1 _09823_ (.A(_04069_),
    .B(\genblk1[2].osc.clkdiv_C.cnt[6] ),
    .X(_04262_));
 sky130_fd_sc_hd__a221o_1 _09824_ (.A1(net315),
    .A2(_04257_),
    .B1(_04259_),
    .B2(net480),
    .C1(_04262_),
    .X(_00306_));
 sky130_fd_sc_hd__and2_1 _09825_ (.A(_04069_),
    .B(\genblk1[2].osc.clkdiv_C.cnt[7] ),
    .X(_04263_));
 sky130_fd_sc_hd__a221o_1 _09826_ (.A1(\genblk2[2].wave_shpr.div.quo[16] ),
    .A2(_04257_),
    .B1(_04259_),
    .B2(net315),
    .C1(_04263_),
    .X(_00307_));
 sky130_fd_sc_hd__nor2_1 _09827_ (.A(_04058_),
    .B(_01412_),
    .Y(_04264_));
 sky130_fd_sc_hd__a221o_1 _09828_ (.A1(net393),
    .A2(_04257_),
    .B1(_04259_),
    .B2(net573),
    .C1(_04264_),
    .X(_00308_));
 sky130_fd_sc_hd__and2_1 _09829_ (.A(_04069_),
    .B(\genblk1[2].osc.clkdiv_C.cnt[9] ),
    .X(_04265_));
 sky130_fd_sc_hd__a221o_1 _09830_ (.A1(net339),
    .A2(_04257_),
    .B1(_04259_),
    .B2(net393),
    .C1(_04265_),
    .X(_00309_));
 sky130_fd_sc_hd__and2_1 _09831_ (.A(_04069_),
    .B(\genblk1[2].osc.clkdiv_C.cnt[10] ),
    .X(_04266_));
 sky130_fd_sc_hd__a221o_1 _09832_ (.A1(net322),
    .A2(_04257_),
    .B1(_04259_),
    .B2(net339),
    .C1(_04266_),
    .X(_00310_));
 sky130_fd_sc_hd__and2_1 _09833_ (.A(_04069_),
    .B(\genblk1[2].osc.clkdiv_C.cnt[11] ),
    .X(_04267_));
 sky130_fd_sc_hd__a221o_1 _09834_ (.A1(\genblk2[2].wave_shpr.div.quo[20] ),
    .A2(_04257_),
    .B1(_04259_),
    .B2(net322),
    .C1(_04267_),
    .X(_00311_));
 sky130_fd_sc_hd__buf_4 _09835_ (.A(_02147_),
    .X(_04268_));
 sky130_fd_sc_hd__buf_2 _09836_ (.A(_04268_),
    .X(_04269_));
 sky130_fd_sc_hd__and2_1 _09837_ (.A(_04269_),
    .B(\genblk1[2].osc.clkdiv_C.cnt[12] ),
    .X(_04270_));
 sky130_fd_sc_hd__a221o_1 _09838_ (.A1(net261),
    .A2(_04257_),
    .B1(_04259_),
    .B2(net656),
    .C1(_04270_),
    .X(_00312_));
 sky130_fd_sc_hd__and2_1 _09839_ (.A(_04269_),
    .B(\genblk1[2].osc.clkdiv_C.cnt[13] ),
    .X(_04271_));
 sky130_fd_sc_hd__a221o_1 _09840_ (.A1(\genblk2[2].wave_shpr.div.quo[22] ),
    .A2(_04247_),
    .B1(_04259_),
    .B2(net261),
    .C1(_04271_),
    .X(_00313_));
 sky130_fd_sc_hd__and2_1 _09841_ (.A(_04269_),
    .B(\genblk1[2].osc.clkdiv_C.cnt[14] ),
    .X(_04272_));
 sky130_fd_sc_hd__a221o_1 _09842_ (.A1(net520),
    .A2(_04247_),
    .B1(_04250_),
    .B2(net639),
    .C1(_04272_),
    .X(_00314_));
 sky130_fd_sc_hd__and2_1 _09843_ (.A(_04269_),
    .B(\genblk1[2].osc.clkdiv_C.cnt[15] ),
    .X(_04273_));
 sky130_fd_sc_hd__a221o_1 _09844_ (.A1(net259),
    .A2(_04247_),
    .B1(_04250_),
    .B2(net520),
    .C1(_04273_),
    .X(_00315_));
 sky130_fd_sc_hd__and2_1 _09845_ (.A(_04269_),
    .B(\genblk1[2].osc.clkdiv_C.cnt[16] ),
    .X(_04274_));
 sky130_fd_sc_hd__a221o_1 _09846_ (.A1(\genblk2[2].wave_shpr.div.acc_next[0] ),
    .A2(_04247_),
    .B1(_04250_),
    .B2(net259),
    .C1(_04274_),
    .X(_00316_));
 sky130_fd_sc_hd__inv_2 _09847_ (.A(_04250_),
    .Y(_04275_));
 sky130_fd_sc_hd__nand2_1 _09848_ (.A(_03702_),
    .B(_01416_),
    .Y(_04276_));
 sky130_fd_sc_hd__o221a_1 _09849_ (.A1(\genblk2[2].wave_shpr.div.acc[0] ),
    .A2(_00008_),
    .B1(_04275_),
    .B2(net914),
    .C1(_04276_),
    .X(_00317_));
 sky130_fd_sc_hd__a21oi_1 _09850_ (.A1(\genblk2[2].wave_shpr.div.b1[0] ),
    .A2(_04214_),
    .B1(\genblk2[2].wave_shpr.div.acc[0] ),
    .Y(_04277_));
 sky130_fd_sc_hd__a31o_1 _09851_ (.A1(\genblk2[2].wave_shpr.div.b1[0] ),
    .A2(\genblk2[2].wave_shpr.div.acc[0] ),
    .A3(_04214_),
    .B1(_04275_),
    .X(_04278_));
 sky130_fd_sc_hd__a2bb2o_1 _09852_ (.A1_N(_04277_),
    .A2_N(_04278_),
    .B1(net782),
    .B2(_04248_),
    .X(_00318_));
 sky130_fd_sc_hd__or2_1 _09853_ (.A(\genblk2[2].wave_shpr.div.acc[1] ),
    .B(_04213_),
    .X(_04279_));
 sky130_fd_sc_hd__xnor2_1 _09854_ (.A(_04174_),
    .B(_04175_),
    .Y(_04280_));
 sky130_fd_sc_hd__nand2_1 _09855_ (.A(_04214_),
    .B(_04280_),
    .Y(_04281_));
 sky130_fd_sc_hd__a32o_1 _09856_ (.A1(_04251_),
    .A2(_04279_),
    .A3(_04281_),
    .B1(_04253_),
    .B2(net1137),
    .X(_00319_));
 sky130_fd_sc_hd__clkbuf_4 _09857_ (.A(_04247_),
    .X(_04282_));
 sky130_fd_sc_hd__xor2_1 _09858_ (.A(\genblk2[2].wave_shpr.div.b1[2] ),
    .B(\genblk2[2].wave_shpr.div.acc[2] ),
    .X(_04283_));
 sky130_fd_sc_hd__xnor2_1 _09859_ (.A(_04176_),
    .B(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__mux2_1 _09860_ (.A0(\genblk2[2].wave_shpr.div.acc[2] ),
    .A1(_04284_),
    .S(_04214_),
    .X(_04285_));
 sky130_fd_sc_hd__a22o_1 _09861_ (.A1(net918),
    .A2(_04282_),
    .B1(_04252_),
    .B2(_04285_),
    .X(_00320_));
 sky130_fd_sc_hd__or2b_1 _09862_ (.A(_04179_),
    .B_N(_04170_),
    .X(_04286_));
 sky130_fd_sc_hd__xnor2_1 _09863_ (.A(_04178_),
    .B(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__mux2_1 _09864_ (.A0(\genblk2[2].wave_shpr.div.acc[3] ),
    .A1(_04287_),
    .S(_04214_),
    .X(_04288_));
 sky130_fd_sc_hd__a22o_1 _09865_ (.A1(net975),
    .A2(_04282_),
    .B1(_04252_),
    .B2(_04288_),
    .X(_00321_));
 sky130_fd_sc_hd__clkbuf_4 _09866_ (.A(_04250_),
    .X(_04289_));
 sky130_fd_sc_hd__or2b_1 _09867_ (.A(_04181_),
    .B_N(_04169_),
    .X(_04290_));
 sky130_fd_sc_hd__xnor2_1 _09868_ (.A(_04290_),
    .B(_04180_),
    .Y(_04291_));
 sky130_fd_sc_hd__mux2_1 _09869_ (.A0(\genblk2[2].wave_shpr.div.acc[4] ),
    .A1(_04291_),
    .S(_04214_),
    .X(_04292_));
 sky130_fd_sc_hd__a22o_1 _09870_ (.A1(net919),
    .A2(_04282_),
    .B1(_04289_),
    .B2(_04292_),
    .X(_00322_));
 sky130_fd_sc_hd__or2b_1 _09871_ (.A(_04183_),
    .B_N(_04168_),
    .X(_04293_));
 sky130_fd_sc_hd__xnor2_1 _09872_ (.A(_04293_),
    .B(_04182_),
    .Y(_04294_));
 sky130_fd_sc_hd__mux2_1 _09873_ (.A0(\genblk2[2].wave_shpr.div.acc[5] ),
    .A1(_04294_),
    .S(_04214_),
    .X(_04295_));
 sky130_fd_sc_hd__a22o_1 _09874_ (.A1(net887),
    .A2(_04282_),
    .B1(_04289_),
    .B2(_04295_),
    .X(_00323_));
 sky130_fd_sc_hd__or2b_1 _09875_ (.A(_04185_),
    .B_N(_04167_),
    .X(_04296_));
 sky130_fd_sc_hd__xnor2_1 _09876_ (.A(_04184_),
    .B(_04296_),
    .Y(_04297_));
 sky130_fd_sc_hd__mux2_1 _09877_ (.A0(\genblk2[2].wave_shpr.div.acc[6] ),
    .A1(_04297_),
    .S(_04214_),
    .X(_04298_));
 sky130_fd_sc_hd__a22o_1 _09878_ (.A1(net836),
    .A2(_04282_),
    .B1(_04289_),
    .B2(_04298_),
    .X(_00324_));
 sky130_fd_sc_hd__or2b_1 _09879_ (.A(_04187_),
    .B_N(_04166_),
    .X(_04299_));
 sky130_fd_sc_hd__xnor2_1 _09880_ (.A(_04186_),
    .B(_04299_),
    .Y(_04300_));
 sky130_fd_sc_hd__clkbuf_4 _09881_ (.A(_04213_),
    .X(_04301_));
 sky130_fd_sc_hd__mux2_1 _09882_ (.A0(\genblk2[2].wave_shpr.div.acc[7] ),
    .A1(_04300_),
    .S(_04301_),
    .X(_04302_));
 sky130_fd_sc_hd__a22o_1 _09883_ (.A1(net903),
    .A2(_04282_),
    .B1(_04289_),
    .B2(_04302_),
    .X(_00325_));
 sky130_fd_sc_hd__or2b_1 _09884_ (.A(_04189_),
    .B_N(_04165_),
    .X(_04303_));
 sky130_fd_sc_hd__xnor2_1 _09885_ (.A(_04188_),
    .B(_04303_),
    .Y(_04304_));
 sky130_fd_sc_hd__mux2_1 _09886_ (.A0(\genblk2[2].wave_shpr.div.acc[8] ),
    .A1(_04304_),
    .S(_04301_),
    .X(_04305_));
 sky130_fd_sc_hd__a22o_1 _09887_ (.A1(net895),
    .A2(_04282_),
    .B1(_04289_),
    .B2(_04305_),
    .X(_00326_));
 sky130_fd_sc_hd__or2b_1 _09888_ (.A(_04191_),
    .B_N(_04164_),
    .X(_04306_));
 sky130_fd_sc_hd__xnor2_1 _09889_ (.A(_04190_),
    .B(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__mux2_1 _09890_ (.A0(\genblk2[2].wave_shpr.div.acc[9] ),
    .A1(_04307_),
    .S(_04301_),
    .X(_04308_));
 sky130_fd_sc_hd__a22o_1 _09891_ (.A1(net952),
    .A2(_04282_),
    .B1(_04289_),
    .B2(_04308_),
    .X(_00327_));
 sky130_fd_sc_hd__or2b_1 _09892_ (.A(_04193_),
    .B_N(_04163_),
    .X(_04309_));
 sky130_fd_sc_hd__xnor2_1 _09893_ (.A(_04192_),
    .B(_04309_),
    .Y(_04310_));
 sky130_fd_sc_hd__mux2_1 _09894_ (.A0(\genblk2[2].wave_shpr.div.acc[10] ),
    .A1(_04310_),
    .S(_04301_),
    .X(_04311_));
 sky130_fd_sc_hd__a22o_1 _09895_ (.A1(net830),
    .A2(_04282_),
    .B1(_04289_),
    .B2(_04311_),
    .X(_00328_));
 sky130_fd_sc_hd__or2b_1 _09896_ (.A(_04195_),
    .B_N(_04162_),
    .X(_04312_));
 sky130_fd_sc_hd__xnor2_1 _09897_ (.A(_04194_),
    .B(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__mux2_1 _09898_ (.A0(\genblk2[2].wave_shpr.div.acc[11] ),
    .A1(_04313_),
    .S(_04301_),
    .X(_04314_));
 sky130_fd_sc_hd__a22o_1 _09899_ (.A1(net857),
    .A2(_04282_),
    .B1(_04289_),
    .B2(_04314_),
    .X(_00329_));
 sky130_fd_sc_hd__clkbuf_4 _09900_ (.A(_04247_),
    .X(_04315_));
 sky130_fd_sc_hd__or2b_1 _09901_ (.A(_04197_),
    .B_N(_04161_),
    .X(_04316_));
 sky130_fd_sc_hd__xnor2_1 _09902_ (.A(_04196_),
    .B(_04316_),
    .Y(_04317_));
 sky130_fd_sc_hd__mux2_1 _09903_ (.A0(\genblk2[2].wave_shpr.div.acc[12] ),
    .A1(_04317_),
    .S(_04301_),
    .X(_04318_));
 sky130_fd_sc_hd__a22o_1 _09904_ (.A1(net953),
    .A2(_04315_),
    .B1(_04289_),
    .B2(_04318_),
    .X(_00330_));
 sky130_fd_sc_hd__or2b_1 _09905_ (.A(_04199_),
    .B_N(_04160_),
    .X(_04319_));
 sky130_fd_sc_hd__xnor2_1 _09906_ (.A(_04198_),
    .B(_04319_),
    .Y(_04320_));
 sky130_fd_sc_hd__mux2_1 _09907_ (.A0(\genblk2[2].wave_shpr.div.acc[13] ),
    .A1(_04320_),
    .S(_04301_),
    .X(_04321_));
 sky130_fd_sc_hd__a22o_1 _09908_ (.A1(net1002),
    .A2(_04315_),
    .B1(_04289_),
    .B2(_04321_),
    .X(_00331_));
 sky130_fd_sc_hd__clkbuf_4 _09909_ (.A(_04250_),
    .X(_04322_));
 sky130_fd_sc_hd__or2b_1 _09910_ (.A(_04201_),
    .B_N(_04159_),
    .X(_04323_));
 sky130_fd_sc_hd__xnor2_1 _09911_ (.A(_04200_),
    .B(_04323_),
    .Y(_04324_));
 sky130_fd_sc_hd__mux2_1 _09912_ (.A0(\genblk2[2].wave_shpr.div.acc[14] ),
    .A1(_04324_),
    .S(_04301_),
    .X(_04325_));
 sky130_fd_sc_hd__a22o_1 _09913_ (.A1(net1036),
    .A2(_04315_),
    .B1(_04322_),
    .B2(_04325_),
    .X(_00332_));
 sky130_fd_sc_hd__or2b_1 _09914_ (.A(_04203_),
    .B_N(_04158_),
    .X(_04326_));
 sky130_fd_sc_hd__xnor2_1 _09915_ (.A(_04202_),
    .B(_04326_),
    .Y(_04327_));
 sky130_fd_sc_hd__mux2_1 _09916_ (.A0(\genblk2[2].wave_shpr.div.acc[15] ),
    .A1(_04327_),
    .S(_04301_),
    .X(_04328_));
 sky130_fd_sc_hd__a22o_1 _09917_ (.A1(net845),
    .A2(_04315_),
    .B1(_04322_),
    .B2(_04328_),
    .X(_00333_));
 sky130_fd_sc_hd__or2b_1 _09918_ (.A(_04205_),
    .B_N(_04157_),
    .X(_04329_));
 sky130_fd_sc_hd__xnor2_1 _09919_ (.A(_04329_),
    .B(_04204_),
    .Y(_04330_));
 sky130_fd_sc_hd__mux2_1 _09920_ (.A0(\genblk2[2].wave_shpr.div.acc[16] ),
    .A1(_04330_),
    .S(_04301_),
    .X(_04331_));
 sky130_fd_sc_hd__a22o_1 _09921_ (.A1(net788),
    .A2(_04315_),
    .B1(_04322_),
    .B2(_04331_),
    .X(_00334_));
 sky130_fd_sc_hd__or2b_1 _09922_ (.A(_04207_),
    .B_N(_04156_),
    .X(_04332_));
 sky130_fd_sc_hd__xnor2_1 _09923_ (.A(_04206_),
    .B(_04332_),
    .Y(_04333_));
 sky130_fd_sc_hd__mux2_1 _09924_ (.A0(\genblk2[2].wave_shpr.div.acc[17] ),
    .A1(_04333_),
    .S(_04213_),
    .X(_04334_));
 sky130_fd_sc_hd__a22o_1 _09925_ (.A1(net580),
    .A2(_04315_),
    .B1(_04322_),
    .B2(_04334_),
    .X(_00335_));
 sky130_fd_sc_hd__nor4_1 _09926_ (.A(\genblk2[2].wave_shpr.div.acc[25] ),
    .B(\genblk2[2].wave_shpr.div.acc[24] ),
    .C(\genblk2[2].wave_shpr.div.acc[26] ),
    .D(_04212_),
    .Y(_04335_));
 sky130_fd_sc_hd__or2_1 _09927_ (.A(_04209_),
    .B(net22),
    .X(_04336_));
 sky130_fd_sc_hd__o21ai_1 _09928_ (.A1(_04208_),
    .A2(net22),
    .B1(\genblk2[2].wave_shpr.div.acc[18] ),
    .Y(_04337_));
 sky130_fd_sc_hd__nand2_1 _09929_ (.A(_04336_),
    .B(_04337_),
    .Y(_04338_));
 sky130_fd_sc_hd__a22o_1 _09930_ (.A1(net605),
    .A2(_04315_),
    .B1(_04322_),
    .B2(_04338_),
    .X(_00336_));
 sky130_fd_sc_hd__nor2_1 _09931_ (.A(_04210_),
    .B(net22),
    .Y(_04339_));
 sky130_fd_sc_hd__a21o_1 _09932_ (.A1(net605),
    .A2(_04336_),
    .B1(_04339_),
    .X(_04340_));
 sky130_fd_sc_hd__a22o_1 _09933_ (.A1(net648),
    .A2(_04315_),
    .B1(_04322_),
    .B2(_04340_),
    .X(_00337_));
 sky130_fd_sc_hd__xor2_1 _09934_ (.A(\genblk2[2].wave_shpr.div.acc[20] ),
    .B(_04339_),
    .X(_04341_));
 sky130_fd_sc_hd__a22o_1 _09935_ (.A1(net1034),
    .A2(_04315_),
    .B1(_04322_),
    .B2(_04341_),
    .X(_00338_));
 sky130_fd_sc_hd__or3_1 _09936_ (.A(\genblk2[2].wave_shpr.div.acc[20] ),
    .B(_04210_),
    .C(net1351),
    .X(_04342_));
 sky130_fd_sc_hd__or4_1 _09937_ (.A(\genblk2[2].wave_shpr.div.acc[21] ),
    .B(\genblk2[2].wave_shpr.div.acc[20] ),
    .C(_04210_),
    .D(net22),
    .X(_04343_));
 sky130_fd_sc_hd__a21bo_1 _09938_ (.A1(\genblk2[2].wave_shpr.div.acc[21] ),
    .A2(_04342_),
    .B1_N(_04343_),
    .X(_04344_));
 sky130_fd_sc_hd__a22o_1 _09939_ (.A1(net968),
    .A2(_04315_),
    .B1(_04322_),
    .B2(_04344_),
    .X(_00339_));
 sky130_fd_sc_hd__xnor2_1 _09940_ (.A(\genblk2[2].wave_shpr.div.acc[22] ),
    .B(_04343_),
    .Y(_04345_));
 sky130_fd_sc_hd__a22o_1 _09941_ (.A1(net707),
    .A2(_04253_),
    .B1(_04322_),
    .B2(_04345_),
    .X(_00340_));
 sky130_fd_sc_hd__nor2_1 _09942_ (.A(_04212_),
    .B(_04335_),
    .Y(_04346_));
 sky130_fd_sc_hd__a21o_1 _09943_ (.A1(\genblk2[2].wave_shpr.div.acc[23] ),
    .A2(_04211_),
    .B1(_04346_),
    .X(_04347_));
 sky130_fd_sc_hd__a22o_1 _09944_ (.A1(\genblk2[2].wave_shpr.div.acc[24] ),
    .A2(_04253_),
    .B1(_04322_),
    .B2(_04347_),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _09945_ (.A0(_04346_),
    .A1(_04212_),
    .S(\genblk2[2].wave_shpr.div.acc[24] ),
    .X(_04348_));
 sky130_fd_sc_hd__a22o_1 _09946_ (.A1(net1094),
    .A2(_04253_),
    .B1(_04251_),
    .B2(_04348_),
    .X(_00342_));
 sky130_fd_sc_hd__o21ai_1 _09947_ (.A1(\genblk2[2].wave_shpr.div.acc[24] ),
    .A2(_04212_),
    .B1(\genblk2[2].wave_shpr.div.acc[25] ),
    .Y(_04349_));
 sky130_fd_sc_hd__or4b_1 _09948_ (.A(\genblk2[2].wave_shpr.div.acc[25] ),
    .B(_04212_),
    .C(\genblk2[2].wave_shpr.div.acc[24] ),
    .D_N(\genblk2[2].wave_shpr.div.acc[26] ),
    .X(_04350_));
 sky130_fd_sc_hd__nand2_1 _09949_ (.A(_04349_),
    .B(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__a22o_1 _09950_ (.A1(net962),
    .A2(_04253_),
    .B1(_04251_),
    .B2(_04351_),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _09951_ (.A0(_04250_),
    .A1(_04247_),
    .S(\genblk2[2].wave_shpr.div.i[0] ),
    .X(_04352_));
 sky130_fd_sc_hd__clkbuf_1 _09952_ (.A(_04352_),
    .X(_00344_));
 sky130_fd_sc_hd__or2_1 _09953_ (.A(\genblk2[2].wave_shpr.div.i[1] ),
    .B(\genblk2[2].wave_shpr.div.i[0] ),
    .X(_04353_));
 sky130_fd_sc_hd__nand2_1 _09954_ (.A(\genblk2[2].wave_shpr.div.i[1] ),
    .B(\genblk2[2].wave_shpr.div.i[0] ),
    .Y(_04354_));
 sky130_fd_sc_hd__a32o_1 _09955_ (.A1(_04251_),
    .A2(_04353_),
    .A3(_04354_),
    .B1(_04253_),
    .B2(net1110),
    .X(_00345_));
 sky130_fd_sc_hd__a21o_1 _09956_ (.A1(\genblk2[2].wave_shpr.div.i[1] ),
    .A2(\genblk2[2].wave_shpr.div.i[0] ),
    .B1(\genblk2[2].wave_shpr.div.i[2] ),
    .X(_04355_));
 sky130_fd_sc_hd__and3_1 _09957_ (.A(\genblk2[2].wave_shpr.div.i[1] ),
    .B(\genblk2[2].wave_shpr.div.i[0] ),
    .C(\genblk2[2].wave_shpr.div.i[2] ),
    .X(_04356_));
 sky130_fd_sc_hd__inv_2 _09958_ (.A(_04356_),
    .Y(_04357_));
 sky130_fd_sc_hd__a32o_1 _09959_ (.A1(_04251_),
    .A2(_04355_),
    .A3(_04357_),
    .B1(_04253_),
    .B2(net711),
    .X(_00346_));
 sky130_fd_sc_hd__a21oi_1 _09960_ (.A1(_00008_),
    .A2(_04356_),
    .B1(net1123),
    .Y(_04358_));
 sky130_fd_sc_hd__and3_1 _09961_ (.A(\genblk2[2].wave_shpr.div.i[3] ),
    .B(_02163_),
    .C(_04356_),
    .X(_04359_));
 sky130_fd_sc_hd__nor3_1 _09962_ (.A(_03690_),
    .B(_04358_),
    .C(_04359_),
    .Y(_00347_));
 sky130_fd_sc_hd__o21ai_1 _09963_ (.A1(net282),
    .A2(_04359_),
    .B1(_03855_),
    .Y(_04360_));
 sky130_fd_sc_hd__a21oi_1 _09964_ (.A1(net282),
    .A2(_04359_),
    .B1(_04360_),
    .Y(_00348_));
 sky130_fd_sc_hd__or2b_1 _09965_ (.A(\genblk2[3].wave_shpr.div.acc[17] ),
    .B_N(\genblk2[3].wave_shpr.div.b1[17] ),
    .X(_04361_));
 sky130_fd_sc_hd__nor2_1 _09966_ (.A(_04245_),
    .B(\genblk2[3].wave_shpr.div.acc[16] ),
    .Y(_04362_));
 sky130_fd_sc_hd__or2b_1 _09967_ (.A(\genblk2[3].wave_shpr.div.acc[15] ),
    .B_N(\genblk2[3].wave_shpr.div.b1[15] ),
    .X(_04363_));
 sky130_fd_sc_hd__or2b_1 _09968_ (.A(\genblk2[3].wave_shpr.div.acc[14] ),
    .B_N(\genblk2[3].wave_shpr.div.b1[14] ),
    .X(_04364_));
 sky130_fd_sc_hd__or2b_1 _09969_ (.A(\genblk2[3].wave_shpr.div.acc[13] ),
    .B_N(\genblk2[3].wave_shpr.div.b1[13] ),
    .X(_04365_));
 sky130_fd_sc_hd__or2b_1 _09970_ (.A(\genblk2[3].wave_shpr.div.acc[12] ),
    .B_N(\genblk2[3].wave_shpr.div.b1[12] ),
    .X(_04366_));
 sky130_fd_sc_hd__or2b_1 _09971_ (.A(\genblk2[3].wave_shpr.div.acc[11] ),
    .B_N(\genblk2[3].wave_shpr.div.b1[11] ),
    .X(_04367_));
 sky130_fd_sc_hd__or2b_1 _09972_ (.A(\genblk2[3].wave_shpr.div.acc[10] ),
    .B_N(\genblk2[3].wave_shpr.div.b1[10] ),
    .X(_04368_));
 sky130_fd_sc_hd__or2b_1 _09973_ (.A(\genblk2[3].wave_shpr.div.acc[9] ),
    .B_N(\genblk2[3].wave_shpr.div.b1[9] ),
    .X(_04369_));
 sky130_fd_sc_hd__or2b_1 _09974_ (.A(\genblk2[3].wave_shpr.div.acc[8] ),
    .B_N(\genblk2[3].wave_shpr.div.b1[8] ),
    .X(_04370_));
 sky130_fd_sc_hd__or2b_1 _09975_ (.A(\genblk2[3].wave_shpr.div.acc[7] ),
    .B_N(\genblk2[3].wave_shpr.div.b1[7] ),
    .X(_04371_));
 sky130_fd_sc_hd__or2b_1 _09976_ (.A(\genblk2[3].wave_shpr.div.acc[6] ),
    .B_N(\genblk2[3].wave_shpr.div.b1[6] ),
    .X(_04372_));
 sky130_fd_sc_hd__or2b_1 _09977_ (.A(\genblk2[3].wave_shpr.div.acc[5] ),
    .B_N(\genblk2[3].wave_shpr.div.b1[5] ),
    .X(_04373_));
 sky130_fd_sc_hd__or2b_1 _09978_ (.A(\genblk2[3].wave_shpr.div.b1[4] ),
    .B_N(\genblk2[3].wave_shpr.div.acc[4] ),
    .X(_04374_));
 sky130_fd_sc_hd__or2b_1 _09979_ (.A(\genblk2[3].wave_shpr.div.acc[4] ),
    .B_N(\genblk2[3].wave_shpr.div.b1[4] ),
    .X(_04375_));
 sky130_fd_sc_hd__nand2_1 _09980_ (.A(_04374_),
    .B(_04375_),
    .Y(_04376_));
 sky130_fd_sc_hd__or2b_1 _09981_ (.A(\genblk2[3].wave_shpr.div.acc[3] ),
    .B_N(\genblk2[3].wave_shpr.div.b1[3] ),
    .X(_04377_));
 sky130_fd_sc_hd__or2b_1 _09982_ (.A(\genblk2[3].wave_shpr.div.acc[2] ),
    .B_N(\genblk2[3].wave_shpr.div.b1[2] ),
    .X(_04378_));
 sky130_fd_sc_hd__inv_2 _09983_ (.A(\genblk2[3].wave_shpr.div.b1[1] ),
    .Y(_04379_));
 sky130_fd_sc_hd__inv_2 _09984_ (.A(\genblk2[3].wave_shpr.div.acc[0] ),
    .Y(_04380_));
 sky130_fd_sc_hd__xor2_1 _09985_ (.A(\genblk2[3].wave_shpr.div.b1[1] ),
    .B(\genblk2[3].wave_shpr.div.acc[1] ),
    .X(_04381_));
 sky130_fd_sc_hd__a21oi_1 _09986_ (.A1(\genblk2[3].wave_shpr.div.b1[0] ),
    .A2(_04380_),
    .B1(_04381_),
    .Y(_04382_));
 sky130_fd_sc_hd__a21o_1 _09987_ (.A1(_04379_),
    .A2(\genblk2[3].wave_shpr.div.acc[1] ),
    .B1(_04382_),
    .X(_04383_));
 sky130_fd_sc_hd__and2b_1 _09988_ (.A_N(\genblk2[3].wave_shpr.div.b1[2] ),
    .B(\genblk2[3].wave_shpr.div.acc[2] ),
    .X(_04384_));
 sky130_fd_sc_hd__a21o_1 _09989_ (.A1(_04378_),
    .A2(_04383_),
    .B1(_04384_),
    .X(_04385_));
 sky130_fd_sc_hd__and2b_1 _09990_ (.A_N(\genblk2[3].wave_shpr.div.b1[3] ),
    .B(\genblk2[3].wave_shpr.div.acc[3] ),
    .X(_04386_));
 sky130_fd_sc_hd__a21oi_1 _09991_ (.A1(_04377_),
    .A2(_04385_),
    .B1(_04386_),
    .Y(_04387_));
 sky130_fd_sc_hd__o21ai_1 _09992_ (.A1(_04376_),
    .A2(_04387_),
    .B1(_04374_),
    .Y(_04388_));
 sky130_fd_sc_hd__and2b_1 _09993_ (.A_N(\genblk2[3].wave_shpr.div.b1[5] ),
    .B(\genblk2[3].wave_shpr.div.acc[5] ),
    .X(_04389_));
 sky130_fd_sc_hd__a21o_1 _09994_ (.A1(_04373_),
    .A2(_04388_),
    .B1(_04389_),
    .X(_04390_));
 sky130_fd_sc_hd__and2b_1 _09995_ (.A_N(\genblk2[3].wave_shpr.div.b1[6] ),
    .B(\genblk2[3].wave_shpr.div.acc[6] ),
    .X(_04391_));
 sky130_fd_sc_hd__a21o_1 _09996_ (.A1(_04372_),
    .A2(_04390_),
    .B1(_04391_),
    .X(_04392_));
 sky130_fd_sc_hd__and2b_1 _09997_ (.A_N(\genblk2[3].wave_shpr.div.b1[7] ),
    .B(\genblk2[3].wave_shpr.div.acc[7] ),
    .X(_04393_));
 sky130_fd_sc_hd__a21o_1 _09998_ (.A1(_04371_),
    .A2(_04392_),
    .B1(_04393_),
    .X(_04394_));
 sky130_fd_sc_hd__and2b_1 _09999_ (.A_N(\genblk2[3].wave_shpr.div.b1[8] ),
    .B(\genblk2[3].wave_shpr.div.acc[8] ),
    .X(_04395_));
 sky130_fd_sc_hd__a21o_1 _10000_ (.A1(_04370_),
    .A2(_04394_),
    .B1(_04395_),
    .X(_04396_));
 sky130_fd_sc_hd__and2b_1 _10001_ (.A_N(\genblk2[3].wave_shpr.div.b1[9] ),
    .B(\genblk2[3].wave_shpr.div.acc[9] ),
    .X(_04397_));
 sky130_fd_sc_hd__a21o_1 _10002_ (.A1(_04369_),
    .A2(_04396_),
    .B1(_04397_),
    .X(_04398_));
 sky130_fd_sc_hd__and2b_1 _10003_ (.A_N(\genblk2[3].wave_shpr.div.b1[10] ),
    .B(\genblk2[3].wave_shpr.div.acc[10] ),
    .X(_04399_));
 sky130_fd_sc_hd__a21o_1 _10004_ (.A1(_04368_),
    .A2(_04398_),
    .B1(_04399_),
    .X(_04400_));
 sky130_fd_sc_hd__and2b_1 _10005_ (.A_N(\genblk2[3].wave_shpr.div.b1[11] ),
    .B(\genblk2[3].wave_shpr.div.acc[11] ),
    .X(_04401_));
 sky130_fd_sc_hd__a21o_1 _10006_ (.A1(_04367_),
    .A2(_04400_),
    .B1(_04401_),
    .X(_04402_));
 sky130_fd_sc_hd__and2b_1 _10007_ (.A_N(\genblk2[3].wave_shpr.div.b1[12] ),
    .B(\genblk2[3].wave_shpr.div.acc[12] ),
    .X(_04403_));
 sky130_fd_sc_hd__a21o_1 _10008_ (.A1(_04366_),
    .A2(_04402_),
    .B1(_04403_),
    .X(_04404_));
 sky130_fd_sc_hd__and2b_1 _10009_ (.A_N(\genblk2[3].wave_shpr.div.b1[13] ),
    .B(\genblk2[3].wave_shpr.div.acc[13] ),
    .X(_04405_));
 sky130_fd_sc_hd__a21o_1 _10010_ (.A1(_04365_),
    .A2(_04404_),
    .B1(_04405_),
    .X(_04406_));
 sky130_fd_sc_hd__and2b_1 _10011_ (.A_N(\genblk2[3].wave_shpr.div.b1[14] ),
    .B(\genblk2[3].wave_shpr.div.acc[14] ),
    .X(_04407_));
 sky130_fd_sc_hd__a21o_1 _10012_ (.A1(_04364_),
    .A2(_04406_),
    .B1(_04407_),
    .X(_04408_));
 sky130_fd_sc_hd__and2b_1 _10013_ (.A_N(\genblk2[3].wave_shpr.div.b1[15] ),
    .B(\genblk2[3].wave_shpr.div.acc[15] ),
    .X(_04409_));
 sky130_fd_sc_hd__a21oi_1 _10014_ (.A1(_04363_),
    .A2(_04408_),
    .B1(_04409_),
    .Y(_04410_));
 sky130_fd_sc_hd__and2_1 _10015_ (.A(_04245_),
    .B(\genblk2[3].wave_shpr.div.acc[16] ),
    .X(_04411_));
 sky130_fd_sc_hd__o21bai_1 _10016_ (.A1(_04362_),
    .A2(_04410_),
    .B1_N(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__and2b_1 _10017_ (.A_N(\genblk2[3].wave_shpr.div.b1[17] ),
    .B(\genblk2[3].wave_shpr.div.acc[17] ),
    .X(_04413_));
 sky130_fd_sc_hd__a21o_1 _10018_ (.A1(_04361_),
    .A2(_04412_),
    .B1(_04413_),
    .X(_04414_));
 sky130_fd_sc_hd__or2_1 _10019_ (.A(\genblk2[3].wave_shpr.div.acc[18] ),
    .B(_04414_),
    .X(_04415_));
 sky130_fd_sc_hd__or4_1 _10020_ (.A(\genblk2[3].wave_shpr.div.acc[21] ),
    .B(\genblk2[3].wave_shpr.div.acc[20] ),
    .C(\genblk2[3].wave_shpr.div.acc[19] ),
    .D(_04415_),
    .X(_04416_));
 sky130_fd_sc_hd__or2_2 _10021_ (.A(\genblk2[3].wave_shpr.div.acc[22] ),
    .B(_04416_),
    .X(_04417_));
 sky130_fd_sc_hd__or4_2 _10022_ (.A(\genblk2[3].wave_shpr.div.acc[23] ),
    .B(\genblk2[3].wave_shpr.div.acc[25] ),
    .C(\genblk2[3].wave_shpr.div.acc[24] ),
    .D(\genblk2[3].wave_shpr.div.acc[26] ),
    .X(_04418_));
 sky130_fd_sc_hd__or2_1 _10023_ (.A(_04417_),
    .B(_04418_),
    .X(_04419_));
 sky130_fd_sc_hd__buf_4 _10024_ (.A(_04419_),
    .X(_04420_));
 sky130_fd_sc_hd__and3_2 _10025_ (.A(_02170_),
    .B(\genblk2[3].wave_shpr.div.busy ),
    .C(_02172_),
    .X(_04421_));
 sky130_fd_sc_hd__clkbuf_4 _10026_ (.A(_04421_),
    .X(_04422_));
 sky130_fd_sc_hd__mux2_1 _10027_ (.A0(\genblk2[3].wave_shpr.div.fin_quo[0] ),
    .A1(_04420_),
    .S(_04422_),
    .X(_04423_));
 sky130_fd_sc_hd__clkbuf_1 _10028_ (.A(_04423_),
    .X(_00349_));
 sky130_fd_sc_hd__mux2_1 _10029_ (.A0(\genblk2[3].wave_shpr.div.fin_quo[1] ),
    .A1(\genblk2[3].wave_shpr.div.quo[0] ),
    .S(_04422_),
    .X(_04424_));
 sky130_fd_sc_hd__clkbuf_1 _10030_ (.A(_04424_),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _10031_ (.A0(\genblk2[3].wave_shpr.div.fin_quo[2] ),
    .A1(net326),
    .S(_04422_),
    .X(_04425_));
 sky130_fd_sc_hd__clkbuf_1 _10032_ (.A(_04425_),
    .X(_00351_));
 sky130_fd_sc_hd__mux2_1 _10033_ (.A0(\genblk2[3].wave_shpr.div.fin_quo[3] ),
    .A1(\genblk2[3].wave_shpr.div.quo[2] ),
    .S(_04422_),
    .X(_04426_));
 sky130_fd_sc_hd__clkbuf_1 _10034_ (.A(_04426_),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _10035_ (.A0(\genblk2[3].wave_shpr.div.fin_quo[4] ),
    .A1(\genblk2[3].wave_shpr.div.quo[3] ),
    .S(_04422_),
    .X(_04427_));
 sky130_fd_sc_hd__clkbuf_1 _10036_ (.A(_04427_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _10037_ (.A0(\genblk2[3].wave_shpr.div.fin_quo[5] ),
    .A1(\genblk2[3].wave_shpr.div.quo[4] ),
    .S(_04422_),
    .X(_04428_));
 sky130_fd_sc_hd__clkbuf_1 _10038_ (.A(_04428_),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_1 _10039_ (.A0(\genblk2[3].wave_shpr.div.fin_quo[6] ),
    .A1(net1346),
    .S(_04422_),
    .X(_04429_));
 sky130_fd_sc_hd__clkbuf_1 _10040_ (.A(_04429_),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_1 _10041_ (.A0(\genblk2[3].wave_shpr.div.fin_quo[7] ),
    .A1(\genblk2[3].wave_shpr.div.quo[6] ),
    .S(_04422_),
    .X(_04430_));
 sky130_fd_sc_hd__clkbuf_1 _10042_ (.A(_04430_),
    .X(_00356_));
 sky130_fd_sc_hd__o21a_1 _10043_ (.A1(_03732_),
    .A2(net1071),
    .B1(_03733_),
    .X(_00357_));
 sky130_fd_sc_hd__inv_2 _10044_ (.A(net1100),
    .Y(_04431_));
 sky130_fd_sc_hd__o21ai_1 _10045_ (.A1(_03714_),
    .A2(_04431_),
    .B1(_03717_),
    .Y(_00358_));
 sky130_fd_sc_hd__nor2_2 _10046_ (.A(_01325_),
    .B(_01996_),
    .Y(_04432_));
 sky130_fd_sc_hd__a2bb2o_1 _10047_ (.A1_N(_03727_),
    .A2_N(_04432_),
    .B1(net1075),
    .B2(_03687_),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_1 _10048_ (.A0(\genblk2[4].wave_shpr.div.b1[3] ),
    .A1(_01223_),
    .S(_04238_),
    .X(_04433_));
 sky130_fd_sc_hd__clkbuf_1 _10049_ (.A(_04433_),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _10050_ (.A0(net1188),
    .A1(_01248_),
    .S(_04238_),
    .X(_04434_));
 sky130_fd_sc_hd__clkbuf_1 _10051_ (.A(_04434_),
    .X(_00361_));
 sky130_fd_sc_hd__mux2_1 _10052_ (.A0(\genblk2[4].wave_shpr.div.b1[5] ),
    .A1(_01870_),
    .S(_04238_),
    .X(_04435_));
 sky130_fd_sc_hd__clkbuf_1 _10053_ (.A(_04435_),
    .X(_00362_));
 sky130_fd_sc_hd__inv_2 _10054_ (.A(_01557_),
    .Y(_04436_));
 sky130_fd_sc_hd__mux2_1 _10055_ (.A0(net1178),
    .A1(_04436_),
    .S(_04238_),
    .X(_04437_));
 sky130_fd_sc_hd__clkbuf_1 _10056_ (.A(_04437_),
    .X(_00363_));
 sky130_fd_sc_hd__mux2_1 _10057_ (.A0(net1225),
    .A1(_01329_),
    .S(_04238_),
    .X(_04438_));
 sky130_fd_sc_hd__clkbuf_1 _10058_ (.A(_04438_),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _10059_ (.A0(net1206),
    .A1(_01263_),
    .S(_04238_),
    .X(_04439_));
 sky130_fd_sc_hd__clkbuf_1 _10060_ (.A(_04439_),
    .X(_00365_));
 sky130_fd_sc_hd__buf_4 _10061_ (.A(_03701_),
    .X(_04440_));
 sky130_fd_sc_hd__mux2_1 _10062_ (.A0(net1186),
    .A1(_01240_),
    .S(_04440_),
    .X(_04441_));
 sky130_fd_sc_hd__clkbuf_1 _10063_ (.A(_04441_),
    .X(_00366_));
 sky130_fd_sc_hd__mux2_1 _10064_ (.A0(net1232),
    .A1(_01589_),
    .S(_04440_),
    .X(_04442_));
 sky130_fd_sc_hd__clkbuf_1 _10065_ (.A(_04442_),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _10066_ (.A0(net1192),
    .A1(_04229_),
    .S(_04440_),
    .X(_04443_));
 sky130_fd_sc_hd__clkbuf_1 _10067_ (.A(_04443_),
    .X(_00368_));
 sky130_fd_sc_hd__nor2_2 _10068_ (.A(_01325_),
    .B(_01226_),
    .Y(_04444_));
 sky130_fd_sc_hd__mux2_1 _10069_ (.A0(net1205),
    .A1(_04444_),
    .S(_04440_),
    .X(_04445_));
 sky130_fd_sc_hd__clkbuf_1 _10070_ (.A(_04445_),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_1 _10071_ (.A0(net1281),
    .A1(_01595_),
    .S(_04440_),
    .X(_04446_));
 sky130_fd_sc_hd__clkbuf_1 _10072_ (.A(_04446_),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _10073_ (.A0(net1262),
    .A1(_04242_),
    .S(_04440_),
    .X(_04447_));
 sky130_fd_sc_hd__clkbuf_1 _10074_ (.A(_04447_),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _10075_ (.A0(\genblk2[4].wave_shpr.div.b1[15] ),
    .A1(_01365_),
    .S(_04440_),
    .X(_04448_));
 sky130_fd_sc_hd__clkbuf_1 _10076_ (.A(_04448_),
    .X(_00372_));
 sky130_fd_sc_hd__inv_2 _10077_ (.A(net667),
    .Y(_04449_));
 sky130_fd_sc_hd__o21ai_1 _10078_ (.A1(_03714_),
    .A2(_04449_),
    .B1(_03736_),
    .Y(_00373_));
 sky130_fd_sc_hd__and2_1 _10079_ (.A(_03833_),
    .B(net1227),
    .X(_04450_));
 sky130_fd_sc_hd__clkbuf_1 _10080_ (.A(_04450_),
    .X(_00374_));
 sky130_fd_sc_hd__buf_4 _10081_ (.A(_02169_),
    .X(_04451_));
 sky130_fd_sc_hd__clkbuf_4 _10082_ (.A(_04451_),
    .X(_04452_));
 sky130_fd_sc_hd__and3_1 _10083_ (.A(_02170_),
    .B(\genblk2[3].wave_shpr.div.busy ),
    .C(_02167_),
    .X(_04453_));
 sky130_fd_sc_hd__buf_4 _10084_ (.A(_04453_),
    .X(_04454_));
 sky130_fd_sc_hd__a22o_1 _10085_ (.A1(net794),
    .A2(_04452_),
    .B1(_04420_),
    .B2(_04454_),
    .X(_00375_));
 sky130_fd_sc_hd__clkbuf_4 _10086_ (.A(_04453_),
    .X(_04455_));
 sky130_fd_sc_hd__clkbuf_4 _10087_ (.A(_04455_),
    .X(_04456_));
 sky130_fd_sc_hd__a22o_1 _10088_ (.A1(net326),
    .A2(_04452_),
    .B1(_04456_),
    .B2(net794),
    .X(_00376_));
 sky130_fd_sc_hd__a22o_1 _10089_ (.A1(\genblk2[3].wave_shpr.div.quo[2] ),
    .A2(_04452_),
    .B1(_04456_),
    .B2(net326),
    .X(_00377_));
 sky130_fd_sc_hd__a22o_1 _10090_ (.A1(\genblk2[3].wave_shpr.div.quo[3] ),
    .A2(_04452_),
    .B1(_04456_),
    .B2(net737),
    .X(_00378_));
 sky130_fd_sc_hd__a22o_1 _10091_ (.A1(\genblk2[3].wave_shpr.div.quo[4] ),
    .A2(_04452_),
    .B1(_04456_),
    .B2(net779),
    .X(_00379_));
 sky130_fd_sc_hd__a22o_1 _10092_ (.A1(net814),
    .A2(_04452_),
    .B1(_04456_),
    .B2(net849),
    .X(_00380_));
 sky130_fd_sc_hd__a22o_1 _10093_ (.A1(\genblk2[3].wave_shpr.div.quo[6] ),
    .A2(_04452_),
    .B1(_04456_),
    .B2(net814),
    .X(_00381_));
 sky130_fd_sc_hd__a22o_1 _10094_ (.A1(net401),
    .A2(_04452_),
    .B1(_04456_),
    .B2(net820),
    .X(_00382_));
 sky130_fd_sc_hd__a22o_1 _10095_ (.A1(\genblk2[3].wave_shpr.div.quo[8] ),
    .A2(_04452_),
    .B1(_04456_),
    .B2(net401),
    .X(_00383_));
 sky130_fd_sc_hd__clkbuf_4 _10096_ (.A(_04451_),
    .X(_04457_));
 sky130_fd_sc_hd__and2_1 _10097_ (.A(_04269_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[0] ),
    .X(_04458_));
 sky130_fd_sc_hd__a221o_1 _10098_ (.A1(net538),
    .A2(_04457_),
    .B1(_04454_),
    .B2(\genblk2[3].wave_shpr.div.quo[8] ),
    .C1(_04458_),
    .X(_00384_));
 sky130_fd_sc_hd__and2_1 _10099_ (.A(_04269_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[1] ),
    .X(_04459_));
 sky130_fd_sc_hd__a221o_1 _10100_ (.A1(net631),
    .A2(_04457_),
    .B1(_04454_),
    .B2(net538),
    .C1(_04459_),
    .X(_00385_));
 sky130_fd_sc_hd__and2_1 _10101_ (.A(_04269_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[2] ),
    .X(_04460_));
 sky130_fd_sc_hd__a221o_1 _10102_ (.A1(net525),
    .A2(_04457_),
    .B1(_04454_),
    .B2(net631),
    .C1(_04460_),
    .X(_00386_));
 sky130_fd_sc_hd__buf_2 _10103_ (.A(_04451_),
    .X(_04461_));
 sky130_fd_sc_hd__buf_2 _10104_ (.A(_04455_),
    .X(_04462_));
 sky130_fd_sc_hd__and2_1 _10105_ (.A(_04269_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[3] ),
    .X(_04463_));
 sky130_fd_sc_hd__a221o_1 _10106_ (.A1(net387),
    .A2(_04461_),
    .B1(_04462_),
    .B2(net525),
    .C1(_04463_),
    .X(_00387_));
 sky130_fd_sc_hd__and2_1 _10107_ (.A(_04269_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[4] ),
    .X(_04464_));
 sky130_fd_sc_hd__a221o_1 _10108_ (.A1(\genblk2[3].wave_shpr.div.quo[13] ),
    .A2(_04461_),
    .B1(_04462_),
    .B2(net387),
    .C1(_04464_),
    .X(_00388_));
 sky130_fd_sc_hd__clkbuf_2 _10109_ (.A(_04268_),
    .X(_04465_));
 sky130_fd_sc_hd__and2_1 _10110_ (.A(_04465_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[5] ),
    .X(_04466_));
 sky130_fd_sc_hd__a221o_1 _10111_ (.A1(net634),
    .A2(_04461_),
    .B1(_04462_),
    .B2(\genblk2[3].wave_shpr.div.quo[13] ),
    .C1(_04466_),
    .X(_00389_));
 sky130_fd_sc_hd__and2_1 _10112_ (.A(_04465_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[6] ),
    .X(_04467_));
 sky130_fd_sc_hd__a221o_1 _10113_ (.A1(net514),
    .A2(_04461_),
    .B1(_04462_),
    .B2(net634),
    .C1(_04467_),
    .X(_00390_));
 sky130_fd_sc_hd__and2_1 _10114_ (.A(_04465_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[7] ),
    .X(_04468_));
 sky130_fd_sc_hd__a221o_1 _10115_ (.A1(net376),
    .A2(_04461_),
    .B1(_04462_),
    .B2(net514),
    .C1(_04468_),
    .X(_00391_));
 sky130_fd_sc_hd__and2_1 _10116_ (.A(_04465_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[8] ),
    .X(_04469_));
 sky130_fd_sc_hd__a221o_1 _10117_ (.A1(\genblk2[3].wave_shpr.div.quo[17] ),
    .A2(_04461_),
    .B1(_04462_),
    .B2(net376),
    .C1(_04469_),
    .X(_00392_));
 sky130_fd_sc_hd__and2_1 _10118_ (.A(_04465_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[9] ),
    .X(_04470_));
 sky130_fd_sc_hd__a221o_1 _10119_ (.A1(net451),
    .A2(_04461_),
    .B1(_04462_),
    .B2(\genblk2[3].wave_shpr.div.quo[17] ),
    .C1(_04470_),
    .X(_00393_));
 sky130_fd_sc_hd__and2_1 _10120_ (.A(_04465_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[10] ),
    .X(_04471_));
 sky130_fd_sc_hd__a221o_1 _10121_ (.A1(net296),
    .A2(_04461_),
    .B1(_04462_),
    .B2(net451),
    .C1(_04471_),
    .X(_00394_));
 sky130_fd_sc_hd__nor2_1 _10122_ (.A(_04058_),
    .B(_01486_),
    .Y(_04472_));
 sky130_fd_sc_hd__a221o_1 _10123_ (.A1(\genblk2[3].wave_shpr.div.quo[20] ),
    .A2(_04461_),
    .B1(_04462_),
    .B2(net296),
    .C1(_04472_),
    .X(_00395_));
 sky130_fd_sc_hd__and2_1 _10124_ (.A(_04465_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[12] ),
    .X(_04473_));
 sky130_fd_sc_hd__a221o_1 _10125_ (.A1(\genblk2[3].wave_shpr.div.quo[21] ),
    .A2(_04461_),
    .B1(_04462_),
    .B2(net545),
    .C1(_04473_),
    .X(_00396_));
 sky130_fd_sc_hd__and2_1 _10126_ (.A(_04465_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[13] ),
    .X(_04474_));
 sky130_fd_sc_hd__a221o_1 _10127_ (.A1(net529),
    .A2(_04451_),
    .B1(_04455_),
    .B2(net607),
    .C1(_04474_),
    .X(_00397_));
 sky130_fd_sc_hd__and2_1 _10128_ (.A(_04465_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[14] ),
    .X(_04475_));
 sky130_fd_sc_hd__a221o_1 _10129_ (.A1(net490),
    .A2(_04451_),
    .B1(_04455_),
    .B2(net529),
    .C1(_04475_),
    .X(_00398_));
 sky130_fd_sc_hd__and2_1 _10130_ (.A(_04465_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[15] ),
    .X(_04476_));
 sky130_fd_sc_hd__a221o_1 _10131_ (.A1(\genblk2[3].wave_shpr.div.quo[24] ),
    .A2(_04451_),
    .B1(_04455_),
    .B2(net490),
    .C1(_04476_),
    .X(_00399_));
 sky130_fd_sc_hd__buf_2 _10132_ (.A(_04268_),
    .X(_04477_));
 sky130_fd_sc_hd__and2_1 _10133_ (.A(_04477_),
    .B(\genblk1[3].osc.clkdiv_C.cnt[16] ),
    .X(_04478_));
 sky130_fd_sc_hd__a221o_1 _10134_ (.A1(\genblk2[3].wave_shpr.div.acc_next[0] ),
    .A2(_04451_),
    .B1(_04455_),
    .B2(net561),
    .C1(_04478_),
    .X(_00400_));
 sky130_fd_sc_hd__or2b_1 _10135_ (.A(\genblk2[3].wave_shpr.div.acc_next[0] ),
    .B_N(_04455_),
    .X(_04479_));
 sky130_fd_sc_hd__o221a_1 _10136_ (.A1(_03819_),
    .A2(net436),
    .B1(_00010_),
    .B2(\genblk2[3].wave_shpr.div.acc[0] ),
    .C1(_04479_),
    .X(_00401_));
 sky130_fd_sc_hd__nor2_2 _10137_ (.A(_04417_),
    .B(_04418_),
    .Y(_04480_));
 sky130_fd_sc_hd__or3b_1 _10138_ (.A(_04480_),
    .B(_04380_),
    .C_N(\genblk2[3].wave_shpr.div.b1[0] ),
    .X(_04481_));
 sky130_fd_sc_hd__a21o_1 _10139_ (.A1(\genblk2[3].wave_shpr.div.b1[0] ),
    .A2(_04420_),
    .B1(\genblk2[3].wave_shpr.div.acc[0] ),
    .X(_04482_));
 sky130_fd_sc_hd__a32o_1 _10140_ (.A1(_04454_),
    .A2(_04481_),
    .A3(_04482_),
    .B1(_04457_),
    .B2(net1067),
    .X(_00402_));
 sky130_fd_sc_hd__and3_1 _10141_ (.A(\genblk2[3].wave_shpr.div.b1[0] ),
    .B(_04380_),
    .C(_04381_),
    .X(_04483_));
 sky130_fd_sc_hd__nor2_1 _10142_ (.A(_04382_),
    .B(_04483_),
    .Y(_04484_));
 sky130_fd_sc_hd__mux2_1 _10143_ (.A0(\genblk2[3].wave_shpr.div.acc[1] ),
    .A1(_04484_),
    .S(_04420_),
    .X(_04485_));
 sky130_fd_sc_hd__a22o_1 _10144_ (.A1(net976),
    .A2(_04452_),
    .B1(_04456_),
    .B2(_04485_),
    .X(_00403_));
 sky130_fd_sc_hd__clkbuf_4 _10145_ (.A(_04451_),
    .X(_04486_));
 sky130_fd_sc_hd__or2b_1 _10146_ (.A(_04384_),
    .B_N(_04378_),
    .X(_04487_));
 sky130_fd_sc_hd__xnor2_1 _10147_ (.A(_04383_),
    .B(_04487_),
    .Y(_04488_));
 sky130_fd_sc_hd__mux2_1 _10148_ (.A0(net976),
    .A1(_04488_),
    .S(_04420_),
    .X(_04489_));
 sky130_fd_sc_hd__a22o_1 _10149_ (.A1(net1057),
    .A2(_04486_),
    .B1(_04456_),
    .B2(_04489_),
    .X(_00404_));
 sky130_fd_sc_hd__clkbuf_4 _10150_ (.A(_04455_),
    .X(_04490_));
 sky130_fd_sc_hd__or2b_1 _10151_ (.A(_04386_),
    .B_N(_04377_),
    .X(_04491_));
 sky130_fd_sc_hd__xnor2_1 _10152_ (.A(_04385_),
    .B(_04491_),
    .Y(_04492_));
 sky130_fd_sc_hd__mux2_1 _10153_ (.A0(\genblk2[3].wave_shpr.div.acc[3] ),
    .A1(_04492_),
    .S(_04420_),
    .X(_04493_));
 sky130_fd_sc_hd__a22o_1 _10154_ (.A1(net979),
    .A2(_04486_),
    .B1(_04490_),
    .B2(_04493_),
    .X(_00405_));
 sky130_fd_sc_hd__xor2_1 _10155_ (.A(_04376_),
    .B(_04387_),
    .X(_04494_));
 sky130_fd_sc_hd__mux2_1 _10156_ (.A0(\genblk2[3].wave_shpr.div.acc[4] ),
    .A1(_04494_),
    .S(_04420_),
    .X(_04495_));
 sky130_fd_sc_hd__a22o_1 _10157_ (.A1(net963),
    .A2(_04486_),
    .B1(_04490_),
    .B2(_04495_),
    .X(_00406_));
 sky130_fd_sc_hd__or2b_1 _10158_ (.A(_04389_),
    .B_N(_04373_),
    .X(_04496_));
 sky130_fd_sc_hd__xnor2_1 _10159_ (.A(_04496_),
    .B(_04388_),
    .Y(_04497_));
 sky130_fd_sc_hd__mux2_1 _10160_ (.A0(\genblk2[3].wave_shpr.div.acc[5] ),
    .A1(_04497_),
    .S(_04420_),
    .X(_04498_));
 sky130_fd_sc_hd__a22o_1 _10161_ (.A1(net941),
    .A2(_04486_),
    .B1(_04490_),
    .B2(_04498_),
    .X(_00407_));
 sky130_fd_sc_hd__or2b_1 _10162_ (.A(_04391_),
    .B_N(_04372_),
    .X(_04499_));
 sky130_fd_sc_hd__xnor2_1 _10163_ (.A(_04390_),
    .B(_04499_),
    .Y(_04500_));
 sky130_fd_sc_hd__mux2_1 _10164_ (.A0(\genblk2[3].wave_shpr.div.acc[6] ),
    .A1(_04500_),
    .S(_04420_),
    .X(_04501_));
 sky130_fd_sc_hd__a22o_1 _10165_ (.A1(net890),
    .A2(_04486_),
    .B1(_04490_),
    .B2(_04501_),
    .X(_00408_));
 sky130_fd_sc_hd__or2b_1 _10166_ (.A(_04393_),
    .B_N(_04371_),
    .X(_04502_));
 sky130_fd_sc_hd__xnor2_1 _10167_ (.A(_04392_),
    .B(_04502_),
    .Y(_04503_));
 sky130_fd_sc_hd__mux2_1 _10168_ (.A0(\genblk2[3].wave_shpr.div.acc[7] ),
    .A1(_04503_),
    .S(_04420_),
    .X(_04504_));
 sky130_fd_sc_hd__a22o_1 _10169_ (.A1(net966),
    .A2(_04486_),
    .B1(_04490_),
    .B2(_04504_),
    .X(_00409_));
 sky130_fd_sc_hd__or2b_1 _10170_ (.A(_04395_),
    .B_N(_04370_),
    .X(_04505_));
 sky130_fd_sc_hd__xnor2_1 _10171_ (.A(_04394_),
    .B(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hd__buf_4 _10172_ (.A(_04419_),
    .X(_04507_));
 sky130_fd_sc_hd__mux2_1 _10173_ (.A0(\genblk2[3].wave_shpr.div.acc[8] ),
    .A1(_04506_),
    .S(_04507_),
    .X(_04508_));
 sky130_fd_sc_hd__a22o_1 _10174_ (.A1(net796),
    .A2(_04486_),
    .B1(_04490_),
    .B2(_04508_),
    .X(_00410_));
 sky130_fd_sc_hd__or2b_1 _10175_ (.A(_04397_),
    .B_N(_04369_),
    .X(_04509_));
 sky130_fd_sc_hd__xnor2_1 _10176_ (.A(_04396_),
    .B(_04509_),
    .Y(_04510_));
 sky130_fd_sc_hd__mux2_1 _10177_ (.A0(\genblk2[3].wave_shpr.div.acc[9] ),
    .A1(_04510_),
    .S(_04507_),
    .X(_04511_));
 sky130_fd_sc_hd__a22o_1 _10178_ (.A1(net790),
    .A2(_04486_),
    .B1(_04490_),
    .B2(_04511_),
    .X(_00411_));
 sky130_fd_sc_hd__or2b_1 _10179_ (.A(_04399_),
    .B_N(_04368_),
    .X(_04512_));
 sky130_fd_sc_hd__xnor2_1 _10180_ (.A(_04398_),
    .B(_04512_),
    .Y(_04513_));
 sky130_fd_sc_hd__mux2_1 _10181_ (.A0(\genblk2[3].wave_shpr.div.acc[10] ),
    .A1(_04513_),
    .S(_04507_),
    .X(_04514_));
 sky130_fd_sc_hd__a22o_1 _10182_ (.A1(net791),
    .A2(_04486_),
    .B1(_04490_),
    .B2(_04514_),
    .X(_00412_));
 sky130_fd_sc_hd__or2b_1 _10183_ (.A(_04401_),
    .B_N(_04367_),
    .X(_04515_));
 sky130_fd_sc_hd__xnor2_1 _10184_ (.A(_04400_),
    .B(_04515_),
    .Y(_04516_));
 sky130_fd_sc_hd__mux2_1 _10185_ (.A0(\genblk2[3].wave_shpr.div.acc[11] ),
    .A1(_04516_),
    .S(_04507_),
    .X(_04517_));
 sky130_fd_sc_hd__a22o_1 _10186_ (.A1(net942),
    .A2(_04486_),
    .B1(_04490_),
    .B2(_04517_),
    .X(_00413_));
 sky130_fd_sc_hd__clkbuf_4 _10187_ (.A(_04451_),
    .X(_04518_));
 sky130_fd_sc_hd__or2b_1 _10188_ (.A(_04403_),
    .B_N(_04366_),
    .X(_04519_));
 sky130_fd_sc_hd__xnor2_1 _10189_ (.A(_04402_),
    .B(_04519_),
    .Y(_04520_));
 sky130_fd_sc_hd__mux2_1 _10190_ (.A0(\genblk2[3].wave_shpr.div.acc[12] ),
    .A1(_04520_),
    .S(_04507_),
    .X(_04521_));
 sky130_fd_sc_hd__a22o_1 _10191_ (.A1(net1017),
    .A2(_04518_),
    .B1(_04490_),
    .B2(_04521_),
    .X(_00414_));
 sky130_fd_sc_hd__clkbuf_4 _10192_ (.A(_04455_),
    .X(_04522_));
 sky130_fd_sc_hd__or2b_1 _10193_ (.A(_04405_),
    .B_N(_04365_),
    .X(_04523_));
 sky130_fd_sc_hd__xnor2_1 _10194_ (.A(_04404_),
    .B(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__mux2_1 _10195_ (.A0(\genblk2[3].wave_shpr.div.acc[13] ),
    .A1(_04524_),
    .S(_04507_),
    .X(_04525_));
 sky130_fd_sc_hd__a22o_1 _10196_ (.A1(net862),
    .A2(_04518_),
    .B1(_04522_),
    .B2(_04525_),
    .X(_00415_));
 sky130_fd_sc_hd__or2b_1 _10197_ (.A(_04407_),
    .B_N(_04364_),
    .X(_04526_));
 sky130_fd_sc_hd__xnor2_1 _10198_ (.A(_04406_),
    .B(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__mux2_1 _10199_ (.A0(\genblk2[3].wave_shpr.div.acc[14] ),
    .A1(_04527_),
    .S(_04507_),
    .X(_04528_));
 sky130_fd_sc_hd__a22o_1 _10200_ (.A1(net930),
    .A2(_04518_),
    .B1(_04522_),
    .B2(_04528_),
    .X(_00416_));
 sky130_fd_sc_hd__or2b_1 _10201_ (.A(_04409_),
    .B_N(_04363_),
    .X(_04529_));
 sky130_fd_sc_hd__xnor2_1 _10202_ (.A(_04408_),
    .B(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__mux2_1 _10203_ (.A0(\genblk2[3].wave_shpr.div.acc[15] ),
    .A1(_04530_),
    .S(_04507_),
    .X(_04531_));
 sky130_fd_sc_hd__a22o_1 _10204_ (.A1(net1016),
    .A2(_04518_),
    .B1(_04522_),
    .B2(_04531_),
    .X(_00417_));
 sky130_fd_sc_hd__nor2_1 _10205_ (.A(_04411_),
    .B(_04362_),
    .Y(_04532_));
 sky130_fd_sc_hd__xnor2_1 _10206_ (.A(_04532_),
    .B(_04410_),
    .Y(_04533_));
 sky130_fd_sc_hd__mux2_1 _10207_ (.A0(\genblk2[3].wave_shpr.div.acc[16] ),
    .A1(_04533_),
    .S(_04507_),
    .X(_04534_));
 sky130_fd_sc_hd__a22o_1 _10208_ (.A1(net948),
    .A2(_04518_),
    .B1(_04522_),
    .B2(_04534_),
    .X(_00418_));
 sky130_fd_sc_hd__or2b_1 _10209_ (.A(_04413_),
    .B_N(_04361_),
    .X(_04535_));
 sky130_fd_sc_hd__xnor2_1 _10210_ (.A(_04412_),
    .B(_04535_),
    .Y(_04536_));
 sky130_fd_sc_hd__mux2_1 _10211_ (.A0(\genblk2[3].wave_shpr.div.acc[17] ),
    .A1(_04536_),
    .S(_04507_),
    .X(_04537_));
 sky130_fd_sc_hd__a22o_1 _10212_ (.A1(net657),
    .A2(_04518_),
    .B1(_04522_),
    .B2(_04537_),
    .X(_00419_));
 sky130_fd_sc_hd__or2_1 _10213_ (.A(_04415_),
    .B(_04480_),
    .X(_04538_));
 sky130_fd_sc_hd__o21ai_1 _10214_ (.A1(_04414_),
    .A2(_04480_),
    .B1(\genblk2[3].wave_shpr.div.acc[18] ),
    .Y(_04539_));
 sky130_fd_sc_hd__nand2_1 _10215_ (.A(_04538_),
    .B(_04539_),
    .Y(_04540_));
 sky130_fd_sc_hd__a22o_1 _10216_ (.A1(net904),
    .A2(_04518_),
    .B1(_04522_),
    .B2(_04540_),
    .X(_00420_));
 sky130_fd_sc_hd__or2_1 _10217_ (.A(\genblk2[3].wave_shpr.div.acc[19] ),
    .B(_04538_),
    .X(_04541_));
 sky130_fd_sc_hd__a21bo_1 _10218_ (.A1(net904),
    .A2(_04415_),
    .B1_N(_04541_),
    .X(_04542_));
 sky130_fd_sc_hd__a22o_1 _10219_ (.A1(net1055),
    .A2(_04518_),
    .B1(_04522_),
    .B2(_04542_),
    .X(_00421_));
 sky130_fd_sc_hd__or2_1 _10220_ (.A(\genblk2[3].wave_shpr.div.acc[20] ),
    .B(_04541_),
    .X(_04543_));
 sky130_fd_sc_hd__nand2_1 _10221_ (.A(\genblk2[3].wave_shpr.div.acc[20] ),
    .B(_04541_),
    .Y(_04544_));
 sky130_fd_sc_hd__nand2_1 _10222_ (.A(_04543_),
    .B(_04544_),
    .Y(_04545_));
 sky130_fd_sc_hd__a22o_1 _10223_ (.A1(net524),
    .A2(_04518_),
    .B1(_04522_),
    .B2(_04545_),
    .X(_00422_));
 sky130_fd_sc_hd__a2bb2o_1 _10224_ (.A1_N(_04416_),
    .A2_N(_04480_),
    .B1(_04543_),
    .B2(net524),
    .X(_04546_));
 sky130_fd_sc_hd__a22o_1 _10225_ (.A1(net710),
    .A2(_04518_),
    .B1(_04522_),
    .B2(_04546_),
    .X(_00423_));
 sky130_fd_sc_hd__and2b_1 _10226_ (.A_N(_04417_),
    .B(_04418_),
    .X(_04547_));
 sky130_fd_sc_hd__a21o_1 _10227_ (.A1(\genblk2[3].wave_shpr.div.acc[22] ),
    .A2(_04416_),
    .B1(_04547_),
    .X(_04548_));
 sky130_fd_sc_hd__a22o_1 _10228_ (.A1(net1000),
    .A2(_04457_),
    .B1(_04522_),
    .B2(_04548_),
    .X(_00424_));
 sky130_fd_sc_hd__nor2_1 _10229_ (.A(\genblk2[3].wave_shpr.div.acc[23] ),
    .B(_04417_),
    .Y(_04549_));
 sky130_fd_sc_hd__and2_1 _10230_ (.A(\genblk2[3].wave_shpr.div.acc[23] ),
    .B(_04417_),
    .X(_04550_));
 sky130_fd_sc_hd__or2_1 _10231_ (.A(_04549_),
    .B(_04550_),
    .X(_04551_));
 sky130_fd_sc_hd__a32o_1 _10232_ (.A1(_04418_),
    .A2(_04454_),
    .A3(_04551_),
    .B1(_04457_),
    .B2(net1064),
    .X(_00425_));
 sky130_fd_sc_hd__inv_2 _10233_ (.A(\genblk2[3].wave_shpr.div.acc[24] ),
    .Y(_04552_));
 sky130_fd_sc_hd__or3b_1 _10234_ (.A(\genblk2[3].wave_shpr.div.acc[24] ),
    .B(_04480_),
    .C_N(_04549_),
    .X(_04553_));
 sky130_fd_sc_hd__o21ai_1 _10235_ (.A1(_04552_),
    .A2(_04549_),
    .B1(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hd__a22o_1 _10236_ (.A1(net1021),
    .A2(_04457_),
    .B1(_04454_),
    .B2(_04554_),
    .X(_00426_));
 sky130_fd_sc_hd__xnor2_1 _10237_ (.A(\genblk2[3].wave_shpr.div.acc[25] ),
    .B(_04553_),
    .Y(_04555_));
 sky130_fd_sc_hd__a22o_1 _10238_ (.A1(net375),
    .A2(_04457_),
    .B1(_04454_),
    .B2(_04555_),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_1 _10239_ (.A0(_04455_),
    .A1(_04451_),
    .S(\genblk2[3].wave_shpr.div.i[0] ),
    .X(_04556_));
 sky130_fd_sc_hd__clkbuf_1 _10240_ (.A(_04556_),
    .X(_00428_));
 sky130_fd_sc_hd__or2_1 _10241_ (.A(\genblk2[3].wave_shpr.div.i[1] ),
    .B(\genblk2[3].wave_shpr.div.i[0] ),
    .X(_04557_));
 sky130_fd_sc_hd__nand2_1 _10242_ (.A(\genblk2[3].wave_shpr.div.i[1] ),
    .B(\genblk2[3].wave_shpr.div.i[0] ),
    .Y(_04558_));
 sky130_fd_sc_hd__a32o_1 _10243_ (.A1(_04454_),
    .A2(_04557_),
    .A3(_04558_),
    .B1(_04457_),
    .B2(net1079),
    .X(_00429_));
 sky130_fd_sc_hd__a21o_1 _10244_ (.A1(\genblk2[3].wave_shpr.div.i[1] ),
    .A2(\genblk2[3].wave_shpr.div.i[0] ),
    .B1(\genblk2[3].wave_shpr.div.i[2] ),
    .X(_04559_));
 sky130_fd_sc_hd__and3_1 _10245_ (.A(\genblk2[3].wave_shpr.div.i[1] ),
    .B(\genblk2[3].wave_shpr.div.i[0] ),
    .C(\genblk2[3].wave_shpr.div.i[2] ),
    .X(_04560_));
 sky130_fd_sc_hd__inv_2 _10246_ (.A(_04560_),
    .Y(_04561_));
 sky130_fd_sc_hd__a32o_1 _10247_ (.A1(_04454_),
    .A2(_04559_),
    .A3(_04561_),
    .B1(_04457_),
    .B2(net725),
    .X(_00430_));
 sky130_fd_sc_hd__a21oi_1 _10248_ (.A1(_00010_),
    .A2(_04560_),
    .B1(net1148),
    .Y(_04562_));
 sky130_fd_sc_hd__and3_1 _10249_ (.A(\genblk2[3].wave_shpr.div.i[3] ),
    .B(_02168_),
    .C(_04560_),
    .X(_04563_));
 sky130_fd_sc_hd__nor3_1 _10250_ (.A(_03690_),
    .B(_04562_),
    .C(_04563_),
    .Y(_00431_));
 sky130_fd_sc_hd__o21ai_1 _10251_ (.A1(net333),
    .A2(_04563_),
    .B1(_03855_),
    .Y(_04564_));
 sky130_fd_sc_hd__a21oi_1 _10252_ (.A1(net333),
    .A2(_04563_),
    .B1(_04564_),
    .Y(_00432_));
 sky130_fd_sc_hd__or2b_1 _10253_ (.A(\genblk2[4].wave_shpr.div.acc[17] ),
    .B_N(\genblk2[4].wave_shpr.div.b1[17] ),
    .X(_04565_));
 sky130_fd_sc_hd__nor2_1 _10254_ (.A(_04449_),
    .B(\genblk2[4].wave_shpr.div.acc[16] ),
    .Y(_04566_));
 sky130_fd_sc_hd__or2b_1 _10255_ (.A(\genblk2[4].wave_shpr.div.acc[15] ),
    .B_N(\genblk2[4].wave_shpr.div.b1[15] ),
    .X(_04567_));
 sky130_fd_sc_hd__or2b_1 _10256_ (.A(\genblk2[4].wave_shpr.div.acc[14] ),
    .B_N(\genblk2[4].wave_shpr.div.b1[14] ),
    .X(_04568_));
 sky130_fd_sc_hd__or2b_1 _10257_ (.A(\genblk2[4].wave_shpr.div.acc[13] ),
    .B_N(\genblk2[4].wave_shpr.div.b1[13] ),
    .X(_04569_));
 sky130_fd_sc_hd__or2b_1 _10258_ (.A(\genblk2[4].wave_shpr.div.acc[12] ),
    .B_N(\genblk2[4].wave_shpr.div.b1[12] ),
    .X(_04570_));
 sky130_fd_sc_hd__or2b_1 _10259_ (.A(\genblk2[4].wave_shpr.div.acc[11] ),
    .B_N(\genblk2[4].wave_shpr.div.b1[11] ),
    .X(_04571_));
 sky130_fd_sc_hd__or2b_1 _10260_ (.A(\genblk2[4].wave_shpr.div.acc[10] ),
    .B_N(\genblk2[4].wave_shpr.div.b1[10] ),
    .X(_04572_));
 sky130_fd_sc_hd__or2b_1 _10261_ (.A(\genblk2[4].wave_shpr.div.acc[9] ),
    .B_N(\genblk2[4].wave_shpr.div.b1[9] ),
    .X(_04573_));
 sky130_fd_sc_hd__or2b_1 _10262_ (.A(\genblk2[4].wave_shpr.div.acc[8] ),
    .B_N(\genblk2[4].wave_shpr.div.b1[8] ),
    .X(_04574_));
 sky130_fd_sc_hd__or2b_1 _10263_ (.A(\genblk2[4].wave_shpr.div.acc[7] ),
    .B_N(\genblk2[4].wave_shpr.div.b1[7] ),
    .X(_04575_));
 sky130_fd_sc_hd__or2b_1 _10264_ (.A(\genblk2[4].wave_shpr.div.acc[6] ),
    .B_N(\genblk2[4].wave_shpr.div.b1[6] ),
    .X(_04576_));
 sky130_fd_sc_hd__or2b_1 _10265_ (.A(\genblk2[4].wave_shpr.div.acc[5] ),
    .B_N(\genblk2[4].wave_shpr.div.b1[5] ),
    .X(_04577_));
 sky130_fd_sc_hd__or2b_1 _10266_ (.A(\genblk2[4].wave_shpr.div.b1[4] ),
    .B_N(\genblk2[4].wave_shpr.div.acc[4] ),
    .X(_04578_));
 sky130_fd_sc_hd__or2b_1 _10267_ (.A(\genblk2[4].wave_shpr.div.acc[4] ),
    .B_N(\genblk2[4].wave_shpr.div.b1[4] ),
    .X(_04579_));
 sky130_fd_sc_hd__nand2_1 _10268_ (.A(_04578_),
    .B(_04579_),
    .Y(_04580_));
 sky130_fd_sc_hd__or2b_1 _10269_ (.A(\genblk2[4].wave_shpr.div.acc[3] ),
    .B_N(\genblk2[4].wave_shpr.div.b1[3] ),
    .X(_04581_));
 sky130_fd_sc_hd__or2b_1 _10270_ (.A(\genblk2[4].wave_shpr.div.acc[2] ),
    .B_N(\genblk2[4].wave_shpr.div.b1[2] ),
    .X(_04582_));
 sky130_fd_sc_hd__inv_2 _10271_ (.A(\genblk2[4].wave_shpr.div.acc[0] ),
    .Y(_04583_));
 sky130_fd_sc_hd__xor2_1 _10272_ (.A(\genblk2[4].wave_shpr.div.b1[1] ),
    .B(\genblk2[4].wave_shpr.div.acc[1] ),
    .X(_04584_));
 sky130_fd_sc_hd__a21oi_1 _10273_ (.A1(\genblk2[4].wave_shpr.div.b1[0] ),
    .A2(_04583_),
    .B1(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__a21o_1 _10274_ (.A1(_04431_),
    .A2(\genblk2[4].wave_shpr.div.acc[1] ),
    .B1(_04585_),
    .X(_04586_));
 sky130_fd_sc_hd__and2b_1 _10275_ (.A_N(\genblk2[4].wave_shpr.div.b1[2] ),
    .B(\genblk2[4].wave_shpr.div.acc[2] ),
    .X(_04587_));
 sky130_fd_sc_hd__a21o_1 _10276_ (.A1(_04582_),
    .A2(_04586_),
    .B1(_04587_),
    .X(_04588_));
 sky130_fd_sc_hd__and2b_1 _10277_ (.A_N(\genblk2[4].wave_shpr.div.b1[3] ),
    .B(\genblk2[4].wave_shpr.div.acc[3] ),
    .X(_04589_));
 sky130_fd_sc_hd__a21oi_1 _10278_ (.A1(_04581_),
    .A2(_04588_),
    .B1(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__o21ai_1 _10279_ (.A1(_04580_),
    .A2(_04590_),
    .B1(_04578_),
    .Y(_04591_));
 sky130_fd_sc_hd__and2b_1 _10280_ (.A_N(\genblk2[4].wave_shpr.div.b1[5] ),
    .B(\genblk2[4].wave_shpr.div.acc[5] ),
    .X(_04592_));
 sky130_fd_sc_hd__a21o_1 _10281_ (.A1(_04577_),
    .A2(_04591_),
    .B1(_04592_),
    .X(_04593_));
 sky130_fd_sc_hd__and2b_1 _10282_ (.A_N(\genblk2[4].wave_shpr.div.b1[6] ),
    .B(\genblk2[4].wave_shpr.div.acc[6] ),
    .X(_04594_));
 sky130_fd_sc_hd__a21o_1 _10283_ (.A1(_04576_),
    .A2(_04593_),
    .B1(_04594_),
    .X(_04595_));
 sky130_fd_sc_hd__and2b_1 _10284_ (.A_N(\genblk2[4].wave_shpr.div.b1[7] ),
    .B(\genblk2[4].wave_shpr.div.acc[7] ),
    .X(_04596_));
 sky130_fd_sc_hd__a21o_1 _10285_ (.A1(_04575_),
    .A2(_04595_),
    .B1(_04596_),
    .X(_04597_));
 sky130_fd_sc_hd__and2b_1 _10286_ (.A_N(\genblk2[4].wave_shpr.div.b1[8] ),
    .B(\genblk2[4].wave_shpr.div.acc[8] ),
    .X(_04598_));
 sky130_fd_sc_hd__a21o_1 _10287_ (.A1(_04574_),
    .A2(_04597_),
    .B1(_04598_),
    .X(_04599_));
 sky130_fd_sc_hd__and2b_1 _10288_ (.A_N(\genblk2[4].wave_shpr.div.b1[9] ),
    .B(\genblk2[4].wave_shpr.div.acc[9] ),
    .X(_04600_));
 sky130_fd_sc_hd__a21o_1 _10289_ (.A1(_04573_),
    .A2(_04599_),
    .B1(_04600_),
    .X(_04601_));
 sky130_fd_sc_hd__and2b_1 _10290_ (.A_N(\genblk2[4].wave_shpr.div.b1[10] ),
    .B(\genblk2[4].wave_shpr.div.acc[10] ),
    .X(_04602_));
 sky130_fd_sc_hd__a21o_1 _10291_ (.A1(_04572_),
    .A2(_04601_),
    .B1(_04602_),
    .X(_04603_));
 sky130_fd_sc_hd__and2b_1 _10292_ (.A_N(\genblk2[4].wave_shpr.div.b1[11] ),
    .B(\genblk2[4].wave_shpr.div.acc[11] ),
    .X(_04604_));
 sky130_fd_sc_hd__a21o_1 _10293_ (.A1(_04571_),
    .A2(_04603_),
    .B1(_04604_),
    .X(_04605_));
 sky130_fd_sc_hd__and2b_1 _10294_ (.A_N(\genblk2[4].wave_shpr.div.b1[12] ),
    .B(\genblk2[4].wave_shpr.div.acc[12] ),
    .X(_04606_));
 sky130_fd_sc_hd__a21o_1 _10295_ (.A1(_04570_),
    .A2(_04605_),
    .B1(_04606_),
    .X(_04607_));
 sky130_fd_sc_hd__and2b_1 _10296_ (.A_N(\genblk2[4].wave_shpr.div.b1[13] ),
    .B(\genblk2[4].wave_shpr.div.acc[13] ),
    .X(_04608_));
 sky130_fd_sc_hd__a21o_1 _10297_ (.A1(_04569_),
    .A2(_04607_),
    .B1(_04608_),
    .X(_04609_));
 sky130_fd_sc_hd__and2b_1 _10298_ (.A_N(\genblk2[4].wave_shpr.div.b1[14] ),
    .B(\genblk2[4].wave_shpr.div.acc[14] ),
    .X(_04610_));
 sky130_fd_sc_hd__a21o_1 _10299_ (.A1(_04568_),
    .A2(_04609_),
    .B1(_04610_),
    .X(_04611_));
 sky130_fd_sc_hd__and2b_1 _10300_ (.A_N(\genblk2[4].wave_shpr.div.b1[15] ),
    .B(\genblk2[4].wave_shpr.div.acc[15] ),
    .X(_04612_));
 sky130_fd_sc_hd__a21oi_1 _10301_ (.A1(_04567_),
    .A2(_04611_),
    .B1(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hd__and2_1 _10302_ (.A(_04449_),
    .B(\genblk2[4].wave_shpr.div.acc[16] ),
    .X(_04614_));
 sky130_fd_sc_hd__o21bai_2 _10303_ (.A1(_04566_),
    .A2(_04613_),
    .B1_N(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__and2b_1 _10304_ (.A_N(\genblk2[4].wave_shpr.div.b1[17] ),
    .B(\genblk2[4].wave_shpr.div.acc[17] ),
    .X(_04616_));
 sky130_fd_sc_hd__a21o_1 _10305_ (.A1(_04565_),
    .A2(_04615_),
    .B1(_04616_),
    .X(_04617_));
 sky130_fd_sc_hd__or2_1 _10306_ (.A(\genblk2[4].wave_shpr.div.acc[19] ),
    .B(\genblk2[4].wave_shpr.div.acc[18] ),
    .X(_04618_));
 sky130_fd_sc_hd__or4_1 _10307_ (.A(\genblk2[4].wave_shpr.div.acc[21] ),
    .B(\genblk2[4].wave_shpr.div.acc[20] ),
    .C(_04617_),
    .D(_04618_),
    .X(_04619_));
 sky130_fd_sc_hd__or2_1 _10308_ (.A(\genblk2[4].wave_shpr.div.acc[22] ),
    .B(_04619_),
    .X(_04620_));
 sky130_fd_sc_hd__nor2_1 _10309_ (.A(\genblk2[4].wave_shpr.div.acc[23] ),
    .B(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hd__or4b_4 _10310_ (.A(\genblk2[4].wave_shpr.div.acc[25] ),
    .B(\genblk2[4].wave_shpr.div.acc[24] ),
    .C(\genblk2[4].wave_shpr.div.acc[26] ),
    .D_N(_04621_),
    .X(_04622_));
 sky130_fd_sc_hd__clkbuf_4 _10311_ (.A(_04622_),
    .X(_04623_));
 sky130_fd_sc_hd__mux2_1 _10312_ (.A0(\genblk2[4].wave_shpr.div.fin_quo[0] ),
    .A1(_04623_),
    .S(_00013_),
    .X(_04624_));
 sky130_fd_sc_hd__clkbuf_1 _10313_ (.A(_04624_),
    .X(_00433_));
 sky130_fd_sc_hd__mux2_1 _10314_ (.A0(\genblk2[4].wave_shpr.div.fin_quo[1] ),
    .A1(net1309),
    .S(_00013_),
    .X(_04625_));
 sky130_fd_sc_hd__clkbuf_1 _10315_ (.A(_04625_),
    .X(_00434_));
 sky130_fd_sc_hd__mux2_1 _10316_ (.A0(\genblk2[4].wave_shpr.div.fin_quo[2] ),
    .A1(\genblk2[4].wave_shpr.div.quo[1] ),
    .S(_00013_),
    .X(_04626_));
 sky130_fd_sc_hd__clkbuf_1 _10317_ (.A(_04626_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _10318_ (.A0(\genblk2[4].wave_shpr.div.fin_quo[3] ),
    .A1(\genblk2[4].wave_shpr.div.quo[2] ),
    .S(_00013_),
    .X(_04627_));
 sky130_fd_sc_hd__clkbuf_1 _10319_ (.A(_04627_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _10320_ (.A0(\genblk2[4].wave_shpr.div.fin_quo[4] ),
    .A1(net1333),
    .S(_00013_),
    .X(_04628_));
 sky130_fd_sc_hd__clkbuf_1 _10321_ (.A(_04628_),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _10322_ (.A0(\genblk2[4].wave_shpr.div.fin_quo[5] ),
    .A1(\genblk2[4].wave_shpr.div.quo[4] ),
    .S(_00013_),
    .X(_04629_));
 sky130_fd_sc_hd__clkbuf_1 _10323_ (.A(_04629_),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _10324_ (.A0(\genblk2[4].wave_shpr.div.fin_quo[6] ),
    .A1(\genblk2[4].wave_shpr.div.quo[5] ),
    .S(_00013_),
    .X(_04630_));
 sky130_fd_sc_hd__clkbuf_1 _10325_ (.A(_04630_),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _10326_ (.A0(\genblk2[4].wave_shpr.div.fin_quo[7] ),
    .A1(net1263),
    .S(_00013_),
    .X(_04631_));
 sky130_fd_sc_hd__clkbuf_1 _10327_ (.A(net1264),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _10328_ (.A0(\genblk2[5].wave_shpr.div.b1[0] ),
    .A1(_01735_),
    .S(_04440_),
    .X(_04632_));
 sky130_fd_sc_hd__clkbuf_1 _10329_ (.A(_04632_),
    .X(_00441_));
 sky130_fd_sc_hd__inv_2 _10330_ (.A(\genblk2[5].wave_shpr.div.b1[1] ),
    .Y(_04633_));
 sky130_fd_sc_hd__mux2_1 _10331_ (.A0(_04633_),
    .A1(_01304_),
    .S(_03689_),
    .X(_04634_));
 sky130_fd_sc_hd__nand2_1 _10332_ (.A(_03717_),
    .B(_04634_),
    .Y(_00442_));
 sky130_fd_sc_hd__o22a_1 _10333_ (.A1(_03714_),
    .A2(net692),
    .B1(_01262_),
    .B2(_03705_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _10334_ (.A0(net1212),
    .A1(_01240_),
    .S(_04440_),
    .X(_04635_));
 sky130_fd_sc_hd__clkbuf_1 _10335_ (.A(_04635_),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _10336_ (.A0(net1287),
    .A1(_01256_),
    .S(_04440_),
    .X(_04636_));
 sky130_fd_sc_hd__clkbuf_1 _10337_ (.A(_04636_),
    .X(_00445_));
 sky130_fd_sc_hd__a21bo_1 _10338_ (.A1(_03831_),
    .A2(net625),
    .B1_N(_03733_),
    .X(_00446_));
 sky130_fd_sc_hd__o21a_1 _10339_ (.A1(_03732_),
    .A2(net708),
    .B1(_03717_),
    .X(_00447_));
 sky130_fd_sc_hd__o22a_1 _10340_ (.A1(_03714_),
    .A2(net1097),
    .B1(_04432_),
    .B2(_03727_),
    .X(_00448_));
 sky130_fd_sc_hd__buf_4 _10341_ (.A(_03701_),
    .X(_04637_));
 sky130_fd_sc_hd__mux2_1 _10342_ (.A0(\genblk2[5].wave_shpr.div.b1[8] ),
    .A1(_01326_),
    .S(_04637_),
    .X(_04638_));
 sky130_fd_sc_hd__clkbuf_1 _10343_ (.A(_04638_),
    .X(_00449_));
 sky130_fd_sc_hd__inv_2 _10344_ (.A(_01678_),
    .Y(_04639_));
 sky130_fd_sc_hd__mux2_1 _10345_ (.A0(net1303),
    .A1(_04639_),
    .S(_04637_),
    .X(_04640_));
 sky130_fd_sc_hd__clkbuf_1 _10346_ (.A(_04640_),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _10347_ (.A0(net1283),
    .A1(_01658_),
    .S(_04637_),
    .X(_04641_));
 sky130_fd_sc_hd__clkbuf_1 _10348_ (.A(_04641_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _10349_ (.A0(net1266),
    .A1(_01757_),
    .S(_04637_),
    .X(_04642_));
 sky130_fd_sc_hd__clkbuf_1 _10350_ (.A(_04642_),
    .X(_00452_));
 sky130_fd_sc_hd__inv_2 _10351_ (.A(_01355_),
    .Y(_04643_));
 sky130_fd_sc_hd__mux2_1 _10352_ (.A0(net1279),
    .A1(_04643_),
    .S(_04637_),
    .X(_04644_));
 sky130_fd_sc_hd__clkbuf_1 _10353_ (.A(_04644_),
    .X(_00453_));
 sky130_fd_sc_hd__nor2_1 _10354_ (.A(_01490_),
    .B(_01242_),
    .Y(_04645_));
 sky130_fd_sc_hd__mux2_1 _10355_ (.A0(\genblk2[5].wave_shpr.div.b1[13] ),
    .A1(_04645_),
    .S(_04637_),
    .X(_04646_));
 sky130_fd_sc_hd__clkbuf_1 _10356_ (.A(_04646_),
    .X(_00454_));
 sky130_fd_sc_hd__and3_4 _10357_ (.A(_03708_),
    .B(_01441_),
    .C(_01367_),
    .X(_04647_));
 sky130_fd_sc_hd__a21o_1 _10358_ (.A1(_03704_),
    .A2(net800),
    .B1(_04647_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _10359_ (.A0(\genblk2[5].wave_shpr.div.b1[15] ),
    .A1(_01365_),
    .S(_04637_),
    .X(_04648_));
 sky130_fd_sc_hd__clkbuf_1 _10360_ (.A(_04648_),
    .X(_00456_));
 sky130_fd_sc_hd__inv_2 _10361_ (.A(net834),
    .Y(_04649_));
 sky130_fd_sc_hd__o21ai_1 _10362_ (.A1(_03726_),
    .A2(_04649_),
    .B1(_03736_),
    .Y(_00457_));
 sky130_fd_sc_hd__and2_1 _10363_ (.A(_03833_),
    .B(net1223),
    .X(_04650_));
 sky130_fd_sc_hd__clkbuf_1 _10364_ (.A(_04650_),
    .X(_00458_));
 sky130_fd_sc_hd__clkbuf_4 _10365_ (.A(_02177_),
    .X(_04651_));
 sky130_fd_sc_hd__buf_2 _10366_ (.A(_04651_),
    .X(_04652_));
 sky130_fd_sc_hd__and3_1 _10367_ (.A(_02152_),
    .B(\genblk2[4].wave_shpr.div.busy ),
    .C(_02175_),
    .X(_04653_));
 sky130_fd_sc_hd__clkbuf_4 _10368_ (.A(_04653_),
    .X(_04654_));
 sky130_fd_sc_hd__clkbuf_4 _10369_ (.A(_04654_),
    .X(_04655_));
 sky130_fd_sc_hd__a22o_1 _10370_ (.A1(net418),
    .A2(_04652_),
    .B1(_04623_),
    .B2(_04655_),
    .X(_00459_));
 sky130_fd_sc_hd__buf_2 _10371_ (.A(_04654_),
    .X(_04656_));
 sky130_fd_sc_hd__a22o_1 _10372_ (.A1(\genblk2[4].wave_shpr.div.quo[1] ),
    .A2(_04652_),
    .B1(_04656_),
    .B2(net418),
    .X(_00460_));
 sky130_fd_sc_hd__a22o_1 _10373_ (.A1(\genblk2[4].wave_shpr.div.quo[2] ),
    .A2(_04652_),
    .B1(_04656_),
    .B2(net464),
    .X(_00461_));
 sky130_fd_sc_hd__a22o_1 _10374_ (.A1(net732),
    .A2(_04652_),
    .B1(_04656_),
    .B2(net793),
    .X(_00462_));
 sky130_fd_sc_hd__a22o_1 _10375_ (.A1(\genblk2[4].wave_shpr.div.quo[4] ),
    .A2(_04652_),
    .B1(_04656_),
    .B2(net732),
    .X(_00463_));
 sky130_fd_sc_hd__a22o_1 _10376_ (.A1(\genblk2[4].wave_shpr.div.quo[5] ),
    .A2(_04652_),
    .B1(_04656_),
    .B2(net749),
    .X(_00464_));
 sky130_fd_sc_hd__a22o_1 _10377_ (.A1(net508),
    .A2(_04652_),
    .B1(_04656_),
    .B2(net781),
    .X(_00465_));
 sky130_fd_sc_hd__a22o_1 _10378_ (.A1(net408),
    .A2(_04652_),
    .B1(_04656_),
    .B2(net508),
    .X(_00466_));
 sky130_fd_sc_hd__a22o_1 _10379_ (.A1(net251),
    .A2(_04652_),
    .B1(_04656_),
    .B2(net408),
    .X(_00467_));
 sky130_fd_sc_hd__clkbuf_4 _10380_ (.A(_04651_),
    .X(_04657_));
 sky130_fd_sc_hd__and2_1 _10381_ (.A(_04477_),
    .B(\genblk1[4].osc.clkdiv_C.cnt[0] ),
    .X(_04658_));
 sky130_fd_sc_hd__a221o_1 _10382_ (.A1(\genblk2[4].wave_shpr.div.quo[9] ),
    .A2(_04657_),
    .B1(_04655_),
    .B2(net251),
    .C1(_04658_),
    .X(_00468_));
 sky130_fd_sc_hd__nor2_1 _10383_ (.A(_04058_),
    .B(_01568_),
    .Y(_04659_));
 sky130_fd_sc_hd__a221o_1 _10384_ (.A1(net672),
    .A2(_04657_),
    .B1(_04655_),
    .B2(\genblk2[4].wave_shpr.div.quo[9] ),
    .C1(_04659_),
    .X(_00469_));
 sky130_fd_sc_hd__and2_1 _10385_ (.A(_04477_),
    .B(\genblk1[4].osc.clkdiv_C.cnt[2] ),
    .X(_04660_));
 sky130_fd_sc_hd__a221o_1 _10386_ (.A1(net602),
    .A2(_04657_),
    .B1(_04655_),
    .B2(\genblk2[4].wave_shpr.div.quo[10] ),
    .C1(_04660_),
    .X(_00470_));
 sky130_fd_sc_hd__buf_2 _10387_ (.A(_04651_),
    .X(_04661_));
 sky130_fd_sc_hd__and2_1 _10388_ (.A(_04477_),
    .B(\genblk1[4].osc.clkdiv_C.cnt[3] ),
    .X(_04662_));
 sky130_fd_sc_hd__a221o_1 _10389_ (.A1(net675),
    .A2(_04661_),
    .B1(_04655_),
    .B2(net602),
    .C1(_04662_),
    .X(_00471_));
 sky130_fd_sc_hd__buf_2 _10390_ (.A(_04654_),
    .X(_04663_));
 sky130_fd_sc_hd__nor2_1 _10391_ (.A(_04058_),
    .B(_01570_),
    .Y(_04664_));
 sky130_fd_sc_hd__a221o_1 _10392_ (.A1(net637),
    .A2(_04661_),
    .B1(_04663_),
    .B2(\genblk2[4].wave_shpr.div.quo[12] ),
    .C1(_04664_),
    .X(_00472_));
 sky130_fd_sc_hd__and2_1 _10393_ (.A(_04477_),
    .B(\genblk1[4].osc.clkdiv_C.cnt[5] ),
    .X(_04665_));
 sky130_fd_sc_hd__a221o_1 _10394_ (.A1(net596),
    .A2(_04661_),
    .B1(_04663_),
    .B2(net637),
    .C1(_04665_),
    .X(_00473_));
 sky130_fd_sc_hd__and2_1 _10395_ (.A(_04477_),
    .B(\genblk1[4].osc.clkdiv_C.cnt[6] ),
    .X(_04666_));
 sky130_fd_sc_hd__a221o_1 _10396_ (.A1(\genblk2[4].wave_shpr.div.quo[15] ),
    .A2(_04661_),
    .B1(_04663_),
    .B2(net596),
    .C1(_04666_),
    .X(_00474_));
 sky130_fd_sc_hd__and2_1 _10397_ (.A(_04477_),
    .B(\genblk1[4].osc.clkdiv_C.cnt[7] ),
    .X(_04667_));
 sky130_fd_sc_hd__a221o_1 _10398_ (.A1(net680),
    .A2(_04661_),
    .B1(_04663_),
    .B2(\genblk2[4].wave_shpr.div.quo[15] ),
    .C1(_04667_),
    .X(_00475_));
 sky130_fd_sc_hd__and2_1 _10399_ (.A(_04477_),
    .B(\genblk1[4].osc.clkdiv_C.cnt[8] ),
    .X(_04668_));
 sky130_fd_sc_hd__a221o_1 _10400_ (.A1(net531),
    .A2(_04661_),
    .B1(_04663_),
    .B2(\genblk2[4].wave_shpr.div.quo[16] ),
    .C1(_04668_),
    .X(_00476_));
 sky130_fd_sc_hd__and2_1 _10401_ (.A(_04477_),
    .B(\genblk1[4].osc.clkdiv_C.cnt[9] ),
    .X(_04669_));
 sky130_fd_sc_hd__a221o_1 _10402_ (.A1(net255),
    .A2(_04661_),
    .B1(_04663_),
    .B2(net531),
    .C1(_04669_),
    .X(_00477_));
 sky130_fd_sc_hd__nor2_1 _10403_ (.A(_04058_),
    .B(_01588_),
    .Y(_04670_));
 sky130_fd_sc_hd__a221o_1 _10404_ (.A1(\genblk2[4].wave_shpr.div.quo[19] ),
    .A2(_04661_),
    .B1(_04663_),
    .B2(net255),
    .C1(_04670_),
    .X(_00478_));
 sky130_fd_sc_hd__and2_1 _10405_ (.A(_04477_),
    .B(\genblk1[4].osc.clkdiv_C.cnt[11] ),
    .X(_04671_));
 sky130_fd_sc_hd__a221o_1 _10406_ (.A1(net626),
    .A2(_04661_),
    .B1(_04663_),
    .B2(net658),
    .C1(_04671_),
    .X(_00479_));
 sky130_fd_sc_hd__buf_2 _10407_ (.A(_04268_),
    .X(_04672_));
 sky130_fd_sc_hd__and2_1 _10408_ (.A(_04672_),
    .B(\genblk1[4].osc.clkdiv_C.cnt[12] ),
    .X(_04673_));
 sky130_fd_sc_hd__a221o_1 _10409_ (.A1(\genblk2[4].wave_shpr.div.quo[21] ),
    .A2(_04661_),
    .B1(_04663_),
    .B2(net626),
    .C1(_04673_),
    .X(_00480_));
 sky130_fd_sc_hd__nor2_1 _10410_ (.A(_04058_),
    .B(_01644_),
    .Y(_04674_));
 sky130_fd_sc_hd__a221o_1 _10411_ (.A1(net665),
    .A2(_04651_),
    .B1(_04663_),
    .B2(\genblk2[4].wave_shpr.div.quo[21] ),
    .C1(_04674_),
    .X(_00481_));
 sky130_fd_sc_hd__and2_1 _10412_ (.A(_04672_),
    .B(\genblk1[4].osc.clkdiv_C.cnt[14] ),
    .X(_04675_));
 sky130_fd_sc_hd__a221o_1 _10413_ (.A1(net698),
    .A2(_04651_),
    .B1(_04654_),
    .B2(net665),
    .C1(_04675_),
    .X(_00482_));
 sky130_fd_sc_hd__buf_6 _10414_ (.A(_03719_),
    .X(_04676_));
 sky130_fd_sc_hd__nor2_1 _10415_ (.A(_04676_),
    .B(_01650_),
    .Y(_04677_));
 sky130_fd_sc_hd__a221o_1 _10416_ (.A1(net714),
    .A2(_04651_),
    .B1(_04654_),
    .B2(net698),
    .C1(_04677_),
    .X(_00483_));
 sky130_fd_sc_hd__and2_1 _10417_ (.A(_04672_),
    .B(\genblk1[4].osc.clkdiv_C.cnt[16] ),
    .X(_04678_));
 sky130_fd_sc_hd__a221o_1 _10418_ (.A1(net643),
    .A2(_04651_),
    .B1(_04654_),
    .B2(\genblk2[4].wave_shpr.div.quo[24] ),
    .C1(_04678_),
    .X(_00484_));
 sky130_fd_sc_hd__inv_2 _10419_ (.A(_04654_),
    .Y(_04679_));
 sky130_fd_sc_hd__or2_1 _10420_ (.A(_03719_),
    .B(\genblk1[4].osc.clkdiv_C.cnt[17] ),
    .X(_04680_));
 sky130_fd_sc_hd__o221a_1 _10421_ (.A1(\genblk2[4].wave_shpr.div.acc[0] ),
    .A2(_00012_),
    .B1(_04679_),
    .B2(net643),
    .C1(_04680_),
    .X(_00485_));
 sky130_fd_sc_hd__a21oi_1 _10422_ (.A1(\genblk2[4].wave_shpr.div.b1[0] ),
    .A2(_04623_),
    .B1(\genblk2[4].wave_shpr.div.acc[0] ),
    .Y(_04681_));
 sky130_fd_sc_hd__a31o_1 _10423_ (.A1(\genblk2[4].wave_shpr.div.b1[0] ),
    .A2(\genblk2[4].wave_shpr.div.acc[0] ),
    .A3(_04623_),
    .B1(_04679_),
    .X(_04682_));
 sky130_fd_sc_hd__a2bb2o_1 _10424_ (.A1_N(_04681_),
    .A2_N(_04682_),
    .B1(net1129),
    .B2(_04652_),
    .X(_00486_));
 sky130_fd_sc_hd__clkbuf_4 _10425_ (.A(_04651_),
    .X(_04683_));
 sky130_fd_sc_hd__and3_1 _10426_ (.A(\genblk2[4].wave_shpr.div.b1[0] ),
    .B(_04583_),
    .C(_04584_),
    .X(_04684_));
 sky130_fd_sc_hd__nor2_1 _10427_ (.A(_04585_),
    .B(_04684_),
    .Y(_04685_));
 sky130_fd_sc_hd__mux2_1 _10428_ (.A0(\genblk2[4].wave_shpr.div.acc[1] ),
    .A1(_04685_),
    .S(_04623_),
    .X(_04686_));
 sky130_fd_sc_hd__a22o_1 _10429_ (.A1(net937),
    .A2(_04683_),
    .B1(_04656_),
    .B2(_04686_),
    .X(_00487_));
 sky130_fd_sc_hd__or2b_1 _10430_ (.A(_04587_),
    .B_N(_04582_),
    .X(_04687_));
 sky130_fd_sc_hd__xnor2_1 _10431_ (.A(_04586_),
    .B(_04687_),
    .Y(_04688_));
 sky130_fd_sc_hd__mux2_1 _10432_ (.A0(\genblk2[4].wave_shpr.div.acc[2] ),
    .A1(_04688_),
    .S(_04623_),
    .X(_04689_));
 sky130_fd_sc_hd__a22o_1 _10433_ (.A1(net1068),
    .A2(_04683_),
    .B1(_04656_),
    .B2(_04689_),
    .X(_00488_));
 sky130_fd_sc_hd__clkbuf_4 _10434_ (.A(_04654_),
    .X(_04690_));
 sky130_fd_sc_hd__or2b_1 _10435_ (.A(_04589_),
    .B_N(_04581_),
    .X(_04691_));
 sky130_fd_sc_hd__xnor2_1 _10436_ (.A(_04588_),
    .B(_04691_),
    .Y(_04692_));
 sky130_fd_sc_hd__mux2_1 _10437_ (.A0(\genblk2[4].wave_shpr.div.acc[3] ),
    .A1(_04692_),
    .S(_04623_),
    .X(_04693_));
 sky130_fd_sc_hd__a22o_1 _10438_ (.A1(net842),
    .A2(_04683_),
    .B1(_04690_),
    .B2(_04693_),
    .X(_00489_));
 sky130_fd_sc_hd__xor2_1 _10439_ (.A(_04580_),
    .B(_04590_),
    .X(_04694_));
 sky130_fd_sc_hd__mux2_1 _10440_ (.A0(\genblk2[4].wave_shpr.div.acc[4] ),
    .A1(_04694_),
    .S(_04623_),
    .X(_04695_));
 sky130_fd_sc_hd__a22o_1 _10441_ (.A1(net970),
    .A2(_04683_),
    .B1(_04690_),
    .B2(_04695_),
    .X(_00490_));
 sky130_fd_sc_hd__or2b_1 _10442_ (.A(_04592_),
    .B_N(_04577_),
    .X(_04696_));
 sky130_fd_sc_hd__xnor2_1 _10443_ (.A(_04696_),
    .B(_04591_),
    .Y(_04697_));
 sky130_fd_sc_hd__mux2_1 _10444_ (.A0(\genblk2[4].wave_shpr.div.acc[5] ),
    .A1(_04697_),
    .S(_04623_),
    .X(_04698_));
 sky130_fd_sc_hd__a22o_1 _10445_ (.A1(net998),
    .A2(_04683_),
    .B1(_04690_),
    .B2(_04698_),
    .X(_00491_));
 sky130_fd_sc_hd__or2b_1 _10446_ (.A(_04594_),
    .B_N(_04576_),
    .X(_04699_));
 sky130_fd_sc_hd__xnor2_1 _10447_ (.A(_04593_),
    .B(_04699_),
    .Y(_04700_));
 sky130_fd_sc_hd__mux2_1 _10448_ (.A0(\genblk2[4].wave_shpr.div.acc[6] ),
    .A1(_04700_),
    .S(_04623_),
    .X(_04701_));
 sky130_fd_sc_hd__a22o_1 _10449_ (.A1(net971),
    .A2(_04683_),
    .B1(_04690_),
    .B2(_04701_),
    .X(_00492_));
 sky130_fd_sc_hd__or2b_1 _10450_ (.A(_04596_),
    .B_N(_04575_),
    .X(_04702_));
 sky130_fd_sc_hd__xnor2_1 _10451_ (.A(_04595_),
    .B(_04702_),
    .Y(_04703_));
 sky130_fd_sc_hd__buf_4 _10452_ (.A(_04622_),
    .X(_04704_));
 sky130_fd_sc_hd__mux2_1 _10453_ (.A0(net1340),
    .A1(_04703_),
    .S(_04704_),
    .X(_04705_));
 sky130_fd_sc_hd__a22o_1 _10454_ (.A1(net891),
    .A2(_04683_),
    .B1(_04690_),
    .B2(_04705_),
    .X(_00493_));
 sky130_fd_sc_hd__or2b_1 _10455_ (.A(_04598_),
    .B_N(_04574_),
    .X(_04706_));
 sky130_fd_sc_hd__xnor2_1 _10456_ (.A(_04597_),
    .B(_04706_),
    .Y(_04707_));
 sky130_fd_sc_hd__mux2_1 _10457_ (.A0(\genblk2[4].wave_shpr.div.acc[8] ),
    .A1(_04707_),
    .S(_04704_),
    .X(_04708_));
 sky130_fd_sc_hd__a22o_1 _10458_ (.A1(net928),
    .A2(_04683_),
    .B1(_04690_),
    .B2(_04708_),
    .X(_00494_));
 sky130_fd_sc_hd__or2b_1 _10459_ (.A(_04600_),
    .B_N(_04573_),
    .X(_04709_));
 sky130_fd_sc_hd__xnor2_1 _10460_ (.A(_04599_),
    .B(_04709_),
    .Y(_04710_));
 sky130_fd_sc_hd__mux2_1 _10461_ (.A0(\genblk2[4].wave_shpr.div.acc[9] ),
    .A1(_04710_),
    .S(_04704_),
    .X(_04711_));
 sky130_fd_sc_hd__a22o_1 _10462_ (.A1(net1024),
    .A2(_04683_),
    .B1(_04690_),
    .B2(_04711_),
    .X(_00495_));
 sky130_fd_sc_hd__or2b_1 _10463_ (.A(_04602_),
    .B_N(_04572_),
    .X(_04712_));
 sky130_fd_sc_hd__xnor2_1 _10464_ (.A(_04601_),
    .B(_04712_),
    .Y(_04713_));
 sky130_fd_sc_hd__mux2_1 _10465_ (.A0(\genblk2[4].wave_shpr.div.acc[10] ),
    .A1(_04713_),
    .S(_04704_),
    .X(_04714_));
 sky130_fd_sc_hd__a22o_1 _10466_ (.A1(net1008),
    .A2(_04683_),
    .B1(_04690_),
    .B2(_04714_),
    .X(_00496_));
 sky130_fd_sc_hd__clkbuf_4 _10467_ (.A(_04651_),
    .X(_04715_));
 sky130_fd_sc_hd__or2b_1 _10468_ (.A(_04604_),
    .B_N(_04571_),
    .X(_04716_));
 sky130_fd_sc_hd__xnor2_1 _10469_ (.A(_04603_),
    .B(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__mux2_1 _10470_ (.A0(\genblk2[4].wave_shpr.div.acc[11] ),
    .A1(_04717_),
    .S(_04704_),
    .X(_04718_));
 sky130_fd_sc_hd__a22o_1 _10471_ (.A1(net778),
    .A2(_04715_),
    .B1(_04690_),
    .B2(_04718_),
    .X(_00497_));
 sky130_fd_sc_hd__or2b_1 _10472_ (.A(_04606_),
    .B_N(_04570_),
    .X(_04719_));
 sky130_fd_sc_hd__xnor2_1 _10473_ (.A(_04605_),
    .B(_04719_),
    .Y(_04720_));
 sky130_fd_sc_hd__mux2_1 _10474_ (.A0(\genblk2[4].wave_shpr.div.acc[12] ),
    .A1(_04720_),
    .S(_04704_),
    .X(_04721_));
 sky130_fd_sc_hd__a22o_1 _10475_ (.A1(net901),
    .A2(_04715_),
    .B1(_04690_),
    .B2(_04721_),
    .X(_00498_));
 sky130_fd_sc_hd__clkbuf_4 _10476_ (.A(_04654_),
    .X(_04722_));
 sky130_fd_sc_hd__or2b_1 _10477_ (.A(_04608_),
    .B_N(_04569_),
    .X(_04723_));
 sky130_fd_sc_hd__xnor2_1 _10478_ (.A(_04607_),
    .B(_04723_),
    .Y(_04724_));
 sky130_fd_sc_hd__mux2_1 _10479_ (.A0(\genblk2[4].wave_shpr.div.acc[13] ),
    .A1(_04724_),
    .S(_04704_),
    .X(_04725_));
 sky130_fd_sc_hd__a22o_1 _10480_ (.A1(net850),
    .A2(_04715_),
    .B1(_04722_),
    .B2(_04725_),
    .X(_00499_));
 sky130_fd_sc_hd__or2b_1 _10481_ (.A(_04610_),
    .B_N(_04568_),
    .X(_04726_));
 sky130_fd_sc_hd__xnor2_1 _10482_ (.A(_04609_),
    .B(_04726_),
    .Y(_04727_));
 sky130_fd_sc_hd__mux2_1 _10483_ (.A0(\genblk2[4].wave_shpr.div.acc[14] ),
    .A1(_04727_),
    .S(_04704_),
    .X(_04728_));
 sky130_fd_sc_hd__a22o_1 _10484_ (.A1(net784),
    .A2(_04715_),
    .B1(_04722_),
    .B2(_04728_),
    .X(_00500_));
 sky130_fd_sc_hd__or2b_1 _10485_ (.A(_04612_),
    .B_N(_04567_),
    .X(_04729_));
 sky130_fd_sc_hd__xnor2_1 _10486_ (.A(_04611_),
    .B(_04729_),
    .Y(_04730_));
 sky130_fd_sc_hd__mux2_1 _10487_ (.A0(\genblk2[4].wave_shpr.div.acc[15] ),
    .A1(_04730_),
    .S(_04704_),
    .X(_04731_));
 sky130_fd_sc_hd__a22o_1 _10488_ (.A1(net881),
    .A2(_04715_),
    .B1(_04722_),
    .B2(_04731_),
    .X(_00501_));
 sky130_fd_sc_hd__nor2_1 _10489_ (.A(_04614_),
    .B(_04566_),
    .Y(_04732_));
 sky130_fd_sc_hd__xnor2_1 _10490_ (.A(_04732_),
    .B(_04613_),
    .Y(_04733_));
 sky130_fd_sc_hd__mux2_1 _10491_ (.A0(\genblk2[4].wave_shpr.div.acc[16] ),
    .A1(_04733_),
    .S(_04704_),
    .X(_04734_));
 sky130_fd_sc_hd__a22o_1 _10492_ (.A1(net926),
    .A2(_04715_),
    .B1(_04722_),
    .B2(_04734_),
    .X(_00502_));
 sky130_fd_sc_hd__or2b_1 _10493_ (.A(_04616_),
    .B_N(_04565_),
    .X(_04735_));
 sky130_fd_sc_hd__xnor2_1 _10494_ (.A(_04615_),
    .B(_04735_),
    .Y(_04736_));
 sky130_fd_sc_hd__mux2_1 _10495_ (.A0(\genblk2[4].wave_shpr.div.acc[17] ),
    .A1(_04736_),
    .S(_04622_),
    .X(_04737_));
 sky130_fd_sc_hd__a22o_1 _10496_ (.A1(net1074),
    .A2(_04715_),
    .B1(_04722_),
    .B2(_04737_),
    .X(_00503_));
 sky130_fd_sc_hd__nand2b_1 _10497_ (.A_N(_04617_),
    .B(_04622_),
    .Y(_04738_));
 sky130_fd_sc_hd__xnor2_1 _10498_ (.A(\genblk2[4].wave_shpr.div.acc[18] ),
    .B(_04738_),
    .Y(_04739_));
 sky130_fd_sc_hd__a22o_1 _10499_ (.A1(net591),
    .A2(_04715_),
    .B1(_04722_),
    .B2(_04739_),
    .X(_00504_));
 sky130_fd_sc_hd__or2_1 _10500_ (.A(_04618_),
    .B(_04738_),
    .X(_04740_));
 sky130_fd_sc_hd__o21ai_1 _10501_ (.A1(\genblk2[4].wave_shpr.div.acc[18] ),
    .A2(_04738_),
    .B1(net591),
    .Y(_04741_));
 sky130_fd_sc_hd__nand2_1 _10502_ (.A(_04740_),
    .B(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__a22o_1 _10503_ (.A1(net694),
    .A2(_04715_),
    .B1(_04722_),
    .B2(_04742_),
    .X(_00505_));
 sky130_fd_sc_hd__xnor2_1 _10504_ (.A(\genblk2[4].wave_shpr.div.acc[20] ),
    .B(_04740_),
    .Y(_04743_));
 sky130_fd_sc_hd__a22o_1 _10505_ (.A1(net472),
    .A2(_04715_),
    .B1(_04722_),
    .B2(_04743_),
    .X(_00506_));
 sky130_fd_sc_hd__or2_1 _10506_ (.A(\genblk2[4].wave_shpr.div.acc[20] ),
    .B(_04740_),
    .X(_04744_));
 sky130_fd_sc_hd__and2b_1 _10507_ (.A_N(_04619_),
    .B(_04622_),
    .X(_04745_));
 sky130_fd_sc_hd__a21o_1 _10508_ (.A1(net472),
    .A2(_04744_),
    .B1(_04745_),
    .X(_04746_));
 sky130_fd_sc_hd__a22o_1 _10509_ (.A1(\genblk2[4].wave_shpr.div.acc[22] ),
    .A2(_04657_),
    .B1(_04722_),
    .B2(_04746_),
    .X(_00507_));
 sky130_fd_sc_hd__mux2_1 _10510_ (.A0(_04745_),
    .A1(_04619_),
    .S(\genblk2[4].wave_shpr.div.acc[22] ),
    .X(_04747_));
 sky130_fd_sc_hd__a22o_1 _10511_ (.A1(net787),
    .A2(_04657_),
    .B1(_04722_),
    .B2(_04747_),
    .X(_00508_));
 sky130_fd_sc_hd__o31a_1 _10512_ (.A1(\genblk2[4].wave_shpr.div.acc[25] ),
    .A2(\genblk2[4].wave_shpr.div.acc[24] ),
    .A3(\genblk2[4].wave_shpr.div.acc[26] ),
    .B1(_04621_),
    .X(_04748_));
 sky130_fd_sc_hd__a21o_1 _10513_ (.A1(\genblk2[4].wave_shpr.div.acc[23] ),
    .A2(_04620_),
    .B1(_04748_),
    .X(_04749_));
 sky130_fd_sc_hd__a22o_1 _10514_ (.A1(net1144),
    .A2(_04657_),
    .B1(_04655_),
    .B2(_04749_),
    .X(_00509_));
 sky130_fd_sc_hd__inv_2 _10515_ (.A(\genblk2[4].wave_shpr.div.acc[24] ),
    .Y(_04750_));
 sky130_fd_sc_hd__nand2_1 _10516_ (.A(_04750_),
    .B(_04748_),
    .Y(_04751_));
 sky130_fd_sc_hd__o21ai_1 _10517_ (.A1(_04750_),
    .A2(_04621_),
    .B1(_04751_),
    .Y(_04752_));
 sky130_fd_sc_hd__a22o_1 _10518_ (.A1(net777),
    .A2(_04657_),
    .B1(_04655_),
    .B2(_04752_),
    .X(_00510_));
 sky130_fd_sc_hd__xnor2_1 _10519_ (.A(\genblk2[4].wave_shpr.div.acc[25] ),
    .B(_04751_),
    .Y(_04753_));
 sky130_fd_sc_hd__a22o_1 _10520_ (.A1(net763),
    .A2(_04657_),
    .B1(_04655_),
    .B2(_04753_),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _10521_ (.A0(_04654_),
    .A1(_04651_),
    .S(\genblk2[4].wave_shpr.div.i[0] ),
    .X(_04754_));
 sky130_fd_sc_hd__clkbuf_1 _10522_ (.A(_04754_),
    .X(_00512_));
 sky130_fd_sc_hd__or2_1 _10523_ (.A(\genblk2[4].wave_shpr.div.i[1] ),
    .B(\genblk2[4].wave_shpr.div.i[0] ),
    .X(_04755_));
 sky130_fd_sc_hd__nand2_1 _10524_ (.A(\genblk2[4].wave_shpr.div.i[1] ),
    .B(\genblk2[4].wave_shpr.div.i[0] ),
    .Y(_04756_));
 sky130_fd_sc_hd__a32o_1 _10525_ (.A1(_04655_),
    .A2(_04755_),
    .A3(_04756_),
    .B1(_04657_),
    .B2(net1108),
    .X(_00513_));
 sky130_fd_sc_hd__a21o_1 _10526_ (.A1(\genblk2[4].wave_shpr.div.i[1] ),
    .A2(\genblk2[4].wave_shpr.div.i[0] ),
    .B1(\genblk2[4].wave_shpr.div.i[2] ),
    .X(_04757_));
 sky130_fd_sc_hd__and3_1 _10527_ (.A(\genblk2[4].wave_shpr.div.i[1] ),
    .B(\genblk2[4].wave_shpr.div.i[0] ),
    .C(\genblk2[4].wave_shpr.div.i[2] ),
    .X(_04758_));
 sky130_fd_sc_hd__inv_2 _10528_ (.A(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hd__a32o_1 _10529_ (.A1(_04655_),
    .A2(_04757_),
    .A3(_04759_),
    .B1(_04657_),
    .B2(net734),
    .X(_00514_));
 sky130_fd_sc_hd__a21oi_1 _10530_ (.A1(_00012_),
    .A2(_04758_),
    .B1(net1160),
    .Y(_04760_));
 sky130_fd_sc_hd__and3_1 _10531_ (.A(\genblk2[4].wave_shpr.div.i[3] ),
    .B(_02176_),
    .C(_04758_),
    .X(_04761_));
 sky130_fd_sc_hd__nor3_1 _10532_ (.A(_03690_),
    .B(_04760_),
    .C(_04761_),
    .Y(_00515_));
 sky130_fd_sc_hd__o21ai_1 _10533_ (.A1(net281),
    .A2(_04761_),
    .B1(_03855_),
    .Y(_04762_));
 sky130_fd_sc_hd__a21oi_1 _10534_ (.A1(net281),
    .A2(_04761_),
    .B1(_04762_),
    .Y(_00516_));
 sky130_fd_sc_hd__or2b_1 _10535_ (.A(\genblk2[5].wave_shpr.div.acc[17] ),
    .B_N(\genblk2[5].wave_shpr.div.b1[17] ),
    .X(_04763_));
 sky130_fd_sc_hd__nor2_1 _10536_ (.A(_04649_),
    .B(\genblk2[5].wave_shpr.div.acc[16] ),
    .Y(_04764_));
 sky130_fd_sc_hd__or2b_1 _10537_ (.A(\genblk2[5].wave_shpr.div.acc[15] ),
    .B_N(\genblk2[5].wave_shpr.div.b1[15] ),
    .X(_04765_));
 sky130_fd_sc_hd__or2b_1 _10538_ (.A(\genblk2[5].wave_shpr.div.acc[14] ),
    .B_N(\genblk2[5].wave_shpr.div.b1[14] ),
    .X(_04766_));
 sky130_fd_sc_hd__or2b_1 _10539_ (.A(\genblk2[5].wave_shpr.div.acc[13] ),
    .B_N(\genblk2[5].wave_shpr.div.b1[13] ),
    .X(_04767_));
 sky130_fd_sc_hd__or2b_1 _10540_ (.A(\genblk2[5].wave_shpr.div.acc[12] ),
    .B_N(\genblk2[5].wave_shpr.div.b1[12] ),
    .X(_04768_));
 sky130_fd_sc_hd__or2b_1 _10541_ (.A(\genblk2[5].wave_shpr.div.acc[11] ),
    .B_N(\genblk2[5].wave_shpr.div.b1[11] ),
    .X(_04769_));
 sky130_fd_sc_hd__or2b_1 _10542_ (.A(\genblk2[5].wave_shpr.div.acc[10] ),
    .B_N(\genblk2[5].wave_shpr.div.b1[10] ),
    .X(_04770_));
 sky130_fd_sc_hd__or2b_1 _10543_ (.A(\genblk2[5].wave_shpr.div.acc[9] ),
    .B_N(\genblk2[5].wave_shpr.div.b1[9] ),
    .X(_04771_));
 sky130_fd_sc_hd__or2b_1 _10544_ (.A(\genblk2[5].wave_shpr.div.acc[8] ),
    .B_N(\genblk2[5].wave_shpr.div.b1[8] ),
    .X(_04772_));
 sky130_fd_sc_hd__or2b_1 _10545_ (.A(\genblk2[5].wave_shpr.div.acc[7] ),
    .B_N(\genblk2[5].wave_shpr.div.b1[7] ),
    .X(_04773_));
 sky130_fd_sc_hd__or2b_1 _10546_ (.A(\genblk2[5].wave_shpr.div.acc[6] ),
    .B_N(\genblk2[5].wave_shpr.div.b1[6] ),
    .X(_04774_));
 sky130_fd_sc_hd__or2b_1 _10547_ (.A(\genblk2[5].wave_shpr.div.acc[5] ),
    .B_N(\genblk2[5].wave_shpr.div.b1[5] ),
    .X(_04775_));
 sky130_fd_sc_hd__or2b_1 _10548_ (.A(\genblk2[5].wave_shpr.div.b1[4] ),
    .B_N(\genblk2[5].wave_shpr.div.acc[4] ),
    .X(_04776_));
 sky130_fd_sc_hd__or2b_1 _10549_ (.A(\genblk2[5].wave_shpr.div.acc[4] ),
    .B_N(\genblk2[5].wave_shpr.div.b1[4] ),
    .X(_04777_));
 sky130_fd_sc_hd__nand2_1 _10550_ (.A(_04776_),
    .B(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__or2b_1 _10551_ (.A(\genblk2[5].wave_shpr.div.acc[3] ),
    .B_N(\genblk2[5].wave_shpr.div.b1[3] ),
    .X(_04779_));
 sky130_fd_sc_hd__or2b_1 _10552_ (.A(\genblk2[5].wave_shpr.div.acc[2] ),
    .B_N(\genblk2[5].wave_shpr.div.b1[2] ),
    .X(_04780_));
 sky130_fd_sc_hd__inv_2 _10553_ (.A(\genblk2[5].wave_shpr.div.acc[0] ),
    .Y(_04781_));
 sky130_fd_sc_hd__xor2_1 _10554_ (.A(\genblk2[5].wave_shpr.div.b1[1] ),
    .B(\genblk2[5].wave_shpr.div.acc[1] ),
    .X(_04782_));
 sky130_fd_sc_hd__a21oi_1 _10555_ (.A1(\genblk2[5].wave_shpr.div.b1[0] ),
    .A2(_04781_),
    .B1(_04782_),
    .Y(_04783_));
 sky130_fd_sc_hd__a21o_1 _10556_ (.A1(_04633_),
    .A2(\genblk2[5].wave_shpr.div.acc[1] ),
    .B1(_04783_),
    .X(_04784_));
 sky130_fd_sc_hd__and2b_1 _10557_ (.A_N(\genblk2[5].wave_shpr.div.b1[2] ),
    .B(\genblk2[5].wave_shpr.div.acc[2] ),
    .X(_04785_));
 sky130_fd_sc_hd__a21o_1 _10558_ (.A1(_04780_),
    .A2(_04784_),
    .B1(_04785_),
    .X(_04786_));
 sky130_fd_sc_hd__and2b_1 _10559_ (.A_N(\genblk2[5].wave_shpr.div.b1[3] ),
    .B(\genblk2[5].wave_shpr.div.acc[3] ),
    .X(_04787_));
 sky130_fd_sc_hd__a21oi_1 _10560_ (.A1(_04779_),
    .A2(_04786_),
    .B1(_04787_),
    .Y(_04788_));
 sky130_fd_sc_hd__o21ai_1 _10561_ (.A1(_04778_),
    .A2(_04788_),
    .B1(_04776_),
    .Y(_04789_));
 sky130_fd_sc_hd__and2b_1 _10562_ (.A_N(\genblk2[5].wave_shpr.div.b1[5] ),
    .B(\genblk2[5].wave_shpr.div.acc[5] ),
    .X(_04790_));
 sky130_fd_sc_hd__a21o_1 _10563_ (.A1(_04775_),
    .A2(_04789_),
    .B1(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__and2b_1 _10564_ (.A_N(\genblk2[5].wave_shpr.div.b1[6] ),
    .B(\genblk2[5].wave_shpr.div.acc[6] ),
    .X(_04792_));
 sky130_fd_sc_hd__a21o_1 _10565_ (.A1(_04774_),
    .A2(_04791_),
    .B1(_04792_),
    .X(_04793_));
 sky130_fd_sc_hd__and2b_1 _10566_ (.A_N(\genblk2[5].wave_shpr.div.b1[7] ),
    .B(\genblk2[5].wave_shpr.div.acc[7] ),
    .X(_04794_));
 sky130_fd_sc_hd__a21o_1 _10567_ (.A1(_04773_),
    .A2(_04793_),
    .B1(_04794_),
    .X(_04795_));
 sky130_fd_sc_hd__and2b_1 _10568_ (.A_N(\genblk2[5].wave_shpr.div.b1[8] ),
    .B(\genblk2[5].wave_shpr.div.acc[8] ),
    .X(_04796_));
 sky130_fd_sc_hd__a21o_1 _10569_ (.A1(_04772_),
    .A2(_04795_),
    .B1(_04796_),
    .X(_04797_));
 sky130_fd_sc_hd__and2b_1 _10570_ (.A_N(\genblk2[5].wave_shpr.div.b1[9] ),
    .B(\genblk2[5].wave_shpr.div.acc[9] ),
    .X(_04798_));
 sky130_fd_sc_hd__a21o_1 _10571_ (.A1(_04771_),
    .A2(_04797_),
    .B1(_04798_),
    .X(_04799_));
 sky130_fd_sc_hd__and2b_1 _10572_ (.A_N(\genblk2[5].wave_shpr.div.b1[10] ),
    .B(\genblk2[5].wave_shpr.div.acc[10] ),
    .X(_04800_));
 sky130_fd_sc_hd__a21o_1 _10573_ (.A1(_04770_),
    .A2(_04799_),
    .B1(_04800_),
    .X(_04801_));
 sky130_fd_sc_hd__and2b_1 _10574_ (.A_N(\genblk2[5].wave_shpr.div.b1[11] ),
    .B(\genblk2[5].wave_shpr.div.acc[11] ),
    .X(_04802_));
 sky130_fd_sc_hd__a21o_1 _10575_ (.A1(_04769_),
    .A2(_04801_),
    .B1(_04802_),
    .X(_04803_));
 sky130_fd_sc_hd__and2b_1 _10576_ (.A_N(\genblk2[5].wave_shpr.div.b1[12] ),
    .B(\genblk2[5].wave_shpr.div.acc[12] ),
    .X(_04804_));
 sky130_fd_sc_hd__a21o_1 _10577_ (.A1(_04768_),
    .A2(_04803_),
    .B1(_04804_),
    .X(_04805_));
 sky130_fd_sc_hd__and2b_1 _10578_ (.A_N(\genblk2[5].wave_shpr.div.b1[13] ),
    .B(\genblk2[5].wave_shpr.div.acc[13] ),
    .X(_04806_));
 sky130_fd_sc_hd__a21o_1 _10579_ (.A1(_04767_),
    .A2(_04805_),
    .B1(_04806_),
    .X(_04807_));
 sky130_fd_sc_hd__and2b_1 _10580_ (.A_N(\genblk2[5].wave_shpr.div.b1[14] ),
    .B(\genblk2[5].wave_shpr.div.acc[14] ),
    .X(_04808_));
 sky130_fd_sc_hd__a21o_1 _10581_ (.A1(_04766_),
    .A2(_04807_),
    .B1(_04808_),
    .X(_04809_));
 sky130_fd_sc_hd__and2b_1 _10582_ (.A_N(\genblk2[5].wave_shpr.div.b1[15] ),
    .B(\genblk2[5].wave_shpr.div.acc[15] ),
    .X(_04810_));
 sky130_fd_sc_hd__a21oi_1 _10583_ (.A1(_04765_),
    .A2(_04809_),
    .B1(_04810_),
    .Y(_04811_));
 sky130_fd_sc_hd__and2_1 _10584_ (.A(_04649_),
    .B(\genblk2[5].wave_shpr.div.acc[16] ),
    .X(_04812_));
 sky130_fd_sc_hd__o21bai_1 _10585_ (.A1(_04764_),
    .A2(_04811_),
    .B1_N(_04812_),
    .Y(_04813_));
 sky130_fd_sc_hd__and2b_1 _10586_ (.A_N(\genblk2[5].wave_shpr.div.b1[17] ),
    .B(\genblk2[5].wave_shpr.div.acc[17] ),
    .X(_04814_));
 sky130_fd_sc_hd__a21o_1 _10587_ (.A1(_04763_),
    .A2(_04813_),
    .B1(_04814_),
    .X(_04815_));
 sky130_fd_sc_hd__or2_1 _10588_ (.A(\genblk2[5].wave_shpr.div.acc[18] ),
    .B(_04815_),
    .X(_04816_));
 sky130_fd_sc_hd__or4_1 _10589_ (.A(\genblk2[5].wave_shpr.div.acc[21] ),
    .B(\genblk2[5].wave_shpr.div.acc[20] ),
    .C(\genblk2[5].wave_shpr.div.acc[19] ),
    .D(_04816_),
    .X(_04817_));
 sky130_fd_sc_hd__or2_2 _10590_ (.A(\genblk2[5].wave_shpr.div.acc[22] ),
    .B(_04817_),
    .X(_04818_));
 sky130_fd_sc_hd__or4_2 _10591_ (.A(\genblk2[5].wave_shpr.div.acc[23] ),
    .B(\genblk2[5].wave_shpr.div.acc[25] ),
    .C(\genblk2[5].wave_shpr.div.acc[24] ),
    .D(\genblk2[5].wave_shpr.div.acc[26] ),
    .X(_04819_));
 sky130_fd_sc_hd__or2_1 _10592_ (.A(_04818_),
    .B(_04819_),
    .X(_04820_));
 sky130_fd_sc_hd__buf_4 _10593_ (.A(_04820_),
    .X(_04821_));
 sky130_fd_sc_hd__mux2_1 _10594_ (.A0(\genblk2[5].wave_shpr.div.fin_quo[0] ),
    .A1(_04821_),
    .S(_00015_),
    .X(_04822_));
 sky130_fd_sc_hd__clkbuf_1 _10595_ (.A(_04822_),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_1 _10596_ (.A0(\genblk2[5].wave_shpr.div.fin_quo[1] ),
    .A1(\genblk2[5].wave_shpr.div.quo[0] ),
    .S(_00015_),
    .X(_04823_));
 sky130_fd_sc_hd__clkbuf_1 _10597_ (.A(_04823_),
    .X(_00518_));
 sky130_fd_sc_hd__mux2_1 _10598_ (.A0(\genblk2[5].wave_shpr.div.fin_quo[2] ),
    .A1(net1336),
    .S(_00015_),
    .X(_04824_));
 sky130_fd_sc_hd__clkbuf_1 _10599_ (.A(_04824_),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_1 _10600_ (.A0(\genblk2[5].wave_shpr.div.fin_quo[3] ),
    .A1(\genblk2[5].wave_shpr.div.quo[2] ),
    .S(_00015_),
    .X(_04825_));
 sky130_fd_sc_hd__clkbuf_1 _10601_ (.A(_04825_),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_1 _10602_ (.A0(\genblk2[5].wave_shpr.div.fin_quo[4] ),
    .A1(net1326),
    .S(_00015_),
    .X(_04826_));
 sky130_fd_sc_hd__clkbuf_1 _10603_ (.A(_04826_),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _10604_ (.A0(\genblk2[5].wave_shpr.div.fin_quo[5] ),
    .A1(net1330),
    .S(_00015_),
    .X(_04827_));
 sky130_fd_sc_hd__clkbuf_1 _10605_ (.A(_04827_),
    .X(_00522_));
 sky130_fd_sc_hd__mux2_1 _10606_ (.A0(\genblk2[5].wave_shpr.div.fin_quo[6] ),
    .A1(net1315),
    .S(_00015_),
    .X(_04828_));
 sky130_fd_sc_hd__clkbuf_1 _10607_ (.A(_04828_),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _10608_ (.A0(\genblk2[5].wave_shpr.div.fin_quo[7] ),
    .A1(net1344),
    .S(_00015_),
    .X(_04829_));
 sky130_fd_sc_hd__clkbuf_1 _10609_ (.A(_04829_),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _10610_ (.A0(\genblk2[6].wave_shpr.div.b1[0] ),
    .A1(_01189_),
    .S(_04637_),
    .X(_04830_));
 sky130_fd_sc_hd__clkbuf_1 _10611_ (.A(_04830_),
    .X(_00525_));
 sky130_fd_sc_hd__inv_2 _10612_ (.A(_01738_),
    .Y(_04831_));
 sky130_fd_sc_hd__mux2_1 _10613_ (.A0(\genblk2[6].wave_shpr.div.b1[1] ),
    .A1(_04831_),
    .S(_04637_),
    .X(_04832_));
 sky130_fd_sc_hd__clkbuf_1 _10614_ (.A(_04832_),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _10615_ (.A0(\genblk2[6].wave_shpr.div.b1[2] ),
    .A1(_01684_),
    .S(_04637_),
    .X(_04833_));
 sky130_fd_sc_hd__clkbuf_1 _10616_ (.A(_04833_),
    .X(_00527_));
 sky130_fd_sc_hd__buf_4 _10617_ (.A(_03701_),
    .X(_04834_));
 sky130_fd_sc_hd__mux2_1 _10618_ (.A0(\genblk2[6].wave_shpr.div.b1[3] ),
    .A1(_01758_),
    .S(_04834_),
    .X(_04835_));
 sky130_fd_sc_hd__clkbuf_1 _10619_ (.A(_04835_),
    .X(_00528_));
 sky130_fd_sc_hd__inv_2 _10620_ (.A(_01730_),
    .Y(_04836_));
 sky130_fd_sc_hd__mux2_1 _10621_ (.A0(\genblk2[6].wave_shpr.div.b1[4] ),
    .A1(_04836_),
    .S(_04834_),
    .X(_04837_));
 sky130_fd_sc_hd__clkbuf_1 _10622_ (.A(_04837_),
    .X(_00529_));
 sky130_fd_sc_hd__inv_2 _10623_ (.A(_01747_),
    .Y(_04838_));
 sky130_fd_sc_hd__mux2_1 _10624_ (.A0(\genblk2[6].wave_shpr.div.b1[5] ),
    .A1(_04838_),
    .S(_04834_),
    .X(_04839_));
 sky130_fd_sc_hd__clkbuf_1 _10625_ (.A(_04839_),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_1 _10626_ (.A0(net1258),
    .A1(net37),
    .S(_04834_),
    .X(_04840_));
 sky130_fd_sc_hd__clkbuf_1 _10627_ (.A(_04840_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _10628_ (.A0(net1211),
    .A1(_01189_),
    .S(_04834_),
    .X(_04841_));
 sky130_fd_sc_hd__clkbuf_1 _10629_ (.A(_04841_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _10630_ (.A0(net1308),
    .A1(_02725_),
    .S(_04834_),
    .X(_04842_));
 sky130_fd_sc_hd__clkbuf_1 _10631_ (.A(_04842_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _10632_ (.A0(\genblk2[6].wave_shpr.div.b1[9] ),
    .A1(_01923_),
    .S(_04834_),
    .X(_04843_));
 sky130_fd_sc_hd__clkbuf_1 _10633_ (.A(_04843_),
    .X(_00534_));
 sky130_fd_sc_hd__inv_2 _10634_ (.A(_01742_),
    .Y(_04844_));
 sky130_fd_sc_hd__mux2_1 _10635_ (.A0(\genblk2[6].wave_shpr.div.b1[10] ),
    .A1(_04844_),
    .S(_04834_),
    .X(_04845_));
 sky130_fd_sc_hd__clkbuf_1 _10636_ (.A(_04845_),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _10637_ (.A0(net1233),
    .A1(_04223_),
    .S(_04834_),
    .X(_04846_));
 sky130_fd_sc_hd__clkbuf_1 _10638_ (.A(_04846_),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_1 _10639_ (.A0(net1248),
    .A1(_04225_),
    .S(_04834_),
    .X(_04847_));
 sky130_fd_sc_hd__clkbuf_1 _10640_ (.A(_04847_),
    .X(_00537_));
 sky130_fd_sc_hd__clkbuf_8 _10641_ (.A(_03707_),
    .X(_04848_));
 sky130_fd_sc_hd__mux2_1 _10642_ (.A0(\genblk2[6].wave_shpr.div.b1[13] ),
    .A1(_04645_),
    .S(_04848_),
    .X(_04849_));
 sky130_fd_sc_hd__clkbuf_1 _10643_ (.A(_04849_),
    .X(_00538_));
 sky130_fd_sc_hd__a21o_1 _10644_ (.A1(_03704_),
    .A2(net747),
    .B1(_04647_),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _10645_ (.A0(\genblk2[6].wave_shpr.div.b1[15] ),
    .A1(_01365_),
    .S(_04848_),
    .X(_04850_));
 sky130_fd_sc_hd__clkbuf_1 _10646_ (.A(_04850_),
    .X(_00540_));
 sky130_fd_sc_hd__inv_2 _10647_ (.A(net1096),
    .Y(_04851_));
 sky130_fd_sc_hd__o21ai_1 _10648_ (.A1(_03726_),
    .A2(_04851_),
    .B1(_03736_),
    .Y(_00541_));
 sky130_fd_sc_hd__and2_1 _10649_ (.A(_02171_),
    .B(\genblk2[6].wave_shpr.div.b1[17] ),
    .X(_04852_));
 sky130_fd_sc_hd__clkbuf_1 _10650_ (.A(_04852_),
    .X(_00542_));
 sky130_fd_sc_hd__clkbuf_4 _10651_ (.A(_02183_),
    .X(_04853_));
 sky130_fd_sc_hd__and3_1 _10652_ (.A(_02170_),
    .B(\genblk2[5].wave_shpr.div.busy ),
    .C(_02180_),
    .X(_04854_));
 sky130_fd_sc_hd__clkbuf_4 _10653_ (.A(_04854_),
    .X(_04855_));
 sky130_fd_sc_hd__a22o_1 _10654_ (.A1(net1342),
    .A2(_04853_),
    .B1(_04821_),
    .B2(_04855_),
    .X(_00543_));
 sky130_fd_sc_hd__clkbuf_4 _10655_ (.A(_04854_),
    .X(_04856_));
 sky130_fd_sc_hd__clkbuf_4 _10656_ (.A(_04856_),
    .X(_04857_));
 sky130_fd_sc_hd__a22o_1 _10657_ (.A1(net879),
    .A2(_04853_),
    .B1(_04857_),
    .B2(net1056),
    .X(_00544_));
 sky130_fd_sc_hd__a22o_1 _10658_ (.A1(\genblk2[5].wave_shpr.div.quo[2] ),
    .A2(_04853_),
    .B1(_04857_),
    .B2(net879),
    .X(_00545_));
 sky130_fd_sc_hd__a22o_1 _10659_ (.A1(net745),
    .A2(_04853_),
    .B1(_04857_),
    .B2(net882),
    .X(_00546_));
 sky130_fd_sc_hd__a22o_1 _10660_ (.A1(net729),
    .A2(_04853_),
    .B1(_04857_),
    .B2(net745),
    .X(_00547_));
 sky130_fd_sc_hd__a22o_1 _10661_ (.A1(net253),
    .A2(_04853_),
    .B1(_04857_),
    .B2(net729),
    .X(_00548_));
 sky130_fd_sc_hd__a22o_1 _10662_ (.A1(\genblk2[5].wave_shpr.div.quo[6] ),
    .A2(_04853_),
    .B1(_04857_),
    .B2(net253),
    .X(_00549_));
 sky130_fd_sc_hd__a22o_1 _10663_ (.A1(net308),
    .A2(_04853_),
    .B1(_04857_),
    .B2(net770),
    .X(_00550_));
 sky130_fd_sc_hd__a22o_1 _10664_ (.A1(\genblk2[5].wave_shpr.div.quo[8] ),
    .A2(_04853_),
    .B1(_04857_),
    .B2(net308),
    .X(_00551_));
 sky130_fd_sc_hd__clkbuf_4 _10665_ (.A(_02182_),
    .X(_04858_));
 sky130_fd_sc_hd__and2_1 _10666_ (.A(_04672_),
    .B(\genblk1[5].osc.clkdiv_C.cnt[0] ),
    .X(_04859_));
 sky130_fd_sc_hd__a221o_1 _10667_ (.A1(net310),
    .A2(_04858_),
    .B1(_04855_),
    .B2(net423),
    .C1(_04859_),
    .X(_00552_));
 sky130_fd_sc_hd__and2_1 _10668_ (.A(_04672_),
    .B(\genblk1[5].osc.clkdiv_C.cnt[1] ),
    .X(_04860_));
 sky130_fd_sc_hd__a221o_1 _10669_ (.A1(\genblk2[5].wave_shpr.div.quo[10] ),
    .A2(_04858_),
    .B1(_04855_),
    .B2(net310),
    .C1(_04860_),
    .X(_00553_));
 sky130_fd_sc_hd__clkbuf_4 _10670_ (.A(_02182_),
    .X(_04861_));
 sky130_fd_sc_hd__clkbuf_4 _10671_ (.A(_04854_),
    .X(_04862_));
 sky130_fd_sc_hd__and2_1 _10672_ (.A(_04672_),
    .B(\genblk1[5].osc.clkdiv_C.cnt[2] ),
    .X(_04863_));
 sky130_fd_sc_hd__a221o_1 _10673_ (.A1(net500),
    .A2(_04861_),
    .B1(_04862_),
    .B2(net572),
    .C1(_04863_),
    .X(_00554_));
 sky130_fd_sc_hd__and2_1 _10674_ (.A(_04672_),
    .B(\genblk1[5].osc.clkdiv_C.cnt[3] ),
    .X(_04864_));
 sky130_fd_sc_hd__a221o_1 _10675_ (.A1(net453),
    .A2(_04861_),
    .B1(_04862_),
    .B2(net500),
    .C1(_04864_),
    .X(_00555_));
 sky130_fd_sc_hd__and2_1 _10676_ (.A(_04672_),
    .B(\genblk1[5].osc.clkdiv_C.cnt[4] ),
    .X(_04865_));
 sky130_fd_sc_hd__a221o_1 _10677_ (.A1(net294),
    .A2(_04861_),
    .B1(_04862_),
    .B2(net453),
    .C1(_04865_),
    .X(_00556_));
 sky130_fd_sc_hd__and2_1 _10678_ (.A(_04672_),
    .B(\genblk1[5].osc.clkdiv_C.cnt[5] ),
    .X(_04866_));
 sky130_fd_sc_hd__a221o_1 _10679_ (.A1(net249),
    .A2(_04861_),
    .B1(_04862_),
    .B2(net294),
    .C1(_04866_),
    .X(_00557_));
 sky130_fd_sc_hd__nor2_1 _10680_ (.A(_04676_),
    .B(_01670_),
    .Y(_04867_));
 sky130_fd_sc_hd__a221o_1 _10681_ (.A1(\genblk2[5].wave_shpr.div.quo[15] ),
    .A2(_04861_),
    .B1(_04862_),
    .B2(net249),
    .C1(_04867_),
    .X(_00558_));
 sky130_fd_sc_hd__and2_1 _10682_ (.A(_04672_),
    .B(\genblk1[5].osc.clkdiv_C.cnt[7] ),
    .X(_04868_));
 sky130_fd_sc_hd__a221o_1 _10683_ (.A1(net378),
    .A2(_04861_),
    .B1(_04862_),
    .B2(net551),
    .C1(_04868_),
    .X(_00559_));
 sky130_fd_sc_hd__clkbuf_2 _10684_ (.A(_04268_),
    .X(_04869_));
 sky130_fd_sc_hd__and2_1 _10685_ (.A(_04869_),
    .B(\genblk1[5].osc.clkdiv_C.cnt[8] ),
    .X(_04870_));
 sky130_fd_sc_hd__a221o_1 _10686_ (.A1(net235),
    .A2(_04861_),
    .B1(_04862_),
    .B2(net378),
    .C1(_04870_),
    .X(_00560_));
 sky130_fd_sc_hd__and2_1 _10687_ (.A(_04869_),
    .B(\genblk1[5].osc.clkdiv_C.cnt[9] ),
    .X(_04871_));
 sky130_fd_sc_hd__a221o_1 _10688_ (.A1(\genblk2[5].wave_shpr.div.quo[18] ),
    .A2(_04861_),
    .B1(_04862_),
    .B2(net235),
    .C1(_04871_),
    .X(_00561_));
 sky130_fd_sc_hd__and2_1 _10689_ (.A(_04869_),
    .B(\genblk1[5].osc.clkdiv_C.cnt[10] ),
    .X(_04872_));
 sky130_fd_sc_hd__a221o_1 _10690_ (.A1(net233),
    .A2(_04861_),
    .B1(_04862_),
    .B2(net507),
    .C1(_04872_),
    .X(_00562_));
 sky130_fd_sc_hd__and2_1 _10691_ (.A(_04869_),
    .B(\genblk1[5].osc.clkdiv_C.cnt[11] ),
    .X(_04873_));
 sky130_fd_sc_hd__a221o_1 _10692_ (.A1(\genblk2[5].wave_shpr.div.quo[20] ),
    .A2(_04861_),
    .B1(_04862_),
    .B2(net233),
    .C1(_04873_),
    .X(_00563_));
 sky130_fd_sc_hd__and2_1 _10693_ (.A(_04869_),
    .B(\genblk1[5].osc.clkdiv_C.cnt[12] ),
    .X(_04874_));
 sky130_fd_sc_hd__a221o_1 _10694_ (.A1(net245),
    .A2(_02183_),
    .B1(_04856_),
    .B2(net503),
    .C1(_04874_),
    .X(_00564_));
 sky130_fd_sc_hd__and2_1 _10695_ (.A(_04869_),
    .B(\genblk1[5].osc.clkdiv_C.cnt[13] ),
    .X(_04875_));
 sky130_fd_sc_hd__a221o_1 _10696_ (.A1(\genblk2[5].wave_shpr.div.quo[22] ),
    .A2(_02183_),
    .B1(_04856_),
    .B2(net245),
    .C1(_04875_),
    .X(_00565_));
 sky130_fd_sc_hd__and2_1 _10697_ (.A(_04869_),
    .B(\genblk1[5].osc.clkdiv_C.cnt[14] ),
    .X(_04876_));
 sky130_fd_sc_hd__a221o_1 _10698_ (.A1(net459),
    .A2(_02183_),
    .B1(_04856_),
    .B2(net471),
    .C1(_04876_),
    .X(_00566_));
 sky130_fd_sc_hd__and2_1 _10699_ (.A(_04869_),
    .B(\genblk1[5].osc.clkdiv_C.cnt[15] ),
    .X(_04877_));
 sky130_fd_sc_hd__a221o_1 _10700_ (.A1(net324),
    .A2(_02183_),
    .B1(_04856_),
    .B2(net459),
    .C1(_04877_),
    .X(_00567_));
 sky130_fd_sc_hd__and2_1 _10701_ (.A(_04869_),
    .B(\genblk1[5].osc.clkdiv_C.cnt[16] ),
    .X(_04878_));
 sky130_fd_sc_hd__a221o_1 _10702_ (.A1(\genblk2[5].wave_shpr.div.acc_next[0] ),
    .A2(_02183_),
    .B1(_04856_),
    .B2(net324),
    .C1(_04878_),
    .X(_00568_));
 sky130_fd_sc_hd__or2b_1 _10703_ (.A(\genblk2[5].wave_shpr.div.acc_next[0] ),
    .B_N(_04856_),
    .X(_04879_));
 sky130_fd_sc_hd__o221a_1 _10704_ (.A1(_03819_),
    .A2(net493),
    .B1(_00014_),
    .B2(\genblk2[5].wave_shpr.div.acc[0] ),
    .C1(_04879_),
    .X(_00569_));
 sky130_fd_sc_hd__nor2_2 _10705_ (.A(_04818_),
    .B(_04819_),
    .Y(_04880_));
 sky130_fd_sc_hd__or3b_1 _10706_ (.A(_04880_),
    .B(_04781_),
    .C_N(\genblk2[5].wave_shpr.div.b1[0] ),
    .X(_04881_));
 sky130_fd_sc_hd__a21o_1 _10707_ (.A1(\genblk2[5].wave_shpr.div.b1[0] ),
    .A2(_04821_),
    .B1(\genblk2[5].wave_shpr.div.acc[0] ),
    .X(_04882_));
 sky130_fd_sc_hd__a32o_1 _10708_ (.A1(_04855_),
    .A2(_04881_),
    .A3(_04882_),
    .B1(_04858_),
    .B2(net1062),
    .X(_00570_));
 sky130_fd_sc_hd__and3_1 _10709_ (.A(\genblk2[5].wave_shpr.div.b1[0] ),
    .B(_04781_),
    .C(_04782_),
    .X(_04883_));
 sky130_fd_sc_hd__nor2_1 _10710_ (.A(_04783_),
    .B(_04883_),
    .Y(_04884_));
 sky130_fd_sc_hd__mux2_1 _10711_ (.A0(\genblk2[5].wave_shpr.div.acc[1] ),
    .A1(_04884_),
    .S(_04821_),
    .X(_04885_));
 sky130_fd_sc_hd__a22o_1 _10712_ (.A1(net910),
    .A2(_04853_),
    .B1(_04857_),
    .B2(_04885_),
    .X(_00571_));
 sky130_fd_sc_hd__clkbuf_4 _10713_ (.A(_02183_),
    .X(_04886_));
 sky130_fd_sc_hd__or2b_1 _10714_ (.A(_04785_),
    .B_N(_04780_),
    .X(_04887_));
 sky130_fd_sc_hd__xnor2_1 _10715_ (.A(_04784_),
    .B(_04887_),
    .Y(_04888_));
 sky130_fd_sc_hd__mux2_1 _10716_ (.A0(\genblk2[5].wave_shpr.div.acc[2] ),
    .A1(_04888_),
    .S(_04821_),
    .X(_04889_));
 sky130_fd_sc_hd__a22o_1 _10717_ (.A1(net961),
    .A2(_04886_),
    .B1(_04857_),
    .B2(_04889_),
    .X(_00572_));
 sky130_fd_sc_hd__clkbuf_4 _10718_ (.A(_04856_),
    .X(_04890_));
 sky130_fd_sc_hd__or2b_1 _10719_ (.A(_04787_),
    .B_N(_04779_),
    .X(_04891_));
 sky130_fd_sc_hd__xnor2_1 _10720_ (.A(_04786_),
    .B(_04891_),
    .Y(_04892_));
 sky130_fd_sc_hd__mux2_1 _10721_ (.A0(\genblk2[5].wave_shpr.div.acc[3] ),
    .A1(_04892_),
    .S(_04821_),
    .X(_04893_));
 sky130_fd_sc_hd__a22o_1 _10722_ (.A1(net888),
    .A2(_04886_),
    .B1(_04890_),
    .B2(_04893_),
    .X(_00573_));
 sky130_fd_sc_hd__xor2_1 _10723_ (.A(_04778_),
    .B(_04788_),
    .X(_04894_));
 sky130_fd_sc_hd__mux2_1 _10724_ (.A0(\genblk2[5].wave_shpr.div.acc[4] ),
    .A1(_04894_),
    .S(_04821_),
    .X(_04895_));
 sky130_fd_sc_hd__a22o_1 _10725_ (.A1(net885),
    .A2(_04886_),
    .B1(_04890_),
    .B2(_04895_),
    .X(_00574_));
 sky130_fd_sc_hd__or2b_1 _10726_ (.A(_04790_),
    .B_N(_04775_),
    .X(_04896_));
 sky130_fd_sc_hd__xnor2_1 _10727_ (.A(_04896_),
    .B(_04789_),
    .Y(_04897_));
 sky130_fd_sc_hd__mux2_1 _10728_ (.A0(\genblk2[5].wave_shpr.div.acc[5] ),
    .A1(_04897_),
    .S(_04821_),
    .X(_04898_));
 sky130_fd_sc_hd__a22o_1 _10729_ (.A1(net863),
    .A2(_04886_),
    .B1(_04890_),
    .B2(_04898_),
    .X(_00575_));
 sky130_fd_sc_hd__or2b_1 _10730_ (.A(_04792_),
    .B_N(_04774_),
    .X(_04899_));
 sky130_fd_sc_hd__xnor2_1 _10731_ (.A(_04791_),
    .B(_04899_),
    .Y(_04900_));
 sky130_fd_sc_hd__mux2_1 _10732_ (.A0(\genblk2[5].wave_shpr.div.acc[6] ),
    .A1(_04900_),
    .S(_04821_),
    .X(_04901_));
 sky130_fd_sc_hd__a22o_1 _10733_ (.A1(net1037),
    .A2(_04886_),
    .B1(_04890_),
    .B2(_04901_),
    .X(_00576_));
 sky130_fd_sc_hd__or2b_1 _10734_ (.A(_04794_),
    .B_N(_04773_),
    .X(_04902_));
 sky130_fd_sc_hd__xnor2_1 _10735_ (.A(_04793_),
    .B(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__mux2_1 _10736_ (.A0(\genblk2[5].wave_shpr.div.acc[7] ),
    .A1(_04903_),
    .S(_04821_),
    .X(_04904_));
 sky130_fd_sc_hd__a22o_1 _10737_ (.A1(net927),
    .A2(_04886_),
    .B1(_04890_),
    .B2(_04904_),
    .X(_00577_));
 sky130_fd_sc_hd__or2b_1 _10738_ (.A(_04796_),
    .B_N(_04772_),
    .X(_04905_));
 sky130_fd_sc_hd__xnor2_1 _10739_ (.A(_04795_),
    .B(_04905_),
    .Y(_04906_));
 sky130_fd_sc_hd__buf_4 _10740_ (.A(_04820_),
    .X(_04907_));
 sky130_fd_sc_hd__mux2_1 _10741_ (.A0(\genblk2[5].wave_shpr.div.acc[8] ),
    .A1(_04906_),
    .S(_04907_),
    .X(_04908_));
 sky130_fd_sc_hd__a22o_1 _10742_ (.A1(net772),
    .A2(_04886_),
    .B1(_04890_),
    .B2(_04908_),
    .X(_00578_));
 sky130_fd_sc_hd__or2b_1 _10743_ (.A(_04798_),
    .B_N(_04771_),
    .X(_04909_));
 sky130_fd_sc_hd__xnor2_1 _10744_ (.A(_04797_),
    .B(_04909_),
    .Y(_04910_));
 sky130_fd_sc_hd__mux2_1 _10745_ (.A0(net772),
    .A1(_04910_),
    .S(_04907_),
    .X(_04911_));
 sky130_fd_sc_hd__a22o_1 _10746_ (.A1(\genblk2[5].wave_shpr.div.acc[10] ),
    .A2(_04886_),
    .B1(_04890_),
    .B2(_04911_),
    .X(_00579_));
 sky130_fd_sc_hd__or2b_1 _10747_ (.A(_04800_),
    .B_N(_04770_),
    .X(_04912_));
 sky130_fd_sc_hd__xnor2_1 _10748_ (.A(_04799_),
    .B(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__mux2_1 _10749_ (.A0(\genblk2[5].wave_shpr.div.acc[10] ),
    .A1(_04913_),
    .S(_04907_),
    .X(_04914_));
 sky130_fd_sc_hd__a22o_1 _10750_ (.A1(net1061),
    .A2(_04886_),
    .B1(_04890_),
    .B2(_04914_),
    .X(_00580_));
 sky130_fd_sc_hd__or2b_1 _10751_ (.A(_04802_),
    .B_N(_04769_),
    .X(_04915_));
 sky130_fd_sc_hd__xnor2_1 _10752_ (.A(_04801_),
    .B(_04915_),
    .Y(_04916_));
 sky130_fd_sc_hd__mux2_1 _10753_ (.A0(\genblk2[5].wave_shpr.div.acc[11] ),
    .A1(_04916_),
    .S(_04907_),
    .X(_04917_));
 sky130_fd_sc_hd__a22o_1 _10754_ (.A1(net1014),
    .A2(_04886_),
    .B1(_04890_),
    .B2(_04917_),
    .X(_00581_));
 sky130_fd_sc_hd__clkbuf_4 _10755_ (.A(_02183_),
    .X(_04918_));
 sky130_fd_sc_hd__or2b_1 _10756_ (.A(_04804_),
    .B_N(_04768_),
    .X(_04919_));
 sky130_fd_sc_hd__xnor2_1 _10757_ (.A(_04803_),
    .B(_04919_),
    .Y(_04920_));
 sky130_fd_sc_hd__mux2_1 _10758_ (.A0(\genblk2[5].wave_shpr.div.acc[12] ),
    .A1(_04920_),
    .S(_04907_),
    .X(_04921_));
 sky130_fd_sc_hd__a22o_1 _10759_ (.A1(net981),
    .A2(_04918_),
    .B1(_04890_),
    .B2(_04921_),
    .X(_00582_));
 sky130_fd_sc_hd__clkbuf_4 _10760_ (.A(_04856_),
    .X(_04922_));
 sky130_fd_sc_hd__or2b_1 _10761_ (.A(_04806_),
    .B_N(_04767_),
    .X(_04923_));
 sky130_fd_sc_hd__xnor2_1 _10762_ (.A(_04805_),
    .B(_04923_),
    .Y(_04924_));
 sky130_fd_sc_hd__mux2_1 _10763_ (.A0(\genblk2[5].wave_shpr.div.acc[13] ),
    .A1(_04924_),
    .S(_04907_),
    .X(_04925_));
 sky130_fd_sc_hd__a22o_1 _10764_ (.A1(net902),
    .A2(_04918_),
    .B1(_04922_),
    .B2(_04925_),
    .X(_00583_));
 sky130_fd_sc_hd__or2b_1 _10765_ (.A(_04808_),
    .B_N(_04766_),
    .X(_04926_));
 sky130_fd_sc_hd__xnor2_1 _10766_ (.A(_04807_),
    .B(_04926_),
    .Y(_04927_));
 sky130_fd_sc_hd__mux2_1 _10767_ (.A0(\genblk2[5].wave_shpr.div.acc[14] ),
    .A1(_04927_),
    .S(_04907_),
    .X(_04928_));
 sky130_fd_sc_hd__a22o_1 _10768_ (.A1(net835),
    .A2(_04918_),
    .B1(_04922_),
    .B2(_04928_),
    .X(_00584_));
 sky130_fd_sc_hd__or2b_1 _10769_ (.A(_04810_),
    .B_N(_04765_),
    .X(_04929_));
 sky130_fd_sc_hd__xnor2_1 _10770_ (.A(_04809_),
    .B(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__mux2_1 _10771_ (.A0(\genblk2[5].wave_shpr.div.acc[15] ),
    .A1(_04930_),
    .S(_04907_),
    .X(_04931_));
 sky130_fd_sc_hd__a22o_1 _10772_ (.A1(net925),
    .A2(_04918_),
    .B1(_04922_),
    .B2(_04931_),
    .X(_00585_));
 sky130_fd_sc_hd__nor2_1 _10773_ (.A(_04812_),
    .B(_04764_),
    .Y(_04932_));
 sky130_fd_sc_hd__xnor2_1 _10774_ (.A(_04932_),
    .B(_04811_),
    .Y(_04933_));
 sky130_fd_sc_hd__mux2_1 _10775_ (.A0(\genblk2[5].wave_shpr.div.acc[16] ),
    .A1(_04933_),
    .S(_04907_),
    .X(_04934_));
 sky130_fd_sc_hd__a22o_1 _10776_ (.A1(net828),
    .A2(_04918_),
    .B1(_04922_),
    .B2(_04934_),
    .X(_00586_));
 sky130_fd_sc_hd__or2b_1 _10777_ (.A(_04814_),
    .B_N(_04763_),
    .X(_04935_));
 sky130_fd_sc_hd__xnor2_1 _10778_ (.A(_04813_),
    .B(_04935_),
    .Y(_04936_));
 sky130_fd_sc_hd__mux2_1 _10779_ (.A0(\genblk2[5].wave_shpr.div.acc[17] ),
    .A1(_04936_),
    .S(_04907_),
    .X(_04937_));
 sky130_fd_sc_hd__a22o_1 _10780_ (.A1(net630),
    .A2(_04918_),
    .B1(_04922_),
    .B2(_04937_),
    .X(_00587_));
 sky130_fd_sc_hd__or2_1 _10781_ (.A(_04816_),
    .B(_04880_),
    .X(_04938_));
 sky130_fd_sc_hd__o21ai_1 _10782_ (.A1(_04815_),
    .A2(_04880_),
    .B1(net630),
    .Y(_04939_));
 sky130_fd_sc_hd__nand2_1 _10783_ (.A(_04938_),
    .B(_04939_),
    .Y(_04940_));
 sky130_fd_sc_hd__a22o_1 _10784_ (.A1(net896),
    .A2(_04918_),
    .B1(_04922_),
    .B2(_04940_),
    .X(_00588_));
 sky130_fd_sc_hd__or2_1 _10785_ (.A(\genblk2[5].wave_shpr.div.acc[19] ),
    .B(_04938_),
    .X(_04941_));
 sky130_fd_sc_hd__a21bo_1 _10786_ (.A1(\genblk2[5].wave_shpr.div.acc[19] ),
    .A2(_04816_),
    .B1_N(_04941_),
    .X(_04942_));
 sky130_fd_sc_hd__a22o_1 _10787_ (.A1(net982),
    .A2(_04918_),
    .B1(_04922_),
    .B2(_04942_),
    .X(_00589_));
 sky130_fd_sc_hd__or2_1 _10788_ (.A(\genblk2[5].wave_shpr.div.acc[20] ),
    .B(_04941_),
    .X(_04943_));
 sky130_fd_sc_hd__nand2_1 _10789_ (.A(net1345),
    .B(_04941_),
    .Y(_04944_));
 sky130_fd_sc_hd__nand2_1 _10790_ (.A(_04943_),
    .B(_04944_),
    .Y(_04945_));
 sky130_fd_sc_hd__a22o_1 _10791_ (.A1(net566),
    .A2(_04918_),
    .B1(_04922_),
    .B2(_04945_),
    .X(_00590_));
 sky130_fd_sc_hd__a2bb2o_1 _10792_ (.A1_N(_04817_),
    .A2_N(_04880_),
    .B1(_04943_),
    .B2(\genblk2[5].wave_shpr.div.acc[21] ),
    .X(_04946_));
 sky130_fd_sc_hd__a22o_1 _10793_ (.A1(net654),
    .A2(_04918_),
    .B1(_04922_),
    .B2(_04946_),
    .X(_00591_));
 sky130_fd_sc_hd__and2b_1 _10794_ (.A_N(_04818_),
    .B(_04819_),
    .X(_04947_));
 sky130_fd_sc_hd__a21o_1 _10795_ (.A1(\genblk2[5].wave_shpr.div.acc[22] ),
    .A2(_04817_),
    .B1(_04947_),
    .X(_04948_));
 sky130_fd_sc_hd__a22o_1 _10796_ (.A1(net1012),
    .A2(_04858_),
    .B1(_04922_),
    .B2(_04948_),
    .X(_00592_));
 sky130_fd_sc_hd__nor2_1 _10797_ (.A(\genblk2[5].wave_shpr.div.acc[23] ),
    .B(_04818_),
    .Y(_04949_));
 sky130_fd_sc_hd__and2_1 _10798_ (.A(\genblk2[5].wave_shpr.div.acc[23] ),
    .B(_04818_),
    .X(_04950_));
 sky130_fd_sc_hd__or2_1 _10799_ (.A(_04949_),
    .B(_04950_),
    .X(_04951_));
 sky130_fd_sc_hd__a32o_1 _10800_ (.A1(_04819_),
    .A2(_04855_),
    .A3(_04951_),
    .B1(_04858_),
    .B2(net1038),
    .X(_00593_));
 sky130_fd_sc_hd__inv_2 _10801_ (.A(\genblk2[5].wave_shpr.div.acc[24] ),
    .Y(_04952_));
 sky130_fd_sc_hd__or3b_1 _10802_ (.A(\genblk2[5].wave_shpr.div.acc[24] ),
    .B(_04880_),
    .C_N(_04949_),
    .X(_04953_));
 sky130_fd_sc_hd__o21ai_1 _10803_ (.A1(_04952_),
    .A2(_04949_),
    .B1(_04953_),
    .Y(_04954_));
 sky130_fd_sc_hd__a22o_1 _10804_ (.A1(net1041),
    .A2(_04858_),
    .B1(_04855_),
    .B2(_04954_),
    .X(_00594_));
 sky130_fd_sc_hd__xnor2_1 _10805_ (.A(\genblk2[5].wave_shpr.div.acc[25] ),
    .B(_04953_),
    .Y(_04955_));
 sky130_fd_sc_hd__a22o_1 _10806_ (.A1(net392),
    .A2(_04858_),
    .B1(_04855_),
    .B2(_04955_),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _10807_ (.A0(_04856_),
    .A1(_02183_),
    .S(\genblk2[5].wave_shpr.div.i[0] ),
    .X(_04956_));
 sky130_fd_sc_hd__clkbuf_1 _10808_ (.A(_04956_),
    .X(_00596_));
 sky130_fd_sc_hd__or2_1 _10809_ (.A(\genblk2[5].wave_shpr.div.i[1] ),
    .B(\genblk2[5].wave_shpr.div.i[0] ),
    .X(_04957_));
 sky130_fd_sc_hd__nand2_1 _10810_ (.A(\genblk2[5].wave_shpr.div.i[1] ),
    .B(\genblk2[5].wave_shpr.div.i[0] ),
    .Y(_04958_));
 sky130_fd_sc_hd__a32o_1 _10811_ (.A1(_04855_),
    .A2(_04957_),
    .A3(_04958_),
    .B1(_04858_),
    .B2(net1117),
    .X(_00597_));
 sky130_fd_sc_hd__a21o_1 _10812_ (.A1(\genblk2[5].wave_shpr.div.i[1] ),
    .A2(\genblk2[5].wave_shpr.div.i[0] ),
    .B1(\genblk2[5].wave_shpr.div.i[2] ),
    .X(_04959_));
 sky130_fd_sc_hd__nand3_1 _10813_ (.A(\genblk2[5].wave_shpr.div.i[1] ),
    .B(\genblk2[5].wave_shpr.div.i[0] ),
    .C(\genblk2[5].wave_shpr.div.i[2] ),
    .Y(_04960_));
 sky130_fd_sc_hd__a32o_1 _10814_ (.A1(_04855_),
    .A2(_04959_),
    .A3(_04960_),
    .B1(_04858_),
    .B2(net1154),
    .X(_00598_));
 sky130_fd_sc_hd__a31o_1 _10815_ (.A1(\genblk2[5].wave_shpr.div.i[1] ),
    .A2(\genblk2[5].wave_shpr.div.i[0] ),
    .A3(\genblk2[5].wave_shpr.div.i[2] ),
    .B1(\genblk2[5].wave_shpr.div.i[3] ),
    .X(_04961_));
 sky130_fd_sc_hd__and4_1 _10816_ (.A(\genblk2[5].wave_shpr.div.i[1] ),
    .B(\genblk2[5].wave_shpr.div.i[0] ),
    .C(\genblk2[5].wave_shpr.div.i[2] ),
    .D(\genblk2[5].wave_shpr.div.i[3] ),
    .X(_04962_));
 sky130_fd_sc_hd__inv_2 _10817_ (.A(_04962_),
    .Y(_04963_));
 sky130_fd_sc_hd__a32o_1 _10818_ (.A1(_04855_),
    .A2(_04961_),
    .A3(_04963_),
    .B1(_04858_),
    .B2(net783),
    .X(_00599_));
 sky130_fd_sc_hd__a21oi_1 _10819_ (.A1(\genblk2[5].wave_shpr.div.busy ),
    .A2(_04962_),
    .B1(net855),
    .Y(_04964_));
 sky130_fd_sc_hd__a31o_1 _10820_ (.A1(net855),
    .A2(_02181_),
    .A3(_04962_),
    .B1(_03708_),
    .X(_04965_));
 sky130_fd_sc_hd__nor2_1 _10821_ (.A(net856),
    .B(_04965_),
    .Y(_00600_));
 sky130_fd_sc_hd__or2b_1 _10822_ (.A(\genblk2[6].wave_shpr.div.acc[17] ),
    .B_N(\genblk2[6].wave_shpr.div.b1[17] ),
    .X(_04966_));
 sky130_fd_sc_hd__xor2_1 _10823_ (.A(\genblk2[6].wave_shpr.div.b1[16] ),
    .B(\genblk2[6].wave_shpr.div.acc[16] ),
    .X(_04967_));
 sky130_fd_sc_hd__or2b_1 _10824_ (.A(\genblk2[6].wave_shpr.div.acc[15] ),
    .B_N(\genblk2[6].wave_shpr.div.b1[15] ),
    .X(_04968_));
 sky130_fd_sc_hd__or2b_1 _10825_ (.A(\genblk2[6].wave_shpr.div.acc[14] ),
    .B_N(\genblk2[6].wave_shpr.div.b1[14] ),
    .X(_04969_));
 sky130_fd_sc_hd__or2b_1 _10826_ (.A(\genblk2[6].wave_shpr.div.acc[13] ),
    .B_N(\genblk2[6].wave_shpr.div.b1[13] ),
    .X(_04970_));
 sky130_fd_sc_hd__or2b_1 _10827_ (.A(\genblk2[6].wave_shpr.div.acc[12] ),
    .B_N(\genblk2[6].wave_shpr.div.b1[12] ),
    .X(_04971_));
 sky130_fd_sc_hd__or2b_1 _10828_ (.A(\genblk2[6].wave_shpr.div.acc[11] ),
    .B_N(\genblk2[6].wave_shpr.div.b1[11] ),
    .X(_04972_));
 sky130_fd_sc_hd__or2b_1 _10829_ (.A(\genblk2[6].wave_shpr.div.acc[10] ),
    .B_N(\genblk2[6].wave_shpr.div.b1[10] ),
    .X(_04973_));
 sky130_fd_sc_hd__or2b_1 _10830_ (.A(\genblk2[6].wave_shpr.div.acc[9] ),
    .B_N(\genblk2[6].wave_shpr.div.b1[9] ),
    .X(_04974_));
 sky130_fd_sc_hd__or2b_1 _10831_ (.A(\genblk2[6].wave_shpr.div.acc[8] ),
    .B_N(\genblk2[6].wave_shpr.div.b1[8] ),
    .X(_04975_));
 sky130_fd_sc_hd__or2b_1 _10832_ (.A(\genblk2[6].wave_shpr.div.acc[7] ),
    .B_N(\genblk2[6].wave_shpr.div.b1[7] ),
    .X(_04976_));
 sky130_fd_sc_hd__or2b_1 _10833_ (.A(\genblk2[6].wave_shpr.div.acc[6] ),
    .B_N(\genblk2[6].wave_shpr.div.b1[6] ),
    .X(_04977_));
 sky130_fd_sc_hd__or2b_1 _10834_ (.A(\genblk2[6].wave_shpr.div.acc[5] ),
    .B_N(\genblk2[6].wave_shpr.div.b1[5] ),
    .X(_04978_));
 sky130_fd_sc_hd__or2b_1 _10835_ (.A(\genblk2[6].wave_shpr.div.acc[4] ),
    .B_N(\genblk2[6].wave_shpr.div.b1[4] ),
    .X(_04979_));
 sky130_fd_sc_hd__or2b_1 _10836_ (.A(\genblk2[6].wave_shpr.div.acc[3] ),
    .B_N(\genblk2[6].wave_shpr.div.b1[3] ),
    .X(_04980_));
 sky130_fd_sc_hd__inv_2 _10837_ (.A(\genblk2[6].wave_shpr.div.b1[2] ),
    .Y(_04981_));
 sky130_fd_sc_hd__xor2_1 _10838_ (.A(\genblk2[6].wave_shpr.div.acc[1] ),
    .B(\genblk2[6].wave_shpr.div.b1[1] ),
    .X(_04982_));
 sky130_fd_sc_hd__and2b_1 _10839_ (.A_N(\genblk2[6].wave_shpr.div.acc[0] ),
    .B(\genblk2[6].wave_shpr.div.b1[0] ),
    .X(_04983_));
 sky130_fd_sc_hd__or2b_1 _10840_ (.A(\genblk2[6].wave_shpr.div.b1[1] ),
    .B_N(\genblk2[6].wave_shpr.div.acc[1] ),
    .X(_04984_));
 sky130_fd_sc_hd__o21ai_1 _10841_ (.A1(_04982_),
    .A2(_04983_),
    .B1(_04984_),
    .Y(_04985_));
 sky130_fd_sc_hd__o21a_1 _10842_ (.A1(_04981_),
    .A2(\genblk2[6].wave_shpr.div.acc[2] ),
    .B1(_04985_),
    .X(_04986_));
 sky130_fd_sc_hd__a21o_1 _10843_ (.A1(_04981_),
    .A2(\genblk2[6].wave_shpr.div.acc[2] ),
    .B1(_04986_),
    .X(_04987_));
 sky130_fd_sc_hd__and2b_1 _10844_ (.A_N(\genblk2[6].wave_shpr.div.b1[3] ),
    .B(\genblk2[6].wave_shpr.div.acc[3] ),
    .X(_04988_));
 sky130_fd_sc_hd__a21o_1 _10845_ (.A1(_04980_),
    .A2(_04987_),
    .B1(_04988_),
    .X(_04989_));
 sky130_fd_sc_hd__and2b_1 _10846_ (.A_N(\genblk2[6].wave_shpr.div.b1[4] ),
    .B(\genblk2[6].wave_shpr.div.acc[4] ),
    .X(_04990_));
 sky130_fd_sc_hd__a21o_1 _10847_ (.A1(_04979_),
    .A2(_04989_),
    .B1(_04990_),
    .X(_04991_));
 sky130_fd_sc_hd__and2b_1 _10848_ (.A_N(\genblk2[6].wave_shpr.div.b1[5] ),
    .B(\genblk2[6].wave_shpr.div.acc[5] ),
    .X(_04992_));
 sky130_fd_sc_hd__a21o_1 _10849_ (.A1(_04978_),
    .A2(_04991_),
    .B1(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__and2b_1 _10850_ (.A_N(\genblk2[6].wave_shpr.div.b1[6] ),
    .B(\genblk2[6].wave_shpr.div.acc[6] ),
    .X(_04994_));
 sky130_fd_sc_hd__a21o_1 _10851_ (.A1(_04977_),
    .A2(_04993_),
    .B1(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__and2b_1 _10852_ (.A_N(\genblk2[6].wave_shpr.div.b1[7] ),
    .B(\genblk2[6].wave_shpr.div.acc[7] ),
    .X(_04996_));
 sky130_fd_sc_hd__a21o_1 _10853_ (.A1(_04976_),
    .A2(_04995_),
    .B1(_04996_),
    .X(_04997_));
 sky130_fd_sc_hd__and2b_1 _10854_ (.A_N(\genblk2[6].wave_shpr.div.b1[8] ),
    .B(\genblk2[6].wave_shpr.div.acc[8] ),
    .X(_04998_));
 sky130_fd_sc_hd__a21o_1 _10855_ (.A1(_04975_),
    .A2(_04997_),
    .B1(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__and2b_1 _10856_ (.A_N(\genblk2[6].wave_shpr.div.b1[9] ),
    .B(\genblk2[6].wave_shpr.div.acc[9] ),
    .X(_05000_));
 sky130_fd_sc_hd__a21o_1 _10857_ (.A1(_04974_),
    .A2(_04999_),
    .B1(_05000_),
    .X(_05001_));
 sky130_fd_sc_hd__and2b_1 _10858_ (.A_N(\genblk2[6].wave_shpr.div.b1[10] ),
    .B(\genblk2[6].wave_shpr.div.acc[10] ),
    .X(_05002_));
 sky130_fd_sc_hd__a21o_1 _10859_ (.A1(_04973_),
    .A2(_05001_),
    .B1(_05002_),
    .X(_05003_));
 sky130_fd_sc_hd__and2b_1 _10860_ (.A_N(\genblk2[6].wave_shpr.div.b1[11] ),
    .B(\genblk2[6].wave_shpr.div.acc[11] ),
    .X(_05004_));
 sky130_fd_sc_hd__a21o_1 _10861_ (.A1(_04972_),
    .A2(_05003_),
    .B1(_05004_),
    .X(_05005_));
 sky130_fd_sc_hd__and2b_1 _10862_ (.A_N(\genblk2[6].wave_shpr.div.b1[12] ),
    .B(\genblk2[6].wave_shpr.div.acc[12] ),
    .X(_05006_));
 sky130_fd_sc_hd__a21o_1 _10863_ (.A1(_04971_),
    .A2(_05005_),
    .B1(_05006_),
    .X(_05007_));
 sky130_fd_sc_hd__and2b_1 _10864_ (.A_N(\genblk2[6].wave_shpr.div.b1[13] ),
    .B(\genblk2[6].wave_shpr.div.acc[13] ),
    .X(_05008_));
 sky130_fd_sc_hd__a21o_1 _10865_ (.A1(_04970_),
    .A2(_05007_),
    .B1(_05008_),
    .X(_05009_));
 sky130_fd_sc_hd__and2b_1 _10866_ (.A_N(\genblk2[6].wave_shpr.div.b1[14] ),
    .B(\genblk2[6].wave_shpr.div.acc[14] ),
    .X(_05010_));
 sky130_fd_sc_hd__a21o_1 _10867_ (.A1(_04969_),
    .A2(_05009_),
    .B1(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__and2b_1 _10868_ (.A_N(\genblk2[6].wave_shpr.div.b1[15] ),
    .B(\genblk2[6].wave_shpr.div.acc[15] ),
    .X(_05012_));
 sky130_fd_sc_hd__a21o_1 _10869_ (.A1(_04968_),
    .A2(_05011_),
    .B1(_05012_),
    .X(_05013_));
 sky130_fd_sc_hd__and2b_1 _10870_ (.A_N(_04967_),
    .B(_05013_),
    .X(_05014_));
 sky130_fd_sc_hd__a21o_1 _10871_ (.A1(_04851_),
    .A2(\genblk2[6].wave_shpr.div.acc[16] ),
    .B1(_05014_),
    .X(_05015_));
 sky130_fd_sc_hd__and2b_1 _10872_ (.A_N(\genblk2[6].wave_shpr.div.b1[17] ),
    .B(\genblk2[6].wave_shpr.div.acc[17] ),
    .X(_05016_));
 sky130_fd_sc_hd__a21o_1 _10873_ (.A1(_04966_),
    .A2(_05015_),
    .B1(_05016_),
    .X(_05017_));
 sky130_fd_sc_hd__or2_1 _10874_ (.A(\genblk2[6].wave_shpr.div.acc[18] ),
    .B(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__or2_1 _10875_ (.A(\genblk2[6].wave_shpr.div.acc[19] ),
    .B(_05018_),
    .X(_05019_));
 sky130_fd_sc_hd__or4_1 _10876_ (.A(\genblk2[6].wave_shpr.div.acc[22] ),
    .B(\genblk2[6].wave_shpr.div.acc[21] ),
    .C(\genblk2[6].wave_shpr.div.acc[20] ),
    .D(_05019_),
    .X(_05020_));
 sky130_fd_sc_hd__or2_2 _10877_ (.A(\genblk2[6].wave_shpr.div.acc[23] ),
    .B(_05020_),
    .X(_05021_));
 sky130_fd_sc_hd__or4_2 _10878_ (.A(\genblk2[6].wave_shpr.div.acc[25] ),
    .B(\genblk2[6].wave_shpr.div.acc[24] ),
    .C(\genblk2[6].wave_shpr.div.acc[26] ),
    .D(_05021_),
    .X(_05022_));
 sky130_fd_sc_hd__buf_4 _10879_ (.A(_05022_),
    .X(_05023_));
 sky130_fd_sc_hd__mux2_1 _10880_ (.A0(\genblk2[6].wave_shpr.div.fin_quo[0] ),
    .A1(_05023_),
    .S(_00017_),
    .X(_05024_));
 sky130_fd_sc_hd__clkbuf_1 _10881_ (.A(_05024_),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _10882_ (.A0(\genblk2[6].wave_shpr.div.fin_quo[1] ),
    .A1(\genblk2[6].wave_shpr.div.quo[0] ),
    .S(_00017_),
    .X(_05025_));
 sky130_fd_sc_hd__clkbuf_1 _10883_ (.A(_05025_),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _10884_ (.A0(\genblk2[6].wave_shpr.div.fin_quo[2] ),
    .A1(net1338),
    .S(_00017_),
    .X(_05026_));
 sky130_fd_sc_hd__clkbuf_1 _10885_ (.A(_05026_),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _10886_ (.A0(\genblk2[6].wave_shpr.div.fin_quo[3] ),
    .A1(net1320),
    .S(_00017_),
    .X(_05027_));
 sky130_fd_sc_hd__clkbuf_1 _10887_ (.A(_05027_),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_1 _10888_ (.A0(\genblk2[6].wave_shpr.div.fin_quo[4] ),
    .A1(net1319),
    .S(_00017_),
    .X(_05028_));
 sky130_fd_sc_hd__clkbuf_1 _10889_ (.A(_05028_),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_1 _10890_ (.A0(\genblk2[6].wave_shpr.div.fin_quo[5] ),
    .A1(net720),
    .S(_00017_),
    .X(_05029_));
 sky130_fd_sc_hd__clkbuf_1 _10891_ (.A(_05029_),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_1 _10892_ (.A0(\genblk2[6].wave_shpr.div.fin_quo[6] ),
    .A1(\genblk2[6].wave_shpr.div.quo[5] ),
    .S(_00017_),
    .X(_05030_));
 sky130_fd_sc_hd__clkbuf_1 _10893_ (.A(_05030_),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _10894_ (.A0(\genblk2[6].wave_shpr.div.fin_quo[7] ),
    .A1(net1349),
    .S(_00017_),
    .X(_05031_));
 sky130_fd_sc_hd__clkbuf_1 _10895_ (.A(_05031_),
    .X(_00608_));
 sky130_fd_sc_hd__mux2_1 _10896_ (.A0(\genblk2[7].wave_shpr.div.b1[0] ),
    .A1(_01514_),
    .S(_04848_),
    .X(_05032_));
 sky130_fd_sc_hd__clkbuf_1 _10897_ (.A(_05032_),
    .X(_00609_));
 sky130_fd_sc_hd__inv_2 _10898_ (.A(net1140),
    .Y(_05033_));
 sky130_fd_sc_hd__a21oi_1 _10899_ (.A1(_03687_),
    .A2(_05033_),
    .B1(_04233_),
    .Y(_00610_));
 sky130_fd_sc_hd__mux2_1 _10900_ (.A0(net1288),
    .A1(_01991_),
    .S(_04848_),
    .X(_05034_));
 sky130_fd_sc_hd__clkbuf_1 _10901_ (.A(_05034_),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _10902_ (.A0(net1250),
    .A1(_01923_),
    .S(_04848_),
    .X(_05035_));
 sky130_fd_sc_hd__clkbuf_1 _10903_ (.A(_05035_),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_1 _10904_ (.A0(net1200),
    .A1(_01799_),
    .S(_04848_),
    .X(_05036_));
 sky130_fd_sc_hd__clkbuf_1 _10905_ (.A(_05036_),
    .X(_00613_));
 sky130_fd_sc_hd__inv_2 _10906_ (.A(_01805_),
    .Y(_05037_));
 sky130_fd_sc_hd__mux2_1 _10907_ (.A0(net1293),
    .A1(_05037_),
    .S(_04848_),
    .X(_05038_));
 sky130_fd_sc_hd__clkbuf_1 _10908_ (.A(_05038_),
    .X(_00614_));
 sky130_fd_sc_hd__mux2_1 _10909_ (.A0(net1202),
    .A1(_04432_),
    .S(_04848_),
    .X(_05039_));
 sky130_fd_sc_hd__clkbuf_1 _10910_ (.A(_05039_),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _10911_ (.A0(\genblk2[7].wave_shpr.div.b1[7] ),
    .A1(_04444_),
    .S(_04848_),
    .X(_05040_));
 sky130_fd_sc_hd__clkbuf_1 _10912_ (.A(_05040_),
    .X(_00616_));
 sky130_fd_sc_hd__mux2_1 _10913_ (.A0(net1201),
    .A1(_01819_),
    .S(_04848_),
    .X(_05041_));
 sky130_fd_sc_hd__clkbuf_1 _10914_ (.A(_05041_),
    .X(_00617_));
 sky130_fd_sc_hd__buf_4 _10915_ (.A(_03707_),
    .X(_05042_));
 sky130_fd_sc_hd__mux2_1 _10916_ (.A0(net1286),
    .A1(_01797_),
    .S(_05042_),
    .X(_05043_));
 sky130_fd_sc_hd__clkbuf_1 _10917_ (.A(_05043_),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _10918_ (.A0(net1253),
    .A1(net34),
    .S(_05042_),
    .X(_05044_));
 sky130_fd_sc_hd__clkbuf_1 _10919_ (.A(_05044_),
    .X(_00619_));
 sky130_fd_sc_hd__mux2_1 _10920_ (.A0(\genblk2[7].wave_shpr.div.b1[11] ),
    .A1(_02433_),
    .S(_05042_),
    .X(_05045_));
 sky130_fd_sc_hd__clkbuf_1 _10921_ (.A(_05045_),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _10922_ (.A0(net1301),
    .A1(_01811_),
    .S(_05042_),
    .X(_05046_));
 sky130_fd_sc_hd__clkbuf_1 _10923_ (.A(_05046_),
    .X(_00621_));
 sky130_fd_sc_hd__mux2_1 _10924_ (.A0(\genblk2[7].wave_shpr.div.b1[13] ),
    .A1(_02374_),
    .S(_05042_),
    .X(_05047_));
 sky130_fd_sc_hd__clkbuf_1 _10925_ (.A(_05047_),
    .X(_00622_));
 sky130_fd_sc_hd__a21o_1 _10926_ (.A1(_03704_),
    .A2(net484),
    .B1(_04647_),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _10927_ (.A0(\genblk2[7].wave_shpr.div.b1[15] ),
    .A1(_01365_),
    .S(_05042_),
    .X(_05048_));
 sky130_fd_sc_hd__clkbuf_1 _10928_ (.A(_05048_),
    .X(_00624_));
 sky130_fd_sc_hd__inv_2 _10929_ (.A(net758),
    .Y(_05049_));
 sky130_fd_sc_hd__o21ai_1 _10930_ (.A1(_03726_),
    .A2(_05049_),
    .B1(_03736_),
    .Y(_00625_));
 sky130_fd_sc_hd__and2_1 _10931_ (.A(_02171_),
    .B(net1234),
    .X(_05050_));
 sky130_fd_sc_hd__clkbuf_1 _10932_ (.A(_05050_),
    .X(_00626_));
 sky130_fd_sc_hd__clkbuf_4 _10933_ (.A(_02188_),
    .X(_05051_));
 sky130_fd_sc_hd__clkbuf_4 _10934_ (.A(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__and3_1 _10935_ (.A(_02152_),
    .B(\genblk2[6].wave_shpr.div.busy ),
    .C(_02186_),
    .X(_05053_));
 sky130_fd_sc_hd__clkbuf_4 _10936_ (.A(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__buf_4 _10937_ (.A(_05054_),
    .X(_05055_));
 sky130_fd_sc_hd__a22o_1 _10938_ (.A1(net792),
    .A2(_05052_),
    .B1(_05023_),
    .B2(_05055_),
    .X(_00627_));
 sky130_fd_sc_hd__buf_4 _10939_ (.A(_05054_),
    .X(_05056_));
 sky130_fd_sc_hd__a22o_1 _10940_ (.A1(net756),
    .A2(_05052_),
    .B1(_05056_),
    .B2(net792),
    .X(_00628_));
 sky130_fd_sc_hd__a22o_1 _10941_ (.A1(net671),
    .A2(_05052_),
    .B1(_05056_),
    .B2(net756),
    .X(_00629_));
 sky130_fd_sc_hd__a22o_1 _10942_ (.A1(net271),
    .A2(_05052_),
    .B1(_05056_),
    .B2(net671),
    .X(_00630_));
 sky130_fd_sc_hd__a22o_1 _10943_ (.A1(\genblk2[6].wave_shpr.div.quo[4] ),
    .A2(_05052_),
    .B1(_05056_),
    .B2(net271),
    .X(_00631_));
 sky130_fd_sc_hd__a22o_1 _10944_ (.A1(\genblk2[6].wave_shpr.div.quo[5] ),
    .A2(_05052_),
    .B1(_05056_),
    .B2(net720),
    .X(_00632_));
 sky130_fd_sc_hd__a22o_1 _10945_ (.A1(net241),
    .A2(_05052_),
    .B1(_05056_),
    .B2(net742),
    .X(_00633_));
 sky130_fd_sc_hd__a22o_1 _10946_ (.A1(\genblk2[6].wave_shpr.div.quo[7] ),
    .A2(_05052_),
    .B1(_05056_),
    .B2(net241),
    .X(_00634_));
 sky130_fd_sc_hd__a22o_1 _10947_ (.A1(net515),
    .A2(_05052_),
    .B1(_05056_),
    .B2(net523),
    .X(_00635_));
 sky130_fd_sc_hd__clkbuf_4 _10948_ (.A(_05051_),
    .X(_05057_));
 sky130_fd_sc_hd__and2_1 _10949_ (.A(_04869_),
    .B(\genblk1[6].osc.clkdiv_C.cnt[0] ),
    .X(_05058_));
 sky130_fd_sc_hd__a221o_1 _10950_ (.A1(net477),
    .A2(_05057_),
    .B1(_05055_),
    .B2(net515),
    .C1(_05058_),
    .X(_00636_));
 sky130_fd_sc_hd__clkbuf_2 _10951_ (.A(_04268_),
    .X(_05059_));
 sky130_fd_sc_hd__and2_1 _10952_ (.A(_05059_),
    .B(\genblk1[6].osc.clkdiv_C.cnt[1] ),
    .X(_05060_));
 sky130_fd_sc_hd__a221o_1 _10953_ (.A1(net344),
    .A2(_05057_),
    .B1(_05055_),
    .B2(net477),
    .C1(_05060_),
    .X(_00637_));
 sky130_fd_sc_hd__nor2_1 _10954_ (.A(_04676_),
    .B(_01729_),
    .Y(_05061_));
 sky130_fd_sc_hd__a221o_1 _10955_ (.A1(\genblk2[6].wave_shpr.div.quo[11] ),
    .A2(_05057_),
    .B1(_05055_),
    .B2(net344),
    .C1(_05061_),
    .X(_00638_));
 sky130_fd_sc_hd__buf_2 _10956_ (.A(_05051_),
    .X(_05062_));
 sky130_fd_sc_hd__and2_1 _10957_ (.A(_05059_),
    .B(\genblk1[6].osc.clkdiv_C.cnt[3] ),
    .X(_05063_));
 sky130_fd_sc_hd__a221o_1 _10958_ (.A1(\genblk2[6].wave_shpr.div.quo[12] ),
    .A2(_05062_),
    .B1(_05055_),
    .B2(net623),
    .C1(_05063_),
    .X(_00639_));
 sky130_fd_sc_hd__buf_2 _10959_ (.A(_05054_),
    .X(_05064_));
 sky130_fd_sc_hd__and2_1 _10960_ (.A(_05059_),
    .B(\genblk1[6].osc.clkdiv_C.cnt[4] ),
    .X(_05065_));
 sky130_fd_sc_hd__a221o_1 _10961_ (.A1(net620),
    .A2(_05062_),
    .B1(_05064_),
    .B2(\genblk2[6].wave_shpr.div.quo[12] ),
    .C1(_05065_),
    .X(_00640_));
 sky130_fd_sc_hd__and2_1 _10962_ (.A(_05059_),
    .B(\genblk1[6].osc.clkdiv_C.cnt[5] ),
    .X(_05066_));
 sky130_fd_sc_hd__a221o_1 _10963_ (.A1(net498),
    .A2(_05062_),
    .B1(_05064_),
    .B2(\genblk2[6].wave_shpr.div.quo[13] ),
    .C1(_05066_),
    .X(_00641_));
 sky130_fd_sc_hd__and2_1 _10964_ (.A(_05059_),
    .B(\genblk1[6].osc.clkdiv_C.cnt[6] ),
    .X(_05067_));
 sky130_fd_sc_hd__a221o_1 _10965_ (.A1(net594),
    .A2(_05062_),
    .B1(_05064_),
    .B2(net498),
    .C1(_05067_),
    .X(_00642_));
 sky130_fd_sc_hd__nor2_1 _10966_ (.A(_04676_),
    .B(_01753_),
    .Y(_05068_));
 sky130_fd_sc_hd__a221o_1 _10967_ (.A1(net595),
    .A2(_05062_),
    .B1(_05064_),
    .B2(net594),
    .C1(_05068_),
    .X(_00643_));
 sky130_fd_sc_hd__and2_1 _10968_ (.A(_05059_),
    .B(\genblk1[6].osc.clkdiv_C.cnt[8] ),
    .X(_05069_));
 sky130_fd_sc_hd__a221o_1 _10969_ (.A1(net582),
    .A2(_05062_),
    .B1(_05064_),
    .B2(net595),
    .C1(_05069_),
    .X(_00644_));
 sky130_fd_sc_hd__and2_1 _10970_ (.A(_05059_),
    .B(\genblk1[6].osc.clkdiv_C.cnt[9] ),
    .X(_05070_));
 sky130_fd_sc_hd__a221o_1 _10971_ (.A1(net486),
    .A2(_05062_),
    .B1(_05064_),
    .B2(net582),
    .C1(_05070_),
    .X(_00645_));
 sky130_fd_sc_hd__and2_1 _10972_ (.A(_05059_),
    .B(\genblk1[6].osc.clkdiv_C.cnt[10] ),
    .X(_05071_));
 sky130_fd_sc_hd__a221o_1 _10973_ (.A1(net313),
    .A2(_05062_),
    .B1(_05064_),
    .B2(net486),
    .C1(_05071_),
    .X(_00646_));
 sky130_fd_sc_hd__and2_1 _10974_ (.A(_05059_),
    .B(\genblk1[6].osc.clkdiv_C.cnt[11] ),
    .X(_05072_));
 sky130_fd_sc_hd__a221o_1 _10975_ (.A1(\genblk2[6].wave_shpr.div.quo[20] ),
    .A2(_05062_),
    .B1(_05064_),
    .B2(net313),
    .C1(_05072_),
    .X(_00647_));
 sky130_fd_sc_hd__and2_1 _10976_ (.A(_05059_),
    .B(\genblk1[6].osc.clkdiv_C.cnt[12] ),
    .X(_05073_));
 sky130_fd_sc_hd__a221o_1 _10977_ (.A1(\genblk2[6].wave_shpr.div.quo[21] ),
    .A2(_05062_),
    .B1(_05064_),
    .B2(net567),
    .C1(_05073_),
    .X(_00648_));
 sky130_fd_sc_hd__clkbuf_4 _10978_ (.A(_04268_),
    .X(_05074_));
 sky130_fd_sc_hd__and2_1 _10979_ (.A(_05074_),
    .B(\genblk1[6].osc.clkdiv_C.cnt[13] ),
    .X(_05075_));
 sky130_fd_sc_hd__a221o_1 _10980_ (.A1(net609),
    .A2(_05051_),
    .B1(_05064_),
    .B2(net616),
    .C1(_05075_),
    .X(_00649_));
 sky130_fd_sc_hd__and2_1 _10981_ (.A(_05074_),
    .B(\genblk1[6].osc.clkdiv_C.cnt[14] ),
    .X(_05076_));
 sky130_fd_sc_hd__a221o_1 _10982_ (.A1(net385),
    .A2(_05051_),
    .B1(_05054_),
    .B2(net609),
    .C1(_05076_),
    .X(_00650_));
 sky130_fd_sc_hd__and2_1 _10983_ (.A(_05074_),
    .B(\genblk1[6].osc.clkdiv_C.cnt[15] ),
    .X(_05077_));
 sky130_fd_sc_hd__a221o_1 _10984_ (.A1(\genblk2[6].wave_shpr.div.quo[24] ),
    .A2(_05051_),
    .B1(_05054_),
    .B2(net385),
    .C1(_05077_),
    .X(_00651_));
 sky130_fd_sc_hd__and2_1 _10985_ (.A(_05074_),
    .B(\genblk1[6].osc.clkdiv_C.cnt[16] ),
    .X(_05078_));
 sky130_fd_sc_hd__a221o_1 _10986_ (.A1(net283),
    .A2(_05051_),
    .B1(_05054_),
    .B2(net668),
    .C1(_05078_),
    .X(_00652_));
 sky130_fd_sc_hd__inv_2 _10987_ (.A(_05054_),
    .Y(_05079_));
 sky130_fd_sc_hd__or2_1 _10988_ (.A(_03719_),
    .B(\genblk1[6].osc.clkdiv_C.cnt[17] ),
    .X(_05080_));
 sky130_fd_sc_hd__o221a_1 _10989_ (.A1(\genblk2[6].wave_shpr.div.acc[0] ),
    .A2(_00016_),
    .B1(_05079_),
    .B2(net283),
    .C1(_05080_),
    .X(_00653_));
 sky130_fd_sc_hd__a21oi_1 _10990_ (.A1(\genblk2[6].wave_shpr.div.b1[0] ),
    .A2(_05023_),
    .B1(\genblk2[6].wave_shpr.div.acc[0] ),
    .Y(_05081_));
 sky130_fd_sc_hd__a31o_1 _10991_ (.A1(\genblk2[6].wave_shpr.div.b1[0] ),
    .A2(\genblk2[6].wave_shpr.div.acc[0] ),
    .A3(_05023_),
    .B1(_05079_),
    .X(_05082_));
 sky130_fd_sc_hd__a2bb2o_1 _10992_ (.A1_N(_05081_),
    .A2_N(_05082_),
    .B1(net1122),
    .B2(_05052_),
    .X(_00654_));
 sky130_fd_sc_hd__or2_1 _10993_ (.A(\genblk2[6].wave_shpr.div.acc[1] ),
    .B(_05022_),
    .X(_05083_));
 sky130_fd_sc_hd__xnor2_1 _10994_ (.A(_04982_),
    .B(_04983_),
    .Y(_05084_));
 sky130_fd_sc_hd__nand2_1 _10995_ (.A(_05023_),
    .B(_05084_),
    .Y(_05085_));
 sky130_fd_sc_hd__a32o_1 _10996_ (.A1(_05055_),
    .A2(_05083_),
    .A3(_05085_),
    .B1(_05057_),
    .B2(net1165),
    .X(_00655_));
 sky130_fd_sc_hd__clkbuf_4 _10997_ (.A(_05051_),
    .X(_05086_));
 sky130_fd_sc_hd__xor2_1 _10998_ (.A(\genblk2[6].wave_shpr.div.b1[2] ),
    .B(\genblk2[6].wave_shpr.div.acc[2] ),
    .X(_05087_));
 sky130_fd_sc_hd__xnor2_1 _10999_ (.A(_04985_),
    .B(_05087_),
    .Y(_05088_));
 sky130_fd_sc_hd__mux2_1 _11000_ (.A0(\genblk2[6].wave_shpr.div.acc[2] ),
    .A1(_05088_),
    .S(_05023_),
    .X(_05089_));
 sky130_fd_sc_hd__a22o_1 _11001_ (.A1(net1015),
    .A2(_05086_),
    .B1(_05056_),
    .B2(_05089_),
    .X(_00656_));
 sky130_fd_sc_hd__or2b_1 _11002_ (.A(_04988_),
    .B_N(_04980_),
    .X(_05090_));
 sky130_fd_sc_hd__xnor2_1 _11003_ (.A(_04987_),
    .B(_05090_),
    .Y(_05091_));
 sky130_fd_sc_hd__mux2_1 _11004_ (.A0(\genblk2[6].wave_shpr.div.acc[3] ),
    .A1(_05091_),
    .S(_05023_),
    .X(_05092_));
 sky130_fd_sc_hd__a22o_1 _11005_ (.A1(net986),
    .A2(_05086_),
    .B1(_05056_),
    .B2(_05092_),
    .X(_00657_));
 sky130_fd_sc_hd__clkbuf_4 _11006_ (.A(_05054_),
    .X(_05093_));
 sky130_fd_sc_hd__or2b_1 _11007_ (.A(_04990_),
    .B_N(_04979_),
    .X(_05094_));
 sky130_fd_sc_hd__xnor2_1 _11008_ (.A(_05094_),
    .B(_04989_),
    .Y(_05095_));
 sky130_fd_sc_hd__mux2_1 _11009_ (.A0(\genblk2[6].wave_shpr.div.acc[4] ),
    .A1(_05095_),
    .S(_05023_),
    .X(_05096_));
 sky130_fd_sc_hd__a22o_1 _11010_ (.A1(net907),
    .A2(_05086_),
    .B1(_05093_),
    .B2(_05096_),
    .X(_00658_));
 sky130_fd_sc_hd__or2b_1 _11011_ (.A(_04992_),
    .B_N(_04978_),
    .X(_05097_));
 sky130_fd_sc_hd__xnor2_1 _11012_ (.A(_05097_),
    .B(_04991_),
    .Y(_05098_));
 sky130_fd_sc_hd__mux2_1 _11013_ (.A0(\genblk2[6].wave_shpr.div.acc[5] ),
    .A1(_05098_),
    .S(_05023_),
    .X(_05099_));
 sky130_fd_sc_hd__a22o_1 _11014_ (.A1(net819),
    .A2(_05086_),
    .B1(_05093_),
    .B2(_05099_),
    .X(_00659_));
 sky130_fd_sc_hd__or2b_1 _11015_ (.A(_04994_),
    .B_N(_04977_),
    .X(_05100_));
 sky130_fd_sc_hd__xnor2_1 _11016_ (.A(_04993_),
    .B(_05100_),
    .Y(_05101_));
 sky130_fd_sc_hd__mux2_1 _11017_ (.A0(\genblk2[6].wave_shpr.div.acc[6] ),
    .A1(_05101_),
    .S(_05023_),
    .X(_05102_));
 sky130_fd_sc_hd__a22o_1 _11018_ (.A1(net826),
    .A2(_05086_),
    .B1(_05093_),
    .B2(_05102_),
    .X(_00660_));
 sky130_fd_sc_hd__or2b_1 _11019_ (.A(_04996_),
    .B_N(_04976_),
    .X(_05103_));
 sky130_fd_sc_hd__xnor2_1 _11020_ (.A(_04995_),
    .B(_05103_),
    .Y(_05104_));
 sky130_fd_sc_hd__clkbuf_4 _11021_ (.A(_05022_),
    .X(_05105_));
 sky130_fd_sc_hd__mux2_1 _11022_ (.A0(\genblk2[6].wave_shpr.div.acc[7] ),
    .A1(_05104_),
    .S(_05105_),
    .X(_05106_));
 sky130_fd_sc_hd__a22o_1 _11023_ (.A1(net867),
    .A2(_05086_),
    .B1(_05093_),
    .B2(_05106_),
    .X(_00661_));
 sky130_fd_sc_hd__or2b_1 _11024_ (.A(_04998_),
    .B_N(_04975_),
    .X(_05107_));
 sky130_fd_sc_hd__xnor2_1 _11025_ (.A(_04997_),
    .B(_05107_),
    .Y(_05108_));
 sky130_fd_sc_hd__mux2_1 _11026_ (.A0(\genblk2[6].wave_shpr.div.acc[8] ),
    .A1(_05108_),
    .S(_05105_),
    .X(_05109_));
 sky130_fd_sc_hd__a22o_1 _11027_ (.A1(net806),
    .A2(_05086_),
    .B1(_05093_),
    .B2(_05109_),
    .X(_00662_));
 sky130_fd_sc_hd__or2b_1 _11028_ (.A(_05000_),
    .B_N(_04974_),
    .X(_05110_));
 sky130_fd_sc_hd__xnor2_1 _11029_ (.A(_04999_),
    .B(_05110_),
    .Y(_05111_));
 sky130_fd_sc_hd__mux2_1 _11030_ (.A0(\genblk2[6].wave_shpr.div.acc[9] ),
    .A1(_05111_),
    .S(_05105_),
    .X(_05112_));
 sky130_fd_sc_hd__a22o_1 _11031_ (.A1(net1003),
    .A2(_05086_),
    .B1(_05093_),
    .B2(_05112_),
    .X(_00663_));
 sky130_fd_sc_hd__or2b_1 _11032_ (.A(_05002_),
    .B_N(_04973_),
    .X(_05113_));
 sky130_fd_sc_hd__xnor2_1 _11033_ (.A(_05001_),
    .B(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__mux2_1 _11034_ (.A0(\genblk2[6].wave_shpr.div.acc[10] ),
    .A1(_05114_),
    .S(_05105_),
    .X(_05115_));
 sky130_fd_sc_hd__a22o_1 _11035_ (.A1(net900),
    .A2(_05086_),
    .B1(_05093_),
    .B2(_05115_),
    .X(_00664_));
 sky130_fd_sc_hd__or2b_1 _11036_ (.A(_05004_),
    .B_N(_04972_),
    .X(_05116_));
 sky130_fd_sc_hd__xnor2_1 _11037_ (.A(_05003_),
    .B(_05116_),
    .Y(_05117_));
 sky130_fd_sc_hd__mux2_1 _11038_ (.A0(\genblk2[6].wave_shpr.div.acc[11] ),
    .A1(_05117_),
    .S(_05105_),
    .X(_05118_));
 sky130_fd_sc_hd__a22o_1 _11039_ (.A1(net838),
    .A2(_05086_),
    .B1(_05093_),
    .B2(_05118_),
    .X(_00665_));
 sky130_fd_sc_hd__clkbuf_4 _11040_ (.A(_05051_),
    .X(_05119_));
 sky130_fd_sc_hd__or2b_1 _11041_ (.A(_05006_),
    .B_N(_04971_),
    .X(_05120_));
 sky130_fd_sc_hd__xnor2_1 _11042_ (.A(_05005_),
    .B(_05120_),
    .Y(_05121_));
 sky130_fd_sc_hd__mux2_1 _11043_ (.A0(\genblk2[6].wave_shpr.div.acc[12] ),
    .A1(_05121_),
    .S(_05105_),
    .X(_05122_));
 sky130_fd_sc_hd__a22o_1 _11044_ (.A1(net883),
    .A2(_05119_),
    .B1(_05093_),
    .B2(_05122_),
    .X(_00666_));
 sky130_fd_sc_hd__or2b_1 _11045_ (.A(_05008_),
    .B_N(_04970_),
    .X(_05123_));
 sky130_fd_sc_hd__xnor2_1 _11046_ (.A(_05007_),
    .B(_05123_),
    .Y(_05124_));
 sky130_fd_sc_hd__mux2_1 _11047_ (.A0(\genblk2[6].wave_shpr.div.acc[13] ),
    .A1(_05124_),
    .S(_05105_),
    .X(_05125_));
 sky130_fd_sc_hd__a22o_1 _11048_ (.A1(net921),
    .A2(_05119_),
    .B1(_05093_),
    .B2(_05125_),
    .X(_00667_));
 sky130_fd_sc_hd__clkbuf_4 _11049_ (.A(_05054_),
    .X(_05126_));
 sky130_fd_sc_hd__or2b_1 _11050_ (.A(_05010_),
    .B_N(_04969_),
    .X(_05127_));
 sky130_fd_sc_hd__xnor2_1 _11051_ (.A(_05009_),
    .B(_05127_),
    .Y(_05128_));
 sky130_fd_sc_hd__mux2_1 _11052_ (.A0(\genblk2[6].wave_shpr.div.acc[14] ),
    .A1(_05128_),
    .S(_05105_),
    .X(_05129_));
 sky130_fd_sc_hd__a22o_1 _11053_ (.A1(net818),
    .A2(_05119_),
    .B1(_05126_),
    .B2(_05129_),
    .X(_00668_));
 sky130_fd_sc_hd__or2b_1 _11054_ (.A(_05012_),
    .B_N(_04968_),
    .X(_05130_));
 sky130_fd_sc_hd__xnor2_1 _11055_ (.A(_05011_),
    .B(_05130_),
    .Y(_05131_));
 sky130_fd_sc_hd__mux2_1 _11056_ (.A0(\genblk2[6].wave_shpr.div.acc[15] ),
    .A1(_05131_),
    .S(_05105_),
    .X(_05132_));
 sky130_fd_sc_hd__a22o_1 _11057_ (.A1(net1093),
    .A2(_05119_),
    .B1(_05126_),
    .B2(_05132_),
    .X(_00669_));
 sky130_fd_sc_hd__xnor2_1 _11058_ (.A(_04967_),
    .B(_05013_),
    .Y(_05133_));
 sky130_fd_sc_hd__mux2_1 _11059_ (.A0(\genblk2[6].wave_shpr.div.acc[16] ),
    .A1(_05133_),
    .S(_05105_),
    .X(_05134_));
 sky130_fd_sc_hd__a22o_1 _11060_ (.A1(net899),
    .A2(_05119_),
    .B1(_05126_),
    .B2(_05134_),
    .X(_00670_));
 sky130_fd_sc_hd__or2b_1 _11061_ (.A(_05016_),
    .B_N(_04966_),
    .X(_05135_));
 sky130_fd_sc_hd__xnor2_1 _11062_ (.A(_05015_),
    .B(_05135_),
    .Y(_05136_));
 sky130_fd_sc_hd__mux2_1 _11063_ (.A0(\genblk2[6].wave_shpr.div.acc[17] ),
    .A1(_05136_),
    .S(_05022_),
    .X(_05137_));
 sky130_fd_sc_hd__a22o_1 _11064_ (.A1(net560),
    .A2(_05119_),
    .B1(_05126_),
    .B2(_05137_),
    .X(_00671_));
 sky130_fd_sc_hd__nor4_1 _11065_ (.A(\genblk2[6].wave_shpr.div.acc[25] ),
    .B(\genblk2[6].wave_shpr.div.acc[24] ),
    .C(\genblk2[6].wave_shpr.div.acc[26] ),
    .D(_05021_),
    .Y(_05138_));
 sky130_fd_sc_hd__or2_1 _11066_ (.A(_05018_),
    .B(net21),
    .X(_05139_));
 sky130_fd_sc_hd__o21ai_1 _11067_ (.A1(_05017_),
    .A2(net21),
    .B1(\genblk2[6].wave_shpr.div.acc[18] ),
    .Y(_05140_));
 sky130_fd_sc_hd__nand2_1 _11068_ (.A(_05139_),
    .B(_05140_),
    .Y(_05141_));
 sky130_fd_sc_hd__a22o_1 _11069_ (.A1(net622),
    .A2(_05119_),
    .B1(_05126_),
    .B2(_05141_),
    .X(_00672_));
 sky130_fd_sc_hd__nor2_1 _11070_ (.A(_05019_),
    .B(net21),
    .Y(_05142_));
 sky130_fd_sc_hd__a21o_1 _11071_ (.A1(net622),
    .A2(_05139_),
    .B1(_05142_),
    .X(_05143_));
 sky130_fd_sc_hd__a22o_1 _11072_ (.A1(net1138),
    .A2(_05119_),
    .B1(_05126_),
    .B2(_05143_),
    .X(_00673_));
 sky130_fd_sc_hd__xor2_1 _11073_ (.A(\genblk2[6].wave_shpr.div.acc[20] ),
    .B(_05142_),
    .X(_05144_));
 sky130_fd_sc_hd__a22o_1 _11074_ (.A1(net1001),
    .A2(_05119_),
    .B1(_05126_),
    .B2(_05144_),
    .X(_00674_));
 sky130_fd_sc_hd__or3_1 _11075_ (.A(\genblk2[6].wave_shpr.div.acc[20] ),
    .B(_05019_),
    .C(net1350),
    .X(_05145_));
 sky130_fd_sc_hd__or4_1 _11076_ (.A(\genblk2[6].wave_shpr.div.acc[21] ),
    .B(\genblk2[6].wave_shpr.div.acc[20] ),
    .C(_05019_),
    .D(net1350),
    .X(_05146_));
 sky130_fd_sc_hd__a21bo_1 _11077_ (.A1(\genblk2[6].wave_shpr.div.acc[21] ),
    .A2(_05145_),
    .B1_N(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__a22o_1 _11078_ (.A1(net1031),
    .A2(_05119_),
    .B1(_05126_),
    .B2(_05147_),
    .X(_00675_));
 sky130_fd_sc_hd__xnor2_1 _11079_ (.A(\genblk2[6].wave_shpr.div.acc[22] ),
    .B(_05146_),
    .Y(_05148_));
 sky130_fd_sc_hd__a22o_1 _11080_ (.A1(net659),
    .A2(_05057_),
    .B1(_05126_),
    .B2(_05148_),
    .X(_00676_));
 sky130_fd_sc_hd__nor2_1 _11081_ (.A(_05021_),
    .B(_05138_),
    .Y(_05149_));
 sky130_fd_sc_hd__a21o_1 _11082_ (.A1(\genblk2[6].wave_shpr.div.acc[23] ),
    .A2(_05020_),
    .B1(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__a22o_1 _11083_ (.A1(\genblk2[6].wave_shpr.div.acc[24] ),
    .A2(_05057_),
    .B1(_05126_),
    .B2(_05150_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _11084_ (.A0(_05149_),
    .A1(_05021_),
    .S(\genblk2[6].wave_shpr.div.acc[24] ),
    .X(_05151_));
 sky130_fd_sc_hd__a22o_1 _11085_ (.A1(net1076),
    .A2(_05057_),
    .B1(_05055_),
    .B2(_05151_),
    .X(_00678_));
 sky130_fd_sc_hd__o21ai_1 _11086_ (.A1(\genblk2[6].wave_shpr.div.acc[24] ),
    .A2(_05021_),
    .B1(\genblk2[6].wave_shpr.div.acc[25] ),
    .Y(_05152_));
 sky130_fd_sc_hd__or4b_1 _11087_ (.A(\genblk2[6].wave_shpr.div.acc[25] ),
    .B(_05021_),
    .C(\genblk2[6].wave_shpr.div.acc[24] ),
    .D_N(\genblk2[6].wave_shpr.div.acc[26] ),
    .X(_05153_));
 sky130_fd_sc_hd__nand2_1 _11088_ (.A(_05152_),
    .B(_05153_),
    .Y(_05154_));
 sky130_fd_sc_hd__a22o_1 _11089_ (.A1(net1043),
    .A2(_05057_),
    .B1(_05055_),
    .B2(_05154_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _11090_ (.A0(_05054_),
    .A1(_05051_),
    .S(\genblk2[6].wave_shpr.div.i[0] ),
    .X(_05155_));
 sky130_fd_sc_hd__clkbuf_1 _11091_ (.A(_05155_),
    .X(_00680_));
 sky130_fd_sc_hd__or2_1 _11092_ (.A(\genblk2[6].wave_shpr.div.i[1] ),
    .B(\genblk2[6].wave_shpr.div.i[0] ),
    .X(_05156_));
 sky130_fd_sc_hd__nand2_1 _11093_ (.A(\genblk2[6].wave_shpr.div.i[1] ),
    .B(\genblk2[6].wave_shpr.div.i[0] ),
    .Y(_05157_));
 sky130_fd_sc_hd__a32o_1 _11094_ (.A1(_05055_),
    .A2(_05156_),
    .A3(_05157_),
    .B1(_05057_),
    .B2(net1130),
    .X(_00681_));
 sky130_fd_sc_hd__a21o_1 _11095_ (.A1(\genblk2[6].wave_shpr.div.i[1] ),
    .A2(\genblk2[6].wave_shpr.div.i[0] ),
    .B1(\genblk2[6].wave_shpr.div.i[2] ),
    .X(_05158_));
 sky130_fd_sc_hd__and3_1 _11096_ (.A(\genblk2[6].wave_shpr.div.i[1] ),
    .B(\genblk2[6].wave_shpr.div.i[0] ),
    .C(\genblk2[6].wave_shpr.div.i[2] ),
    .X(_05159_));
 sky130_fd_sc_hd__inv_2 _11097_ (.A(_05159_),
    .Y(_05160_));
 sky130_fd_sc_hd__a32o_1 _11098_ (.A1(_05055_),
    .A2(_05158_),
    .A3(_05160_),
    .B1(_05057_),
    .B2(net739),
    .X(_00682_));
 sky130_fd_sc_hd__a21oi_1 _11099_ (.A1(_00016_),
    .A2(_05159_),
    .B1(net1177),
    .Y(_05161_));
 sky130_fd_sc_hd__and3_1 _11100_ (.A(\genblk2[6].wave_shpr.div.i[3] ),
    .B(_02187_),
    .C(_05159_),
    .X(_05162_));
 sky130_fd_sc_hd__nor3_1 _11101_ (.A(_03690_),
    .B(_05161_),
    .C(_05162_),
    .Y(_00683_));
 sky130_fd_sc_hd__o21ai_1 _11102_ (.A1(net280),
    .A2(_05162_),
    .B1(_03855_),
    .Y(_05163_));
 sky130_fd_sc_hd__a21oi_1 _11103_ (.A1(net280),
    .A2(_05162_),
    .B1(_05163_),
    .Y(_00684_));
 sky130_fd_sc_hd__or2b_1 _11104_ (.A(\genblk2[7].wave_shpr.div.acc[17] ),
    .B_N(\genblk2[7].wave_shpr.div.b1[17] ),
    .X(_05164_));
 sky130_fd_sc_hd__nor2_1 _11105_ (.A(_05049_),
    .B(\genblk2[7].wave_shpr.div.acc[16] ),
    .Y(_05165_));
 sky130_fd_sc_hd__or2b_1 _11106_ (.A(\genblk2[7].wave_shpr.div.acc[15] ),
    .B_N(\genblk2[7].wave_shpr.div.b1[15] ),
    .X(_05166_));
 sky130_fd_sc_hd__or2b_1 _11107_ (.A(\genblk2[7].wave_shpr.div.acc[14] ),
    .B_N(\genblk2[7].wave_shpr.div.b1[14] ),
    .X(_05167_));
 sky130_fd_sc_hd__or2b_1 _11108_ (.A(\genblk2[7].wave_shpr.div.acc[13] ),
    .B_N(\genblk2[7].wave_shpr.div.b1[13] ),
    .X(_05168_));
 sky130_fd_sc_hd__or2b_1 _11109_ (.A(\genblk2[7].wave_shpr.div.acc[12] ),
    .B_N(\genblk2[7].wave_shpr.div.b1[12] ),
    .X(_05169_));
 sky130_fd_sc_hd__or2b_1 _11110_ (.A(\genblk2[7].wave_shpr.div.acc[11] ),
    .B_N(\genblk2[7].wave_shpr.div.b1[11] ),
    .X(_05170_));
 sky130_fd_sc_hd__or2b_1 _11111_ (.A(\genblk2[7].wave_shpr.div.acc[10] ),
    .B_N(\genblk2[7].wave_shpr.div.b1[10] ),
    .X(_05171_));
 sky130_fd_sc_hd__or2b_1 _11112_ (.A(\genblk2[7].wave_shpr.div.acc[9] ),
    .B_N(\genblk2[7].wave_shpr.div.b1[9] ),
    .X(_05172_));
 sky130_fd_sc_hd__or2b_1 _11113_ (.A(\genblk2[7].wave_shpr.div.acc[8] ),
    .B_N(\genblk2[7].wave_shpr.div.b1[8] ),
    .X(_05173_));
 sky130_fd_sc_hd__or2b_1 _11114_ (.A(\genblk2[7].wave_shpr.div.acc[7] ),
    .B_N(\genblk2[7].wave_shpr.div.b1[7] ),
    .X(_05174_));
 sky130_fd_sc_hd__or2b_1 _11115_ (.A(\genblk2[7].wave_shpr.div.acc[6] ),
    .B_N(\genblk2[7].wave_shpr.div.b1[6] ),
    .X(_05175_));
 sky130_fd_sc_hd__or2b_1 _11116_ (.A(\genblk2[7].wave_shpr.div.acc[5] ),
    .B_N(\genblk2[7].wave_shpr.div.b1[5] ),
    .X(_05176_));
 sky130_fd_sc_hd__or2b_1 _11117_ (.A(\genblk2[7].wave_shpr.div.b1[4] ),
    .B_N(\genblk2[7].wave_shpr.div.acc[4] ),
    .X(_05177_));
 sky130_fd_sc_hd__or2b_1 _11118_ (.A(\genblk2[7].wave_shpr.div.acc[4] ),
    .B_N(\genblk2[7].wave_shpr.div.b1[4] ),
    .X(_05178_));
 sky130_fd_sc_hd__nand2_1 _11119_ (.A(_05177_),
    .B(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hd__or2b_1 _11120_ (.A(\genblk2[7].wave_shpr.div.acc[3] ),
    .B_N(\genblk2[7].wave_shpr.div.b1[3] ),
    .X(_05180_));
 sky130_fd_sc_hd__or2b_1 _11121_ (.A(\genblk2[7].wave_shpr.div.acc[2] ),
    .B_N(\genblk2[7].wave_shpr.div.b1[2] ),
    .X(_05181_));
 sky130_fd_sc_hd__inv_2 _11122_ (.A(\genblk2[7].wave_shpr.div.acc[0] ),
    .Y(_05182_));
 sky130_fd_sc_hd__xor2_1 _11123_ (.A(\genblk2[7].wave_shpr.div.b1[1] ),
    .B(\genblk2[7].wave_shpr.div.acc[1] ),
    .X(_05183_));
 sky130_fd_sc_hd__a21oi_1 _11124_ (.A1(\genblk2[7].wave_shpr.div.b1[0] ),
    .A2(_05182_),
    .B1(_05183_),
    .Y(_05184_));
 sky130_fd_sc_hd__a21o_1 _11125_ (.A1(_05033_),
    .A2(\genblk2[7].wave_shpr.div.acc[1] ),
    .B1(_05184_),
    .X(_05185_));
 sky130_fd_sc_hd__and2b_1 _11126_ (.A_N(\genblk2[7].wave_shpr.div.b1[2] ),
    .B(\genblk2[7].wave_shpr.div.acc[2] ),
    .X(_05186_));
 sky130_fd_sc_hd__a21o_1 _11127_ (.A1(_05181_),
    .A2(_05185_),
    .B1(_05186_),
    .X(_05187_));
 sky130_fd_sc_hd__and2b_1 _11128_ (.A_N(\genblk2[7].wave_shpr.div.b1[3] ),
    .B(\genblk2[7].wave_shpr.div.acc[3] ),
    .X(_05188_));
 sky130_fd_sc_hd__a21oi_1 _11129_ (.A1(_05180_),
    .A2(_05187_),
    .B1(_05188_),
    .Y(_05189_));
 sky130_fd_sc_hd__o21ai_1 _11130_ (.A1(_05179_),
    .A2(_05189_),
    .B1(_05177_),
    .Y(_05190_));
 sky130_fd_sc_hd__and2b_1 _11131_ (.A_N(\genblk2[7].wave_shpr.div.b1[5] ),
    .B(\genblk2[7].wave_shpr.div.acc[5] ),
    .X(_05191_));
 sky130_fd_sc_hd__a21o_1 _11132_ (.A1(_05176_),
    .A2(_05190_),
    .B1(_05191_),
    .X(_05192_));
 sky130_fd_sc_hd__and2b_1 _11133_ (.A_N(\genblk2[7].wave_shpr.div.b1[6] ),
    .B(\genblk2[7].wave_shpr.div.acc[6] ),
    .X(_05193_));
 sky130_fd_sc_hd__a21o_1 _11134_ (.A1(_05175_),
    .A2(_05192_),
    .B1(_05193_),
    .X(_05194_));
 sky130_fd_sc_hd__and2b_1 _11135_ (.A_N(\genblk2[7].wave_shpr.div.b1[7] ),
    .B(\genblk2[7].wave_shpr.div.acc[7] ),
    .X(_05195_));
 sky130_fd_sc_hd__a21o_1 _11136_ (.A1(_05174_),
    .A2(_05194_),
    .B1(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__and2b_1 _11137_ (.A_N(\genblk2[7].wave_shpr.div.b1[8] ),
    .B(\genblk2[7].wave_shpr.div.acc[8] ),
    .X(_05197_));
 sky130_fd_sc_hd__a21o_1 _11138_ (.A1(_05173_),
    .A2(_05196_),
    .B1(_05197_),
    .X(_05198_));
 sky130_fd_sc_hd__and2b_1 _11139_ (.A_N(\genblk2[7].wave_shpr.div.b1[9] ),
    .B(\genblk2[7].wave_shpr.div.acc[9] ),
    .X(_05199_));
 sky130_fd_sc_hd__a21o_1 _11140_ (.A1(_05172_),
    .A2(_05198_),
    .B1(_05199_),
    .X(_05200_));
 sky130_fd_sc_hd__and2b_1 _11141_ (.A_N(\genblk2[7].wave_shpr.div.b1[10] ),
    .B(\genblk2[7].wave_shpr.div.acc[10] ),
    .X(_05201_));
 sky130_fd_sc_hd__a21o_1 _11142_ (.A1(_05171_),
    .A2(_05200_),
    .B1(_05201_),
    .X(_05202_));
 sky130_fd_sc_hd__and2b_1 _11143_ (.A_N(\genblk2[7].wave_shpr.div.b1[11] ),
    .B(\genblk2[7].wave_shpr.div.acc[11] ),
    .X(_05203_));
 sky130_fd_sc_hd__a21o_1 _11144_ (.A1(_05170_),
    .A2(_05202_),
    .B1(_05203_),
    .X(_05204_));
 sky130_fd_sc_hd__and2b_1 _11145_ (.A_N(\genblk2[7].wave_shpr.div.b1[12] ),
    .B(\genblk2[7].wave_shpr.div.acc[12] ),
    .X(_05205_));
 sky130_fd_sc_hd__a21o_1 _11146_ (.A1(_05169_),
    .A2(_05204_),
    .B1(_05205_),
    .X(_05206_));
 sky130_fd_sc_hd__and2b_1 _11147_ (.A_N(\genblk2[7].wave_shpr.div.b1[13] ),
    .B(\genblk2[7].wave_shpr.div.acc[13] ),
    .X(_05207_));
 sky130_fd_sc_hd__a21o_1 _11148_ (.A1(_05168_),
    .A2(_05206_),
    .B1(_05207_),
    .X(_05208_));
 sky130_fd_sc_hd__and2b_1 _11149_ (.A_N(\genblk2[7].wave_shpr.div.b1[14] ),
    .B(\genblk2[7].wave_shpr.div.acc[14] ),
    .X(_05209_));
 sky130_fd_sc_hd__a21o_1 _11150_ (.A1(_05167_),
    .A2(_05208_),
    .B1(_05209_),
    .X(_05210_));
 sky130_fd_sc_hd__and2b_1 _11151_ (.A_N(\genblk2[7].wave_shpr.div.b1[15] ),
    .B(\genblk2[7].wave_shpr.div.acc[15] ),
    .X(_05211_));
 sky130_fd_sc_hd__a21oi_1 _11152_ (.A1(_05166_),
    .A2(_05210_),
    .B1(_05211_),
    .Y(_05212_));
 sky130_fd_sc_hd__and2_1 _11153_ (.A(_05049_),
    .B(\genblk2[7].wave_shpr.div.acc[16] ),
    .X(_05213_));
 sky130_fd_sc_hd__o21bai_2 _11154_ (.A1(_05165_),
    .A2(_05212_),
    .B1_N(_05213_),
    .Y(_05214_));
 sky130_fd_sc_hd__and2b_1 _11155_ (.A_N(\genblk2[7].wave_shpr.div.b1[17] ),
    .B(\genblk2[7].wave_shpr.div.acc[17] ),
    .X(_05215_));
 sky130_fd_sc_hd__a21o_1 _11156_ (.A1(_05164_),
    .A2(_05214_),
    .B1(_05215_),
    .X(_05216_));
 sky130_fd_sc_hd__or2_1 _11157_ (.A(\genblk2[7].wave_shpr.div.acc[18] ),
    .B(_05216_),
    .X(_05217_));
 sky130_fd_sc_hd__or4_1 _11158_ (.A(\genblk2[7].wave_shpr.div.acc[21] ),
    .B(\genblk2[7].wave_shpr.div.acc[20] ),
    .C(\genblk2[7].wave_shpr.div.acc[19] ),
    .D(_05217_),
    .X(_05218_));
 sky130_fd_sc_hd__or2_2 _11159_ (.A(\genblk2[7].wave_shpr.div.acc[22] ),
    .B(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__or4_2 _11160_ (.A(\genblk2[7].wave_shpr.div.acc[23] ),
    .B(\genblk2[7].wave_shpr.div.acc[25] ),
    .C(\genblk2[7].wave_shpr.div.acc[24] ),
    .D(\genblk2[7].wave_shpr.div.acc[26] ),
    .X(_05220_));
 sky130_fd_sc_hd__or2_1 _11161_ (.A(_05219_),
    .B(_05220_),
    .X(_05221_));
 sky130_fd_sc_hd__clkbuf_4 _11162_ (.A(_05221_),
    .X(_05222_));
 sky130_fd_sc_hd__mux2_1 _11163_ (.A0(\genblk2[7].wave_shpr.div.fin_quo[0] ),
    .A1(_05222_),
    .S(_00019_),
    .X(_05223_));
 sky130_fd_sc_hd__clkbuf_1 _11164_ (.A(_05223_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _11165_ (.A0(\genblk2[7].wave_shpr.div.fin_quo[1] ),
    .A1(net1347),
    .S(_00019_),
    .X(_05224_));
 sky130_fd_sc_hd__clkbuf_1 _11166_ (.A(_05224_),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _11167_ (.A0(\genblk2[7].wave_shpr.div.fin_quo[2] ),
    .A1(net1311),
    .S(_00019_),
    .X(_05225_));
 sky130_fd_sc_hd__clkbuf_1 _11168_ (.A(_05225_),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _11169_ (.A0(\genblk2[7].wave_shpr.div.fin_quo[3] ),
    .A1(\genblk2[7].wave_shpr.div.quo[2] ),
    .S(_00019_),
    .X(_05226_));
 sky130_fd_sc_hd__clkbuf_1 _11170_ (.A(_05226_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _11171_ (.A0(\genblk2[7].wave_shpr.div.fin_quo[4] ),
    .A1(net1318),
    .S(_00019_),
    .X(_05227_));
 sky130_fd_sc_hd__clkbuf_1 _11172_ (.A(_05227_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _11173_ (.A0(\genblk2[7].wave_shpr.div.fin_quo[5] ),
    .A1(\genblk2[7].wave_shpr.div.quo[4] ),
    .S(_00019_),
    .X(_05228_));
 sky130_fd_sc_hd__clkbuf_1 _11174_ (.A(_05228_),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _11175_ (.A0(\genblk2[7].wave_shpr.div.fin_quo[6] ),
    .A1(net754),
    .S(_00019_),
    .X(_05229_));
 sky130_fd_sc_hd__clkbuf_1 _11176_ (.A(_05229_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _11177_ (.A0(net1215),
    .A1(\genblk2[7].wave_shpr.div.quo[6] ),
    .S(_00019_),
    .X(_05230_));
 sky130_fd_sc_hd__clkbuf_1 _11178_ (.A(net1216),
    .X(_00692_));
 sky130_fd_sc_hd__a21bo_1 _11179_ (.A1(_03831_),
    .A2(net864),
    .B1_N(_03705_),
    .X(_00693_));
 sky130_fd_sc_hd__or2_1 _11180_ (.A(_03708_),
    .B(\genblk2[8].wave_shpr.div.b1[1] ),
    .X(_05231_));
 sky130_fd_sc_hd__o31a_1 _11181_ (.A1(_03819_),
    .A2(_01242_),
    .A3(_02064_),
    .B1(_05231_),
    .X(_00694_));
 sky130_fd_sc_hd__o21a_1 _11182_ (.A1(_03732_),
    .A2(net389),
    .B1(_04241_),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _11183_ (.A0(net1214),
    .A1(_04242_),
    .S(_05042_),
    .X(_05232_));
 sky130_fd_sc_hd__clkbuf_1 _11184_ (.A(_05232_),
    .X(_00696_));
 sky130_fd_sc_hd__a2bb2o_1 _11185_ (.A1_N(_03727_),
    .A2_N(_01432_),
    .B1(net593),
    .B2(_03687_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _11186_ (.A0(\genblk2[8].wave_shpr.div.b1[5] ),
    .A1(_01508_),
    .S(_05042_),
    .X(_05233_));
 sky130_fd_sc_hd__clkbuf_1 _11187_ (.A(_05233_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _11188_ (.A0(\genblk2[8].wave_shpr.div.b1[6] ),
    .A1(_01507_),
    .S(_05042_),
    .X(_05234_));
 sky130_fd_sc_hd__clkbuf_1 _11189_ (.A(_05234_),
    .X(_00699_));
 sky130_fd_sc_hd__a21bo_1 _11190_ (.A1(_03831_),
    .A2(net768),
    .B1_N(_04241_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _11191_ (.A0(net1280),
    .A1(_01556_),
    .S(_05042_),
    .X(_05235_));
 sky130_fd_sc_hd__clkbuf_1 _11192_ (.A(_05235_),
    .X(_00701_));
 sky130_fd_sc_hd__inv_2 _11193_ (.A(_01865_),
    .Y(_05236_));
 sky130_fd_sc_hd__clkbuf_4 _11194_ (.A(_03707_),
    .X(_05237_));
 sky130_fd_sc_hd__mux2_1 _11195_ (.A0(net1246),
    .A1(_05236_),
    .S(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__clkbuf_1 _11196_ (.A(_05238_),
    .X(_00702_));
 sky130_fd_sc_hd__inv_2 _11197_ (.A(_01859_),
    .Y(_05239_));
 sky130_fd_sc_hd__mux2_1 _11198_ (.A0(\genblk2[8].wave_shpr.div.b1[10] ),
    .A1(_05239_),
    .S(_05237_),
    .X(_05240_));
 sky130_fd_sc_hd__clkbuf_1 _11199_ (.A(_05240_),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _11200_ (.A0(\genblk2[8].wave_shpr.div.b1[11] ),
    .A1(_01565_),
    .S(_05237_),
    .X(_05241_));
 sky130_fd_sc_hd__clkbuf_1 _11201_ (.A(_05241_),
    .X(_00704_));
 sky130_fd_sc_hd__nor2_1 _11202_ (.A(_03702_),
    .B(net1147),
    .Y(_05242_));
 sky130_fd_sc_hd__a21oi_1 _11203_ (.A1(_03726_),
    .A2(_01869_),
    .B1(_05242_),
    .Y(_00705_));
 sky130_fd_sc_hd__a2bb2o_1 _11204_ (.A1_N(_03727_),
    .A2_N(_01490_),
    .B1(_03687_),
    .B2(net1005),
    .X(_00706_));
 sky130_fd_sc_hd__a21bo_1 _11205_ (.A1(_03831_),
    .A2(net722),
    .B1_N(_03728_),
    .X(_00707_));
 sky130_fd_sc_hd__a21bo_1 _11206_ (.A1(_03831_),
    .A2(net391),
    .B1_N(_03717_),
    .X(_00708_));
 sky130_fd_sc_hd__inv_2 _11207_ (.A(net703),
    .Y(_05243_));
 sky130_fd_sc_hd__o21ai_1 _11208_ (.A1(_03726_),
    .A2(_05243_),
    .B1(_03736_),
    .Y(_00709_));
 sky130_fd_sc_hd__and2_1 _11209_ (.A(_02171_),
    .B(net1191),
    .X(_05244_));
 sky130_fd_sc_hd__clkbuf_1 _11210_ (.A(_05244_),
    .X(_00710_));
 sky130_fd_sc_hd__clkbuf_4 _11211_ (.A(_02193_),
    .X(_05245_));
 sky130_fd_sc_hd__clkbuf_4 _11212_ (.A(_05245_),
    .X(_05246_));
 sky130_fd_sc_hd__and3_1 _11213_ (.A(_02170_),
    .B(\genblk2[7].wave_shpr.div.busy ),
    .C(_02191_),
    .X(_05247_));
 sky130_fd_sc_hd__clkbuf_4 _11214_ (.A(_05247_),
    .X(_05248_));
 sky130_fd_sc_hd__a22o_1 _11215_ (.A1(net822),
    .A2(_05246_),
    .B1(_05222_),
    .B2(_05248_),
    .X(_00711_));
 sky130_fd_sc_hd__clkbuf_4 _11216_ (.A(_05247_),
    .X(_05249_));
 sky130_fd_sc_hd__clkbuf_4 _11217_ (.A(_05249_),
    .X(_05250_));
 sky130_fd_sc_hd__a22o_1 _11218_ (.A1(net563),
    .A2(_05246_),
    .B1(_05250_),
    .B2(net822),
    .X(_00712_));
 sky130_fd_sc_hd__a22o_1 _11219_ (.A1(\genblk2[7].wave_shpr.div.quo[2] ),
    .A2(_05246_),
    .B1(_05250_),
    .B2(net563),
    .X(_00713_));
 sky130_fd_sc_hd__a22o_1 _11220_ (.A1(net331),
    .A2(_05246_),
    .B1(_05250_),
    .B2(net693),
    .X(_00714_));
 sky130_fd_sc_hd__a22o_1 _11221_ (.A1(\genblk2[7].wave_shpr.div.quo[4] ),
    .A2(_05246_),
    .B1(_05250_),
    .B2(net331),
    .X(_00715_));
 sky130_fd_sc_hd__a22o_1 _11222_ (.A1(\genblk2[7].wave_shpr.div.quo[5] ),
    .A2(_05246_),
    .B1(_05250_),
    .B2(net661),
    .X(_00716_));
 sky130_fd_sc_hd__a22o_1 _11223_ (.A1(net317),
    .A2(_05246_),
    .B1(_05250_),
    .B2(net754),
    .X(_00717_));
 sky130_fd_sc_hd__a22o_1 _11224_ (.A1(\genblk2[7].wave_shpr.div.quo[7] ),
    .A2(_05246_),
    .B1(_05250_),
    .B2(net317),
    .X(_00718_));
 sky130_fd_sc_hd__a22o_1 _11225_ (.A1(\genblk2[7].wave_shpr.div.quo[8] ),
    .A2(_05246_),
    .B1(_05250_),
    .B2(net421),
    .X(_00719_));
 sky130_fd_sc_hd__clkbuf_4 _11226_ (.A(_05245_),
    .X(_05251_));
 sky130_fd_sc_hd__and2_1 _11227_ (.A(_05074_),
    .B(\genblk1[7].osc.clkdiv_C.cnt[0] ),
    .X(_05252_));
 sky130_fd_sc_hd__a221o_1 _11228_ (.A1(net302),
    .A2(_05251_),
    .B1(_05248_),
    .B2(net492),
    .C1(_05252_),
    .X(_00720_));
 sky130_fd_sc_hd__and2_1 _11229_ (.A(_05074_),
    .B(\genblk1[7].osc.clkdiv_C.cnt[1] ),
    .X(_05253_));
 sky130_fd_sc_hd__a221o_1 _11230_ (.A1(\genblk2[7].wave_shpr.div.quo[10] ),
    .A2(_05251_),
    .B1(_05248_),
    .B2(net302),
    .C1(_05253_),
    .X(_00721_));
 sky130_fd_sc_hd__and2_1 _11231_ (.A(_05074_),
    .B(\genblk1[7].osc.clkdiv_C.cnt[2] ),
    .X(_05254_));
 sky130_fd_sc_hd__a221o_1 _11232_ (.A1(net370),
    .A2(_05251_),
    .B1(_05248_),
    .B2(net736),
    .C1(_05254_),
    .X(_00722_));
 sky130_fd_sc_hd__buf_2 _11233_ (.A(_05245_),
    .X(_05255_));
 sky130_fd_sc_hd__buf_2 _11234_ (.A(_05249_),
    .X(_05256_));
 sky130_fd_sc_hd__and2_1 _11235_ (.A(_05074_),
    .B(\genblk1[7].osc.clkdiv_C.cnt[3] ),
    .X(_05257_));
 sky130_fd_sc_hd__a221o_1 _11236_ (.A1(\genblk2[7].wave_shpr.div.quo[12] ),
    .A2(_05255_),
    .B1(_05256_),
    .B2(net370),
    .C1(_05257_),
    .X(_00723_));
 sky130_fd_sc_hd__and2_1 _11237_ (.A(_05074_),
    .B(\genblk1[7].osc.clkdiv_C.cnt[4] ),
    .X(_05258_));
 sky130_fd_sc_hd__a221o_1 _11238_ (.A1(net640),
    .A2(_05255_),
    .B1(_05256_),
    .B2(net670),
    .C1(_05258_),
    .X(_00724_));
 sky130_fd_sc_hd__and2_1 _11239_ (.A(_05074_),
    .B(\genblk1[7].osc.clkdiv_C.cnt[5] ),
    .X(_05259_));
 sky130_fd_sc_hd__a221o_1 _11240_ (.A1(net613),
    .A2(_05255_),
    .B1(_05256_),
    .B2(net640),
    .C1(_05259_),
    .X(_00725_));
 sky130_fd_sc_hd__clkbuf_2 _11241_ (.A(_04268_),
    .X(_05260_));
 sky130_fd_sc_hd__and2_1 _11242_ (.A(_05260_),
    .B(\genblk1[7].osc.clkdiv_C.cnt[6] ),
    .X(_05261_));
 sky130_fd_sc_hd__a221o_1 _11243_ (.A1(net550),
    .A2(_05255_),
    .B1(_05256_),
    .B2(net613),
    .C1(_05261_),
    .X(_00726_));
 sky130_fd_sc_hd__and2_1 _11244_ (.A(_05260_),
    .B(\genblk1[7].osc.clkdiv_C.cnt[7] ),
    .X(_05262_));
 sky130_fd_sc_hd__a221o_1 _11245_ (.A1(net548),
    .A2(_05255_),
    .B1(_05256_),
    .B2(net550),
    .C1(_05262_),
    .X(_00727_));
 sky130_fd_sc_hd__and2_1 _11246_ (.A(_05260_),
    .B(\genblk1[7].osc.clkdiv_C.cnt[8] ),
    .X(_05263_));
 sky130_fd_sc_hd__a221o_1 _11247_ (.A1(\genblk2[7].wave_shpr.div.quo[17] ),
    .A2(_05255_),
    .B1(_05256_),
    .B2(net548),
    .C1(_05263_),
    .X(_00728_));
 sky130_fd_sc_hd__and2_1 _11248_ (.A(_05260_),
    .B(\genblk1[7].osc.clkdiv_C.cnt[9] ),
    .X(_05264_));
 sky130_fd_sc_hd__a221o_1 _11249_ (.A1(net400),
    .A2(_05255_),
    .B1(_05256_),
    .B2(net585),
    .C1(_05264_),
    .X(_00729_));
 sky130_fd_sc_hd__and2_1 _11250_ (.A(_05260_),
    .B(\genblk1[7].osc.clkdiv_C.cnt[10] ),
    .X(_05265_));
 sky130_fd_sc_hd__a221o_1 _11251_ (.A1(net231),
    .A2(_05255_),
    .B1(_05256_),
    .B2(net400),
    .C1(_05265_),
    .X(_00730_));
 sky130_fd_sc_hd__and2_1 _11252_ (.A(_05260_),
    .B(\genblk1[7].osc.clkdiv_C.cnt[11] ),
    .X(_05266_));
 sky130_fd_sc_hd__a221o_1 _11253_ (.A1(\genblk2[7].wave_shpr.div.quo[20] ),
    .A2(_05255_),
    .B1(_05256_),
    .B2(net231),
    .C1(_05266_),
    .X(_00731_));
 sky130_fd_sc_hd__and2_1 _11254_ (.A(_05260_),
    .B(\genblk1[7].osc.clkdiv_C.cnt[12] ),
    .X(_05267_));
 sky130_fd_sc_hd__a221o_1 _11255_ (.A1(\genblk2[7].wave_shpr.div.quo[21] ),
    .A2(_05255_),
    .B1(_05256_),
    .B2(net527),
    .C1(_05267_),
    .X(_00732_));
 sky130_fd_sc_hd__and2_1 _11256_ (.A(_05260_),
    .B(\genblk1[7].osc.clkdiv_C.cnt[13] ),
    .X(_05268_));
 sky130_fd_sc_hd__a221o_1 _11257_ (.A1(net487),
    .A2(_05245_),
    .B1(_05249_),
    .B2(net542),
    .C1(_05268_),
    .X(_00733_));
 sky130_fd_sc_hd__and2_1 _11258_ (.A(_05260_),
    .B(\genblk1[7].osc.clkdiv_C.cnt[14] ),
    .X(_05269_));
 sky130_fd_sc_hd__a221o_1 _11259_ (.A1(\genblk2[7].wave_shpr.div.quo[23] ),
    .A2(_05245_),
    .B1(_05249_),
    .B2(net487),
    .C1(_05269_),
    .X(_00734_));
 sky130_fd_sc_hd__and2_1 _11260_ (.A(_05260_),
    .B(\genblk1[7].osc.clkdiv_C.cnt[15] ),
    .X(_05270_));
 sky130_fd_sc_hd__a221o_1 _11261_ (.A1(net534),
    .A2(_05245_),
    .B1(_05249_),
    .B2(\genblk2[7].wave_shpr.div.quo[23] ),
    .C1(_05270_),
    .X(_00735_));
 sky130_fd_sc_hd__nor2_1 _11262_ (.A(_04676_),
    .B(_01813_),
    .Y(_05271_));
 sky130_fd_sc_hd__a221o_1 _11263_ (.A1(net540),
    .A2(_05245_),
    .B1(_05249_),
    .B2(net534),
    .C1(_05271_),
    .X(_00736_));
 sky130_fd_sc_hd__or2b_1 _11264_ (.A(net540),
    .B_N(_05249_),
    .X(_05272_));
 sky130_fd_sc_hd__o221a_1 _11265_ (.A1(_03819_),
    .A2(net1255),
    .B1(_00018_),
    .B2(\genblk2[7].wave_shpr.div.acc[0] ),
    .C1(_05272_),
    .X(_00737_));
 sky130_fd_sc_hd__nor2_2 _11266_ (.A(_05219_),
    .B(_05220_),
    .Y(_05273_));
 sky130_fd_sc_hd__or3b_1 _11267_ (.A(_05273_),
    .B(_05182_),
    .C_N(\genblk2[7].wave_shpr.div.b1[0] ),
    .X(_05274_));
 sky130_fd_sc_hd__a21o_1 _11268_ (.A1(\genblk2[7].wave_shpr.div.b1[0] ),
    .A2(_05222_),
    .B1(\genblk2[7].wave_shpr.div.acc[0] ),
    .X(_05275_));
 sky130_fd_sc_hd__a32o_1 _11269_ (.A1(_05248_),
    .A2(_05274_),
    .A3(_05275_),
    .B1(_05251_),
    .B2(net1070),
    .X(_00738_));
 sky130_fd_sc_hd__and3_1 _11270_ (.A(\genblk2[7].wave_shpr.div.b1[0] ),
    .B(_05182_),
    .C(_05183_),
    .X(_05276_));
 sky130_fd_sc_hd__nor2_1 _11271_ (.A(_05184_),
    .B(_05276_),
    .Y(_05277_));
 sky130_fd_sc_hd__mux2_1 _11272_ (.A0(\genblk2[7].wave_shpr.div.acc[1] ),
    .A1(_05277_),
    .S(_05222_),
    .X(_05278_));
 sky130_fd_sc_hd__a22o_1 _11273_ (.A1(net1013),
    .A2(_05246_),
    .B1(_05250_),
    .B2(_05278_),
    .X(_00739_));
 sky130_fd_sc_hd__clkbuf_4 _11274_ (.A(_05245_),
    .X(_05279_));
 sky130_fd_sc_hd__or2b_1 _11275_ (.A(_05186_),
    .B_N(_05181_),
    .X(_05280_));
 sky130_fd_sc_hd__xnor2_1 _11276_ (.A(_05185_),
    .B(_05280_),
    .Y(_05281_));
 sky130_fd_sc_hd__mux2_1 _11277_ (.A0(\genblk2[7].wave_shpr.div.acc[2] ),
    .A1(_05281_),
    .S(_05222_),
    .X(_05282_));
 sky130_fd_sc_hd__a22o_1 _11278_ (.A1(net992),
    .A2(_05279_),
    .B1(_05250_),
    .B2(_05282_),
    .X(_00740_));
 sky130_fd_sc_hd__clkbuf_4 _11279_ (.A(_05249_),
    .X(_05283_));
 sky130_fd_sc_hd__or2b_1 _11280_ (.A(_05188_),
    .B_N(_05180_),
    .X(_05284_));
 sky130_fd_sc_hd__xnor2_1 _11281_ (.A(_05187_),
    .B(_05284_),
    .Y(_05285_));
 sky130_fd_sc_hd__mux2_1 _11282_ (.A0(\genblk2[7].wave_shpr.div.acc[3] ),
    .A1(_05285_),
    .S(_05222_),
    .X(_05286_));
 sky130_fd_sc_hd__a22o_1 _11283_ (.A1(net877),
    .A2(_05279_),
    .B1(_05283_),
    .B2(_05286_),
    .X(_00741_));
 sky130_fd_sc_hd__xor2_1 _11284_ (.A(_05179_),
    .B(_05189_),
    .X(_05287_));
 sky130_fd_sc_hd__mux2_1 _11285_ (.A0(net877),
    .A1(_05287_),
    .S(_05222_),
    .X(_05288_));
 sky130_fd_sc_hd__a22o_1 _11286_ (.A1(net1030),
    .A2(_05279_),
    .B1(_05283_),
    .B2(_05288_),
    .X(_00742_));
 sky130_fd_sc_hd__or2b_1 _11287_ (.A(_05191_),
    .B_N(_05176_),
    .X(_05289_));
 sky130_fd_sc_hd__xnor2_1 _11288_ (.A(_05289_),
    .B(_05190_),
    .Y(_05290_));
 sky130_fd_sc_hd__mux2_1 _11289_ (.A0(\genblk2[7].wave_shpr.div.acc[5] ),
    .A1(_05290_),
    .S(_05222_),
    .X(_05291_));
 sky130_fd_sc_hd__a22o_1 _11290_ (.A1(net988),
    .A2(_05279_),
    .B1(_05283_),
    .B2(_05291_),
    .X(_00743_));
 sky130_fd_sc_hd__or2b_1 _11291_ (.A(_05193_),
    .B_N(_05175_),
    .X(_05292_));
 sky130_fd_sc_hd__xnor2_1 _11292_ (.A(_05192_),
    .B(_05292_),
    .Y(_05293_));
 sky130_fd_sc_hd__mux2_1 _11293_ (.A0(\genblk2[7].wave_shpr.div.acc[6] ),
    .A1(_05293_),
    .S(_05222_),
    .X(_05294_));
 sky130_fd_sc_hd__a22o_1 _11294_ (.A1(net893),
    .A2(_05279_),
    .B1(_05283_),
    .B2(_05294_),
    .X(_00744_));
 sky130_fd_sc_hd__or2b_1 _11295_ (.A(_05195_),
    .B_N(_05174_),
    .X(_05295_));
 sky130_fd_sc_hd__xnor2_1 _11296_ (.A(_05194_),
    .B(_05295_),
    .Y(_05296_));
 sky130_fd_sc_hd__mux2_1 _11297_ (.A0(net893),
    .A1(_05296_),
    .S(_05222_),
    .X(_05297_));
 sky130_fd_sc_hd__a22o_1 _11298_ (.A1(net1009),
    .A2(_05279_),
    .B1(_05283_),
    .B2(_05297_),
    .X(_00745_));
 sky130_fd_sc_hd__or2b_1 _11299_ (.A(_05197_),
    .B_N(_05173_),
    .X(_05298_));
 sky130_fd_sc_hd__xnor2_1 _11300_ (.A(_05196_),
    .B(_05298_),
    .Y(_05299_));
 sky130_fd_sc_hd__clkbuf_4 _11301_ (.A(_05221_),
    .X(_05300_));
 sky130_fd_sc_hd__mux2_1 _11302_ (.A0(\genblk2[7].wave_shpr.div.acc[8] ),
    .A1(_05299_),
    .S(_05300_),
    .X(_05301_));
 sky130_fd_sc_hd__a22o_1 _11303_ (.A1(net916),
    .A2(_05279_),
    .B1(_05283_),
    .B2(_05301_),
    .X(_00746_));
 sky130_fd_sc_hd__or2b_1 _11304_ (.A(_05199_),
    .B_N(_05172_),
    .X(_05302_));
 sky130_fd_sc_hd__xnor2_1 _11305_ (.A(_05198_),
    .B(_05302_),
    .Y(_05303_));
 sky130_fd_sc_hd__mux2_1 _11306_ (.A0(\genblk2[7].wave_shpr.div.acc[9] ),
    .A1(_05303_),
    .S(_05300_),
    .X(_05304_));
 sky130_fd_sc_hd__a22o_1 _11307_ (.A1(net797),
    .A2(_05279_),
    .B1(_05283_),
    .B2(_05304_),
    .X(_00747_));
 sky130_fd_sc_hd__or2b_1 _11308_ (.A(_05201_),
    .B_N(_05171_),
    .X(_05305_));
 sky130_fd_sc_hd__xnor2_1 _11309_ (.A(_05200_),
    .B(_05305_),
    .Y(_05306_));
 sky130_fd_sc_hd__mux2_1 _11310_ (.A0(\genblk2[7].wave_shpr.div.acc[10] ),
    .A1(_05306_),
    .S(_05300_),
    .X(_05307_));
 sky130_fd_sc_hd__a22o_1 _11311_ (.A1(net894),
    .A2(_05279_),
    .B1(_05283_),
    .B2(_05307_),
    .X(_00748_));
 sky130_fd_sc_hd__or2b_1 _11312_ (.A(_05203_),
    .B_N(_05170_),
    .X(_05308_));
 sky130_fd_sc_hd__xnor2_1 _11313_ (.A(_05202_),
    .B(_05308_),
    .Y(_05309_));
 sky130_fd_sc_hd__mux2_1 _11314_ (.A0(\genblk2[7].wave_shpr.div.acc[11] ),
    .A1(_05309_),
    .S(_05300_),
    .X(_05310_));
 sky130_fd_sc_hd__a22o_1 _11315_ (.A1(net852),
    .A2(_05279_),
    .B1(_05283_),
    .B2(_05310_),
    .X(_00749_));
 sky130_fd_sc_hd__clkbuf_4 _11316_ (.A(_05245_),
    .X(_05311_));
 sky130_fd_sc_hd__or2b_1 _11317_ (.A(_05205_),
    .B_N(_05169_),
    .X(_05312_));
 sky130_fd_sc_hd__xnor2_1 _11318_ (.A(_05204_),
    .B(_05312_),
    .Y(_05313_));
 sky130_fd_sc_hd__mux2_1 _11319_ (.A0(\genblk2[7].wave_shpr.div.acc[12] ),
    .A1(_05313_),
    .S(_05300_),
    .X(_05314_));
 sky130_fd_sc_hd__a22o_1 _11320_ (.A1(net808),
    .A2(_05311_),
    .B1(_05283_),
    .B2(_05314_),
    .X(_00750_));
 sky130_fd_sc_hd__clkbuf_4 _11321_ (.A(_05249_),
    .X(_05315_));
 sky130_fd_sc_hd__or2b_1 _11322_ (.A(_05207_),
    .B_N(_05168_),
    .X(_05316_));
 sky130_fd_sc_hd__xnor2_1 _11323_ (.A(_05206_),
    .B(_05316_),
    .Y(_05317_));
 sky130_fd_sc_hd__mux2_1 _11324_ (.A0(\genblk2[7].wave_shpr.div.acc[13] ),
    .A1(_05317_),
    .S(_05300_),
    .X(_05318_));
 sky130_fd_sc_hd__a22o_1 _11325_ (.A1(net805),
    .A2(_05311_),
    .B1(_05315_),
    .B2(_05318_),
    .X(_00751_));
 sky130_fd_sc_hd__or2b_1 _11326_ (.A(_05209_),
    .B_N(_05167_),
    .X(_05319_));
 sky130_fd_sc_hd__xnor2_1 _11327_ (.A(_05208_),
    .B(_05319_),
    .Y(_05320_));
 sky130_fd_sc_hd__mux2_1 _11328_ (.A0(\genblk2[7].wave_shpr.div.acc[14] ),
    .A1(_05320_),
    .S(_05300_),
    .X(_05321_));
 sky130_fd_sc_hd__a22o_1 _11329_ (.A1(net809),
    .A2(_05311_),
    .B1(_05315_),
    .B2(_05321_),
    .X(_00752_));
 sky130_fd_sc_hd__or2b_1 _11330_ (.A(_05211_),
    .B_N(_05166_),
    .X(_05322_));
 sky130_fd_sc_hd__xnor2_1 _11331_ (.A(_05210_),
    .B(_05322_),
    .Y(_05323_));
 sky130_fd_sc_hd__mux2_1 _11332_ (.A0(\genblk2[7].wave_shpr.div.acc[15] ),
    .A1(_05323_),
    .S(_05300_),
    .X(_05324_));
 sky130_fd_sc_hd__a22o_1 _11333_ (.A1(net1010),
    .A2(_05311_),
    .B1(_05315_),
    .B2(_05324_),
    .X(_00753_));
 sky130_fd_sc_hd__nor2_1 _11334_ (.A(_05213_),
    .B(_05165_),
    .Y(_05325_));
 sky130_fd_sc_hd__xnor2_1 _11335_ (.A(_05325_),
    .B(_05212_),
    .Y(_05326_));
 sky130_fd_sc_hd__mux2_1 _11336_ (.A0(\genblk2[7].wave_shpr.div.acc[16] ),
    .A1(_05326_),
    .S(_05300_),
    .X(_05327_));
 sky130_fd_sc_hd__a22o_1 _11337_ (.A1(net924),
    .A2(_05311_),
    .B1(_05315_),
    .B2(_05327_),
    .X(_00754_));
 sky130_fd_sc_hd__or2b_1 _11338_ (.A(_05215_),
    .B_N(_05164_),
    .X(_05328_));
 sky130_fd_sc_hd__xnor2_1 _11339_ (.A(_05214_),
    .B(_05328_),
    .Y(_05329_));
 sky130_fd_sc_hd__mux2_1 _11340_ (.A0(\genblk2[7].wave_shpr.div.acc[17] ),
    .A1(_05329_),
    .S(_05300_),
    .X(_05330_));
 sky130_fd_sc_hd__a22o_1 _11341_ (.A1(net628),
    .A2(_05311_),
    .B1(_05315_),
    .B2(_05330_),
    .X(_00755_));
 sky130_fd_sc_hd__or2_1 _11342_ (.A(_05217_),
    .B(_05273_),
    .X(_05331_));
 sky130_fd_sc_hd__o21ai_1 _11343_ (.A1(_05216_),
    .A2(_05273_),
    .B1(\genblk2[7].wave_shpr.div.acc[18] ),
    .Y(_05332_));
 sky130_fd_sc_hd__nand2_1 _11344_ (.A(_05331_),
    .B(_05332_),
    .Y(_05333_));
 sky130_fd_sc_hd__a22o_1 _11345_ (.A1(net1048),
    .A2(_05311_),
    .B1(_05315_),
    .B2(_05333_),
    .X(_00756_));
 sky130_fd_sc_hd__or2_1 _11346_ (.A(\genblk2[7].wave_shpr.div.acc[19] ),
    .B(_05331_),
    .X(_05334_));
 sky130_fd_sc_hd__a21bo_1 _11347_ (.A1(\genblk2[7].wave_shpr.div.acc[19] ),
    .A2(_05217_),
    .B1_N(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__a22o_1 _11348_ (.A1(net923),
    .A2(_05311_),
    .B1(_05315_),
    .B2(_05335_),
    .X(_00757_));
 sky130_fd_sc_hd__or2_1 _11349_ (.A(\genblk2[7].wave_shpr.div.acc[20] ),
    .B(_05334_),
    .X(_05336_));
 sky130_fd_sc_hd__nand2_1 _11350_ (.A(\genblk2[7].wave_shpr.div.acc[20] ),
    .B(_05334_),
    .Y(_05337_));
 sky130_fd_sc_hd__nand2_1 _11351_ (.A(_05336_),
    .B(_05337_),
    .Y(_05338_));
 sky130_fd_sc_hd__a22o_1 _11352_ (.A1(net679),
    .A2(_05311_),
    .B1(_05315_),
    .B2(_05338_),
    .X(_00758_));
 sky130_fd_sc_hd__a2bb2o_1 _11353_ (.A1_N(_05218_),
    .A2_N(_05273_),
    .B1(_05336_),
    .B2(\genblk2[7].wave_shpr.div.acc[21] ),
    .X(_05339_));
 sky130_fd_sc_hd__a22o_1 _11354_ (.A1(net706),
    .A2(_05311_),
    .B1(_05315_),
    .B2(_05339_),
    .X(_00759_));
 sky130_fd_sc_hd__and2b_1 _11355_ (.A_N(_05219_),
    .B(_05220_),
    .X(_05340_));
 sky130_fd_sc_hd__a21o_1 _11356_ (.A1(\genblk2[7].wave_shpr.div.acc[22] ),
    .A2(_05218_),
    .B1(_05340_),
    .X(_05341_));
 sky130_fd_sc_hd__a22o_1 _11357_ (.A1(net873),
    .A2(_05251_),
    .B1(_05315_),
    .B2(_05341_),
    .X(_00760_));
 sky130_fd_sc_hd__nor2_1 _11358_ (.A(\genblk2[7].wave_shpr.div.acc[23] ),
    .B(_05219_),
    .Y(_05342_));
 sky130_fd_sc_hd__and2_1 _11359_ (.A(\genblk2[7].wave_shpr.div.acc[23] ),
    .B(_05219_),
    .X(_05343_));
 sky130_fd_sc_hd__or2_1 _11360_ (.A(_05342_),
    .B(_05343_),
    .X(_05344_));
 sky130_fd_sc_hd__a32o_1 _11361_ (.A1(_05220_),
    .A2(_05248_),
    .A3(_05344_),
    .B1(_05251_),
    .B2(net1029),
    .X(_00761_));
 sky130_fd_sc_hd__inv_2 _11362_ (.A(\genblk2[7].wave_shpr.div.acc[24] ),
    .Y(_05345_));
 sky130_fd_sc_hd__or3b_1 _11363_ (.A(\genblk2[7].wave_shpr.div.acc[24] ),
    .B(_05273_),
    .C_N(_05342_),
    .X(_05346_));
 sky130_fd_sc_hd__o21ai_1 _11364_ (.A1(_05345_),
    .A2(_05342_),
    .B1(_05346_),
    .Y(_05347_));
 sky130_fd_sc_hd__a22o_1 _11365_ (.A1(net1053),
    .A2(_05251_),
    .B1(_05248_),
    .B2(_05347_),
    .X(_00762_));
 sky130_fd_sc_hd__xnor2_1 _11366_ (.A(\genblk2[7].wave_shpr.div.acc[25] ),
    .B(_05346_),
    .Y(_05348_));
 sky130_fd_sc_hd__a22o_1 _11367_ (.A1(net381),
    .A2(_05251_),
    .B1(_05248_),
    .B2(_05348_),
    .X(_00763_));
 sky130_fd_sc_hd__mux2_1 _11368_ (.A0(_05249_),
    .A1(_05245_),
    .S(\genblk2[7].wave_shpr.div.i[0] ),
    .X(_05349_));
 sky130_fd_sc_hd__clkbuf_1 _11369_ (.A(_05349_),
    .X(_00764_));
 sky130_fd_sc_hd__or2_1 _11370_ (.A(\genblk2[7].wave_shpr.div.i[1] ),
    .B(\genblk2[7].wave_shpr.div.i[0] ),
    .X(_05350_));
 sky130_fd_sc_hd__nand2_1 _11371_ (.A(\genblk2[7].wave_shpr.div.i[1] ),
    .B(\genblk2[7].wave_shpr.div.i[0] ),
    .Y(_05351_));
 sky130_fd_sc_hd__a32o_1 _11372_ (.A1(_05248_),
    .A2(_05350_),
    .A3(_05351_),
    .B1(_05251_),
    .B2(net1113),
    .X(_00765_));
 sky130_fd_sc_hd__a21o_1 _11373_ (.A1(\genblk2[7].wave_shpr.div.i[1] ),
    .A2(\genblk2[7].wave_shpr.div.i[0] ),
    .B1(\genblk2[7].wave_shpr.div.i[2] ),
    .X(_05352_));
 sky130_fd_sc_hd__and3_1 _11374_ (.A(\genblk2[7].wave_shpr.div.i[1] ),
    .B(\genblk2[7].wave_shpr.div.i[0] ),
    .C(\genblk2[7].wave_shpr.div.i[2] ),
    .X(_05353_));
 sky130_fd_sc_hd__inv_2 _11375_ (.A(_05353_),
    .Y(_05354_));
 sky130_fd_sc_hd__a32o_1 _11376_ (.A1(_05248_),
    .A2(_05352_),
    .A3(_05354_),
    .B1(_05251_),
    .B2(net801),
    .X(_00766_));
 sky130_fd_sc_hd__a21oi_1 _11377_ (.A1(_00018_),
    .A2(_05353_),
    .B1(net1181),
    .Y(_05355_));
 sky130_fd_sc_hd__and3_1 _11378_ (.A(\genblk2[7].wave_shpr.div.i[3] ),
    .B(_02192_),
    .C(_05353_),
    .X(_05356_));
 sky130_fd_sc_hd__nor3_1 _11379_ (.A(_03690_),
    .B(_05355_),
    .C(_05356_),
    .Y(_00767_));
 sky130_fd_sc_hd__o21ai_1 _11380_ (.A1(net328),
    .A2(_05356_),
    .B1(_03855_),
    .Y(_05357_));
 sky130_fd_sc_hd__a21oi_1 _11381_ (.A1(net328),
    .A2(_05356_),
    .B1(_05357_),
    .Y(_00768_));
 sky130_fd_sc_hd__or2b_1 _11382_ (.A(\genblk2[8].wave_shpr.div.acc[17] ),
    .B_N(\genblk2[8].wave_shpr.div.b1[17] ),
    .X(_05358_));
 sky130_fd_sc_hd__or2_1 _11383_ (.A(_05243_),
    .B(\genblk2[8].wave_shpr.div.acc[16] ),
    .X(_05359_));
 sky130_fd_sc_hd__or2b_1 _11384_ (.A(\genblk2[8].wave_shpr.div.acc[15] ),
    .B_N(\genblk2[8].wave_shpr.div.b1[15] ),
    .X(_05360_));
 sky130_fd_sc_hd__or2b_1 _11385_ (.A(\genblk2[8].wave_shpr.div.acc[14] ),
    .B_N(\genblk2[8].wave_shpr.div.b1[14] ),
    .X(_05361_));
 sky130_fd_sc_hd__or2b_1 _11386_ (.A(\genblk2[8].wave_shpr.div.acc[13] ),
    .B_N(\genblk2[8].wave_shpr.div.b1[13] ),
    .X(_05362_));
 sky130_fd_sc_hd__or2b_1 _11387_ (.A(\genblk2[8].wave_shpr.div.acc[12] ),
    .B_N(\genblk2[8].wave_shpr.div.b1[12] ),
    .X(_05363_));
 sky130_fd_sc_hd__or2b_1 _11388_ (.A(\genblk2[8].wave_shpr.div.acc[11] ),
    .B_N(\genblk2[8].wave_shpr.div.b1[11] ),
    .X(_05364_));
 sky130_fd_sc_hd__or2b_1 _11389_ (.A(\genblk2[8].wave_shpr.div.acc[10] ),
    .B_N(\genblk2[8].wave_shpr.div.b1[10] ),
    .X(_05365_));
 sky130_fd_sc_hd__or2b_1 _11390_ (.A(\genblk2[8].wave_shpr.div.acc[9] ),
    .B_N(\genblk2[8].wave_shpr.div.b1[9] ),
    .X(_05366_));
 sky130_fd_sc_hd__or2b_1 _11391_ (.A(\genblk2[8].wave_shpr.div.acc[8] ),
    .B_N(\genblk2[8].wave_shpr.div.b1[8] ),
    .X(_05367_));
 sky130_fd_sc_hd__or2b_1 _11392_ (.A(\genblk2[8].wave_shpr.div.acc[7] ),
    .B_N(\genblk2[8].wave_shpr.div.b1[7] ),
    .X(_05368_));
 sky130_fd_sc_hd__or2b_1 _11393_ (.A(\genblk2[8].wave_shpr.div.acc[6] ),
    .B_N(\genblk2[8].wave_shpr.div.b1[6] ),
    .X(_05369_));
 sky130_fd_sc_hd__or2b_1 _11394_ (.A(\genblk2[8].wave_shpr.div.acc[5] ),
    .B_N(\genblk2[8].wave_shpr.div.b1[5] ),
    .X(_05370_));
 sky130_fd_sc_hd__or2b_1 _11395_ (.A(\genblk2[8].wave_shpr.div.acc[4] ),
    .B_N(\genblk2[8].wave_shpr.div.b1[4] ),
    .X(_05371_));
 sky130_fd_sc_hd__or2b_1 _11396_ (.A(\genblk2[8].wave_shpr.div.acc[3] ),
    .B_N(\genblk2[8].wave_shpr.div.b1[3] ),
    .X(_05372_));
 sky130_fd_sc_hd__or2b_1 _11397_ (.A(\genblk2[8].wave_shpr.div.acc[2] ),
    .B_N(\genblk2[8].wave_shpr.div.b1[2] ),
    .X(_05373_));
 sky130_fd_sc_hd__xor2_1 _11398_ (.A(\genblk2[8].wave_shpr.div.acc[1] ),
    .B(\genblk2[8].wave_shpr.div.b1[1] ),
    .X(_05374_));
 sky130_fd_sc_hd__and2b_1 _11399_ (.A_N(\genblk2[8].wave_shpr.div.acc[0] ),
    .B(\genblk2[8].wave_shpr.div.b1[0] ),
    .X(_05375_));
 sky130_fd_sc_hd__or2b_1 _11400_ (.A(\genblk2[8].wave_shpr.div.b1[1] ),
    .B_N(\genblk2[8].wave_shpr.div.acc[1] ),
    .X(_05376_));
 sky130_fd_sc_hd__o21ai_1 _11401_ (.A1(_05374_),
    .A2(_05375_),
    .B1(_05376_),
    .Y(_05377_));
 sky130_fd_sc_hd__and2b_1 _11402_ (.A_N(\genblk2[8].wave_shpr.div.b1[2] ),
    .B(\genblk2[8].wave_shpr.div.acc[2] ),
    .X(_05378_));
 sky130_fd_sc_hd__a21o_1 _11403_ (.A1(_05373_),
    .A2(_05377_),
    .B1(_05378_),
    .X(_05379_));
 sky130_fd_sc_hd__and2b_1 _11404_ (.A_N(\genblk2[8].wave_shpr.div.b1[3] ),
    .B(\genblk2[8].wave_shpr.div.acc[3] ),
    .X(_05380_));
 sky130_fd_sc_hd__a21o_1 _11405_ (.A1(_05372_),
    .A2(_05379_),
    .B1(_05380_),
    .X(_05381_));
 sky130_fd_sc_hd__and2b_1 _11406_ (.A_N(\genblk2[8].wave_shpr.div.b1[4] ),
    .B(\genblk2[8].wave_shpr.div.acc[4] ),
    .X(_05382_));
 sky130_fd_sc_hd__a21o_1 _11407_ (.A1(_05371_),
    .A2(_05381_),
    .B1(_05382_),
    .X(_05383_));
 sky130_fd_sc_hd__and2b_1 _11408_ (.A_N(\genblk2[8].wave_shpr.div.b1[5] ),
    .B(\genblk2[8].wave_shpr.div.acc[5] ),
    .X(_05384_));
 sky130_fd_sc_hd__a21o_1 _11409_ (.A1(_05370_),
    .A2(_05383_),
    .B1(_05384_),
    .X(_05385_));
 sky130_fd_sc_hd__and2b_1 _11410_ (.A_N(\genblk2[8].wave_shpr.div.b1[6] ),
    .B(\genblk2[8].wave_shpr.div.acc[6] ),
    .X(_05386_));
 sky130_fd_sc_hd__a21o_1 _11411_ (.A1(_05369_),
    .A2(_05385_),
    .B1(_05386_),
    .X(_05387_));
 sky130_fd_sc_hd__and2b_1 _11412_ (.A_N(\genblk2[8].wave_shpr.div.b1[7] ),
    .B(\genblk2[8].wave_shpr.div.acc[7] ),
    .X(_05388_));
 sky130_fd_sc_hd__a21o_1 _11413_ (.A1(_05368_),
    .A2(_05387_),
    .B1(_05388_),
    .X(_05389_));
 sky130_fd_sc_hd__and2b_1 _11414_ (.A_N(\genblk2[8].wave_shpr.div.b1[8] ),
    .B(\genblk2[8].wave_shpr.div.acc[8] ),
    .X(_05390_));
 sky130_fd_sc_hd__a21o_1 _11415_ (.A1(_05367_),
    .A2(_05389_),
    .B1(_05390_),
    .X(_05391_));
 sky130_fd_sc_hd__and2b_1 _11416_ (.A_N(\genblk2[8].wave_shpr.div.b1[9] ),
    .B(\genblk2[8].wave_shpr.div.acc[9] ),
    .X(_05392_));
 sky130_fd_sc_hd__a21o_1 _11417_ (.A1(_05366_),
    .A2(_05391_),
    .B1(_05392_),
    .X(_05393_));
 sky130_fd_sc_hd__and2b_1 _11418_ (.A_N(\genblk2[8].wave_shpr.div.b1[10] ),
    .B(\genblk2[8].wave_shpr.div.acc[10] ),
    .X(_05394_));
 sky130_fd_sc_hd__a21o_1 _11419_ (.A1(_05365_),
    .A2(_05393_),
    .B1(_05394_),
    .X(_05395_));
 sky130_fd_sc_hd__and2b_1 _11420_ (.A_N(\genblk2[8].wave_shpr.div.b1[11] ),
    .B(\genblk2[8].wave_shpr.div.acc[11] ),
    .X(_05396_));
 sky130_fd_sc_hd__a21o_1 _11421_ (.A1(_05364_),
    .A2(_05395_),
    .B1(_05396_),
    .X(_05397_));
 sky130_fd_sc_hd__and2b_1 _11422_ (.A_N(\genblk2[8].wave_shpr.div.b1[12] ),
    .B(\genblk2[8].wave_shpr.div.acc[12] ),
    .X(_05398_));
 sky130_fd_sc_hd__a21o_1 _11423_ (.A1(_05363_),
    .A2(_05397_),
    .B1(_05398_),
    .X(_05399_));
 sky130_fd_sc_hd__and2b_1 _11424_ (.A_N(\genblk2[8].wave_shpr.div.b1[13] ),
    .B(\genblk2[8].wave_shpr.div.acc[13] ),
    .X(_05400_));
 sky130_fd_sc_hd__a21o_1 _11425_ (.A1(_05362_),
    .A2(_05399_),
    .B1(_05400_),
    .X(_05401_));
 sky130_fd_sc_hd__and2b_1 _11426_ (.A_N(\genblk2[8].wave_shpr.div.b1[14] ),
    .B(\genblk2[8].wave_shpr.div.acc[14] ),
    .X(_05402_));
 sky130_fd_sc_hd__a21o_1 _11427_ (.A1(_05361_),
    .A2(_05401_),
    .B1(_05402_),
    .X(_05403_));
 sky130_fd_sc_hd__and2b_1 _11428_ (.A_N(\genblk2[8].wave_shpr.div.b1[15] ),
    .B(\genblk2[8].wave_shpr.div.acc[15] ),
    .X(_05404_));
 sky130_fd_sc_hd__a21o_1 _11429_ (.A1(_05360_),
    .A2(_05403_),
    .B1(_05404_),
    .X(_05405_));
 sky130_fd_sc_hd__and2_1 _11430_ (.A(_05243_),
    .B(\genblk2[8].wave_shpr.div.acc[16] ),
    .X(_05406_));
 sky130_fd_sc_hd__a21o_1 _11431_ (.A1(_05359_),
    .A2(_05405_),
    .B1(_05406_),
    .X(_05407_));
 sky130_fd_sc_hd__and2b_1 _11432_ (.A_N(\genblk2[8].wave_shpr.div.b1[17] ),
    .B(\genblk2[8].wave_shpr.div.acc[17] ),
    .X(_05408_));
 sky130_fd_sc_hd__a21o_1 _11433_ (.A1(_05358_),
    .A2(_05407_),
    .B1(_05408_),
    .X(_05409_));
 sky130_fd_sc_hd__or4_1 _11434_ (.A(\genblk2[8].wave_shpr.div.acc[20] ),
    .B(\genblk2[8].wave_shpr.div.acc[18] ),
    .C(\genblk2[8].wave_shpr.div.acc[19] ),
    .D(_05409_),
    .X(_05410_));
 sky130_fd_sc_hd__or2_1 _11435_ (.A(\genblk2[8].wave_shpr.div.acc[21] ),
    .B(_05410_),
    .X(_05411_));
 sky130_fd_sc_hd__or2_1 _11436_ (.A(\genblk2[8].wave_shpr.div.acc[22] ),
    .B(_05411_),
    .X(_05412_));
 sky130_fd_sc_hd__or2_1 _11437_ (.A(\genblk2[8].wave_shpr.div.acc[23] ),
    .B(_05412_),
    .X(_05413_));
 sky130_fd_sc_hd__or2_1 _11438_ (.A(\genblk2[8].wave_shpr.div.acc[24] ),
    .B(_05413_),
    .X(_05414_));
 sky130_fd_sc_hd__or3_1 _11439_ (.A(\genblk2[8].wave_shpr.div.acc[25] ),
    .B(\genblk2[8].wave_shpr.div.acc[26] ),
    .C(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__buf_2 _11440_ (.A(_05415_),
    .X(_05416_));
 sky130_fd_sc_hd__clkbuf_4 _11441_ (.A(_05416_),
    .X(_05417_));
 sky130_fd_sc_hd__mux2_1 _11442_ (.A0(\genblk2[8].wave_shpr.div.fin_quo[0] ),
    .A1(_05417_),
    .S(_00021_),
    .X(_05418_));
 sky130_fd_sc_hd__clkbuf_1 _11443_ (.A(_05418_),
    .X(_00769_));
 sky130_fd_sc_hd__mux2_1 _11444_ (.A0(\genblk2[8].wave_shpr.div.fin_quo[1] ),
    .A1(net1331),
    .S(_00021_),
    .X(_05419_));
 sky130_fd_sc_hd__clkbuf_1 _11445_ (.A(_05419_),
    .X(_00770_));
 sky130_fd_sc_hd__mux2_1 _11446_ (.A0(\genblk2[8].wave_shpr.div.fin_quo[2] ),
    .A1(\genblk2[8].wave_shpr.div.quo[1] ),
    .S(_00021_),
    .X(_05420_));
 sky130_fd_sc_hd__clkbuf_1 _11447_ (.A(_05420_),
    .X(_00771_));
 sky130_fd_sc_hd__mux2_1 _11448_ (.A0(\genblk2[8].wave_shpr.div.fin_quo[3] ),
    .A1(net1337),
    .S(_00021_),
    .X(_05421_));
 sky130_fd_sc_hd__clkbuf_1 _11449_ (.A(_05421_),
    .X(_00772_));
 sky130_fd_sc_hd__mux2_1 _11450_ (.A0(\genblk2[8].wave_shpr.div.fin_quo[4] ),
    .A1(net1321),
    .S(_00021_),
    .X(_05422_));
 sky130_fd_sc_hd__clkbuf_1 _11451_ (.A(_05422_),
    .X(_00773_));
 sky130_fd_sc_hd__mux2_1 _11452_ (.A0(\genblk2[8].wave_shpr.div.fin_quo[5] ),
    .A1(\genblk2[8].wave_shpr.div.quo[4] ),
    .S(_00021_),
    .X(_05423_));
 sky130_fd_sc_hd__clkbuf_1 _11453_ (.A(_05423_),
    .X(_00774_));
 sky130_fd_sc_hd__mux2_1 _11454_ (.A0(\genblk2[8].wave_shpr.div.fin_quo[6] ),
    .A1(net1325),
    .S(_00021_),
    .X(_05424_));
 sky130_fd_sc_hd__clkbuf_1 _11455_ (.A(_05424_),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _11456_ (.A0(\genblk2[8].wave_shpr.div.fin_quo[7] ),
    .A1(net1335),
    .S(_00021_),
    .X(_05425_));
 sky130_fd_sc_hd__clkbuf_1 _11457_ (.A(_05425_),
    .X(_00776_));
 sky130_fd_sc_hd__mux2_1 _11458_ (.A0(\genblk2[9].wave_shpr.div.b1[0] ),
    .A1(_02064_),
    .S(_05237_),
    .X(_05426_));
 sky130_fd_sc_hd__clkbuf_1 _11459_ (.A(_05426_),
    .X(_00777_));
 sky130_fd_sc_hd__mux2_1 _11460_ (.A0(\genblk2[9].wave_shpr.div.b1[1] ),
    .A1(_01819_),
    .S(_05237_),
    .X(_05427_));
 sky130_fd_sc_hd__clkbuf_1 _11461_ (.A(_05427_),
    .X(_00778_));
 sky130_fd_sc_hd__mux2_1 _11462_ (.A0(net1294),
    .A1(_01797_),
    .S(_05237_),
    .X(_05428_));
 sky130_fd_sc_hd__clkbuf_1 _11463_ (.A(_05428_),
    .X(_00779_));
 sky130_fd_sc_hd__mux2_1 _11464_ (.A0(net1230),
    .A1(net34),
    .S(_05237_),
    .X(_05429_));
 sky130_fd_sc_hd__clkbuf_1 _11465_ (.A(_05429_),
    .X(_00780_));
 sky130_fd_sc_hd__mux2_1 _11466_ (.A0(net1268),
    .A1(_02433_),
    .S(_05237_),
    .X(_05430_));
 sky130_fd_sc_hd__clkbuf_1 _11467_ (.A(_05430_),
    .X(_00781_));
 sky130_fd_sc_hd__mux2_1 _11468_ (.A0(net1208),
    .A1(_01811_),
    .S(_05237_),
    .X(_05431_));
 sky130_fd_sc_hd__clkbuf_1 _11469_ (.A(_05431_),
    .X(_00782_));
 sky130_fd_sc_hd__mux2_1 _11470_ (.A0(net1187),
    .A1(_01946_),
    .S(_05237_),
    .X(_05432_));
 sky130_fd_sc_hd__clkbuf_1 _11471_ (.A(_05432_),
    .X(_00783_));
 sky130_fd_sc_hd__clkbuf_4 _11472_ (.A(_03707_),
    .X(_05433_));
 sky130_fd_sc_hd__mux2_1 _11473_ (.A0(\genblk2[9].wave_shpr.div.b1[7] ),
    .A1(_04230_),
    .S(_05433_),
    .X(_05434_));
 sky130_fd_sc_hd__clkbuf_1 _11474_ (.A(_05434_),
    .X(_00784_));
 sky130_fd_sc_hd__mux2_1 _11475_ (.A0(net1236),
    .A1(net34),
    .S(_05433_),
    .X(_05435_));
 sky130_fd_sc_hd__clkbuf_1 _11476_ (.A(_05435_),
    .X(_00785_));
 sky130_fd_sc_hd__a21o_1 _11477_ (.A1(_03704_),
    .A2(net1042),
    .B1(_04233_),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _11478_ (.A0(net1231),
    .A1(_01227_),
    .S(_05433_),
    .X(_05436_));
 sky130_fd_sc_hd__clkbuf_1 _11479_ (.A(_05436_),
    .X(_00787_));
 sky130_fd_sc_hd__mux2_1 _11480_ (.A0(\genblk2[9].wave_shpr.div.b1[11] ),
    .A1(_01732_),
    .S(_05433_),
    .X(_05437_));
 sky130_fd_sc_hd__clkbuf_1 _11481_ (.A(_05437_),
    .X(_00788_));
 sky130_fd_sc_hd__mux2_1 _11482_ (.A0(\genblk2[9].wave_shpr.div.b1[12] ),
    .A1(_02656_),
    .S(_05433_),
    .X(_05438_));
 sky130_fd_sc_hd__clkbuf_1 _11483_ (.A(_05438_),
    .X(_00789_));
 sky130_fd_sc_hd__a2bb2o_1 _11484_ (.A1_N(_03727_),
    .A2_N(_01490_),
    .B1(_03687_),
    .B2(net478),
    .X(_00790_));
 sky130_fd_sc_hd__a21bo_1 _11485_ (.A1(_03831_),
    .A2(net374),
    .B1_N(_03728_),
    .X(_00791_));
 sky130_fd_sc_hd__a21bo_1 _11486_ (.A1(_03831_),
    .A2(net390),
    .B1_N(_03717_),
    .X(_00792_));
 sky130_fd_sc_hd__inv_2 _11487_ (.A(net713),
    .Y(_05439_));
 sky130_fd_sc_hd__o21ai_1 _11488_ (.A1(_03726_),
    .A2(_05439_),
    .B1(_03736_),
    .Y(_00793_));
 sky130_fd_sc_hd__and2_1 _11489_ (.A(_02171_),
    .B(net1239),
    .X(_05440_));
 sky130_fd_sc_hd__clkbuf_1 _11490_ (.A(_05440_),
    .X(_00794_));
 sky130_fd_sc_hd__clkbuf_4 _11491_ (.A(_02198_),
    .X(_05441_));
 sky130_fd_sc_hd__clkbuf_4 _11492_ (.A(_05441_),
    .X(_05442_));
 sky130_fd_sc_hd__and3_1 _11493_ (.A(_02152_),
    .B(\genblk2[8].wave_shpr.div.busy ),
    .C(_02196_),
    .X(_05443_));
 sky130_fd_sc_hd__buf_2 _11494_ (.A(_05443_),
    .X(_05444_));
 sky130_fd_sc_hd__clkbuf_4 _11495_ (.A(_05444_),
    .X(_05445_));
 sky130_fd_sc_hd__a22o_1 _11496_ (.A1(net743),
    .A2(_05442_),
    .B1(_05417_),
    .B2(_05445_),
    .X(_00795_));
 sky130_fd_sc_hd__clkbuf_4 _11497_ (.A(_05444_),
    .X(_05446_));
 sky130_fd_sc_hd__a22o_1 _11498_ (.A1(\genblk2[8].wave_shpr.div.quo[1] ),
    .A2(_05442_),
    .B1(_05446_),
    .B2(net743),
    .X(_00796_));
 sky130_fd_sc_hd__a22o_1 _11499_ (.A1(net709),
    .A2(_05442_),
    .B1(_05446_),
    .B2(net871),
    .X(_00797_));
 sky130_fd_sc_hd__a22o_1 _11500_ (.A1(net346),
    .A2(_05442_),
    .B1(_05446_),
    .B2(net709),
    .X(_00798_));
 sky130_fd_sc_hd__a22o_1 _11501_ (.A1(\genblk2[8].wave_shpr.div.quo[4] ),
    .A2(_05442_),
    .B1(_05446_),
    .B2(net346),
    .X(_00799_));
 sky130_fd_sc_hd__a22o_1 _11502_ (.A1(net751),
    .A2(_05442_),
    .B1(_05446_),
    .B2(net795),
    .X(_00800_));
 sky130_fd_sc_hd__a22o_1 _11503_ (.A1(net676),
    .A2(_05442_),
    .B1(_05446_),
    .B2(net751),
    .X(_00801_));
 sky130_fd_sc_hd__a22o_1 _11504_ (.A1(net404),
    .A2(_05442_),
    .B1(_05446_),
    .B2(net676),
    .X(_00802_));
 sky130_fd_sc_hd__clkbuf_4 _11505_ (.A(_05441_),
    .X(_05447_));
 sky130_fd_sc_hd__a22o_1 _11506_ (.A1(\genblk2[8].wave_shpr.div.quo[8] ),
    .A2(_05447_),
    .B1(_05446_),
    .B2(net404),
    .X(_00803_));
 sky130_fd_sc_hd__clkbuf_4 _11507_ (.A(_05441_),
    .X(_05448_));
 sky130_fd_sc_hd__clkbuf_4 _11508_ (.A(_05444_),
    .X(_05449_));
 sky130_fd_sc_hd__clkbuf_2 _11509_ (.A(_04268_),
    .X(_05450_));
 sky130_fd_sc_hd__and2_1 _11510_ (.A(_05450_),
    .B(\genblk1[8].osc.clkdiv_C.cnt[0] ),
    .X(_05451_));
 sky130_fd_sc_hd__a221o_1 _11511_ (.A1(net329),
    .A2(_05448_),
    .B1(_05449_),
    .B2(net450),
    .C1(_05451_),
    .X(_00804_));
 sky130_fd_sc_hd__and2_1 _11512_ (.A(_05450_),
    .B(\genblk1[8].osc.clkdiv_C.cnt[1] ),
    .X(_05452_));
 sky130_fd_sc_hd__a221o_1 _11513_ (.A1(\genblk2[8].wave_shpr.div.quo[10] ),
    .A2(_05448_),
    .B1(_05449_),
    .B2(net329),
    .C1(_05452_),
    .X(_00805_));
 sky130_fd_sc_hd__nor2_1 _11514_ (.A(_04676_),
    .B(_01879_),
    .Y(_05453_));
 sky130_fd_sc_hd__a221o_1 _11515_ (.A1(\genblk2[8].wave_shpr.div.quo[11] ),
    .A2(_05448_),
    .B1(_05449_),
    .B2(net469),
    .C1(_05453_),
    .X(_00806_));
 sky130_fd_sc_hd__buf_2 _11516_ (.A(_05441_),
    .X(_05454_));
 sky130_fd_sc_hd__and2_1 _11517_ (.A(_05450_),
    .B(\genblk1[8].osc.clkdiv_C.cnt[3] ),
    .X(_05455_));
 sky130_fd_sc_hd__a221o_1 _11518_ (.A1(net482),
    .A2(_05454_),
    .B1(_05449_),
    .B2(net506),
    .C1(_05455_),
    .X(_00807_));
 sky130_fd_sc_hd__and2_1 _11519_ (.A(_05450_),
    .B(\genblk1[8].osc.clkdiv_C.cnt[4] ),
    .X(_05456_));
 sky130_fd_sc_hd__a221o_1 _11520_ (.A1(net312),
    .A2(_05454_),
    .B1(_05449_),
    .B2(net482),
    .C1(_05456_),
    .X(_00808_));
 sky130_fd_sc_hd__and2_1 _11521_ (.A(_05450_),
    .B(\genblk1[8].osc.clkdiv_C.cnt[5] ),
    .X(_05457_));
 sky130_fd_sc_hd__a221o_1 _11522_ (.A1(net237),
    .A2(_05454_),
    .B1(_05449_),
    .B2(net312),
    .C1(_05457_),
    .X(_00809_));
 sky130_fd_sc_hd__clkbuf_4 _11523_ (.A(_05444_),
    .X(_05458_));
 sky130_fd_sc_hd__and2_1 _11524_ (.A(_05450_),
    .B(\genblk1[8].osc.clkdiv_C.cnt[6] ),
    .X(_05459_));
 sky130_fd_sc_hd__a221o_1 _11525_ (.A1(\genblk2[8].wave_shpr.div.quo[15] ),
    .A2(_05454_),
    .B1(_05458_),
    .B2(net237),
    .C1(_05459_),
    .X(_00810_));
 sky130_fd_sc_hd__and2_1 _11526_ (.A(_05450_),
    .B(\genblk1[8].osc.clkdiv_C.cnt[7] ),
    .X(_05460_));
 sky130_fd_sc_hd__a221o_1 _11527_ (.A1(net502),
    .A2(_05454_),
    .B1(_05458_),
    .B2(net611),
    .C1(_05460_),
    .X(_00811_));
 sky130_fd_sc_hd__and2_1 _11528_ (.A(_05450_),
    .B(\genblk1[8].osc.clkdiv_C.cnt[8] ),
    .X(_05461_));
 sky130_fd_sc_hd__a221o_1 _11529_ (.A1(net263),
    .A2(_05454_),
    .B1(_05458_),
    .B2(net502),
    .C1(_05461_),
    .X(_00812_));
 sky130_fd_sc_hd__and2_1 _11530_ (.A(_05450_),
    .B(\genblk1[8].osc.clkdiv_C.cnt[9] ),
    .X(_05462_));
 sky130_fd_sc_hd__a221o_1 _11531_ (.A1(\genblk2[8].wave_shpr.div.quo[18] ),
    .A2(_05454_),
    .B1(_05458_),
    .B2(net263),
    .C1(_05462_),
    .X(_00813_));
 sky130_fd_sc_hd__and2_1 _11532_ (.A(_05450_),
    .B(\genblk1[8].osc.clkdiv_C.cnt[10] ),
    .X(_05463_));
 sky130_fd_sc_hd__a221o_1 _11533_ (.A1(\genblk2[8].wave_shpr.div.quo[19] ),
    .A2(_05454_),
    .B1(_05458_),
    .B2(net617),
    .C1(_05463_),
    .X(_00814_));
 sky130_fd_sc_hd__buf_2 _11534_ (.A(_04268_),
    .X(_05464_));
 sky130_fd_sc_hd__and2_1 _11535_ (.A(_05464_),
    .B(\genblk1[8].osc.clkdiv_C.cnt[11] ),
    .X(_05465_));
 sky130_fd_sc_hd__a221o_1 _11536_ (.A1(net660),
    .A2(_05454_),
    .B1(_05458_),
    .B2(net677),
    .C1(_05465_),
    .X(_00815_));
 sky130_fd_sc_hd__and2_1 _11537_ (.A(_05464_),
    .B(\genblk1[8].osc.clkdiv_C.cnt[12] ),
    .X(_05466_));
 sky130_fd_sc_hd__a221o_1 _11538_ (.A1(net575),
    .A2(_05454_),
    .B1(_05458_),
    .B2(net660),
    .C1(_05466_),
    .X(_00816_));
 sky130_fd_sc_hd__and2_1 _11539_ (.A(_05464_),
    .B(\genblk1[8].osc.clkdiv_C.cnt[13] ),
    .X(_05467_));
 sky130_fd_sc_hd__a221o_1 _11540_ (.A1(net229),
    .A2(_05441_),
    .B1(_05458_),
    .B2(net575),
    .C1(_05467_),
    .X(_00817_));
 sky130_fd_sc_hd__and2_1 _11541_ (.A(_05464_),
    .B(\genblk1[8].osc.clkdiv_C.cnt[14] ),
    .X(_05468_));
 sky130_fd_sc_hd__a221o_1 _11542_ (.A1(\genblk2[8].wave_shpr.div.quo[23] ),
    .A2(_05441_),
    .B1(_05458_),
    .B2(net229),
    .C1(_05468_),
    .X(_00818_));
 sky130_fd_sc_hd__and2_1 _11543_ (.A(_05464_),
    .B(\genblk1[8].osc.clkdiv_C.cnt[15] ),
    .X(_05469_));
 sky130_fd_sc_hd__a221o_1 _11544_ (.A1(net445),
    .A2(_05441_),
    .B1(_05458_),
    .B2(net505),
    .C1(_05469_),
    .X(_00819_));
 sky130_fd_sc_hd__and2_1 _11545_ (.A(_05464_),
    .B(\genblk1[8].osc.clkdiv_C.cnt[16] ),
    .X(_05470_));
 sky130_fd_sc_hd__a221o_1 _11546_ (.A1(net274),
    .A2(_05441_),
    .B1(_05444_),
    .B2(net445),
    .C1(_05470_),
    .X(_00820_));
 sky130_fd_sc_hd__inv_2 _11547_ (.A(_05444_),
    .Y(_05471_));
 sky130_fd_sc_hd__or2_1 _11548_ (.A(_03719_),
    .B(\genblk1[8].osc.clkdiv_C.cnt[17] ),
    .X(_05472_));
 sky130_fd_sc_hd__o221a_1 _11549_ (.A1(\genblk2[8].wave_shpr.div.acc[0] ),
    .A2(_00020_),
    .B1(_05471_),
    .B2(net274),
    .C1(_05472_),
    .X(_00821_));
 sky130_fd_sc_hd__a21oi_1 _11550_ (.A1(\genblk2[8].wave_shpr.div.b1[0] ),
    .A2(_05417_),
    .B1(\genblk2[8].wave_shpr.div.acc[0] ),
    .Y(_05473_));
 sky130_fd_sc_hd__a31o_1 _11551_ (.A1(\genblk2[8].wave_shpr.div.b1[0] ),
    .A2(\genblk2[8].wave_shpr.div.acc[0] ),
    .A3(_05417_),
    .B1(_05471_),
    .X(_05474_));
 sky130_fd_sc_hd__a2bb2o_1 _11552_ (.A1_N(_05473_),
    .A2_N(_05474_),
    .B1(net1116),
    .B2(_05442_),
    .X(_00822_));
 sky130_fd_sc_hd__or2_1 _11553_ (.A(\genblk2[8].wave_shpr.div.acc[1] ),
    .B(_05416_),
    .X(_05475_));
 sky130_fd_sc_hd__xnor2_1 _11554_ (.A(_05374_),
    .B(_05375_),
    .Y(_05476_));
 sky130_fd_sc_hd__nand2_1 _11555_ (.A(_05417_),
    .B(_05476_),
    .Y(_05477_));
 sky130_fd_sc_hd__a32o_1 _11556_ (.A1(_05449_),
    .A2(_05475_),
    .A3(_05477_),
    .B1(_05448_),
    .B2(net699),
    .X(_00823_));
 sky130_fd_sc_hd__or2b_1 _11557_ (.A(_05378_),
    .B_N(_05373_),
    .X(_05478_));
 sky130_fd_sc_hd__xnor2_1 _11558_ (.A(_05377_),
    .B(_05478_),
    .Y(_05479_));
 sky130_fd_sc_hd__mux2_1 _11559_ (.A0(\genblk2[8].wave_shpr.div.acc[2] ),
    .A1(_05479_),
    .S(_05417_),
    .X(_05480_));
 sky130_fd_sc_hd__a22o_1 _11560_ (.A1(net872),
    .A2(_05447_),
    .B1(_05446_),
    .B2(_05480_),
    .X(_00824_));
 sky130_fd_sc_hd__or2b_1 _11561_ (.A(_05380_),
    .B_N(_05372_),
    .X(_05481_));
 sky130_fd_sc_hd__xnor2_1 _11562_ (.A(_05379_),
    .B(_05481_),
    .Y(_05482_));
 sky130_fd_sc_hd__mux2_1 _11563_ (.A0(\genblk2[8].wave_shpr.div.acc[3] ),
    .A1(_05482_),
    .S(_05417_),
    .X(_05483_));
 sky130_fd_sc_hd__a22o_1 _11564_ (.A1(net980),
    .A2(_05447_),
    .B1(_05446_),
    .B2(_05483_),
    .X(_00825_));
 sky130_fd_sc_hd__clkbuf_4 _11565_ (.A(_05444_),
    .X(_05484_));
 sky130_fd_sc_hd__or2b_1 _11566_ (.A(_05382_),
    .B_N(_05371_),
    .X(_05485_));
 sky130_fd_sc_hd__xnor2_1 _11567_ (.A(_05485_),
    .B(_05381_),
    .Y(_05486_));
 sky130_fd_sc_hd__mux2_1 _11568_ (.A0(\genblk2[8].wave_shpr.div.acc[4] ),
    .A1(_05486_),
    .S(_05417_),
    .X(_05487_));
 sky130_fd_sc_hd__a22o_1 _11569_ (.A1(net898),
    .A2(_05447_),
    .B1(_05484_),
    .B2(_05487_),
    .X(_00826_));
 sky130_fd_sc_hd__or2b_1 _11570_ (.A(_05384_),
    .B_N(_05370_),
    .X(_05488_));
 sky130_fd_sc_hd__xnor2_1 _11571_ (.A(_05488_),
    .B(_05383_),
    .Y(_05489_));
 sky130_fd_sc_hd__mux2_1 _11572_ (.A0(\genblk2[8].wave_shpr.div.acc[5] ),
    .A1(_05489_),
    .S(_05417_),
    .X(_05490_));
 sky130_fd_sc_hd__a22o_1 _11573_ (.A1(net932),
    .A2(_05447_),
    .B1(_05484_),
    .B2(_05490_),
    .X(_00827_));
 sky130_fd_sc_hd__or2b_1 _11574_ (.A(_05386_),
    .B_N(_05369_),
    .X(_05491_));
 sky130_fd_sc_hd__xnor2_1 _11575_ (.A(_05385_),
    .B(_05491_),
    .Y(_05492_));
 sky130_fd_sc_hd__clkbuf_4 _11576_ (.A(_05416_),
    .X(_05493_));
 sky130_fd_sc_hd__mux2_1 _11577_ (.A0(\genblk2[8].wave_shpr.div.acc[6] ),
    .A1(_05492_),
    .S(_05493_),
    .X(_05494_));
 sky130_fd_sc_hd__a22o_1 _11578_ (.A1(net950),
    .A2(_05447_),
    .B1(_05484_),
    .B2(_05494_),
    .X(_00828_));
 sky130_fd_sc_hd__or2b_1 _11579_ (.A(_05388_),
    .B_N(_05368_),
    .X(_05495_));
 sky130_fd_sc_hd__xnor2_1 _11580_ (.A(_05387_),
    .B(_05495_),
    .Y(_05496_));
 sky130_fd_sc_hd__mux2_1 _11581_ (.A0(\genblk2[8].wave_shpr.div.acc[7] ),
    .A1(_05496_),
    .S(_05493_),
    .X(_05497_));
 sky130_fd_sc_hd__a22o_1 _11582_ (.A1(net978),
    .A2(_05447_),
    .B1(_05484_),
    .B2(_05497_),
    .X(_00829_));
 sky130_fd_sc_hd__or2b_1 _11583_ (.A(_05390_),
    .B_N(_05367_),
    .X(_05498_));
 sky130_fd_sc_hd__xnor2_1 _11584_ (.A(_05389_),
    .B(_05498_),
    .Y(_05499_));
 sky130_fd_sc_hd__mux2_1 _11585_ (.A0(\genblk2[8].wave_shpr.div.acc[8] ),
    .A1(_05499_),
    .S(_05493_),
    .X(_05500_));
 sky130_fd_sc_hd__a22o_1 _11586_ (.A1(net922),
    .A2(_05447_),
    .B1(_05484_),
    .B2(_05500_),
    .X(_00830_));
 sky130_fd_sc_hd__or2b_1 _11587_ (.A(_05392_),
    .B_N(_05366_),
    .X(_05501_));
 sky130_fd_sc_hd__xnor2_1 _11588_ (.A(_05391_),
    .B(_05501_),
    .Y(_05502_));
 sky130_fd_sc_hd__mux2_1 _11589_ (.A0(\genblk2[8].wave_shpr.div.acc[9] ),
    .A1(_05502_),
    .S(_05493_),
    .X(_05503_));
 sky130_fd_sc_hd__a22o_1 _11590_ (.A1(net908),
    .A2(_05447_),
    .B1(_05484_),
    .B2(_05503_),
    .X(_00831_));
 sky130_fd_sc_hd__or2b_1 _11591_ (.A(_05394_),
    .B_N(_05365_),
    .X(_05504_));
 sky130_fd_sc_hd__xnor2_1 _11592_ (.A(_05393_),
    .B(_05504_),
    .Y(_05505_));
 sky130_fd_sc_hd__mux2_1 _11593_ (.A0(\genblk2[8].wave_shpr.div.acc[10] ),
    .A1(_05505_),
    .S(_05493_),
    .X(_05506_));
 sky130_fd_sc_hd__a22o_1 _11594_ (.A1(net917),
    .A2(_05447_),
    .B1(_05484_),
    .B2(_05506_),
    .X(_00832_));
 sky130_fd_sc_hd__clkbuf_4 _11595_ (.A(_05441_),
    .X(_05507_));
 sky130_fd_sc_hd__or2b_1 _11596_ (.A(_05396_),
    .B_N(_05364_),
    .X(_05508_));
 sky130_fd_sc_hd__xnor2_1 _11597_ (.A(_05395_),
    .B(_05508_),
    .Y(_05509_));
 sky130_fd_sc_hd__mux2_1 _11598_ (.A0(\genblk2[8].wave_shpr.div.acc[11] ),
    .A1(_05509_),
    .S(_05493_),
    .X(_05510_));
 sky130_fd_sc_hd__a22o_1 _11599_ (.A1(net909),
    .A2(_05507_),
    .B1(_05484_),
    .B2(_05510_),
    .X(_00833_));
 sky130_fd_sc_hd__or2b_1 _11600_ (.A(_05398_),
    .B_N(_05363_),
    .X(_05511_));
 sky130_fd_sc_hd__xnor2_1 _11601_ (.A(_05397_),
    .B(_05511_),
    .Y(_05512_));
 sky130_fd_sc_hd__mux2_1 _11602_ (.A0(\genblk2[8].wave_shpr.div.acc[12] ),
    .A1(_05512_),
    .S(_05493_),
    .X(_05513_));
 sky130_fd_sc_hd__a22o_1 _11603_ (.A1(net833),
    .A2(_05507_),
    .B1(_05484_),
    .B2(_05513_),
    .X(_00834_));
 sky130_fd_sc_hd__or2b_1 _11604_ (.A(_05400_),
    .B_N(_05362_),
    .X(_05514_));
 sky130_fd_sc_hd__xnor2_1 _11605_ (.A(_05399_),
    .B(_05514_),
    .Y(_05515_));
 sky130_fd_sc_hd__mux2_1 _11606_ (.A0(\genblk2[8].wave_shpr.div.acc[13] ),
    .A1(_05515_),
    .S(_05493_),
    .X(_05516_));
 sky130_fd_sc_hd__a22o_1 _11607_ (.A1(net846),
    .A2(_05507_),
    .B1(_05484_),
    .B2(_05516_),
    .X(_00835_));
 sky130_fd_sc_hd__or2b_1 _11608_ (.A(_05402_),
    .B_N(_05361_),
    .X(_05517_));
 sky130_fd_sc_hd__xnor2_1 _11609_ (.A(_05401_),
    .B(_05517_),
    .Y(_05518_));
 sky130_fd_sc_hd__mux2_1 _11610_ (.A0(net846),
    .A1(_05518_),
    .S(_05493_),
    .X(_05519_));
 sky130_fd_sc_hd__a22o_1 _11611_ (.A1(net947),
    .A2(_05507_),
    .B1(_05445_),
    .B2(_05519_),
    .X(_00836_));
 sky130_fd_sc_hd__or2b_1 _11612_ (.A(_05404_),
    .B_N(_05360_),
    .X(_05520_));
 sky130_fd_sc_hd__xnor2_1 _11613_ (.A(_05403_),
    .B(_05520_),
    .Y(_05521_));
 sky130_fd_sc_hd__mux2_1 _11614_ (.A0(\genblk2[8].wave_shpr.div.acc[15] ),
    .A1(_05521_),
    .S(_05493_),
    .X(_05522_));
 sky130_fd_sc_hd__a22o_1 _11615_ (.A1(net802),
    .A2(_05507_),
    .B1(_05445_),
    .B2(_05522_),
    .X(_00837_));
 sky130_fd_sc_hd__or2b_1 _11616_ (.A(_05406_),
    .B_N(_05359_),
    .X(_05523_));
 sky130_fd_sc_hd__xnor2_1 _11617_ (.A(_05523_),
    .B(_05405_),
    .Y(_05524_));
 sky130_fd_sc_hd__mux2_1 _11618_ (.A0(\genblk2[8].wave_shpr.div.acc[16] ),
    .A1(_05524_),
    .S(_05416_),
    .X(_05525_));
 sky130_fd_sc_hd__a22o_1 _11619_ (.A1(net991),
    .A2(_05507_),
    .B1(_05445_),
    .B2(_05525_),
    .X(_00838_));
 sky130_fd_sc_hd__or2b_1 _11620_ (.A(_05408_),
    .B_N(_05358_),
    .X(_05526_));
 sky130_fd_sc_hd__xnor2_1 _11621_ (.A(_05407_),
    .B(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hd__mux2_1 _11622_ (.A0(\genblk2[8].wave_shpr.div.acc[17] ),
    .A1(_05527_),
    .S(_05416_),
    .X(_05528_));
 sky130_fd_sc_hd__a22o_1 _11623_ (.A1(net1222),
    .A2(_05507_),
    .B1(_05445_),
    .B2(_05528_),
    .X(_00839_));
 sky130_fd_sc_hd__nand2b_1 _11624_ (.A_N(_05409_),
    .B(_05416_),
    .Y(_05529_));
 sky130_fd_sc_hd__xnor2_1 _11625_ (.A(\genblk2[8].wave_shpr.div.acc[18] ),
    .B(_05529_),
    .Y(_05530_));
 sky130_fd_sc_hd__a22o_1 _11626_ (.A1(net1114),
    .A2(_05507_),
    .B1(_05445_),
    .B2(_05530_),
    .X(_00840_));
 sky130_fd_sc_hd__nor2_1 _11627_ (.A(\genblk2[8].wave_shpr.div.acc[18] ),
    .B(_05529_),
    .Y(_05531_));
 sky130_fd_sc_hd__xnor2_1 _11628_ (.A(\genblk2[8].wave_shpr.div.acc[19] ),
    .B(_05531_),
    .Y(_05532_));
 sky130_fd_sc_hd__a2bb2o_1 _11629_ (.A1_N(_05471_),
    .A2_N(_05532_),
    .B1(net690),
    .B2(_05442_),
    .X(_00841_));
 sky130_fd_sc_hd__or3_1 _11630_ (.A(\genblk2[8].wave_shpr.div.acc[18] ),
    .B(\genblk2[8].wave_shpr.div.acc[19] ),
    .C(_05529_),
    .X(_05533_));
 sky130_fd_sc_hd__and2b_1 _11631_ (.A_N(_05410_),
    .B(_05416_),
    .X(_05534_));
 sky130_fd_sc_hd__a21o_1 _11632_ (.A1(\genblk2[8].wave_shpr.div.acc[20] ),
    .A2(_05533_),
    .B1(_05534_),
    .X(_05535_));
 sky130_fd_sc_hd__a22o_1 _11633_ (.A1(net1018),
    .A2(_05507_),
    .B1(_05445_),
    .B2(_05535_),
    .X(_00842_));
 sky130_fd_sc_hd__nand2_1 _11634_ (.A(\genblk2[8].wave_shpr.div.acc[21] ),
    .B(_05534_),
    .Y(_05536_));
 sky130_fd_sc_hd__or2_1 _11635_ (.A(\genblk2[8].wave_shpr.div.acc[21] ),
    .B(_05534_),
    .X(_05537_));
 sky130_fd_sc_hd__a32o_1 _11636_ (.A1(_05449_),
    .A2(_05536_),
    .A3(_05537_),
    .B1(_05448_),
    .B2(net456),
    .X(_00843_));
 sky130_fd_sc_hd__nand2_1 _11637_ (.A(\genblk2[8].wave_shpr.div.acc[22] ),
    .B(_05411_),
    .Y(_05538_));
 sky130_fd_sc_hd__a21oi_1 _11638_ (.A1(_05412_),
    .A2(_05538_),
    .B1(_05471_),
    .Y(_05539_));
 sky130_fd_sc_hd__a22o_1 _11639_ (.A1(net704),
    .A2(_05507_),
    .B1(_05417_),
    .B2(_05539_),
    .X(_00844_));
 sky130_fd_sc_hd__and2b_1 _11640_ (.A_N(_05413_),
    .B(_05416_),
    .X(_05540_));
 sky130_fd_sc_hd__a21o_1 _11641_ (.A1(\genblk2[8].wave_shpr.div.acc[23] ),
    .A2(_05412_),
    .B1(_05540_),
    .X(_05541_));
 sky130_fd_sc_hd__a22o_1 _11642_ (.A1(net946),
    .A2(_05448_),
    .B1(_05445_),
    .B2(_05541_),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _11643_ (.A0(_05540_),
    .A1(_05413_),
    .S(\genblk2[8].wave_shpr.div.acc[24] ),
    .X(_05542_));
 sky130_fd_sc_hd__a22o_1 _11644_ (.A1(net1052),
    .A2(_05448_),
    .B1(_05445_),
    .B2(_05542_),
    .X(_00846_));
 sky130_fd_sc_hd__or3b_1 _11645_ (.A(_05414_),
    .B(\genblk2[8].wave_shpr.div.acc[25] ),
    .C_N(\genblk2[8].wave_shpr.div.acc[26] ),
    .X(_05543_));
 sky130_fd_sc_hd__a21bo_1 _11646_ (.A1(\genblk2[8].wave_shpr.div.acc[25] ),
    .A2(_05414_),
    .B1_N(_05543_),
    .X(_05544_));
 sky130_fd_sc_hd__a22o_1 _11647_ (.A1(net615),
    .A2(_05448_),
    .B1(_05445_),
    .B2(_05544_),
    .X(_00847_));
 sky130_fd_sc_hd__mux2_1 _11648_ (.A0(_05444_),
    .A1(_05441_),
    .S(\genblk2[8].wave_shpr.div.i[0] ),
    .X(_05545_));
 sky130_fd_sc_hd__clkbuf_1 _11649_ (.A(_05545_),
    .X(_00848_));
 sky130_fd_sc_hd__or2_1 _11650_ (.A(\genblk2[8].wave_shpr.div.i[1] ),
    .B(\genblk2[8].wave_shpr.div.i[0] ),
    .X(_05546_));
 sky130_fd_sc_hd__nand2_1 _11651_ (.A(\genblk2[8].wave_shpr.div.i[1] ),
    .B(\genblk2[8].wave_shpr.div.i[0] ),
    .Y(_05547_));
 sky130_fd_sc_hd__a32o_1 _11652_ (.A1(_05449_),
    .A2(_05546_),
    .A3(_05547_),
    .B1(_05448_),
    .B2(net1098),
    .X(_00849_));
 sky130_fd_sc_hd__a21o_1 _11653_ (.A1(\genblk2[8].wave_shpr.div.i[1] ),
    .A2(\genblk2[8].wave_shpr.div.i[0] ),
    .B1(\genblk2[8].wave_shpr.div.i[2] ),
    .X(_05548_));
 sky130_fd_sc_hd__and3_1 _11654_ (.A(\genblk2[8].wave_shpr.div.i[1] ),
    .B(\genblk2[8].wave_shpr.div.i[0] ),
    .C(\genblk2[8].wave_shpr.div.i[2] ),
    .X(_05549_));
 sky130_fd_sc_hd__inv_2 _11655_ (.A(_05549_),
    .Y(_05550_));
 sky130_fd_sc_hd__a32o_1 _11656_ (.A1(_05449_),
    .A2(_05548_),
    .A3(_05550_),
    .B1(_05448_),
    .B2(net726),
    .X(_00850_));
 sky130_fd_sc_hd__a21oi_1 _11657_ (.A1(_00020_),
    .A2(_05549_),
    .B1(net1164),
    .Y(_05551_));
 sky130_fd_sc_hd__and3_1 _11658_ (.A(\genblk2[8].wave_shpr.div.i[3] ),
    .B(_02197_),
    .C(_05549_),
    .X(_05552_));
 sky130_fd_sc_hd__nor3_1 _11659_ (.A(_03690_),
    .B(_05551_),
    .C(_05552_),
    .Y(_00851_));
 sky130_fd_sc_hd__o21ai_1 _11660_ (.A1(net319),
    .A2(_05552_),
    .B1(_03855_),
    .Y(_05553_));
 sky130_fd_sc_hd__a21oi_1 _11661_ (.A1(net319),
    .A2(_05552_),
    .B1(_05553_),
    .Y(_00852_));
 sky130_fd_sc_hd__or2b_1 _11662_ (.A(\genblk2[9].wave_shpr.div.acc[17] ),
    .B_N(\genblk2[9].wave_shpr.div.b1[17] ),
    .X(_05554_));
 sky130_fd_sc_hd__nor2_1 _11663_ (.A(_05439_),
    .B(\genblk2[9].wave_shpr.div.acc[16] ),
    .Y(_05555_));
 sky130_fd_sc_hd__or2b_1 _11664_ (.A(\genblk2[9].wave_shpr.div.acc[15] ),
    .B_N(\genblk2[9].wave_shpr.div.b1[15] ),
    .X(_05556_));
 sky130_fd_sc_hd__or2b_1 _11665_ (.A(\genblk2[9].wave_shpr.div.acc[14] ),
    .B_N(\genblk2[9].wave_shpr.div.b1[14] ),
    .X(_05557_));
 sky130_fd_sc_hd__or2b_1 _11666_ (.A(\genblk2[9].wave_shpr.div.acc[13] ),
    .B_N(\genblk2[9].wave_shpr.div.b1[13] ),
    .X(_05558_));
 sky130_fd_sc_hd__or2b_1 _11667_ (.A(\genblk2[9].wave_shpr.div.acc[12] ),
    .B_N(\genblk2[9].wave_shpr.div.b1[12] ),
    .X(_05559_));
 sky130_fd_sc_hd__or2b_1 _11668_ (.A(\genblk2[9].wave_shpr.div.acc[11] ),
    .B_N(\genblk2[9].wave_shpr.div.b1[11] ),
    .X(_05560_));
 sky130_fd_sc_hd__or2b_1 _11669_ (.A(\genblk2[9].wave_shpr.div.acc[10] ),
    .B_N(\genblk2[9].wave_shpr.div.b1[10] ),
    .X(_05561_));
 sky130_fd_sc_hd__or2b_1 _11670_ (.A(\genblk2[9].wave_shpr.div.acc[9] ),
    .B_N(\genblk2[9].wave_shpr.div.b1[9] ),
    .X(_05562_));
 sky130_fd_sc_hd__or2b_1 _11671_ (.A(\genblk2[9].wave_shpr.div.acc[8] ),
    .B_N(\genblk2[9].wave_shpr.div.b1[8] ),
    .X(_05563_));
 sky130_fd_sc_hd__or2b_1 _11672_ (.A(\genblk2[9].wave_shpr.div.acc[7] ),
    .B_N(\genblk2[9].wave_shpr.div.b1[7] ),
    .X(_05564_));
 sky130_fd_sc_hd__or2b_1 _11673_ (.A(\genblk2[9].wave_shpr.div.acc[6] ),
    .B_N(\genblk2[9].wave_shpr.div.b1[6] ),
    .X(_05565_));
 sky130_fd_sc_hd__or2b_1 _11674_ (.A(\genblk2[9].wave_shpr.div.acc[5] ),
    .B_N(\genblk2[9].wave_shpr.div.b1[5] ),
    .X(_05566_));
 sky130_fd_sc_hd__or2b_1 _11675_ (.A(\genblk2[9].wave_shpr.div.b1[4] ),
    .B_N(\genblk2[9].wave_shpr.div.acc[4] ),
    .X(_05567_));
 sky130_fd_sc_hd__or2b_1 _11676_ (.A(\genblk2[9].wave_shpr.div.acc[4] ),
    .B_N(\genblk2[9].wave_shpr.div.b1[4] ),
    .X(_05568_));
 sky130_fd_sc_hd__nand2_1 _11677_ (.A(_05567_),
    .B(_05568_),
    .Y(_05569_));
 sky130_fd_sc_hd__or2b_1 _11678_ (.A(\genblk2[9].wave_shpr.div.acc[3] ),
    .B_N(\genblk2[9].wave_shpr.div.b1[3] ),
    .X(_05570_));
 sky130_fd_sc_hd__or2b_1 _11679_ (.A(\genblk2[9].wave_shpr.div.acc[2] ),
    .B_N(\genblk2[9].wave_shpr.div.b1[2] ),
    .X(_05571_));
 sky130_fd_sc_hd__inv_2 _11680_ (.A(\genblk2[9].wave_shpr.div.b1[1] ),
    .Y(_05572_));
 sky130_fd_sc_hd__inv_2 _11681_ (.A(\genblk2[9].wave_shpr.div.acc[0] ),
    .Y(_05573_));
 sky130_fd_sc_hd__xor2_1 _11682_ (.A(\genblk2[9].wave_shpr.div.b1[1] ),
    .B(\genblk2[9].wave_shpr.div.acc[1] ),
    .X(_05574_));
 sky130_fd_sc_hd__a21oi_1 _11683_ (.A1(\genblk2[9].wave_shpr.div.b1[0] ),
    .A2(_05573_),
    .B1(_05574_),
    .Y(_05575_));
 sky130_fd_sc_hd__a21o_1 _11684_ (.A1(_05572_),
    .A2(\genblk2[9].wave_shpr.div.acc[1] ),
    .B1(_05575_),
    .X(_05576_));
 sky130_fd_sc_hd__and2b_1 _11685_ (.A_N(\genblk2[9].wave_shpr.div.b1[2] ),
    .B(\genblk2[9].wave_shpr.div.acc[2] ),
    .X(_05577_));
 sky130_fd_sc_hd__a21o_1 _11686_ (.A1(_05571_),
    .A2(_05576_),
    .B1(_05577_),
    .X(_05578_));
 sky130_fd_sc_hd__and2b_1 _11687_ (.A_N(\genblk2[9].wave_shpr.div.b1[3] ),
    .B(\genblk2[9].wave_shpr.div.acc[3] ),
    .X(_05579_));
 sky130_fd_sc_hd__a21oi_1 _11688_ (.A1(_05570_),
    .A2(_05578_),
    .B1(_05579_),
    .Y(_05580_));
 sky130_fd_sc_hd__o21ai_1 _11689_ (.A1(_05569_),
    .A2(_05580_),
    .B1(_05567_),
    .Y(_05581_));
 sky130_fd_sc_hd__and2b_1 _11690_ (.A_N(\genblk2[9].wave_shpr.div.b1[5] ),
    .B(\genblk2[9].wave_shpr.div.acc[5] ),
    .X(_05582_));
 sky130_fd_sc_hd__a21o_1 _11691_ (.A1(_05566_),
    .A2(_05581_),
    .B1(_05582_),
    .X(_05583_));
 sky130_fd_sc_hd__and2b_1 _11692_ (.A_N(\genblk2[9].wave_shpr.div.b1[6] ),
    .B(\genblk2[9].wave_shpr.div.acc[6] ),
    .X(_05584_));
 sky130_fd_sc_hd__a21o_1 _11693_ (.A1(_05565_),
    .A2(_05583_),
    .B1(_05584_),
    .X(_05585_));
 sky130_fd_sc_hd__and2b_1 _11694_ (.A_N(\genblk2[9].wave_shpr.div.b1[7] ),
    .B(\genblk2[9].wave_shpr.div.acc[7] ),
    .X(_05586_));
 sky130_fd_sc_hd__a21o_1 _11695_ (.A1(_05564_),
    .A2(_05585_),
    .B1(_05586_),
    .X(_05587_));
 sky130_fd_sc_hd__and2b_1 _11696_ (.A_N(\genblk2[9].wave_shpr.div.b1[8] ),
    .B(\genblk2[9].wave_shpr.div.acc[8] ),
    .X(_05588_));
 sky130_fd_sc_hd__a21o_1 _11697_ (.A1(_05563_),
    .A2(_05587_),
    .B1(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__and2b_1 _11698_ (.A_N(\genblk2[9].wave_shpr.div.b1[9] ),
    .B(\genblk2[9].wave_shpr.div.acc[9] ),
    .X(_05590_));
 sky130_fd_sc_hd__a21o_1 _11699_ (.A1(_05562_),
    .A2(_05589_),
    .B1(_05590_),
    .X(_05591_));
 sky130_fd_sc_hd__and2b_1 _11700_ (.A_N(\genblk2[9].wave_shpr.div.b1[10] ),
    .B(\genblk2[9].wave_shpr.div.acc[10] ),
    .X(_05592_));
 sky130_fd_sc_hd__a21o_1 _11701_ (.A1(_05561_),
    .A2(_05591_),
    .B1(_05592_),
    .X(_05593_));
 sky130_fd_sc_hd__and2b_1 _11702_ (.A_N(\genblk2[9].wave_shpr.div.b1[11] ),
    .B(\genblk2[9].wave_shpr.div.acc[11] ),
    .X(_05594_));
 sky130_fd_sc_hd__a21o_1 _11703_ (.A1(_05560_),
    .A2(_05593_),
    .B1(_05594_),
    .X(_05595_));
 sky130_fd_sc_hd__and2b_1 _11704_ (.A_N(\genblk2[9].wave_shpr.div.b1[12] ),
    .B(\genblk2[9].wave_shpr.div.acc[12] ),
    .X(_05596_));
 sky130_fd_sc_hd__a21o_1 _11705_ (.A1(_05559_),
    .A2(_05595_),
    .B1(_05596_),
    .X(_05597_));
 sky130_fd_sc_hd__and2b_1 _11706_ (.A_N(\genblk2[9].wave_shpr.div.b1[13] ),
    .B(\genblk2[9].wave_shpr.div.acc[13] ),
    .X(_05598_));
 sky130_fd_sc_hd__a21o_1 _11707_ (.A1(_05558_),
    .A2(_05597_),
    .B1(_05598_),
    .X(_05599_));
 sky130_fd_sc_hd__and2b_1 _11708_ (.A_N(\genblk2[9].wave_shpr.div.b1[14] ),
    .B(\genblk2[9].wave_shpr.div.acc[14] ),
    .X(_05600_));
 sky130_fd_sc_hd__a21o_1 _11709_ (.A1(_05557_),
    .A2(_05599_),
    .B1(_05600_),
    .X(_05601_));
 sky130_fd_sc_hd__and2b_1 _11710_ (.A_N(\genblk2[9].wave_shpr.div.b1[15] ),
    .B(\genblk2[9].wave_shpr.div.acc[15] ),
    .X(_05602_));
 sky130_fd_sc_hd__a21oi_2 _11711_ (.A1(_05556_),
    .A2(_05601_),
    .B1(_05602_),
    .Y(_05603_));
 sky130_fd_sc_hd__and2_1 _11712_ (.A(_05439_),
    .B(\genblk2[9].wave_shpr.div.acc[16] ),
    .X(_05604_));
 sky130_fd_sc_hd__o21bai_2 _11713_ (.A1(_05555_),
    .A2(_05603_),
    .B1_N(_05604_),
    .Y(_05605_));
 sky130_fd_sc_hd__and2b_1 _11714_ (.A_N(\genblk2[9].wave_shpr.div.b1[17] ),
    .B(\genblk2[9].wave_shpr.div.acc[17] ),
    .X(_05606_));
 sky130_fd_sc_hd__a21o_1 _11715_ (.A1(_05554_),
    .A2(_05605_),
    .B1(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__or2_1 _11716_ (.A(\genblk2[9].wave_shpr.div.acc[18] ),
    .B(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__or4_1 _11717_ (.A(\genblk2[9].wave_shpr.div.acc[21] ),
    .B(\genblk2[9].wave_shpr.div.acc[20] ),
    .C(\genblk2[9].wave_shpr.div.acc[19] ),
    .D(_05608_),
    .X(_05609_));
 sky130_fd_sc_hd__or2_1 _11718_ (.A(\genblk2[9].wave_shpr.div.acc[22] ),
    .B(_05609_),
    .X(_05610_));
 sky130_fd_sc_hd__or4_2 _11719_ (.A(\genblk2[9].wave_shpr.div.acc[23] ),
    .B(\genblk2[9].wave_shpr.div.acc[25] ),
    .C(\genblk2[9].wave_shpr.div.acc[24] ),
    .D(\genblk2[9].wave_shpr.div.acc[26] ),
    .X(_05611_));
 sky130_fd_sc_hd__or2_1 _11720_ (.A(_05610_),
    .B(_05611_),
    .X(_05612_));
 sky130_fd_sc_hd__buf_4 _11721_ (.A(_05612_),
    .X(_05613_));
 sky130_fd_sc_hd__mux2_1 _11722_ (.A0(\genblk2[9].wave_shpr.div.fin_quo[0] ),
    .A1(_05613_),
    .S(_00023_),
    .X(_05614_));
 sky130_fd_sc_hd__clkbuf_1 _11723_ (.A(_05614_),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _11724_ (.A0(\genblk2[9].wave_shpr.div.fin_quo[1] ),
    .A1(net1328),
    .S(_00023_),
    .X(_05615_));
 sky130_fd_sc_hd__clkbuf_1 _11725_ (.A(_05615_),
    .X(_00854_));
 sky130_fd_sc_hd__mux2_1 _11726_ (.A0(\genblk2[9].wave_shpr.div.fin_quo[2] ),
    .A1(net1313),
    .S(_00023_),
    .X(_05616_));
 sky130_fd_sc_hd__clkbuf_1 _11727_ (.A(_05616_),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_1 _11728_ (.A0(\genblk2[9].wave_shpr.div.fin_quo[3] ),
    .A1(\genblk2[9].wave_shpr.div.quo[2] ),
    .S(_00023_),
    .X(_05617_));
 sky130_fd_sc_hd__clkbuf_1 _11729_ (.A(_05617_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _11730_ (.A0(\genblk2[9].wave_shpr.div.fin_quo[4] ),
    .A1(\genblk2[9].wave_shpr.div.quo[3] ),
    .S(_00023_),
    .X(_05618_));
 sky130_fd_sc_hd__clkbuf_1 _11731_ (.A(_05618_),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_1 _11732_ (.A0(\genblk2[9].wave_shpr.div.fin_quo[5] ),
    .A1(net1317),
    .S(_00023_),
    .X(_05619_));
 sky130_fd_sc_hd__clkbuf_1 _11733_ (.A(_05619_),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_1 _11734_ (.A0(\genblk2[9].wave_shpr.div.fin_quo[6] ),
    .A1(\genblk2[9].wave_shpr.div.quo[5] ),
    .S(_00023_),
    .X(_05620_));
 sky130_fd_sc_hd__clkbuf_1 _11735_ (.A(_05620_),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _11736_ (.A0(net1259),
    .A1(\genblk2[9].wave_shpr.div.quo[6] ),
    .S(_00023_),
    .X(_05621_));
 sky130_fd_sc_hd__clkbuf_1 _11737_ (.A(_05621_),
    .X(_00860_));
 sky130_fd_sc_hd__nand2_1 _11738_ (.A(_02248_),
    .B(_01150_),
    .Y(_05622_));
 sky130_fd_sc_hd__a2bb2o_1 _11739_ (.A1_N(_01099_),
    .A2_N(_01147_),
    .B1(_05622_),
    .B2(net1161),
    .X(_00861_));
 sky130_fd_sc_hd__a2bb2o_1 _11740_ (.A1_N(_01099_),
    .A2_N(_01149_),
    .B1(_05622_),
    .B2(net497),
    .X(_00862_));
 sky130_fd_sc_hd__a22o_1 _11741_ (.A1(_02248_),
    .A2(_01145_),
    .B1(_05622_),
    .B2(net1073),
    .X(_00863_));
 sky130_fd_sc_hd__a22o_1 _11742_ (.A1(_02248_),
    .A2(_01144_),
    .B1(_05622_),
    .B2(net1088),
    .X(_00864_));
 sky130_fd_sc_hd__clkbuf_4 _11743_ (.A(_02203_),
    .X(_05623_));
 sky130_fd_sc_hd__clkbuf_4 _11744_ (.A(_03693_),
    .X(_05624_));
 sky130_fd_sc_hd__a22o_1 _11745_ (.A1(net746),
    .A2(_05623_),
    .B1(_05624_),
    .B2(_05613_),
    .X(_00865_));
 sky130_fd_sc_hd__a22o_1 _11746_ (.A1(net649),
    .A2(_05623_),
    .B1(_05624_),
    .B2(net746),
    .X(_00866_));
 sky130_fd_sc_hd__a22o_1 _11747_ (.A1(\genblk2[9].wave_shpr.div.quo[2] ),
    .A2(_05623_),
    .B1(_05624_),
    .B2(net649),
    .X(_00867_));
 sky130_fd_sc_hd__a22o_1 _11748_ (.A1(\genblk2[9].wave_shpr.div.quo[3] ),
    .A2(_05623_),
    .B1(_05624_),
    .B2(net686),
    .X(_00868_));
 sky130_fd_sc_hd__a22o_1 _11749_ (.A1(net586),
    .A2(_05623_),
    .B1(_05624_),
    .B2(net700),
    .X(_00869_));
 sky130_fd_sc_hd__a22o_1 _11750_ (.A1(\genblk2[9].wave_shpr.div.quo[5] ),
    .A2(_05623_),
    .B1(_05624_),
    .B2(net586),
    .X(_00870_));
 sky130_fd_sc_hd__a22o_1 _11751_ (.A1(net267),
    .A2(_05623_),
    .B1(_05624_),
    .B2(net712),
    .X(_00871_));
 sky130_fd_sc_hd__a22o_1 _11752_ (.A1(\genblk2[9].wave_shpr.div.quo[7] ),
    .A2(_05623_),
    .B1(_05624_),
    .B2(net267),
    .X(_00872_));
 sky130_fd_sc_hd__a22o_1 _11753_ (.A1(net526),
    .A2(_05623_),
    .B1(_05624_),
    .B2(net1085),
    .X(_00873_));
 sky130_fd_sc_hd__and2_1 _11754_ (.A(_05464_),
    .B(\genblk1[9].osc.clkdiv_C.cnt[0] ),
    .X(_05625_));
 sky130_fd_sc_hd__a221o_1 _11755_ (.A1(net290),
    .A2(_03696_),
    .B1(_03694_),
    .B2(net526),
    .C1(_05625_),
    .X(_00874_));
 sky130_fd_sc_hd__and2_1 _11756_ (.A(_05464_),
    .B(\genblk1[9].osc.clkdiv_C.cnt[1] ),
    .X(_05626_));
 sky130_fd_sc_hd__a221o_1 _11757_ (.A1(\genblk2[9].wave_shpr.div.quo[10] ),
    .A2(_03696_),
    .B1(_03694_),
    .B2(net290),
    .C1(_05626_),
    .X(_00875_));
 sky130_fd_sc_hd__and2_1 _11758_ (.A(_05464_),
    .B(\genblk1[9].osc.clkdiv_C.cnt[2] ),
    .X(_05627_));
 sky130_fd_sc_hd__a221o_1 _11759_ (.A1(net481),
    .A2(_03696_),
    .B1(_03694_),
    .B2(net557),
    .C1(_05627_),
    .X(_00876_));
 sky130_fd_sc_hd__clkbuf_4 _11760_ (.A(_02203_),
    .X(_05628_));
 sky130_fd_sc_hd__clkbuf_4 _11761_ (.A(_03693_),
    .X(_05629_));
 sky130_fd_sc_hd__and2_1 _11762_ (.A(_05464_),
    .B(\genblk1[9].osc.clkdiv_C.cnt[3] ),
    .X(_05630_));
 sky130_fd_sc_hd__a221o_1 _11763_ (.A1(net243),
    .A2(_05628_),
    .B1(_05629_),
    .B2(net481),
    .C1(_05630_),
    .X(_00877_));
 sky130_fd_sc_hd__clkbuf_2 _11764_ (.A(_02155_),
    .X(_05631_));
 sky130_fd_sc_hd__and2_1 _11765_ (.A(_05631_),
    .B(\genblk1[9].osc.clkdiv_C.cnt[4] ),
    .X(_05632_));
 sky130_fd_sc_hd__a221o_1 _11766_ (.A1(\genblk2[9].wave_shpr.div.quo[13] ),
    .A2(_05628_),
    .B1(_05629_),
    .B2(net243),
    .C1(_05632_),
    .X(_00878_));
 sky130_fd_sc_hd__and2_1 _11767_ (.A(_05631_),
    .B(\genblk1[9].osc.clkdiv_C.cnt[5] ),
    .X(_05633_));
 sky130_fd_sc_hd__a221o_1 _11768_ (.A1(net485),
    .A2(_05628_),
    .B1(_05629_),
    .B2(net541),
    .C1(_05633_),
    .X(_00879_));
 sky130_fd_sc_hd__and2_1 _11769_ (.A(_05631_),
    .B(\genblk1[9].osc.clkdiv_C.cnt[6] ),
    .X(_05634_));
 sky130_fd_sc_hd__a221o_1 _11770_ (.A1(net304),
    .A2(_05628_),
    .B1(_05629_),
    .B2(net485),
    .C1(_05634_),
    .X(_00880_));
 sky130_fd_sc_hd__and2_1 _11771_ (.A(_05631_),
    .B(\genblk1[9].osc.clkdiv_C.cnt[7] ),
    .X(_05635_));
 sky130_fd_sc_hd__a221o_1 _11772_ (.A1(\genblk2[9].wave_shpr.div.quo[16] ),
    .A2(_05628_),
    .B1(_05629_),
    .B2(net304),
    .C1(_05635_),
    .X(_00881_));
 sky130_fd_sc_hd__nor2_1 _11773_ (.A(_04676_),
    .B(_01928_),
    .Y(_05636_));
 sky130_fd_sc_hd__a221o_1 _11774_ (.A1(\genblk2[9].wave_shpr.div.quo[17] ),
    .A2(_05628_),
    .B1(_05629_),
    .B2(net349),
    .C1(_05636_),
    .X(_00882_));
 sky130_fd_sc_hd__nor2_1 _11775_ (.A(_04676_),
    .B(_01930_),
    .Y(_05637_));
 sky130_fd_sc_hd__a221o_1 _11776_ (.A1(net513),
    .A2(_05628_),
    .B1(_05629_),
    .B2(net530),
    .C1(_05637_),
    .X(_00883_));
 sky130_fd_sc_hd__nor2_1 _11777_ (.A(_04676_),
    .B(_02268_),
    .Y(_05638_));
 sky130_fd_sc_hd__a221o_1 _11778_ (.A1(net362),
    .A2(_05628_),
    .B1(_05629_),
    .B2(net513),
    .C1(_05638_),
    .X(_00884_));
 sky130_fd_sc_hd__and2_1 _11779_ (.A(_05631_),
    .B(\genblk1[9].osc.clkdiv_C.cnt[11] ),
    .X(_05639_));
 sky130_fd_sc_hd__a221o_1 _11780_ (.A1(\genblk2[9].wave_shpr.div.quo[20] ),
    .A2(_05628_),
    .B1(_05629_),
    .B2(net362),
    .C1(_05639_),
    .X(_00885_));
 sky130_fd_sc_hd__and2_1 _11781_ (.A(_05631_),
    .B(\genblk1[9].osc.clkdiv_C.cnt[12] ),
    .X(_05640_));
 sky130_fd_sc_hd__a221o_1 _11782_ (.A1(net416),
    .A2(_05628_),
    .B1(_05629_),
    .B2(net533),
    .C1(_05640_),
    .X(_00886_));
 sky130_fd_sc_hd__and2_1 _11783_ (.A(_05631_),
    .B(\genblk1[9].osc.clkdiv_C.cnt[13] ),
    .X(_05641_));
 sky130_fd_sc_hd__a221o_1 _11784_ (.A1(net226),
    .A2(_02203_),
    .B1(_03693_),
    .B2(net416),
    .C1(_05641_),
    .X(_00887_));
 sky130_fd_sc_hd__and2_1 _11785_ (.A(_05631_),
    .B(\genblk1[9].osc.clkdiv_C.cnt[14] ),
    .X(_05642_));
 sky130_fd_sc_hd__a221o_1 _11786_ (.A1(\genblk2[9].wave_shpr.div.quo[23] ),
    .A2(_02203_),
    .B1(_03693_),
    .B2(net226),
    .C1(_05642_),
    .X(_00888_));
 sky130_fd_sc_hd__and2_1 _11787_ (.A(_05631_),
    .B(\genblk1[9].osc.clkdiv_C.cnt[15] ),
    .X(_05643_));
 sky130_fd_sc_hd__a221o_1 _11788_ (.A1(net306),
    .A2(_02203_),
    .B1(_03693_),
    .B2(net565),
    .C1(_05643_),
    .X(_00889_));
 sky130_fd_sc_hd__and2_1 _11789_ (.A(_05631_),
    .B(\genblk1[9].osc.clkdiv_C.cnt[16] ),
    .X(_05644_));
 sky130_fd_sc_hd__a221o_1 _11790_ (.A1(\genblk2[9].wave_shpr.div.acc_next[0] ),
    .A2(_02203_),
    .B1(_03693_),
    .B2(net306),
    .C1(_05644_),
    .X(_00890_));
 sky130_fd_sc_hd__or2b_1 _11791_ (.A(\genblk2[9].wave_shpr.div.acc_next[0] ),
    .B_N(_03693_),
    .X(_05645_));
 sky130_fd_sc_hd__o221a_1 _11792_ (.A1(_03819_),
    .A2(\genblk1[9].osc.clkdiv_C.cnt[17] ),
    .B1(_00022_),
    .B2(net1209),
    .C1(_05645_),
    .X(_00891_));
 sky130_fd_sc_hd__nor2_1 _11793_ (.A(_05610_),
    .B(_05611_),
    .Y(_05646_));
 sky130_fd_sc_hd__or3b_1 _11794_ (.A(_05646_),
    .B(_05573_),
    .C_N(\genblk2[9].wave_shpr.div.b1[0] ),
    .X(_05647_));
 sky130_fd_sc_hd__a21o_1 _11795_ (.A1(\genblk2[9].wave_shpr.div.b1[0] ),
    .A2(_05613_),
    .B1(\genblk2[9].wave_shpr.div.acc[0] ),
    .X(_05648_));
 sky130_fd_sc_hd__a32o_1 _11796_ (.A1(_03694_),
    .A2(_05647_),
    .A3(_05648_),
    .B1(_03696_),
    .B2(net1059),
    .X(_00892_));
 sky130_fd_sc_hd__and3_1 _11797_ (.A(\genblk2[9].wave_shpr.div.b1[0] ),
    .B(_05573_),
    .C(_05574_),
    .X(_05649_));
 sky130_fd_sc_hd__nor2_1 _11798_ (.A(_05575_),
    .B(_05649_),
    .Y(_05650_));
 sky130_fd_sc_hd__mux2_1 _11799_ (.A0(\genblk2[9].wave_shpr.div.acc[1] ),
    .A1(_05650_),
    .S(_05613_),
    .X(_05651_));
 sky130_fd_sc_hd__a22o_1 _11800_ (.A1(net1022),
    .A2(_05623_),
    .B1(_05624_),
    .B2(_05651_),
    .X(_00893_));
 sky130_fd_sc_hd__clkbuf_4 _11801_ (.A(_02203_),
    .X(_05652_));
 sky130_fd_sc_hd__clkbuf_4 _11802_ (.A(_03693_),
    .X(_05653_));
 sky130_fd_sc_hd__or2b_1 _11803_ (.A(_05577_),
    .B_N(_05571_),
    .X(_05654_));
 sky130_fd_sc_hd__xnor2_1 _11804_ (.A(_05576_),
    .B(_05654_),
    .Y(_05655_));
 sky130_fd_sc_hd__mux2_1 _11805_ (.A0(\genblk2[9].wave_shpr.div.acc[2] ),
    .A1(_05655_),
    .S(_05613_),
    .X(_05656_));
 sky130_fd_sc_hd__a22o_1 _11806_ (.A1(net1006),
    .A2(_05652_),
    .B1(_05653_),
    .B2(_05656_),
    .X(_00894_));
 sky130_fd_sc_hd__or2b_1 _11807_ (.A(_05579_),
    .B_N(_05570_),
    .X(_05657_));
 sky130_fd_sc_hd__xnor2_1 _11808_ (.A(_05578_),
    .B(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hd__mux2_1 _11809_ (.A0(\genblk2[9].wave_shpr.div.acc[3] ),
    .A1(_05658_),
    .S(_05613_),
    .X(_05659_));
 sky130_fd_sc_hd__a22o_1 _11810_ (.A1(net886),
    .A2(_05652_),
    .B1(_05653_),
    .B2(_05659_),
    .X(_00895_));
 sky130_fd_sc_hd__xor2_1 _11811_ (.A(_05569_),
    .B(_05580_),
    .X(_05660_));
 sky130_fd_sc_hd__mux2_1 _11812_ (.A0(\genblk2[9].wave_shpr.div.acc[4] ),
    .A1(_05660_),
    .S(_05613_),
    .X(_05661_));
 sky130_fd_sc_hd__a22o_1 _11813_ (.A1(net999),
    .A2(_05652_),
    .B1(_05653_),
    .B2(_05661_),
    .X(_00896_));
 sky130_fd_sc_hd__or2b_1 _11814_ (.A(_05582_),
    .B_N(_05566_),
    .X(_05662_));
 sky130_fd_sc_hd__xnor2_1 _11815_ (.A(_05662_),
    .B(_05581_),
    .Y(_05663_));
 sky130_fd_sc_hd__mux2_1 _11816_ (.A0(\genblk2[9].wave_shpr.div.acc[5] ),
    .A1(_05663_),
    .S(_05613_),
    .X(_05664_));
 sky130_fd_sc_hd__a22o_1 _11817_ (.A1(net938),
    .A2(_05652_),
    .B1(_05653_),
    .B2(_05664_),
    .X(_00897_));
 sky130_fd_sc_hd__or2b_1 _11818_ (.A(_05584_),
    .B_N(_05565_),
    .X(_05665_));
 sky130_fd_sc_hd__xnor2_1 _11819_ (.A(_05583_),
    .B(_05665_),
    .Y(_05666_));
 sky130_fd_sc_hd__mux2_1 _11820_ (.A0(\genblk2[9].wave_shpr.div.acc[6] ),
    .A1(_05666_),
    .S(_05613_),
    .X(_05667_));
 sky130_fd_sc_hd__a22o_1 _11821_ (.A1(net984),
    .A2(_05652_),
    .B1(_05653_),
    .B2(_05667_),
    .X(_00898_));
 sky130_fd_sc_hd__or2b_1 _11822_ (.A(_05586_),
    .B_N(_05564_),
    .X(_05668_));
 sky130_fd_sc_hd__xnor2_1 _11823_ (.A(_05585_),
    .B(_05668_),
    .Y(_05669_));
 sky130_fd_sc_hd__mux2_1 _11824_ (.A0(\genblk2[9].wave_shpr.div.acc[7] ),
    .A1(_05669_),
    .S(_05613_),
    .X(_05670_));
 sky130_fd_sc_hd__a22o_1 _11825_ (.A1(net839),
    .A2(_05652_),
    .B1(_05653_),
    .B2(_05670_),
    .X(_00899_));
 sky130_fd_sc_hd__or2b_1 _11826_ (.A(_05588_),
    .B_N(_05563_),
    .X(_05671_));
 sky130_fd_sc_hd__xnor2_1 _11827_ (.A(_05587_),
    .B(_05671_),
    .Y(_05672_));
 sky130_fd_sc_hd__buf_4 _11828_ (.A(_05612_),
    .X(_05673_));
 sky130_fd_sc_hd__mux2_1 _11829_ (.A0(\genblk2[9].wave_shpr.div.acc[8] ),
    .A1(_05672_),
    .S(_05673_),
    .X(_05674_));
 sky130_fd_sc_hd__a22o_1 _11830_ (.A1(net974),
    .A2(_05652_),
    .B1(_05653_),
    .B2(_05674_),
    .X(_00900_));
 sky130_fd_sc_hd__or2b_1 _11831_ (.A(_05590_),
    .B_N(_05562_),
    .X(_05675_));
 sky130_fd_sc_hd__xnor2_1 _11832_ (.A(_05589_),
    .B(_05675_),
    .Y(_05676_));
 sky130_fd_sc_hd__mux2_1 _11833_ (.A0(\genblk2[9].wave_shpr.div.acc[9] ),
    .A1(_05676_),
    .S(_05673_),
    .X(_05677_));
 sky130_fd_sc_hd__a22o_1 _11834_ (.A1(net884),
    .A2(_05652_),
    .B1(_05653_),
    .B2(_05677_),
    .X(_00901_));
 sky130_fd_sc_hd__or2b_1 _11835_ (.A(_05592_),
    .B_N(_05561_),
    .X(_05678_));
 sky130_fd_sc_hd__xnor2_1 _11836_ (.A(_05591_),
    .B(_05678_),
    .Y(_05679_));
 sky130_fd_sc_hd__mux2_1 _11837_ (.A0(\genblk2[9].wave_shpr.div.acc[10] ),
    .A1(_05679_),
    .S(_05673_),
    .X(_05680_));
 sky130_fd_sc_hd__a22o_1 _11838_ (.A1(net807),
    .A2(_05652_),
    .B1(_05653_),
    .B2(_05680_),
    .X(_00902_));
 sky130_fd_sc_hd__or2b_1 _11839_ (.A(_05594_),
    .B_N(_05560_),
    .X(_05681_));
 sky130_fd_sc_hd__xnor2_1 _11840_ (.A(_05593_),
    .B(_05681_),
    .Y(_05682_));
 sky130_fd_sc_hd__mux2_1 _11841_ (.A0(\genblk2[9].wave_shpr.div.acc[11] ),
    .A1(_05682_),
    .S(_05673_),
    .X(_05683_));
 sky130_fd_sc_hd__a22o_1 _11842_ (.A1(net1046),
    .A2(_05652_),
    .B1(_05653_),
    .B2(_05683_),
    .X(_00903_));
 sky130_fd_sc_hd__clkbuf_4 _11843_ (.A(_02203_),
    .X(_05684_));
 sky130_fd_sc_hd__clkbuf_4 _11844_ (.A(_03693_),
    .X(_05685_));
 sky130_fd_sc_hd__or2b_1 _11845_ (.A(_05596_),
    .B_N(_05559_),
    .X(_05686_));
 sky130_fd_sc_hd__xnor2_1 _11846_ (.A(_05595_),
    .B(_05686_),
    .Y(_05687_));
 sky130_fd_sc_hd__mux2_1 _11847_ (.A0(\genblk2[9].wave_shpr.div.acc[12] ),
    .A1(_05687_),
    .S(_05673_),
    .X(_05688_));
 sky130_fd_sc_hd__a22o_1 _11848_ (.A1(net967),
    .A2(_05684_),
    .B1(_05685_),
    .B2(_05688_),
    .X(_00904_));
 sky130_fd_sc_hd__or2b_1 _11849_ (.A(_05598_),
    .B_N(_05558_),
    .X(_05689_));
 sky130_fd_sc_hd__xnor2_1 _11850_ (.A(_05597_),
    .B(_05689_),
    .Y(_05690_));
 sky130_fd_sc_hd__mux2_1 _11851_ (.A0(\genblk2[9].wave_shpr.div.acc[13] ),
    .A1(_05690_),
    .S(_05673_),
    .X(_05691_));
 sky130_fd_sc_hd__a22o_1 _11852_ (.A1(net799),
    .A2(_05684_),
    .B1(_05685_),
    .B2(_05691_),
    .X(_00905_));
 sky130_fd_sc_hd__or2b_1 _11853_ (.A(_05600_),
    .B_N(_05557_),
    .X(_05692_));
 sky130_fd_sc_hd__xnor2_1 _11854_ (.A(_05599_),
    .B(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hd__mux2_1 _11855_ (.A0(\genblk2[9].wave_shpr.div.acc[14] ),
    .A1(_05693_),
    .S(_05673_),
    .X(_05694_));
 sky130_fd_sc_hd__a22o_1 _11856_ (.A1(net912),
    .A2(_05684_),
    .B1(_05685_),
    .B2(_05694_),
    .X(_00906_));
 sky130_fd_sc_hd__or2b_1 _11857_ (.A(_05602_),
    .B_N(_05556_),
    .X(_05695_));
 sky130_fd_sc_hd__xnor2_1 _11858_ (.A(_05601_),
    .B(_05695_),
    .Y(_05696_));
 sky130_fd_sc_hd__mux2_1 _11859_ (.A0(\genblk2[9].wave_shpr.div.acc[15] ),
    .A1(_05696_),
    .S(_05673_),
    .X(_05697_));
 sky130_fd_sc_hd__a22o_1 _11860_ (.A1(net1060),
    .A2(_05684_),
    .B1(_05685_),
    .B2(_05697_),
    .X(_00907_));
 sky130_fd_sc_hd__nor2_1 _11861_ (.A(_05604_),
    .B(_05555_),
    .Y(_05698_));
 sky130_fd_sc_hd__xnor2_1 _11862_ (.A(_05698_),
    .B(_05603_),
    .Y(_05699_));
 sky130_fd_sc_hd__mux2_1 _11863_ (.A0(\genblk2[9].wave_shpr.div.acc[16] ),
    .A1(_05699_),
    .S(_05673_),
    .X(_05700_));
 sky130_fd_sc_hd__a22o_1 _11864_ (.A1(net987),
    .A2(_05684_),
    .B1(_05685_),
    .B2(_05700_),
    .X(_00908_));
 sky130_fd_sc_hd__or2b_1 _11865_ (.A(_05606_),
    .B_N(_05554_),
    .X(_05701_));
 sky130_fd_sc_hd__xnor2_1 _11866_ (.A(_05605_),
    .B(_05701_),
    .Y(_05702_));
 sky130_fd_sc_hd__mux2_1 _11867_ (.A0(\genblk2[9].wave_shpr.div.acc[17] ),
    .A1(_05702_),
    .S(_05673_),
    .X(_05703_));
 sky130_fd_sc_hd__a22o_1 _11868_ (.A1(net669),
    .A2(_05684_),
    .B1(_05685_),
    .B2(_05703_),
    .X(_00909_));
 sky130_fd_sc_hd__or2_1 _11869_ (.A(_05608_),
    .B(_05646_),
    .X(_05704_));
 sky130_fd_sc_hd__o21ai_1 _11870_ (.A1(_05607_),
    .A2(_05646_),
    .B1(\genblk2[9].wave_shpr.div.acc[18] ),
    .Y(_05705_));
 sky130_fd_sc_hd__nand2_1 _11871_ (.A(_05704_),
    .B(_05705_),
    .Y(_05706_));
 sky130_fd_sc_hd__a22o_1 _11872_ (.A1(net1023),
    .A2(_05684_),
    .B1(_05685_),
    .B2(_05706_),
    .X(_00910_));
 sky130_fd_sc_hd__or2_1 _11873_ (.A(\genblk2[9].wave_shpr.div.acc[19] ),
    .B(_05704_),
    .X(_05707_));
 sky130_fd_sc_hd__a21bo_1 _11874_ (.A1(\genblk2[9].wave_shpr.div.acc[19] ),
    .A2(_05608_),
    .B1_N(_05707_),
    .X(_05708_));
 sky130_fd_sc_hd__a22o_1 _11875_ (.A1(net935),
    .A2(_05684_),
    .B1(_05685_),
    .B2(_05708_),
    .X(_00911_));
 sky130_fd_sc_hd__or2_1 _11876_ (.A(\genblk2[9].wave_shpr.div.acc[20] ),
    .B(_05707_),
    .X(_05709_));
 sky130_fd_sc_hd__nand2_1 _11877_ (.A(\genblk2[9].wave_shpr.div.acc[20] ),
    .B(_05707_),
    .Y(_05710_));
 sky130_fd_sc_hd__nand2_1 _11878_ (.A(_05709_),
    .B(_05710_),
    .Y(_05711_));
 sky130_fd_sc_hd__a22o_1 _11879_ (.A1(net556),
    .A2(_05684_),
    .B1(_05685_),
    .B2(_05711_),
    .X(_00912_));
 sky130_fd_sc_hd__a2bb2o_1 _11880_ (.A1_N(_05609_),
    .A2_N(_05646_),
    .B1(_05709_),
    .B2(\genblk2[9].wave_shpr.div.acc[21] ),
    .X(_05712_));
 sky130_fd_sc_hd__a22o_1 _11881_ (.A1(net646),
    .A2(_05684_),
    .B1(_05685_),
    .B2(_05712_),
    .X(_00913_));
 sky130_fd_sc_hd__and2b_1 _11882_ (.A_N(_05610_),
    .B(_05611_),
    .X(_05713_));
 sky130_fd_sc_hd__a21o_1 _11883_ (.A1(net646),
    .A2(_05609_),
    .B1(_05713_),
    .X(_05714_));
 sky130_fd_sc_hd__a22o_1 _11884_ (.A1(net892),
    .A2(_03696_),
    .B1(_03694_),
    .B2(_05714_),
    .X(_00914_));
 sky130_fd_sc_hd__nor2_1 _11885_ (.A(\genblk2[9].wave_shpr.div.acc[23] ),
    .B(_05610_),
    .Y(_05715_));
 sky130_fd_sc_hd__and2_1 _11886_ (.A(\genblk2[9].wave_shpr.div.acc[23] ),
    .B(_05610_),
    .X(_05716_));
 sky130_fd_sc_hd__or2_1 _11887_ (.A(_05715_),
    .B(_05716_),
    .X(_05717_));
 sky130_fd_sc_hd__a32o_1 _11888_ (.A1(_03694_),
    .A2(_05611_),
    .A3(_05717_),
    .B1(_03696_),
    .B2(net1026),
    .X(_00915_));
 sky130_fd_sc_hd__inv_2 _11889_ (.A(\genblk2[9].wave_shpr.div.acc[24] ),
    .Y(_05718_));
 sky130_fd_sc_hd__or3b_1 _11890_ (.A(\genblk2[9].wave_shpr.div.acc[24] ),
    .B(_05646_),
    .C_N(_05715_),
    .X(_05719_));
 sky130_fd_sc_hd__o21ai_1 _11891_ (.A1(_05718_),
    .A2(_05715_),
    .B1(_05719_),
    .Y(_05720_));
 sky130_fd_sc_hd__a22o_1 _11892_ (.A1(net1045),
    .A2(_03696_),
    .B1(_03694_),
    .B2(_05720_),
    .X(_00916_));
 sky130_fd_sc_hd__xnor2_1 _11893_ (.A(\genblk2[9].wave_shpr.div.acc[25] ),
    .B(_05719_),
    .Y(_05721_));
 sky130_fd_sc_hd__a22o_1 _11894_ (.A1(net348),
    .A2(_03696_),
    .B1(_03694_),
    .B2(_05721_),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _11895_ (.A0(_03838_),
    .A1(_03835_),
    .S(\genblk2[0].wave_shpr.div.i[0] ),
    .X(_05722_));
 sky130_fd_sc_hd__clkbuf_1 _11896_ (.A(_05722_),
    .X(_00918_));
 sky130_fd_sc_hd__or2_1 _11897_ (.A(\genblk2[0].wave_shpr.div.i[1] ),
    .B(\genblk2[0].wave_shpr.div.i[0] ),
    .X(_05723_));
 sky130_fd_sc_hd__nand2_1 _11898_ (.A(\genblk2[0].wave_shpr.div.i[1] ),
    .B(\genblk2[0].wave_shpr.div.i[0] ),
    .Y(_05724_));
 sky130_fd_sc_hd__a32o_1 _11899_ (.A1(_03839_),
    .A2(_05723_),
    .A3(_05724_),
    .B1(_03841_),
    .B2(net1106),
    .X(_00919_));
 sky130_fd_sc_hd__a21o_1 _11900_ (.A1(\genblk2[0].wave_shpr.div.i[1] ),
    .A2(\genblk2[0].wave_shpr.div.i[0] ),
    .B1(\genblk2[0].wave_shpr.div.i[2] ),
    .X(_05725_));
 sky130_fd_sc_hd__and3_1 _11901_ (.A(\genblk2[0].wave_shpr.div.i[1] ),
    .B(\genblk2[0].wave_shpr.div.i[0] ),
    .C(\genblk2[0].wave_shpr.div.i[2] ),
    .X(_05726_));
 sky130_fd_sc_hd__inv_2 _11902_ (.A(_05726_),
    .Y(_05727_));
 sky130_fd_sc_hd__a32o_1 _11903_ (.A1(_03839_),
    .A2(_05725_),
    .A3(_05727_),
    .B1(_03841_),
    .B2(net775),
    .X(_00920_));
 sky130_fd_sc_hd__a21oi_1 _11904_ (.A1(_00000_),
    .A2(_05726_),
    .B1(net1158),
    .Y(_05728_));
 sky130_fd_sc_hd__and3_1 _11905_ (.A(\genblk2[0].wave_shpr.div.i[3] ),
    .B(_02150_),
    .C(_05726_),
    .X(_05729_));
 sky130_fd_sc_hd__nor3_1 _11906_ (.A(_03690_),
    .B(_05728_),
    .C(_05729_),
    .Y(_00921_));
 sky130_fd_sc_hd__o21ai_1 _11907_ (.A1(net273),
    .A2(_05729_),
    .B1(_03855_),
    .Y(_05730_));
 sky130_fd_sc_hd__a21oi_1 _11908_ (.A1(net273),
    .A2(_05729_),
    .B1(_05730_),
    .Y(_00922_));
 sky130_fd_sc_hd__or2b_1 _11909_ (.A(\genblk2[10].wave_shpr.div.acc[17] ),
    .B_N(\genblk2[10].wave_shpr.div.b1[17] ),
    .X(_05731_));
 sky130_fd_sc_hd__nor2_1 _11910_ (.A(_03832_),
    .B(\genblk2[10].wave_shpr.div.acc[16] ),
    .Y(_05732_));
 sky130_fd_sc_hd__or2b_1 _11911_ (.A(\genblk2[10].wave_shpr.div.acc[15] ),
    .B_N(\genblk2[10].wave_shpr.div.b1[15] ),
    .X(_05733_));
 sky130_fd_sc_hd__or2b_1 _11912_ (.A(\genblk2[10].wave_shpr.div.acc[14] ),
    .B_N(\genblk2[10].wave_shpr.div.b1[14] ),
    .X(_05734_));
 sky130_fd_sc_hd__or2b_1 _11913_ (.A(\genblk2[10].wave_shpr.div.acc[13] ),
    .B_N(\genblk2[10].wave_shpr.div.b1[13] ),
    .X(_05735_));
 sky130_fd_sc_hd__or2b_1 _11914_ (.A(\genblk2[10].wave_shpr.div.acc[12] ),
    .B_N(\genblk2[10].wave_shpr.div.b1[12] ),
    .X(_05736_));
 sky130_fd_sc_hd__or2b_1 _11915_ (.A(\genblk2[10].wave_shpr.div.acc[11] ),
    .B_N(\genblk2[10].wave_shpr.div.b1[11] ),
    .X(_05737_));
 sky130_fd_sc_hd__or2b_1 _11916_ (.A(\genblk2[10].wave_shpr.div.acc[10] ),
    .B_N(\genblk2[10].wave_shpr.div.b1[10] ),
    .X(_05738_));
 sky130_fd_sc_hd__or2b_1 _11917_ (.A(\genblk2[10].wave_shpr.div.acc[9] ),
    .B_N(\genblk2[10].wave_shpr.div.b1[9] ),
    .X(_05739_));
 sky130_fd_sc_hd__or2b_1 _11918_ (.A(\genblk2[10].wave_shpr.div.acc[8] ),
    .B_N(\genblk2[10].wave_shpr.div.b1[8] ),
    .X(_05740_));
 sky130_fd_sc_hd__or2b_1 _11919_ (.A(\genblk2[10].wave_shpr.div.acc[7] ),
    .B_N(\genblk2[10].wave_shpr.div.b1[7] ),
    .X(_05741_));
 sky130_fd_sc_hd__and2b_1 _11920_ (.A_N(\genblk2[10].wave_shpr.div.acc[5] ),
    .B(\genblk2[10].wave_shpr.div.b1[5] ),
    .X(_05742_));
 sky130_fd_sc_hd__and2b_1 _11921_ (.A_N(\genblk2[10].wave_shpr.div.acc[4] ),
    .B(\genblk2[10].wave_shpr.div.b1[4] ),
    .X(_05743_));
 sky130_fd_sc_hd__or2b_1 _11922_ (.A(\genblk2[10].wave_shpr.div.acc[3] ),
    .B_N(\genblk2[10].wave_shpr.div.b1[3] ),
    .X(_05744_));
 sky130_fd_sc_hd__or2b_1 _11923_ (.A(\genblk2[10].wave_shpr.div.acc[2] ),
    .B_N(\genblk2[10].wave_shpr.div.b1[2] ),
    .X(_05745_));
 sky130_fd_sc_hd__xnor2_1 _11924_ (.A(\genblk2[10].wave_shpr.div.acc[1] ),
    .B(\genblk2[10].wave_shpr.div.b1[1] ),
    .Y(_05746_));
 sky130_fd_sc_hd__or2b_1 _11925_ (.A(\genblk2[10].wave_shpr.div.acc[0] ),
    .B_N(\genblk2[10].wave_shpr.div.b1[0] ),
    .X(_05747_));
 sky130_fd_sc_hd__and2b_1 _11926_ (.A_N(\genblk2[10].wave_shpr.div.b1[1] ),
    .B(\genblk2[10].wave_shpr.div.acc[1] ),
    .X(_05748_));
 sky130_fd_sc_hd__a21o_1 _11927_ (.A1(_05746_),
    .A2(_05747_),
    .B1(_05748_),
    .X(_05749_));
 sky130_fd_sc_hd__and2b_1 _11928_ (.A_N(\genblk2[10].wave_shpr.div.b1[2] ),
    .B(\genblk2[10].wave_shpr.div.acc[2] ),
    .X(_05750_));
 sky130_fd_sc_hd__a21o_1 _11929_ (.A1(_05745_),
    .A2(_05749_),
    .B1(_05750_),
    .X(_05751_));
 sky130_fd_sc_hd__and2b_1 _11930_ (.A_N(\genblk2[10].wave_shpr.div.b1[3] ),
    .B(\genblk2[10].wave_shpr.div.acc[3] ),
    .X(_05752_));
 sky130_fd_sc_hd__a21oi_1 _11931_ (.A1(_05744_),
    .A2(_05751_),
    .B1(_05752_),
    .Y(_05753_));
 sky130_fd_sc_hd__and2b_1 _11932_ (.A_N(\genblk2[10].wave_shpr.div.b1[4] ),
    .B(\genblk2[10].wave_shpr.div.acc[4] ),
    .X(_05754_));
 sky130_fd_sc_hd__o21ba_1 _11933_ (.A1(_05743_),
    .A2(_05753_),
    .B1_N(_05754_),
    .X(_05755_));
 sky130_fd_sc_hd__and2b_1 _11934_ (.A_N(\genblk2[10].wave_shpr.div.b1[5] ),
    .B(\genblk2[10].wave_shpr.div.acc[5] ),
    .X(_05756_));
 sky130_fd_sc_hd__o21bai_1 _11935_ (.A1(_05742_),
    .A2(_05755_),
    .B1_N(_05756_),
    .Y(_05757_));
 sky130_fd_sc_hd__o21a_1 _11936_ (.A1(_03821_),
    .A2(\genblk2[10].wave_shpr.div.acc[6] ),
    .B1(_05757_),
    .X(_05758_));
 sky130_fd_sc_hd__a21o_1 _11937_ (.A1(_03821_),
    .A2(\genblk2[10].wave_shpr.div.acc[6] ),
    .B1(_05758_),
    .X(_05759_));
 sky130_fd_sc_hd__and2b_1 _11938_ (.A_N(\genblk2[10].wave_shpr.div.b1[7] ),
    .B(\genblk2[10].wave_shpr.div.acc[7] ),
    .X(_05760_));
 sky130_fd_sc_hd__a21o_1 _11939_ (.A1(_05741_),
    .A2(_05759_),
    .B1(_05760_),
    .X(_05761_));
 sky130_fd_sc_hd__and2b_1 _11940_ (.A_N(\genblk2[10].wave_shpr.div.b1[8] ),
    .B(\genblk2[10].wave_shpr.div.acc[8] ),
    .X(_05762_));
 sky130_fd_sc_hd__a21o_1 _11941_ (.A1(_05740_),
    .A2(_05761_),
    .B1(_05762_),
    .X(_05763_));
 sky130_fd_sc_hd__and2b_1 _11942_ (.A_N(\genblk2[10].wave_shpr.div.b1[9] ),
    .B(\genblk2[10].wave_shpr.div.acc[9] ),
    .X(_05764_));
 sky130_fd_sc_hd__a21o_1 _11943_ (.A1(_05739_),
    .A2(_05763_),
    .B1(_05764_),
    .X(_05765_));
 sky130_fd_sc_hd__and2b_1 _11944_ (.A_N(\genblk2[10].wave_shpr.div.b1[10] ),
    .B(\genblk2[10].wave_shpr.div.acc[10] ),
    .X(_05766_));
 sky130_fd_sc_hd__a21o_1 _11945_ (.A1(_05738_),
    .A2(_05765_),
    .B1(_05766_),
    .X(_05767_));
 sky130_fd_sc_hd__and2b_1 _11946_ (.A_N(\genblk2[10].wave_shpr.div.b1[11] ),
    .B(\genblk2[10].wave_shpr.div.acc[11] ),
    .X(_05768_));
 sky130_fd_sc_hd__a21o_1 _11947_ (.A1(_05737_),
    .A2(_05767_),
    .B1(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__and2b_1 _11948_ (.A_N(\genblk2[10].wave_shpr.div.b1[12] ),
    .B(\genblk2[10].wave_shpr.div.acc[12] ),
    .X(_05770_));
 sky130_fd_sc_hd__a21o_1 _11949_ (.A1(_05736_),
    .A2(_05769_),
    .B1(_05770_),
    .X(_05771_));
 sky130_fd_sc_hd__and2b_1 _11950_ (.A_N(\genblk2[10].wave_shpr.div.b1[13] ),
    .B(\genblk2[10].wave_shpr.div.acc[13] ),
    .X(_05772_));
 sky130_fd_sc_hd__a21o_1 _11951_ (.A1(_05735_),
    .A2(_05771_),
    .B1(_05772_),
    .X(_05773_));
 sky130_fd_sc_hd__and2b_1 _11952_ (.A_N(\genblk2[10].wave_shpr.div.b1[14] ),
    .B(\genblk2[10].wave_shpr.div.acc[14] ),
    .X(_05774_));
 sky130_fd_sc_hd__a21o_1 _11953_ (.A1(_05734_),
    .A2(_05773_),
    .B1(_05774_),
    .X(_05775_));
 sky130_fd_sc_hd__and2b_1 _11954_ (.A_N(\genblk2[10].wave_shpr.div.b1[15] ),
    .B(\genblk2[10].wave_shpr.div.acc[15] ),
    .X(_05776_));
 sky130_fd_sc_hd__a21oi_1 _11955_ (.A1(_05733_),
    .A2(_05775_),
    .B1(_05776_),
    .Y(_05777_));
 sky130_fd_sc_hd__and2_1 _11956_ (.A(_03832_),
    .B(\genblk2[10].wave_shpr.div.acc[16] ),
    .X(_05778_));
 sky130_fd_sc_hd__o21bai_1 _11957_ (.A1(_05732_),
    .A2(_05777_),
    .B1_N(_05778_),
    .Y(_05779_));
 sky130_fd_sc_hd__and2b_1 _11958_ (.A_N(\genblk2[10].wave_shpr.div.b1[17] ),
    .B(\genblk2[10].wave_shpr.div.acc[17] ),
    .X(_05780_));
 sky130_fd_sc_hd__a21o_1 _11959_ (.A1(_05731_),
    .A2(_05779_),
    .B1(_05780_),
    .X(_05781_));
 sky130_fd_sc_hd__or2_1 _11960_ (.A(\genblk2[10].wave_shpr.div.acc[18] ),
    .B(_05781_),
    .X(_05782_));
 sky130_fd_sc_hd__or3_1 _11961_ (.A(\genblk2[10].wave_shpr.div.acc[20] ),
    .B(\genblk2[10].wave_shpr.div.acc[19] ),
    .C(_05782_),
    .X(_05783_));
 sky130_fd_sc_hd__or4_1 _11962_ (.A(\genblk2[10].wave_shpr.div.acc[23] ),
    .B(\genblk2[10].wave_shpr.div.acc[22] ),
    .C(\genblk2[10].wave_shpr.div.acc[21] ),
    .D(_05783_),
    .X(_05784_));
 sky130_fd_sc_hd__or2_2 _11963_ (.A(\genblk2[10].wave_shpr.div.acc[24] ),
    .B(_05784_),
    .X(_05785_));
 sky130_fd_sc_hd__or3_2 _11964_ (.A(\genblk2[10].wave_shpr.div.acc[25] ),
    .B(\genblk2[10].wave_shpr.div.acc[26] ),
    .C(_05785_),
    .X(_05786_));
 sky130_fd_sc_hd__clkbuf_8 _11965_ (.A(_05786_),
    .X(_05787_));
 sky130_fd_sc_hd__mux2_1 _11966_ (.A0(\genblk2[10].wave_shpr.div.fin_quo[0] ),
    .A1(_05787_),
    .S(_00003_),
    .X(_05788_));
 sky130_fd_sc_hd__clkbuf_1 _11967_ (.A(_05788_),
    .X(_00923_));
 sky130_fd_sc_hd__mux2_1 _11968_ (.A0(\genblk2[10].wave_shpr.div.fin_quo[1] ),
    .A1(\genblk2[10].wave_shpr.div.quo[0] ),
    .S(_00003_),
    .X(_05789_));
 sky130_fd_sc_hd__clkbuf_1 _11969_ (.A(_05789_),
    .X(_00924_));
 sky130_fd_sc_hd__mux2_1 _11970_ (.A0(\genblk2[10].wave_shpr.div.fin_quo[2] ),
    .A1(net220),
    .S(_00003_),
    .X(_05790_));
 sky130_fd_sc_hd__clkbuf_1 _11971_ (.A(_05790_),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _11972_ (.A0(\genblk2[10].wave_shpr.div.fin_quo[3] ),
    .A1(\genblk2[10].wave_shpr.div.quo[2] ),
    .S(_00003_),
    .X(_05791_));
 sky130_fd_sc_hd__clkbuf_1 _11973_ (.A(_05791_),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _11974_ (.A0(\genblk2[10].wave_shpr.div.fin_quo[4] ),
    .A1(net1323),
    .S(_00003_),
    .X(_05792_));
 sky130_fd_sc_hd__clkbuf_1 _11975_ (.A(_05792_),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _11976_ (.A0(\genblk2[10].wave_shpr.div.fin_quo[5] ),
    .A1(\genblk2[10].wave_shpr.div.quo[4] ),
    .S(_00003_),
    .X(_05793_));
 sky130_fd_sc_hd__clkbuf_1 _11977_ (.A(_05793_),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _11978_ (.A0(\genblk2[10].wave_shpr.div.fin_quo[6] ),
    .A1(net1324),
    .S(_00003_),
    .X(_05794_));
 sky130_fd_sc_hd__clkbuf_1 _11979_ (.A(_05794_),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _11980_ (.A0(\genblk2[10].wave_shpr.div.fin_quo[7] ),
    .A1(\genblk2[10].wave_shpr.div.quo[6] ),
    .S(_00003_),
    .X(_05795_));
 sky130_fd_sc_hd__clkbuf_1 _11981_ (.A(_05795_),
    .X(_00930_));
 sky130_fd_sc_hd__o21ai_4 _11982_ (.A1(_01441_),
    .A2(_01320_),
    .B1(_03702_),
    .Y(_05796_));
 sky130_fd_sc_hd__o21a_1 _11983_ (.A1(_03732_),
    .A2(net1007),
    .B1(_05796_),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _11984_ (.A0(\genblk2[11].wave_shpr.div.b1[1] ),
    .A1(_03813_),
    .S(_05433_),
    .X(_05797_));
 sky130_fd_sc_hd__clkbuf_1 _11985_ (.A(_05797_),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _11986_ (.A0(\genblk2[11].wave_shpr.div.b1[2] ),
    .A1(_01811_),
    .S(_05433_),
    .X(_05798_));
 sky130_fd_sc_hd__clkbuf_1 _11987_ (.A(_05798_),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _11988_ (.A0(net1265),
    .A1(_01946_),
    .S(_05433_),
    .X(_05799_));
 sky130_fd_sc_hd__clkbuf_1 _11989_ (.A(_05799_),
    .X(_00934_));
 sky130_fd_sc_hd__mux2_1 _11990_ (.A0(\genblk2[11].wave_shpr.div.b1[4] ),
    .A1(_04230_),
    .S(_05433_),
    .X(_05800_));
 sky130_fd_sc_hd__clkbuf_1 _11991_ (.A(_05800_),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_1 _11992_ (.A0(\genblk2[11].wave_shpr.div.b1[5] ),
    .A1(_01855_),
    .S(_05433_),
    .X(_05801_));
 sky130_fd_sc_hd__clkbuf_1 _11993_ (.A(_05801_),
    .X(_00936_));
 sky130_fd_sc_hd__clkbuf_8 _11994_ (.A(_03707_),
    .X(_05802_));
 sky130_fd_sc_hd__mux2_1 _11995_ (.A0(net1242),
    .A1(_02805_),
    .S(_05802_),
    .X(_05803_));
 sky130_fd_sc_hd__clkbuf_1 _11996_ (.A(_05803_),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _11997_ (.A0(net1275),
    .A1(_01556_),
    .S(_05802_),
    .X(_05804_));
 sky130_fd_sc_hd__clkbuf_1 _11998_ (.A(_05804_),
    .X(_00938_));
 sky130_fd_sc_hd__a21bo_1 _11999_ (.A1(_03687_),
    .A2(net420),
    .B1_N(_03705_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _12000_ (.A0(net1217),
    .A1(_03706_),
    .S(_05802_),
    .X(_05805_));
 sky130_fd_sc_hd__clkbuf_1 _12001_ (.A(_05805_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _12002_ (.A0(net1204),
    .A1(_02002_),
    .S(_05802_),
    .X(_05806_));
 sky130_fd_sc_hd__clkbuf_1 _12003_ (.A(_05806_),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _12004_ (.A0(\genblk2[11].wave_shpr.div.b1[11] ),
    .A1(_01500_),
    .S(_05802_),
    .X(_05807_));
 sky130_fd_sc_hd__clkbuf_1 _12005_ (.A(_05807_),
    .X(_00942_));
 sky130_fd_sc_hd__mux2_1 _12006_ (.A0(\genblk2[11].wave_shpr.div.b1[12] ),
    .A1(_01494_),
    .S(_05802_),
    .X(_05808_));
 sky130_fd_sc_hd__clkbuf_1 _12007_ (.A(_05808_),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _12008_ (.A0(\genblk2[11].wave_shpr.div.b1[13] ),
    .A1(_01483_),
    .S(_05802_),
    .X(_05809_));
 sky130_fd_sc_hd__clkbuf_1 _12009_ (.A(_05809_),
    .X(_00944_));
 sky130_fd_sc_hd__o21a_1 _12010_ (.A1(_03732_),
    .A2(net384),
    .B1(_03733_),
    .X(_00945_));
 sky130_fd_sc_hd__a21bo_1 _12011_ (.A1(_03687_),
    .A2(net424),
    .B1_N(_03717_),
    .X(_00946_));
 sky130_fd_sc_hd__inv_2 _12012_ (.A(net1086),
    .Y(_05810_));
 sky130_fd_sc_hd__o21ai_1 _12013_ (.A1(_03726_),
    .A2(_05810_),
    .B1(_03735_),
    .Y(_00947_));
 sky130_fd_sc_hd__and2_1 _12014_ (.A(_02171_),
    .B(net1278),
    .X(_05811_));
 sky130_fd_sc_hd__clkbuf_1 _12015_ (.A(_05811_),
    .X(_00948_));
 sky130_fd_sc_hd__clkbuf_4 _12016_ (.A(_02208_),
    .X(_05812_));
 sky130_fd_sc_hd__buf_4 _12017_ (.A(_05812_),
    .X(_05813_));
 sky130_fd_sc_hd__and3_1 _12018_ (.A(_02152_),
    .B(\genblk2[10].wave_shpr.div.busy ),
    .C(_02206_),
    .X(_05814_));
 sky130_fd_sc_hd__clkbuf_4 _12019_ (.A(_05814_),
    .X(_05815_));
 sky130_fd_sc_hd__buf_4 _12020_ (.A(_05815_),
    .X(_05816_));
 sky130_fd_sc_hd__a22o_1 _12021_ (.A1(\genblk2[10].wave_shpr.div.quo[0] ),
    .A2(_05813_),
    .B1(_05787_),
    .B2(_05816_),
    .X(_00949_));
 sky130_fd_sc_hd__buf_4 _12022_ (.A(_05815_),
    .X(_05817_));
 sky130_fd_sc_hd__a22o_1 _12023_ (.A1(net220),
    .A2(_05813_),
    .B1(_05817_),
    .B2(net740),
    .X(_00950_));
 sky130_fd_sc_hd__a22o_1 _12024_ (.A1(\genblk2[10].wave_shpr.div.quo[2] ),
    .A2(_05813_),
    .B1(_05817_),
    .B2(net220),
    .X(_00951_));
 sky130_fd_sc_hd__a22o_1 _12025_ (.A1(net682),
    .A2(_05813_),
    .B1(_05817_),
    .B2(net724),
    .X(_00952_));
 sky130_fd_sc_hd__a22o_1 _12026_ (.A1(\genblk2[10].wave_shpr.div.quo[4] ),
    .A2(_05813_),
    .B1(_05817_),
    .B2(net682),
    .X(_00953_));
 sky130_fd_sc_hd__a22o_1 _12027_ (.A1(net555),
    .A2(_05813_),
    .B1(_05817_),
    .B2(net723),
    .X(_00954_));
 sky130_fd_sc_hd__a22o_1 _12028_ (.A1(\genblk2[10].wave_shpr.div.quo[6] ),
    .A2(_05813_),
    .B1(_05817_),
    .B2(net555),
    .X(_00955_));
 sky130_fd_sc_hd__a22o_1 _12029_ (.A1(net320),
    .A2(_05813_),
    .B1(_05817_),
    .B2(\genblk2[10].wave_shpr.div.quo[6] ),
    .X(_00956_));
 sky130_fd_sc_hd__a22o_1 _12030_ (.A1(\genblk2[10].wave_shpr.div.quo[8] ),
    .A2(_05813_),
    .B1(_05817_),
    .B2(net320),
    .X(_00957_));
 sky130_fd_sc_hd__clkbuf_4 _12031_ (.A(_05812_),
    .X(_05818_));
 sky130_fd_sc_hd__clkbuf_2 _12032_ (.A(_02155_),
    .X(_05819_));
 sky130_fd_sc_hd__and2_1 _12033_ (.A(_05819_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[0] ),
    .X(_05820_));
 sky130_fd_sc_hd__a221o_1 _12034_ (.A1(net432),
    .A2(_05818_),
    .B1(_05816_),
    .B2(\genblk2[10].wave_shpr.div.quo[8] ),
    .C1(_05820_),
    .X(_00958_));
 sky130_fd_sc_hd__and2_1 _12035_ (.A(_05819_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[1] ),
    .X(_05821_));
 sky130_fd_sc_hd__a221o_1 _12036_ (.A1(net398),
    .A2(_05818_),
    .B1(_05816_),
    .B2(net432),
    .C1(_05821_),
    .X(_00959_));
 sky130_fd_sc_hd__and2_1 _12037_ (.A(_05819_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[2] ),
    .X(_05822_));
 sky130_fd_sc_hd__a221o_1 _12038_ (.A1(net223),
    .A2(_05818_),
    .B1(_05816_),
    .B2(net398),
    .C1(_05822_),
    .X(_00960_));
 sky130_fd_sc_hd__clkbuf_4 _12039_ (.A(_05812_),
    .X(_05823_));
 sky130_fd_sc_hd__and2_1 _12040_ (.A(_05819_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[3] ),
    .X(_05824_));
 sky130_fd_sc_hd__a221o_1 _12041_ (.A1(\genblk2[10].wave_shpr.div.quo[12] ),
    .A2(_05823_),
    .B1(_05816_),
    .B2(net223),
    .C1(_05824_),
    .X(_00961_));
 sky130_fd_sc_hd__clkbuf_4 _12042_ (.A(_05815_),
    .X(_05825_));
 sky130_fd_sc_hd__nor2_1 _12043_ (.A(_04676_),
    .B(_01993_),
    .Y(_05826_));
 sky130_fd_sc_hd__a221o_1 _12044_ (.A1(net521),
    .A2(_05823_),
    .B1(_05825_),
    .B2(net583),
    .C1(_05826_),
    .X(_00962_));
 sky130_fd_sc_hd__and2_1 _12045_ (.A(_05819_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[5] ),
    .X(_05827_));
 sky130_fd_sc_hd__a221o_1 _12046_ (.A1(net373),
    .A2(_05823_),
    .B1(_05825_),
    .B2(net521),
    .C1(_05827_),
    .X(_00963_));
 sky130_fd_sc_hd__and2_1 _12047_ (.A(_05819_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[6] ),
    .X(_05828_));
 sky130_fd_sc_hd__a221o_1 _12048_ (.A1(net357),
    .A2(_05823_),
    .B1(_05825_),
    .B2(net373),
    .C1(_05828_),
    .X(_00964_));
 sky130_fd_sc_hd__and2_1 _12049_ (.A(_05819_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[7] ),
    .X(_05829_));
 sky130_fd_sc_hd__a221o_1 _12050_ (.A1(net353),
    .A2(_05823_),
    .B1(_05825_),
    .B2(net357),
    .C1(_05829_),
    .X(_00965_));
 sky130_fd_sc_hd__nor2_1 _12051_ (.A(_03833_),
    .B(_02003_),
    .Y(_05830_));
 sky130_fd_sc_hd__a221o_1 _12052_ (.A1(\genblk2[10].wave_shpr.div.quo[17] ),
    .A2(_05823_),
    .B1(_05825_),
    .B2(net353),
    .C1(_05830_),
    .X(_00966_));
 sky130_fd_sc_hd__and2_1 _12053_ (.A(_05819_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[9] ),
    .X(_05831_));
 sky130_fd_sc_hd__a221o_1 _12054_ (.A1(net518),
    .A2(_05823_),
    .B1(_05825_),
    .B2(net547),
    .C1(_05831_),
    .X(_00967_));
 sky130_fd_sc_hd__and2_1 _12055_ (.A(_05819_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[10] ),
    .X(_05832_));
 sky130_fd_sc_hd__a221o_1 _12056_ (.A1(net440),
    .A2(_05823_),
    .B1(_05825_),
    .B2(net518),
    .C1(_05832_),
    .X(_00968_));
 sky130_fd_sc_hd__and2_1 _12057_ (.A(_05819_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[11] ),
    .X(_05833_));
 sky130_fd_sc_hd__a221o_1 _12058_ (.A1(net383),
    .A2(_05823_),
    .B1(_05825_),
    .B2(net440),
    .C1(_05833_),
    .X(_00969_));
 sky130_fd_sc_hd__nor2_1 _12059_ (.A(_03833_),
    .B(_02023_),
    .Y(_05834_));
 sky130_fd_sc_hd__a221o_1 _12060_ (.A1(net334),
    .A2(_05823_),
    .B1(_05825_),
    .B2(net383),
    .C1(_05834_),
    .X(_00970_));
 sky130_fd_sc_hd__clkbuf_2 _12061_ (.A(_02155_),
    .X(_05835_));
 sky130_fd_sc_hd__and2_1 _12062_ (.A(_05835_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[13] ),
    .X(_05836_));
 sky130_fd_sc_hd__a221o_1 _12063_ (.A1(\genblk2[10].wave_shpr.div.quo[22] ),
    .A2(_05812_),
    .B1(_05825_),
    .B2(net334),
    .C1(_05836_),
    .X(_00971_));
 sky130_fd_sc_hd__nor2_1 _12064_ (.A(_03833_),
    .B(_01995_),
    .Y(_05837_));
 sky130_fd_sc_hd__a221o_1 _12065_ (.A1(\genblk2[10].wave_shpr.div.quo[23] ),
    .A2(_05812_),
    .B1(_05815_),
    .B2(net474),
    .C1(_05837_),
    .X(_00972_));
 sky130_fd_sc_hd__and2_1 _12066_ (.A(_05835_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[15] ),
    .X(_05838_));
 sky130_fd_sc_hd__a221o_1 _12067_ (.A1(net446),
    .A2(_05812_),
    .B1(_05815_),
    .B2(\genblk2[10].wave_shpr.div.quo[23] ),
    .C1(_05838_),
    .X(_00973_));
 sky130_fd_sc_hd__and2_1 _12068_ (.A(_05835_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[16] ),
    .X(_05839_));
 sky130_fd_sc_hd__a221o_1 _12069_ (.A1(net247),
    .A2(_05812_),
    .B1(_05815_),
    .B2(net446),
    .C1(_05839_),
    .X(_00974_));
 sky130_fd_sc_hd__inv_2 _12070_ (.A(_05815_),
    .Y(_05840_));
 sky130_fd_sc_hd__or2_1 _12071_ (.A(_03719_),
    .B(\genblk1[10].osc.clkdiv_C.cnt[17] ),
    .X(_05841_));
 sky130_fd_sc_hd__o221a_1 _12072_ (.A1(\genblk2[10].wave_shpr.div.acc[0] ),
    .A2(_00002_),
    .B1(_05840_),
    .B2(net247),
    .C1(_05841_),
    .X(_00975_));
 sky130_fd_sc_hd__a21oi_1 _12073_ (.A1(\genblk2[10].wave_shpr.div.b1[0] ),
    .A2(_05787_),
    .B1(\genblk2[10].wave_shpr.div.acc[0] ),
    .Y(_05842_));
 sky130_fd_sc_hd__a31o_1 _12074_ (.A1(\genblk2[10].wave_shpr.div.b1[0] ),
    .A2(\genblk2[10].wave_shpr.div.acc[0] ),
    .A3(_05787_),
    .B1(_05840_),
    .X(_05843_));
 sky130_fd_sc_hd__a2bb2o_1 _12075_ (.A1_N(_05842_),
    .A2_N(_05843_),
    .B1(net1118),
    .B2(_05813_),
    .X(_00976_));
 sky130_fd_sc_hd__clkbuf_4 _12076_ (.A(_05812_),
    .X(_05844_));
 sky130_fd_sc_hd__xor2_1 _12077_ (.A(_05746_),
    .B(_05747_),
    .X(_05845_));
 sky130_fd_sc_hd__mux2_1 _12078_ (.A0(\genblk2[10].wave_shpr.div.acc[1] ),
    .A1(_05845_),
    .S(_05787_),
    .X(_05846_));
 sky130_fd_sc_hd__a22o_1 _12079_ (.A1(net989),
    .A2(_05844_),
    .B1(_05817_),
    .B2(_05846_),
    .X(_00977_));
 sky130_fd_sc_hd__or2b_1 _12080_ (.A(_05750_),
    .B_N(_05745_),
    .X(_05847_));
 sky130_fd_sc_hd__xnor2_1 _12081_ (.A(_05749_),
    .B(_05847_),
    .Y(_05848_));
 sky130_fd_sc_hd__mux2_1 _12082_ (.A0(\genblk2[10].wave_shpr.div.acc[2] ),
    .A1(_05848_),
    .S(_05787_),
    .X(_05849_));
 sky130_fd_sc_hd__a22o_1 _12083_ (.A1(net969),
    .A2(_05844_),
    .B1(_05817_),
    .B2(_05849_),
    .X(_00978_));
 sky130_fd_sc_hd__clkbuf_4 _12084_ (.A(_05815_),
    .X(_05850_));
 sky130_fd_sc_hd__or2b_1 _12085_ (.A(_05752_),
    .B_N(_05744_),
    .X(_05851_));
 sky130_fd_sc_hd__xnor2_1 _12086_ (.A(_05751_),
    .B(_05851_),
    .Y(_05852_));
 sky130_fd_sc_hd__mux2_1 _12087_ (.A0(\genblk2[10].wave_shpr.div.acc[3] ),
    .A1(_05852_),
    .S(_05787_),
    .X(_05853_));
 sky130_fd_sc_hd__a22o_1 _12088_ (.A1(net868),
    .A2(_05844_),
    .B1(_05850_),
    .B2(_05853_),
    .X(_00979_));
 sky130_fd_sc_hd__nor2_1 _12089_ (.A(_05754_),
    .B(_05743_),
    .Y(_05854_));
 sky130_fd_sc_hd__xnor2_1 _12090_ (.A(_05854_),
    .B(_05753_),
    .Y(_05855_));
 sky130_fd_sc_hd__mux2_1 _12091_ (.A0(\genblk2[10].wave_shpr.div.acc[4] ),
    .A1(_05855_),
    .S(_05787_),
    .X(_05856_));
 sky130_fd_sc_hd__a22o_1 _12092_ (.A1(net977),
    .A2(_05844_),
    .B1(_05850_),
    .B2(_05856_),
    .X(_00980_));
 sky130_fd_sc_hd__nor2_1 _12093_ (.A(_05756_),
    .B(_05742_),
    .Y(_05857_));
 sky130_fd_sc_hd__xnor2_1 _12094_ (.A(_05857_),
    .B(_05755_),
    .Y(_05858_));
 sky130_fd_sc_hd__mux2_1 _12095_ (.A0(\genblk2[10].wave_shpr.div.acc[5] ),
    .A1(_05858_),
    .S(_05787_),
    .X(_05859_));
 sky130_fd_sc_hd__a22o_1 _12096_ (.A1(net1241),
    .A2(_05844_),
    .B1(_05850_),
    .B2(_05859_),
    .X(_00981_));
 sky130_fd_sc_hd__xor2_1 _12097_ (.A(\genblk2[10].wave_shpr.div.b1[6] ),
    .B(\genblk2[10].wave_shpr.div.acc[6] ),
    .X(_05860_));
 sky130_fd_sc_hd__xnor2_1 _12098_ (.A(_05757_),
    .B(_05860_),
    .Y(_05861_));
 sky130_fd_sc_hd__mux2_1 _12099_ (.A0(\genblk2[10].wave_shpr.div.acc[6] ),
    .A1(_05861_),
    .S(_05787_),
    .X(_05862_));
 sky130_fd_sc_hd__a22o_1 _12100_ (.A1(net929),
    .A2(_05844_),
    .B1(_05850_),
    .B2(_05862_),
    .X(_00982_));
 sky130_fd_sc_hd__or2b_1 _12101_ (.A(_05760_),
    .B_N(_05741_),
    .X(_05863_));
 sky130_fd_sc_hd__xnor2_1 _12102_ (.A(_05759_),
    .B(_05863_),
    .Y(_05864_));
 sky130_fd_sc_hd__buf_4 _12103_ (.A(_05786_),
    .X(_05865_));
 sky130_fd_sc_hd__mux2_1 _12104_ (.A0(\genblk2[10].wave_shpr.div.acc[7] ),
    .A1(_05864_),
    .S(_05865_),
    .X(_05866_));
 sky130_fd_sc_hd__a22o_1 _12105_ (.A1(net954),
    .A2(_05844_),
    .B1(_05850_),
    .B2(_05866_),
    .X(_00983_));
 sky130_fd_sc_hd__or2b_1 _12106_ (.A(_05762_),
    .B_N(_05740_),
    .X(_05867_));
 sky130_fd_sc_hd__xnor2_1 _12107_ (.A(_05761_),
    .B(_05867_),
    .Y(_05868_));
 sky130_fd_sc_hd__mux2_1 _12108_ (.A0(\genblk2[10].wave_shpr.div.acc[8] ),
    .A1(_05868_),
    .S(_05865_),
    .X(_05869_));
 sky130_fd_sc_hd__a22o_1 _12109_ (.A1(net1035),
    .A2(_05844_),
    .B1(_05850_),
    .B2(_05869_),
    .X(_00984_));
 sky130_fd_sc_hd__or2b_1 _12110_ (.A(_05764_),
    .B_N(_05739_),
    .X(_05870_));
 sky130_fd_sc_hd__xnor2_1 _12111_ (.A(_05763_),
    .B(_05870_),
    .Y(_05871_));
 sky130_fd_sc_hd__mux2_1 _12112_ (.A0(\genblk2[10].wave_shpr.div.acc[9] ),
    .A1(_05871_),
    .S(_05865_),
    .X(_05872_));
 sky130_fd_sc_hd__a22o_1 _12113_ (.A1(net951),
    .A2(_05844_),
    .B1(_05850_),
    .B2(_05872_),
    .X(_00985_));
 sky130_fd_sc_hd__or2b_1 _12114_ (.A(_05766_),
    .B_N(_05738_),
    .X(_05873_));
 sky130_fd_sc_hd__xnor2_1 _12115_ (.A(_05765_),
    .B(_05873_),
    .Y(_05874_));
 sky130_fd_sc_hd__mux2_1 _12116_ (.A0(\genblk2[10].wave_shpr.div.acc[10] ),
    .A1(_05874_),
    .S(_05865_),
    .X(_05875_));
 sky130_fd_sc_hd__a22o_1 _12117_ (.A1(net844),
    .A2(_05844_),
    .B1(_05850_),
    .B2(_05875_),
    .X(_00986_));
 sky130_fd_sc_hd__clkbuf_4 _12118_ (.A(_05812_),
    .X(_05876_));
 sky130_fd_sc_hd__or2b_1 _12119_ (.A(_05768_),
    .B_N(_05737_),
    .X(_05877_));
 sky130_fd_sc_hd__xnor2_1 _12120_ (.A(_05767_),
    .B(_05877_),
    .Y(_05878_));
 sky130_fd_sc_hd__mux2_1 _12121_ (.A0(\genblk2[10].wave_shpr.div.acc[11] ),
    .A1(_05878_),
    .S(_05865_),
    .X(_05879_));
 sky130_fd_sc_hd__a22o_1 _12122_ (.A1(net957),
    .A2(_05876_),
    .B1(_05850_),
    .B2(_05879_),
    .X(_00987_));
 sky130_fd_sc_hd__or2b_1 _12123_ (.A(_05770_),
    .B_N(_05736_),
    .X(_05880_));
 sky130_fd_sc_hd__xnor2_1 _12124_ (.A(_05769_),
    .B(_05880_),
    .Y(_05881_));
 sky130_fd_sc_hd__mux2_1 _12125_ (.A0(\genblk2[10].wave_shpr.div.acc[12] ),
    .A1(_05881_),
    .S(_05865_),
    .X(_05882_));
 sky130_fd_sc_hd__a22o_1 _12126_ (.A1(net858),
    .A2(_05876_),
    .B1(_05850_),
    .B2(_05882_),
    .X(_00988_));
 sky130_fd_sc_hd__clkbuf_4 _12127_ (.A(_05815_),
    .X(_05883_));
 sky130_fd_sc_hd__or2b_1 _12128_ (.A(_05772_),
    .B_N(_05735_),
    .X(_05884_));
 sky130_fd_sc_hd__xnor2_1 _12129_ (.A(_05771_),
    .B(_05884_),
    .Y(_05885_));
 sky130_fd_sc_hd__mux2_1 _12130_ (.A0(\genblk2[10].wave_shpr.div.acc[13] ),
    .A1(_05885_),
    .S(_05865_),
    .X(_05886_));
 sky130_fd_sc_hd__a22o_1 _12131_ (.A1(net945),
    .A2(_05876_),
    .B1(_05883_),
    .B2(_05886_),
    .X(_00989_));
 sky130_fd_sc_hd__or2b_1 _12132_ (.A(_05774_),
    .B_N(_05734_),
    .X(_05887_));
 sky130_fd_sc_hd__xnor2_1 _12133_ (.A(_05773_),
    .B(_05887_),
    .Y(_05888_));
 sky130_fd_sc_hd__mux2_1 _12134_ (.A0(\genblk2[10].wave_shpr.div.acc[14] ),
    .A1(_05888_),
    .S(_05865_),
    .X(_05889_));
 sky130_fd_sc_hd__a22o_1 _12135_ (.A1(net944),
    .A2(_05876_),
    .B1(_05883_),
    .B2(_05889_),
    .X(_00990_));
 sky130_fd_sc_hd__or2b_1 _12136_ (.A(_05776_),
    .B_N(_05733_),
    .X(_05890_));
 sky130_fd_sc_hd__xnor2_1 _12137_ (.A(_05775_),
    .B(_05890_),
    .Y(_05891_));
 sky130_fd_sc_hd__mux2_1 _12138_ (.A0(\genblk2[10].wave_shpr.div.acc[15] ),
    .A1(_05891_),
    .S(_05865_),
    .X(_05892_));
 sky130_fd_sc_hd__a22o_1 _12139_ (.A1(net870),
    .A2(_05876_),
    .B1(_05883_),
    .B2(_05892_),
    .X(_00991_));
 sky130_fd_sc_hd__nor2_1 _12140_ (.A(_05778_),
    .B(_05732_),
    .Y(_05893_));
 sky130_fd_sc_hd__xnor2_1 _12141_ (.A(_05893_),
    .B(_05777_),
    .Y(_05894_));
 sky130_fd_sc_hd__mux2_1 _12142_ (.A0(\genblk2[10].wave_shpr.div.acc[16] ),
    .A1(_05894_),
    .S(_05865_),
    .X(_05895_));
 sky130_fd_sc_hd__a22o_1 _12143_ (.A1(net859),
    .A2(_05876_),
    .B1(_05883_),
    .B2(_05895_),
    .X(_00992_));
 sky130_fd_sc_hd__or2b_1 _12144_ (.A(_05780_),
    .B_N(_05731_),
    .X(_05896_));
 sky130_fd_sc_hd__xnor2_1 _12145_ (.A(_05779_),
    .B(_05896_),
    .Y(_05897_));
 sky130_fd_sc_hd__mux2_1 _12146_ (.A0(\genblk2[10].wave_shpr.div.acc[17] ),
    .A1(_05897_),
    .S(_05786_),
    .X(_05898_));
 sky130_fd_sc_hd__a22o_1 _12147_ (.A1(net590),
    .A2(_05876_),
    .B1(_05883_),
    .B2(_05898_),
    .X(_00993_));
 sky130_fd_sc_hd__nor3_2 _12148_ (.A(\genblk2[10].wave_shpr.div.acc[25] ),
    .B(\genblk2[10].wave_shpr.div.acc[26] ),
    .C(_05785_),
    .Y(_05899_));
 sky130_fd_sc_hd__or2_1 _12149_ (.A(_05782_),
    .B(_05899_),
    .X(_05900_));
 sky130_fd_sc_hd__o21ai_1 _12150_ (.A1(_05781_),
    .A2(_05899_),
    .B1(\genblk2[10].wave_shpr.div.acc[18] ),
    .Y(_05901_));
 sky130_fd_sc_hd__nand2_1 _12151_ (.A(_05900_),
    .B(_05901_),
    .Y(_05902_));
 sky130_fd_sc_hd__a22o_1 _12152_ (.A1(net1135),
    .A2(_05876_),
    .B1(_05883_),
    .B2(_05902_),
    .X(_00994_));
 sky130_fd_sc_hd__xnor2_1 _12153_ (.A(\genblk2[10].wave_shpr.div.acc[19] ),
    .B(_05900_),
    .Y(_05903_));
 sky130_fd_sc_hd__a22o_1 _12154_ (.A1(net705),
    .A2(_05876_),
    .B1(_05883_),
    .B2(_05903_),
    .X(_00995_));
 sky130_fd_sc_hd__nor2_1 _12155_ (.A(_05783_),
    .B(_05899_),
    .Y(_05904_));
 sky130_fd_sc_hd__o21a_1 _12156_ (.A1(\genblk2[10].wave_shpr.div.acc[19] ),
    .A2(_05900_),
    .B1(\genblk2[10].wave_shpr.div.acc[20] ),
    .X(_05905_));
 sky130_fd_sc_hd__or2_1 _12157_ (.A(_05904_),
    .B(_05905_),
    .X(_05906_));
 sky130_fd_sc_hd__a22o_1 _12158_ (.A1(net1087),
    .A2(_05876_),
    .B1(_05883_),
    .B2(_05906_),
    .X(_00996_));
 sky130_fd_sc_hd__xor2_1 _12159_ (.A(\genblk2[10].wave_shpr.div.acc[21] ),
    .B(_05904_),
    .X(_05907_));
 sky130_fd_sc_hd__a22o_1 _12160_ (.A1(net1257),
    .A2(_05818_),
    .B1(_05883_),
    .B2(_05907_),
    .X(_00997_));
 sky130_fd_sc_hd__or3_1 _12161_ (.A(\genblk2[10].wave_shpr.div.acc[21] ),
    .B(_05783_),
    .C(_05899_),
    .X(_05908_));
 sky130_fd_sc_hd__xnor2_1 _12162_ (.A(\genblk2[10].wave_shpr.div.acc[22] ),
    .B(_05908_),
    .Y(_05909_));
 sky130_fd_sc_hd__a22o_1 _12163_ (.A1(net906),
    .A2(_05818_),
    .B1(_05883_),
    .B2(_05909_),
    .X(_00998_));
 sky130_fd_sc_hd__or3b_1 _12164_ (.A(\genblk2[10].wave_shpr.div.acc[22] ),
    .B(_05908_),
    .C_N(\genblk2[10].wave_shpr.div.acc[23] ),
    .X(_05910_));
 sky130_fd_sc_hd__o21bai_1 _12165_ (.A1(\genblk2[10].wave_shpr.div.acc[22] ),
    .A2(_05908_),
    .B1_N(\genblk2[10].wave_shpr.div.acc[23] ),
    .Y(_05911_));
 sky130_fd_sc_hd__a32o_1 _12166_ (.A1(_05816_),
    .A2(_05910_),
    .A3(_05911_),
    .B1(_05818_),
    .B2(net536),
    .X(_00999_));
 sky130_fd_sc_hd__nand2_1 _12167_ (.A(\genblk2[10].wave_shpr.div.acc[24] ),
    .B(_05784_),
    .Y(_05912_));
 sky130_fd_sc_hd__o21ai_1 _12168_ (.A1(_05785_),
    .A2(_05899_),
    .B1(_05912_),
    .Y(_05913_));
 sky130_fd_sc_hd__a22o_1 _12169_ (.A1(net1226),
    .A2(_05818_),
    .B1(_05816_),
    .B2(_05913_),
    .X(_01000_));
 sky130_fd_sc_hd__or3b_1 _12170_ (.A(_05785_),
    .B(\genblk2[10].wave_shpr.div.acc[25] ),
    .C_N(\genblk2[10].wave_shpr.div.acc[26] ),
    .X(_05914_));
 sky130_fd_sc_hd__a21bo_1 _12171_ (.A1(\genblk2[10].wave_shpr.div.acc[25] ),
    .A2(_05785_),
    .B1_N(_05914_),
    .X(_05915_));
 sky130_fd_sc_hd__a22o_1 _12172_ (.A1(net1081),
    .A2(_05818_),
    .B1(_05816_),
    .B2(_05915_),
    .X(_01001_));
 sky130_fd_sc_hd__mux2_1 _12173_ (.A0(_05815_),
    .A1(_05812_),
    .S(\genblk2[10].wave_shpr.div.i[0] ),
    .X(_05916_));
 sky130_fd_sc_hd__clkbuf_1 _12174_ (.A(_05916_),
    .X(_01002_));
 sky130_fd_sc_hd__or2_1 _12175_ (.A(\genblk2[10].wave_shpr.div.i[1] ),
    .B(\genblk2[10].wave_shpr.div.i[0] ),
    .X(_05917_));
 sky130_fd_sc_hd__nand2_1 _12176_ (.A(\genblk2[10].wave_shpr.div.i[1] ),
    .B(\genblk2[10].wave_shpr.div.i[0] ),
    .Y(_05918_));
 sky130_fd_sc_hd__a32o_1 _12177_ (.A1(_05816_),
    .A2(_05917_),
    .A3(_05918_),
    .B1(_05818_),
    .B2(net1090),
    .X(_01003_));
 sky130_fd_sc_hd__a21o_1 _12178_ (.A1(\genblk2[10].wave_shpr.div.i[1] ),
    .A2(\genblk2[10].wave_shpr.div.i[0] ),
    .B1(\genblk2[10].wave_shpr.div.i[2] ),
    .X(_05919_));
 sky130_fd_sc_hd__and3_1 _12179_ (.A(\genblk2[10].wave_shpr.div.i[1] ),
    .B(\genblk2[10].wave_shpr.div.i[0] ),
    .C(\genblk2[10].wave_shpr.div.i[2] ),
    .X(_05920_));
 sky130_fd_sc_hd__inv_2 _12180_ (.A(_05920_),
    .Y(_05921_));
 sky130_fd_sc_hd__a32o_1 _12181_ (.A1(_05816_),
    .A2(_05919_),
    .A3(_05921_),
    .B1(_05818_),
    .B2(net748),
    .X(_01004_));
 sky130_fd_sc_hd__a21oi_1 _12182_ (.A1(_00002_),
    .A2(_05920_),
    .B1(net1153),
    .Y(_05922_));
 sky130_fd_sc_hd__and3_1 _12183_ (.A(\genblk2[10].wave_shpr.div.i[3] ),
    .B(_02207_),
    .C(_05920_),
    .X(_05923_));
 sky130_fd_sc_hd__nor3_1 _12184_ (.A(_03690_),
    .B(_05922_),
    .C(_05923_),
    .Y(_01005_));
 sky130_fd_sc_hd__o21ai_1 _12185_ (.A1(net289),
    .A2(_05923_),
    .B1(_03855_),
    .Y(_05924_));
 sky130_fd_sc_hd__a21oi_1 _12186_ (.A1(net289),
    .A2(_05923_),
    .B1(_05924_),
    .Y(_01006_));
 sky130_fd_sc_hd__or2b_1 _12187_ (.A(\genblk2[11].wave_shpr.div.acc[17] ),
    .B_N(\genblk2[11].wave_shpr.div.b1[17] ),
    .X(_05925_));
 sky130_fd_sc_hd__xor2_1 _12188_ (.A(\genblk2[11].wave_shpr.div.b1[16] ),
    .B(\genblk2[11].wave_shpr.div.acc[16] ),
    .X(_05926_));
 sky130_fd_sc_hd__or2b_1 _12189_ (.A(\genblk2[11].wave_shpr.div.acc[15] ),
    .B_N(\genblk2[11].wave_shpr.div.b1[15] ),
    .X(_05927_));
 sky130_fd_sc_hd__or2b_1 _12190_ (.A(\genblk2[11].wave_shpr.div.acc[14] ),
    .B_N(\genblk2[11].wave_shpr.div.b1[14] ),
    .X(_05928_));
 sky130_fd_sc_hd__or2b_1 _12191_ (.A(\genblk2[11].wave_shpr.div.acc[13] ),
    .B_N(\genblk2[11].wave_shpr.div.b1[13] ),
    .X(_05929_));
 sky130_fd_sc_hd__or2b_1 _12192_ (.A(\genblk2[11].wave_shpr.div.acc[12] ),
    .B_N(\genblk2[11].wave_shpr.div.b1[12] ),
    .X(_05930_));
 sky130_fd_sc_hd__or2b_1 _12193_ (.A(\genblk2[11].wave_shpr.div.acc[11] ),
    .B_N(\genblk2[11].wave_shpr.div.b1[11] ),
    .X(_05931_));
 sky130_fd_sc_hd__or2b_1 _12194_ (.A(\genblk2[11].wave_shpr.div.acc[10] ),
    .B_N(\genblk2[11].wave_shpr.div.b1[10] ),
    .X(_05932_));
 sky130_fd_sc_hd__or2b_1 _12195_ (.A(\genblk2[11].wave_shpr.div.acc[9] ),
    .B_N(\genblk2[11].wave_shpr.div.b1[9] ),
    .X(_05933_));
 sky130_fd_sc_hd__or2b_1 _12196_ (.A(\genblk2[11].wave_shpr.div.acc[8] ),
    .B_N(\genblk2[11].wave_shpr.div.b1[8] ),
    .X(_05934_));
 sky130_fd_sc_hd__or2b_1 _12197_ (.A(\genblk2[11].wave_shpr.div.acc[7] ),
    .B_N(\genblk2[11].wave_shpr.div.b1[7] ),
    .X(_05935_));
 sky130_fd_sc_hd__or2b_1 _12198_ (.A(\genblk2[11].wave_shpr.div.acc[6] ),
    .B_N(\genblk2[11].wave_shpr.div.b1[6] ),
    .X(_05936_));
 sky130_fd_sc_hd__or2b_1 _12199_ (.A(\genblk2[11].wave_shpr.div.acc[5] ),
    .B_N(\genblk2[11].wave_shpr.div.b1[5] ),
    .X(_05937_));
 sky130_fd_sc_hd__or2b_1 _12200_ (.A(\genblk2[11].wave_shpr.div.acc[4] ),
    .B_N(\genblk2[11].wave_shpr.div.b1[4] ),
    .X(_05938_));
 sky130_fd_sc_hd__or2b_1 _12201_ (.A(\genblk2[11].wave_shpr.div.acc[3] ),
    .B_N(\genblk2[11].wave_shpr.div.b1[3] ),
    .X(_05939_));
 sky130_fd_sc_hd__inv_2 _12202_ (.A(\genblk2[11].wave_shpr.div.b1[2] ),
    .Y(_05940_));
 sky130_fd_sc_hd__xor2_1 _12203_ (.A(\genblk2[11].wave_shpr.div.acc[1] ),
    .B(\genblk2[11].wave_shpr.div.b1[1] ),
    .X(_05941_));
 sky130_fd_sc_hd__and2b_1 _12204_ (.A_N(\genblk2[11].wave_shpr.div.acc[0] ),
    .B(\genblk2[11].wave_shpr.div.b1[0] ),
    .X(_05942_));
 sky130_fd_sc_hd__or2b_1 _12205_ (.A(\genblk2[11].wave_shpr.div.b1[1] ),
    .B_N(\genblk2[11].wave_shpr.div.acc[1] ),
    .X(_05943_));
 sky130_fd_sc_hd__o21ai_1 _12206_ (.A1(_05941_),
    .A2(_05942_),
    .B1(_05943_),
    .Y(_05944_));
 sky130_fd_sc_hd__o21a_1 _12207_ (.A1(_05940_),
    .A2(\genblk2[11].wave_shpr.div.acc[2] ),
    .B1(_05944_),
    .X(_05945_));
 sky130_fd_sc_hd__a21o_1 _12208_ (.A1(_05940_),
    .A2(\genblk2[11].wave_shpr.div.acc[2] ),
    .B1(_05945_),
    .X(_05946_));
 sky130_fd_sc_hd__and2b_1 _12209_ (.A_N(\genblk2[11].wave_shpr.div.b1[3] ),
    .B(\genblk2[11].wave_shpr.div.acc[3] ),
    .X(_05947_));
 sky130_fd_sc_hd__a21o_1 _12210_ (.A1(_05939_),
    .A2(_05946_),
    .B1(_05947_),
    .X(_05948_));
 sky130_fd_sc_hd__and2b_1 _12211_ (.A_N(\genblk2[11].wave_shpr.div.b1[4] ),
    .B(\genblk2[11].wave_shpr.div.acc[4] ),
    .X(_05949_));
 sky130_fd_sc_hd__a21o_1 _12212_ (.A1(_05938_),
    .A2(_05948_),
    .B1(_05949_),
    .X(_05950_));
 sky130_fd_sc_hd__and2b_1 _12213_ (.A_N(\genblk2[11].wave_shpr.div.b1[5] ),
    .B(\genblk2[11].wave_shpr.div.acc[5] ),
    .X(_05951_));
 sky130_fd_sc_hd__a21o_1 _12214_ (.A1(_05937_),
    .A2(_05950_),
    .B1(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__and2b_1 _12215_ (.A_N(\genblk2[11].wave_shpr.div.b1[6] ),
    .B(\genblk2[11].wave_shpr.div.acc[6] ),
    .X(_05953_));
 sky130_fd_sc_hd__a21o_1 _12216_ (.A1(_05936_),
    .A2(_05952_),
    .B1(_05953_),
    .X(_05954_));
 sky130_fd_sc_hd__and2b_1 _12217_ (.A_N(\genblk2[11].wave_shpr.div.b1[7] ),
    .B(\genblk2[11].wave_shpr.div.acc[7] ),
    .X(_05955_));
 sky130_fd_sc_hd__a21o_1 _12218_ (.A1(_05935_),
    .A2(_05954_),
    .B1(_05955_),
    .X(_05956_));
 sky130_fd_sc_hd__and2b_1 _12219_ (.A_N(\genblk2[11].wave_shpr.div.b1[8] ),
    .B(\genblk2[11].wave_shpr.div.acc[8] ),
    .X(_05957_));
 sky130_fd_sc_hd__a21o_1 _12220_ (.A1(_05934_),
    .A2(_05956_),
    .B1(_05957_),
    .X(_05958_));
 sky130_fd_sc_hd__and2b_1 _12221_ (.A_N(\genblk2[11].wave_shpr.div.b1[9] ),
    .B(\genblk2[11].wave_shpr.div.acc[9] ),
    .X(_05959_));
 sky130_fd_sc_hd__a21o_1 _12222_ (.A1(_05933_),
    .A2(_05958_),
    .B1(_05959_),
    .X(_05960_));
 sky130_fd_sc_hd__and2b_1 _12223_ (.A_N(\genblk2[11].wave_shpr.div.b1[10] ),
    .B(\genblk2[11].wave_shpr.div.acc[10] ),
    .X(_05961_));
 sky130_fd_sc_hd__a21o_1 _12224_ (.A1(_05932_),
    .A2(_05960_),
    .B1(_05961_),
    .X(_05962_));
 sky130_fd_sc_hd__and2b_1 _12225_ (.A_N(\genblk2[11].wave_shpr.div.b1[11] ),
    .B(\genblk2[11].wave_shpr.div.acc[11] ),
    .X(_05963_));
 sky130_fd_sc_hd__a21o_1 _12226_ (.A1(_05931_),
    .A2(_05962_),
    .B1(_05963_),
    .X(_05964_));
 sky130_fd_sc_hd__and2b_1 _12227_ (.A_N(\genblk2[11].wave_shpr.div.b1[12] ),
    .B(\genblk2[11].wave_shpr.div.acc[12] ),
    .X(_05965_));
 sky130_fd_sc_hd__a21o_1 _12228_ (.A1(_05930_),
    .A2(_05964_),
    .B1(_05965_),
    .X(_05966_));
 sky130_fd_sc_hd__and2b_1 _12229_ (.A_N(\genblk2[11].wave_shpr.div.b1[13] ),
    .B(\genblk2[11].wave_shpr.div.acc[13] ),
    .X(_05967_));
 sky130_fd_sc_hd__a21o_1 _12230_ (.A1(_05929_),
    .A2(_05966_),
    .B1(_05967_),
    .X(_05968_));
 sky130_fd_sc_hd__and2b_1 _12231_ (.A_N(\genblk2[11].wave_shpr.div.b1[14] ),
    .B(\genblk2[11].wave_shpr.div.acc[14] ),
    .X(_05969_));
 sky130_fd_sc_hd__a21o_1 _12232_ (.A1(_05928_),
    .A2(_05968_),
    .B1(_05969_),
    .X(_05970_));
 sky130_fd_sc_hd__and2b_1 _12233_ (.A_N(\genblk2[11].wave_shpr.div.b1[15] ),
    .B(\genblk2[11].wave_shpr.div.acc[15] ),
    .X(_05971_));
 sky130_fd_sc_hd__a21o_1 _12234_ (.A1(_05927_),
    .A2(_05970_),
    .B1(_05971_),
    .X(_05972_));
 sky130_fd_sc_hd__and2b_1 _12235_ (.A_N(_05926_),
    .B(_05972_),
    .X(_05973_));
 sky130_fd_sc_hd__a21o_1 _12236_ (.A1(_05810_),
    .A2(\genblk2[11].wave_shpr.div.acc[16] ),
    .B1(_05973_),
    .X(_05974_));
 sky130_fd_sc_hd__and2b_1 _12237_ (.A_N(\genblk2[11].wave_shpr.div.b1[17] ),
    .B(\genblk2[11].wave_shpr.div.acc[17] ),
    .X(_05975_));
 sky130_fd_sc_hd__a21o_1 _12238_ (.A1(_05925_),
    .A2(_05974_),
    .B1(_05975_),
    .X(_05976_));
 sky130_fd_sc_hd__or2_1 _12239_ (.A(\genblk2[11].wave_shpr.div.acc[18] ),
    .B(_05976_),
    .X(_05977_));
 sky130_fd_sc_hd__or2_1 _12240_ (.A(\genblk2[11].wave_shpr.div.acc[19] ),
    .B(_05977_),
    .X(_05978_));
 sky130_fd_sc_hd__or4_1 _12241_ (.A(\genblk2[11].wave_shpr.div.acc[22] ),
    .B(\genblk2[11].wave_shpr.div.acc[21] ),
    .C(\genblk2[11].wave_shpr.div.acc[20] ),
    .D(_05978_),
    .X(_05979_));
 sky130_fd_sc_hd__or2_2 _12242_ (.A(\genblk2[11].wave_shpr.div.acc[23] ),
    .B(_05979_),
    .X(_05980_));
 sky130_fd_sc_hd__or4_2 _12243_ (.A(\genblk2[11].wave_shpr.div.acc[25] ),
    .B(\genblk2[11].wave_shpr.div.acc[24] ),
    .C(\genblk2[11].wave_shpr.div.acc[26] ),
    .D(_05980_),
    .X(_05981_));
 sky130_fd_sc_hd__buf_4 _12244_ (.A(_05981_),
    .X(_05982_));
 sky130_fd_sc_hd__mux2_1 _12245_ (.A0(\genblk2[11].wave_shpr.div.fin_quo[0] ),
    .A1(_05982_),
    .S(_00005_),
    .X(_05983_));
 sky130_fd_sc_hd__clkbuf_1 _12246_ (.A(_05983_),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _12247_ (.A0(\genblk2[11].wave_shpr.div.fin_quo[1] ),
    .A1(net1310),
    .S(_00005_),
    .X(_05984_));
 sky130_fd_sc_hd__clkbuf_1 _12248_ (.A(_05984_),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_1 _12249_ (.A0(\genblk2[11].wave_shpr.div.fin_quo[2] ),
    .A1(net769),
    .S(_00005_),
    .X(_05985_));
 sky130_fd_sc_hd__clkbuf_1 _12250_ (.A(_05985_),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_1 _12251_ (.A0(\genblk2[11].wave_shpr.div.fin_quo[3] ),
    .A1(net402),
    .S(_00005_),
    .X(_05986_));
 sky130_fd_sc_hd__clkbuf_1 _12252_ (.A(_05986_),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_1 _12253_ (.A0(\genblk2[11].wave_shpr.div.fin_quo[4] ),
    .A1(\genblk2[11].wave_shpr.div.quo[3] ),
    .S(_00005_),
    .X(_05987_));
 sky130_fd_sc_hd__clkbuf_1 _12254_ (.A(_05987_),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _12255_ (.A0(\genblk2[11].wave_shpr.div.fin_quo[5] ),
    .A1(net767),
    .S(_00005_),
    .X(_05988_));
 sky130_fd_sc_hd__clkbuf_1 _12256_ (.A(_05988_),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _12257_ (.A0(\genblk2[11].wave_shpr.div.fin_quo[6] ),
    .A1(net1332),
    .S(_00005_),
    .X(_05989_));
 sky130_fd_sc_hd__clkbuf_1 _12258_ (.A(_05989_),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_1 _12259_ (.A0(\genblk2[11].wave_shpr.div.fin_quo[7] ),
    .A1(net1341),
    .S(_00005_),
    .X(_05990_));
 sky130_fd_sc_hd__clkbuf_1 _12260_ (.A(_05990_),
    .X(_01014_));
 sky130_fd_sc_hd__mux2_1 _12261_ (.A0(\genblk2[1].wave_shpr.div.b1[0] ),
    .A1(_01329_),
    .S(_05802_),
    .X(_05991_));
 sky130_fd_sc_hd__clkbuf_1 _12262_ (.A(_05991_),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_1 _12263_ (.A0(\genblk2[1].wave_shpr.div.b1[1] ),
    .A1(_01263_),
    .S(_05802_),
    .X(_05992_));
 sky130_fd_sc_hd__clkbuf_1 _12264_ (.A(_05992_),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_1 _12265_ (.A0(net1295),
    .A1(_01240_),
    .S(_05802_),
    .X(_05993_));
 sky130_fd_sc_hd__clkbuf_1 _12266_ (.A(_05993_),
    .X(_01017_));
 sky130_fd_sc_hd__buf_4 _12267_ (.A(_03707_),
    .X(_05994_));
 sky130_fd_sc_hd__mux2_1 _12268_ (.A0(net1235),
    .A1(_01589_),
    .S(_05994_),
    .X(_05995_));
 sky130_fd_sc_hd__clkbuf_1 _12269_ (.A(_05995_),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_1 _12270_ (.A0(net1267),
    .A1(_04229_),
    .S(_05994_),
    .X(_05996_));
 sky130_fd_sc_hd__clkbuf_1 _12271_ (.A(_05996_),
    .X(_01019_));
 sky130_fd_sc_hd__inv_2 _12272_ (.A(_01305_),
    .Y(_05997_));
 sky130_fd_sc_hd__mux2_1 _12273_ (.A0(net1272),
    .A1(_05997_),
    .S(_05994_),
    .X(_05998_));
 sky130_fd_sc_hd__clkbuf_1 _12274_ (.A(_05998_),
    .X(_01020_));
 sky130_fd_sc_hd__mux2_1 _12275_ (.A0(\genblk2[1].wave_shpr.div.b1[6] ),
    .A1(_01311_),
    .S(_05994_),
    .X(_05999_));
 sky130_fd_sc_hd__clkbuf_1 _12276_ (.A(_05999_),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_1 _12277_ (.A0(net1274),
    .A1(_02001_),
    .S(_05994_),
    .X(_06000_));
 sky130_fd_sc_hd__clkbuf_1 _12278_ (.A(_06000_),
    .X(_01022_));
 sky130_fd_sc_hd__mux2_1 _12279_ (.A0(_01308_),
    .A1(\genblk2[1].wave_shpr.div.b1[8] ),
    .S(_03719_),
    .X(_06001_));
 sky130_fd_sc_hd__clkbuf_1 _12280_ (.A(_06001_),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_1 _12281_ (.A0(\genblk2[1].wave_shpr.div.b1[9] ),
    .A1(_02013_),
    .S(_05994_),
    .X(_06002_));
 sky130_fd_sc_hd__clkbuf_1 _12282_ (.A(_06002_),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_1 _12283_ (.A0(\genblk2[1].wave_shpr.div.b1[10] ),
    .A1(_01946_),
    .S(_05994_),
    .X(_06003_));
 sky130_fd_sc_hd__clkbuf_1 _12284_ (.A(_06003_),
    .X(_01025_));
 sky130_fd_sc_hd__nor2_1 _12285_ (.A(_03702_),
    .B(net1121),
    .Y(_06004_));
 sky130_fd_sc_hd__a21oi_1 _12286_ (.A1(_03726_),
    .A2(_01312_),
    .B1(_06004_),
    .Y(_01026_));
 sky130_fd_sc_hd__inv_2 _12287_ (.A(_01337_),
    .Y(_06005_));
 sky130_fd_sc_hd__mux2_1 _12288_ (.A0(\genblk2[1].wave_shpr.div.b1[12] ),
    .A1(_06005_),
    .S(_05994_),
    .X(_06006_));
 sky130_fd_sc_hd__clkbuf_1 _12289_ (.A(_06006_),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _12290_ (.A0(net1299),
    .A1(_01249_),
    .S(_05994_),
    .X(_06007_));
 sky130_fd_sc_hd__clkbuf_1 _12291_ (.A(_06007_),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_1 _12292_ (.A0(net1270),
    .A1(_01327_),
    .S(_05994_),
    .X(_06008_));
 sky130_fd_sc_hd__clkbuf_1 _12293_ (.A(_06008_),
    .X(_01029_));
 sky130_fd_sc_hd__o21a_1 _12294_ (.A1(_03732_),
    .A2(net406),
    .B1(_03733_),
    .X(_01030_));
 sky130_fd_sc_hd__a21bo_1 _12295_ (.A1(_03687_),
    .A2(net425),
    .B1_N(_03716_),
    .X(_01031_));
 sky130_fd_sc_hd__a21bo_1 _12296_ (.A1(_03687_),
    .A2(net409),
    .B1_N(_03735_),
    .X(_01032_));
 sky130_fd_sc_hd__buf_4 _12297_ (.A(_03942_),
    .X(_06009_));
 sky130_fd_sc_hd__buf_4 _12298_ (.A(_03941_),
    .X(_06010_));
 sky130_fd_sc_hd__a22o_1 _12299_ (.A1(net430),
    .A2(_06009_),
    .B1(_06010_),
    .B2(_05982_),
    .X(_01033_));
 sky130_fd_sc_hd__a22o_1 _12300_ (.A1(\genblk2[11].wave_shpr.div.quo[1] ),
    .A2(_06009_),
    .B1(_06010_),
    .B2(net430),
    .X(_01034_));
 sky130_fd_sc_hd__a22o_1 _12301_ (.A1(net402),
    .A2(_06009_),
    .B1(_06010_),
    .B2(net769),
    .X(_01035_));
 sky130_fd_sc_hd__a22o_1 _12302_ (.A1(\genblk2[11].wave_shpr.div.quo[3] ),
    .A2(_06009_),
    .B1(_06010_),
    .B2(net402),
    .X(_01036_));
 sky130_fd_sc_hd__a22o_1 _12303_ (.A1(net767),
    .A2(_06009_),
    .B1(_06010_),
    .B2(net776),
    .X(_01037_));
 sky130_fd_sc_hd__a22o_1 _12304_ (.A1(net731),
    .A2(_06009_),
    .B1(_06010_),
    .B2(net767),
    .X(_01038_));
 sky130_fd_sc_hd__a22o_1 _12305_ (.A1(net397),
    .A2(_06009_),
    .B1(_06010_),
    .B2(net731),
    .X(_01039_));
 sky130_fd_sc_hd__a22o_1 _12306_ (.A1(net358),
    .A2(_06009_),
    .B1(_06010_),
    .B2(net397),
    .X(_01040_));
 sky130_fd_sc_hd__a22o_1 _12307_ (.A1(net355),
    .A2(_06009_),
    .B1(_06010_),
    .B2(net358),
    .X(_01041_));
 sky130_fd_sc_hd__and2_1 _12308_ (.A(_05835_),
    .B(\genblk1[11].osc.clkdiv_C.cnt[0] ),
    .X(_06011_));
 sky130_fd_sc_hd__a221o_1 _12309_ (.A1(\genblk2[11].wave_shpr.div.quo[9] ),
    .A2(_03947_),
    .B1(_03944_),
    .B2(net355),
    .C1(_06011_),
    .X(_01042_));
 sky130_fd_sc_hd__and2_1 _12310_ (.A(_05835_),
    .B(\genblk1[11].osc.clkdiv_C.cnt[1] ),
    .X(_06012_));
 sky130_fd_sc_hd__a221o_1 _12311_ (.A1(net467),
    .A2(_03947_),
    .B1(_03944_),
    .B2(net479),
    .C1(_06012_),
    .X(_01043_));
 sky130_fd_sc_hd__and2_1 _12312_ (.A(_05835_),
    .B(\genblk1[11].osc.clkdiv_C.cnt[2] ),
    .X(_06013_));
 sky130_fd_sc_hd__a221o_1 _12313_ (.A1(\genblk2[11].wave_shpr.div.quo[11] ),
    .A2(_03947_),
    .B1(_03944_),
    .B2(net467),
    .C1(_06013_),
    .X(_01044_));
 sky130_fd_sc_hd__clkbuf_4 _12314_ (.A(_03942_),
    .X(_06014_));
 sky130_fd_sc_hd__clkbuf_4 _12315_ (.A(_03941_),
    .X(_06015_));
 sky130_fd_sc_hd__and2_1 _12316_ (.A(_05835_),
    .B(\genblk1[11].osc.clkdiv_C.cnt[3] ),
    .X(_06016_));
 sky130_fd_sc_hd__a221o_1 _12317_ (.A1(net443),
    .A2(_06014_),
    .B1(_06015_),
    .B2(\genblk2[11].wave_shpr.div.quo[11] ),
    .C1(_06016_),
    .X(_01045_));
 sky130_fd_sc_hd__and2_1 _12318_ (.A(_05835_),
    .B(\genblk1[11].osc.clkdiv_C.cnt[4] ),
    .X(_06017_));
 sky130_fd_sc_hd__a221o_1 _12319_ (.A1(net342),
    .A2(_06014_),
    .B1(_06015_),
    .B2(net443),
    .C1(_06017_),
    .X(_01046_));
 sky130_fd_sc_hd__and2_1 _12320_ (.A(_05835_),
    .B(\genblk1[11].osc.clkdiv_C.cnt[5] ),
    .X(_06018_));
 sky130_fd_sc_hd__a221o_1 _12321_ (.A1(\genblk2[11].wave_shpr.div.quo[14] ),
    .A2(_06014_),
    .B1(_06015_),
    .B2(net342),
    .C1(_06018_),
    .X(_01047_));
 sky130_fd_sc_hd__and2_1 _12322_ (.A(_05835_),
    .B(\genblk1[11].osc.clkdiv_C.cnt[6] ),
    .X(_06019_));
 sky130_fd_sc_hd__a221o_1 _12323_ (.A1(net351),
    .A2(_06014_),
    .B1(_06015_),
    .B2(net489),
    .C1(_06019_),
    .X(_01048_));
 sky130_fd_sc_hd__and2_1 _12324_ (.A(_03689_),
    .B(\genblk1[11].osc.clkdiv_C.cnt[7] ),
    .X(_06020_));
 sky130_fd_sc_hd__a221o_1 _12325_ (.A1(\genblk2[11].wave_shpr.div.quo[16] ),
    .A2(_06014_),
    .B1(_06015_),
    .B2(net351),
    .C1(_06020_),
    .X(_01049_));
 sky130_fd_sc_hd__and2_1 _12326_ (.A(_03689_),
    .B(\genblk1[11].osc.clkdiv_C.cnt[8] ),
    .X(_06021_));
 sky130_fd_sc_hd__a221o_1 _12327_ (.A1(net510),
    .A2(_06014_),
    .B1(_06015_),
    .B2(net571),
    .C1(_06021_),
    .X(_01050_));
 sky130_fd_sc_hd__and2_1 _12328_ (.A(_03689_),
    .B(\genblk1[11].osc.clkdiv_C.cnt[9] ),
    .X(_06022_));
 sky130_fd_sc_hd__a221o_1 _12329_ (.A1(net509),
    .A2(_06014_),
    .B1(_06015_),
    .B2(net510),
    .C1(_06022_),
    .X(_01051_));
 sky130_fd_sc_hd__and2_1 _12330_ (.A(_03689_),
    .B(\genblk1[11].osc.clkdiv_C.cnt[10] ),
    .X(_06023_));
 sky130_fd_sc_hd__a221o_1 _12331_ (.A1(net483),
    .A2(_06014_),
    .B1(_06015_),
    .B2(net509),
    .C1(_06023_),
    .X(_01052_));
 sky130_fd_sc_hd__nor2_1 _12332_ (.A(_03833_),
    .B(_02128_),
    .Y(_06024_));
 sky130_fd_sc_hd__a221o_1 _12333_ (.A1(net239),
    .A2(_06014_),
    .B1(_06015_),
    .B2(net483),
    .C1(_06024_),
    .X(_01053_));
 sky130_fd_sc_hd__and2_1 _12334_ (.A(_03689_),
    .B(\genblk1[11].osc.clkdiv_C.cnt[12] ),
    .X(_06025_));
 sky130_fd_sc_hd__a221o_1 _12335_ (.A1(\genblk2[11].wave_shpr.div.quo[21] ),
    .A2(_06014_),
    .B1(_06015_),
    .B2(net239),
    .C1(_06025_),
    .X(_01054_));
 sky130_fd_sc_hd__and2_1 _12336_ (.A(_03689_),
    .B(\genblk1[11].osc.clkdiv_C.cnt[13] ),
    .X(_06026_));
 sky130_fd_sc_hd__a221o_1 _12337_ (.A1(net438),
    .A2(_03942_),
    .B1(_03941_),
    .B2(net504),
    .C1(_06026_),
    .X(_01055_));
 sky130_fd_sc_hd__nor2_1 _12338_ (.A(_03833_),
    .B(_02081_),
    .Y(_06027_));
 sky130_fd_sc_hd__a221o_1 _12339_ (.A1(net434),
    .A2(_03942_),
    .B1(_03941_),
    .B2(net438),
    .C1(_06027_),
    .X(_01056_));
 sky130_fd_sc_hd__nor2_1 _12340_ (.A(_03833_),
    .B(_02080_),
    .Y(_06028_));
 sky130_fd_sc_hd__a221o_1 _12341_ (.A1(net412),
    .A2(_03942_),
    .B1(_03941_),
    .B2(net434),
    .C1(_06028_),
    .X(_01057_));
 sky130_fd_sc_hd__and2_1 _12342_ (.A(_03689_),
    .B(\genblk1[11].osc.clkdiv_C.cnt[16] ),
    .X(_06029_));
 sky130_fd_sc_hd__a221o_1 _12343_ (.A1(\genblk2[11].wave_shpr.div.acc_next[0] ),
    .A2(_03942_),
    .B1(_03941_),
    .B2(net412),
    .C1(_06029_),
    .X(_01058_));
 sky130_fd_sc_hd__or2b_1 _12344_ (.A(\genblk2[11].wave_shpr.div.acc_next[0] ),
    .B_N(_03941_),
    .X(_06030_));
 sky130_fd_sc_hd__o221a_1 _12345_ (.A1(_03819_),
    .A2(net1220),
    .B1(_00004_),
    .B2(\genblk2[11].wave_shpr.div.acc[0] ),
    .C1(_06030_),
    .X(_01059_));
 sky130_fd_sc_hd__nand3_1 _12346_ (.A(\genblk2[11].wave_shpr.div.b1[0] ),
    .B(\genblk2[11].wave_shpr.div.acc[0] ),
    .C(_05982_),
    .Y(_06031_));
 sky130_fd_sc_hd__a21o_1 _12347_ (.A1(\genblk2[11].wave_shpr.div.b1[0] ),
    .A2(_05982_),
    .B1(\genblk2[11].wave_shpr.div.acc[0] ),
    .X(_06032_));
 sky130_fd_sc_hd__a32o_1 _12348_ (.A1(_03944_),
    .A2(_06031_),
    .A3(_06032_),
    .B1(_03947_),
    .B2(net1044),
    .X(_01060_));
 sky130_fd_sc_hd__or2_1 _12349_ (.A(\genblk2[11].wave_shpr.div.acc[1] ),
    .B(_05981_),
    .X(_06033_));
 sky130_fd_sc_hd__xnor2_1 _12350_ (.A(_05941_),
    .B(_05942_),
    .Y(_06034_));
 sky130_fd_sc_hd__nand2_1 _12351_ (.A(_05982_),
    .B(_06034_),
    .Y(_06035_));
 sky130_fd_sc_hd__a32o_1 _12352_ (.A1(_03944_),
    .A2(_06033_),
    .A3(_06035_),
    .B1(_03947_),
    .B2(net1127),
    .X(_01061_));
 sky130_fd_sc_hd__xor2_1 _12353_ (.A(\genblk2[11].wave_shpr.div.b1[2] ),
    .B(\genblk2[11].wave_shpr.div.acc[2] ),
    .X(_06036_));
 sky130_fd_sc_hd__xnor2_1 _12354_ (.A(_05944_),
    .B(_06036_),
    .Y(_06037_));
 sky130_fd_sc_hd__mux2_1 _12355_ (.A0(\genblk2[11].wave_shpr.div.acc[2] ),
    .A1(_06037_),
    .S(_05982_),
    .X(_06038_));
 sky130_fd_sc_hd__a22o_1 _12356_ (.A1(net1020),
    .A2(_06009_),
    .B1(_06010_),
    .B2(_06038_),
    .X(_01062_));
 sky130_fd_sc_hd__clkbuf_4 _12357_ (.A(_03942_),
    .X(_06039_));
 sky130_fd_sc_hd__clkbuf_4 _12358_ (.A(_03941_),
    .X(_06040_));
 sky130_fd_sc_hd__or2b_1 _12359_ (.A(_05947_),
    .B_N(_05939_),
    .X(_06041_));
 sky130_fd_sc_hd__xnor2_1 _12360_ (.A(_05946_),
    .B(_06041_),
    .Y(_06042_));
 sky130_fd_sc_hd__mux2_1 _12361_ (.A0(\genblk2[11].wave_shpr.div.acc[3] ),
    .A1(_06042_),
    .S(_05982_),
    .X(_06043_));
 sky130_fd_sc_hd__a22o_1 _12362_ (.A1(net985),
    .A2(_06039_),
    .B1(_06040_),
    .B2(_06043_),
    .X(_01063_));
 sky130_fd_sc_hd__or2b_1 _12363_ (.A(_05949_),
    .B_N(_05938_),
    .X(_06044_));
 sky130_fd_sc_hd__xnor2_1 _12364_ (.A(_06044_),
    .B(_05948_),
    .Y(_06045_));
 sky130_fd_sc_hd__mux2_1 _12365_ (.A0(\genblk2[11].wave_shpr.div.acc[4] ),
    .A1(_06045_),
    .S(_05982_),
    .X(_06046_));
 sky130_fd_sc_hd__a22o_1 _12366_ (.A1(net958),
    .A2(_06039_),
    .B1(_06040_),
    .B2(_06046_),
    .X(_01064_));
 sky130_fd_sc_hd__or2b_1 _12367_ (.A(_05951_),
    .B_N(_05937_),
    .X(_06047_));
 sky130_fd_sc_hd__xnor2_1 _12368_ (.A(_06047_),
    .B(_05950_),
    .Y(_06048_));
 sky130_fd_sc_hd__mux2_1 _12369_ (.A0(\genblk2[11].wave_shpr.div.acc[5] ),
    .A1(_06048_),
    .S(_05982_),
    .X(_06049_));
 sky130_fd_sc_hd__a22o_1 _12370_ (.A1(net841),
    .A2(_06039_),
    .B1(_06040_),
    .B2(_06049_),
    .X(_01065_));
 sky130_fd_sc_hd__or2b_1 _12371_ (.A(_05953_),
    .B_N(_05936_),
    .X(_06050_));
 sky130_fd_sc_hd__xnor2_1 _12372_ (.A(_05952_),
    .B(_06050_),
    .Y(_06051_));
 sky130_fd_sc_hd__mux2_1 _12373_ (.A0(\genblk2[11].wave_shpr.div.acc[6] ),
    .A1(_06051_),
    .S(_05982_),
    .X(_06052_));
 sky130_fd_sc_hd__a22o_1 _12374_ (.A1(net997),
    .A2(_06039_),
    .B1(_06040_),
    .B2(_06052_),
    .X(_01066_));
 sky130_fd_sc_hd__or2b_1 _12375_ (.A(_05955_),
    .B_N(_05935_),
    .X(_06053_));
 sky130_fd_sc_hd__xnor2_1 _12376_ (.A(_05954_),
    .B(_06053_),
    .Y(_06054_));
 sky130_fd_sc_hd__clkbuf_4 _12377_ (.A(_05981_),
    .X(_06055_));
 sky130_fd_sc_hd__mux2_1 _12378_ (.A0(\genblk2[11].wave_shpr.div.acc[7] ),
    .A1(_06054_),
    .S(_06055_),
    .X(_06056_));
 sky130_fd_sc_hd__a22o_1 _12379_ (.A1(net876),
    .A2(_06039_),
    .B1(_06040_),
    .B2(_06056_),
    .X(_01067_));
 sky130_fd_sc_hd__or2b_1 _12380_ (.A(_05957_),
    .B_N(_05934_),
    .X(_06057_));
 sky130_fd_sc_hd__xnor2_1 _12381_ (.A(_05956_),
    .B(_06057_),
    .Y(_06058_));
 sky130_fd_sc_hd__mux2_1 _12382_ (.A0(\genblk2[11].wave_shpr.div.acc[8] ),
    .A1(_06058_),
    .S(_06055_),
    .X(_06059_));
 sky130_fd_sc_hd__a22o_1 _12383_ (.A1(net762),
    .A2(_06039_),
    .B1(_06040_),
    .B2(_06059_),
    .X(_01068_));
 sky130_fd_sc_hd__or2b_1 _12384_ (.A(_05959_),
    .B_N(_05933_),
    .X(_06060_));
 sky130_fd_sc_hd__xnor2_1 _12385_ (.A(_05958_),
    .B(_06060_),
    .Y(_06061_));
 sky130_fd_sc_hd__mux2_1 _12386_ (.A0(\genblk2[11].wave_shpr.div.acc[9] ),
    .A1(_06061_),
    .S(_06055_),
    .X(_06062_));
 sky130_fd_sc_hd__a22o_1 _12387_ (.A1(net816),
    .A2(_06039_),
    .B1(_06040_),
    .B2(_06062_),
    .X(_01069_));
 sky130_fd_sc_hd__or2b_1 _12388_ (.A(_05961_),
    .B_N(_05932_),
    .X(_06063_));
 sky130_fd_sc_hd__xnor2_1 _12389_ (.A(_05960_),
    .B(_06063_),
    .Y(_06064_));
 sky130_fd_sc_hd__mux2_1 _12390_ (.A0(\genblk2[11].wave_shpr.div.acc[10] ),
    .A1(_06064_),
    .S(_06055_),
    .X(_06065_));
 sky130_fd_sc_hd__a22o_1 _12391_ (.A1(net785),
    .A2(_06039_),
    .B1(_06040_),
    .B2(_06065_),
    .X(_01070_));
 sky130_fd_sc_hd__or2b_1 _12392_ (.A(_05963_),
    .B_N(_05931_),
    .X(_06066_));
 sky130_fd_sc_hd__xnor2_1 _12393_ (.A(_05962_),
    .B(_06066_),
    .Y(_06067_));
 sky130_fd_sc_hd__mux2_1 _12394_ (.A0(\genblk2[11].wave_shpr.div.acc[11] ),
    .A1(_06067_),
    .S(_06055_),
    .X(_06068_));
 sky130_fd_sc_hd__a22o_1 _12395_ (.A1(net875),
    .A2(_06039_),
    .B1(_06040_),
    .B2(_06068_),
    .X(_01071_));
 sky130_fd_sc_hd__or2b_1 _12396_ (.A(_05965_),
    .B_N(_05930_),
    .X(_06069_));
 sky130_fd_sc_hd__xnor2_1 _12397_ (.A(_05964_),
    .B(_06069_),
    .Y(_06070_));
 sky130_fd_sc_hd__mux2_1 _12398_ (.A0(\genblk2[11].wave_shpr.div.acc[12] ),
    .A1(_06070_),
    .S(_06055_),
    .X(_06071_));
 sky130_fd_sc_hd__a22o_1 _12399_ (.A1(net949),
    .A2(_06039_),
    .B1(_06040_),
    .B2(_06071_),
    .X(_01072_));
 sky130_fd_sc_hd__clkbuf_4 _12400_ (.A(_03942_),
    .X(_06072_));
 sky130_fd_sc_hd__clkbuf_4 _12401_ (.A(_03941_),
    .X(_06073_));
 sky130_fd_sc_hd__or2b_1 _12402_ (.A(_05967_),
    .B_N(_05929_),
    .X(_06074_));
 sky130_fd_sc_hd__xnor2_1 _12403_ (.A(_05966_),
    .B(_06074_),
    .Y(_06075_));
 sky130_fd_sc_hd__mux2_1 _12404_ (.A0(\genblk2[11].wave_shpr.div.acc[13] ),
    .A1(_06075_),
    .S(_06055_),
    .X(_06076_));
 sky130_fd_sc_hd__a22o_1 _12405_ (.A1(net993),
    .A2(_06072_),
    .B1(_06073_),
    .B2(_06076_),
    .X(_01073_));
 sky130_fd_sc_hd__or2b_1 _12406_ (.A(_05969_),
    .B_N(_05928_),
    .X(_06077_));
 sky130_fd_sc_hd__xnor2_1 _12407_ (.A(_05968_),
    .B(_06077_),
    .Y(_06078_));
 sky130_fd_sc_hd__mux2_1 _12408_ (.A0(\genblk2[11].wave_shpr.div.acc[14] ),
    .A1(_06078_),
    .S(_06055_),
    .X(_06079_));
 sky130_fd_sc_hd__a22o_1 _12409_ (.A1(net897),
    .A2(_06072_),
    .B1(_06073_),
    .B2(_06079_),
    .X(_01074_));
 sky130_fd_sc_hd__or2b_1 _12410_ (.A(_05971_),
    .B_N(_05927_),
    .X(_06080_));
 sky130_fd_sc_hd__xnor2_1 _12411_ (.A(_05970_),
    .B(_06080_),
    .Y(_06081_));
 sky130_fd_sc_hd__mux2_1 _12412_ (.A0(\genblk2[11].wave_shpr.div.acc[15] ),
    .A1(_06081_),
    .S(_06055_),
    .X(_06082_));
 sky130_fd_sc_hd__a22o_1 _12413_ (.A1(net1125),
    .A2(_06072_),
    .B1(_06073_),
    .B2(_06082_),
    .X(_01075_));
 sky130_fd_sc_hd__xnor2_1 _12414_ (.A(_05926_),
    .B(_05972_),
    .Y(_06083_));
 sky130_fd_sc_hd__mux2_1 _12415_ (.A0(\genblk2[11].wave_shpr.div.acc[16] ),
    .A1(_06083_),
    .S(_06055_),
    .X(_06084_));
 sky130_fd_sc_hd__a22o_1 _12416_ (.A1(net878),
    .A2(_06072_),
    .B1(_06073_),
    .B2(_06084_),
    .X(_01076_));
 sky130_fd_sc_hd__or2b_1 _12417_ (.A(_05975_),
    .B_N(_05925_),
    .X(_06085_));
 sky130_fd_sc_hd__xnor2_1 _12418_ (.A(_05974_),
    .B(_06085_),
    .Y(_06086_));
 sky130_fd_sc_hd__mux2_1 _12419_ (.A0(\genblk2[11].wave_shpr.div.acc[17] ),
    .A1(_06086_),
    .S(_05981_),
    .X(_06087_));
 sky130_fd_sc_hd__a22o_1 _12420_ (.A1(net576),
    .A2(_06072_),
    .B1(_06073_),
    .B2(_06087_),
    .X(_01077_));
 sky130_fd_sc_hd__nor4_1 _12421_ (.A(\genblk2[11].wave_shpr.div.acc[25] ),
    .B(\genblk2[11].wave_shpr.div.acc[24] ),
    .C(\genblk2[11].wave_shpr.div.acc[26] ),
    .D(_05980_),
    .Y(_06088_));
 sky130_fd_sc_hd__or2_1 _12422_ (.A(_05977_),
    .B(net20),
    .X(_06089_));
 sky130_fd_sc_hd__o21ai_1 _12423_ (.A1(_05976_),
    .A2(net20),
    .B1(\genblk2[11].wave_shpr.div.acc[18] ),
    .Y(_06090_));
 sky130_fd_sc_hd__nand2_1 _12424_ (.A(_06089_),
    .B(_06090_),
    .Y(_06091_));
 sky130_fd_sc_hd__a22o_1 _12425_ (.A1(net641),
    .A2(_06072_),
    .B1(_06073_),
    .B2(_06091_),
    .X(_01078_));
 sky130_fd_sc_hd__nor2_1 _12426_ (.A(_05978_),
    .B(net20),
    .Y(_06092_));
 sky130_fd_sc_hd__a21o_1 _12427_ (.A1(\genblk2[11].wave_shpr.div.acc[19] ),
    .A2(_06089_),
    .B1(_06092_),
    .X(_06093_));
 sky130_fd_sc_hd__a22o_1 _12428_ (.A1(net1203),
    .A2(_06072_),
    .B1(_06073_),
    .B2(_06093_),
    .X(_01079_));
 sky130_fd_sc_hd__xor2_1 _12429_ (.A(\genblk2[11].wave_shpr.div.acc[20] ),
    .B(_06092_),
    .X(_06094_));
 sky130_fd_sc_hd__a22o_1 _12430_ (.A1(net931),
    .A2(_06072_),
    .B1(_06073_),
    .B2(_06094_),
    .X(_01080_));
 sky130_fd_sc_hd__or3_1 _12431_ (.A(\genblk2[11].wave_shpr.div.acc[20] ),
    .B(_05978_),
    .C(net20),
    .X(_06095_));
 sky130_fd_sc_hd__or4_1 _12432_ (.A(\genblk2[11].wave_shpr.div.acc[21] ),
    .B(\genblk2[11].wave_shpr.div.acc[20] ),
    .C(_05978_),
    .D(net20),
    .X(_06096_));
 sky130_fd_sc_hd__a21bo_1 _12433_ (.A1(\genblk2[11].wave_shpr.div.acc[21] ),
    .A2(_06095_),
    .B1_N(_06096_),
    .X(_06097_));
 sky130_fd_sc_hd__a22o_1 _12434_ (.A1(net955),
    .A2(_06072_),
    .B1(_06073_),
    .B2(_06097_),
    .X(_01081_));
 sky130_fd_sc_hd__xnor2_1 _12435_ (.A(\genblk2[11].wave_shpr.div.acc[22] ),
    .B(_06096_),
    .Y(_06098_));
 sky130_fd_sc_hd__a22o_1 _12436_ (.A1(net619),
    .A2(_06072_),
    .B1(_06073_),
    .B2(_06098_),
    .X(_01082_));
 sky130_fd_sc_hd__nor2_1 _12437_ (.A(_05980_),
    .B(_06088_),
    .Y(_06099_));
 sky130_fd_sc_hd__a21o_1 _12438_ (.A1(\genblk2[11].wave_shpr.div.acc[23] ),
    .A2(_05979_),
    .B1(_06099_),
    .X(_06100_));
 sky130_fd_sc_hd__a22o_1 _12439_ (.A1(\genblk2[11].wave_shpr.div.acc[24] ),
    .A2(_03947_),
    .B1(_03944_),
    .B2(_06100_),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_1 _12440_ (.A0(_06099_),
    .A1(_05980_),
    .S(\genblk2[11].wave_shpr.div.acc[24] ),
    .X(_06101_));
 sky130_fd_sc_hd__a22o_1 _12441_ (.A1(net1078),
    .A2(_03947_),
    .B1(_03944_),
    .B2(_06101_),
    .X(_01084_));
 sky130_fd_sc_hd__o21ai_1 _12442_ (.A1(\genblk2[11].wave_shpr.div.acc[24] ),
    .A2(_05980_),
    .B1(\genblk2[11].wave_shpr.div.acc[25] ),
    .Y(_06102_));
 sky130_fd_sc_hd__or4b_1 _12443_ (.A(\genblk2[11].wave_shpr.div.acc[25] ),
    .B(_05980_),
    .C(\genblk2[11].wave_shpr.div.acc[24] ),
    .D_N(\genblk2[11].wave_shpr.div.acc[26] ),
    .X(_06103_));
 sky130_fd_sc_hd__nand2_1 _12444_ (.A(_06102_),
    .B(_06103_),
    .Y(_06104_));
 sky130_fd_sc_hd__a22o_1 _12445_ (.A1(net960),
    .A2(_03947_),
    .B1(_03944_),
    .B2(_06104_),
    .X(_01085_));
 sky130_fd_sc_hd__dfrtp_1 _12446_ (.CLK(clknet_leaf_99_clk),
    .D(net219),
    .RESET_B(net168),
    .Q(net19));
 sky130_fd_sc_hd__dfrtp_1 _12447_ (.CLK(clknet_leaf_106_clk),
    .D(net940),
    .RESET_B(net153),
    .Q(\sig_norm.i[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12448_ (.CLK(clknet_leaf_105_clk),
    .D(_00027_),
    .RESET_B(net153),
    .Q(\sig_norm.i[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12449_ (.CLK(clknet_leaf_106_clk),
    .D(net766),
    .RESET_B(net153),
    .Q(\sig_norm.i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12450_ (.CLK(clknet_leaf_107_clk),
    .D(_00029_),
    .RESET_B(net153),
    .Q(\sig_norm.i[3] ));
 sky130_fd_sc_hd__dfrtp_4 _12451_ (.CLK(clknet_4_0_0_clk),
    .D(net6),
    .RESET_B(net38),
    .Q(\modein.delay_in[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12452_ (.CLK(clknet_leaf_116_clk),
    .D(net222),
    .RESET_B(net150),
    .Q(\modein.delay_in[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12453_ (.CLK(clknet_leaf_42_clk),
    .D(net5),
    .RESET_B(net123),
    .Q(\modein.delay_octave_up_in[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12454_ (.CLK(clknet_leaf_39_clk),
    .D(net228),
    .RESET_B(net115),
    .Q(\modein.delay_octave_up_in[1] ));
 sky130_fd_sc_hd__dfrtp_2 _12455_ (.CLK(clknet_leaf_33_clk),
    .D(net4),
    .RESET_B(net101),
    .Q(\modein.delay_octave_down_in[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12456_ (.CLK(clknet_leaf_20_clk),
    .D(net225),
    .RESET_B(net108),
    .Q(\modein.delay_octave_down_in[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12457_ (.CLK(clknet_leaf_106_clk),
    .D(_00030_),
    .RESET_B(net155),
    .Q(\PWM.final_sample_in[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12458_ (.CLK(clknet_leaf_104_clk),
    .D(_00031_),
    .RESET_B(net155),
    .Q(\PWM.final_sample_in[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12459_ (.CLK(clknet_leaf_104_clk),
    .D(_00032_),
    .RESET_B(net153),
    .Q(\PWM.final_sample_in[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12460_ (.CLK(clknet_leaf_104_clk),
    .D(_00033_),
    .RESET_B(net155),
    .Q(\PWM.final_sample_in[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12461_ (.CLK(clknet_leaf_104_clk),
    .D(_00034_),
    .RESET_B(net155),
    .Q(\PWM.final_sample_in[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12462_ (.CLK(clknet_leaf_104_clk),
    .D(_00035_),
    .RESET_B(net155),
    .Q(\PWM.final_sample_in[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12463_ (.CLK(clknet_leaf_103_clk),
    .D(_00036_),
    .RESET_B(net156),
    .Q(\PWM.final_sample_in[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12464_ (.CLK(clknet_leaf_103_clk),
    .D(_00037_),
    .RESET_B(net156),
    .Q(\PWM.final_sample_in[7] ));
 sky130_fd_sc_hd__dfrtp_4 _12465_ (.CLK(clknet_leaf_31_clk),
    .D(\smpl_rt_clkdiv.clkDiv_inst.next_hzX ),
    .RESET_B(net99),
    .Q(\genblk2[0].wave_shpr.div.start ));
 sky130_fd_sc_hd__dfrtp_1 _12466_ (.CLK(clknet_leaf_33_clk),
    .D(\smpl_rt_clkdiv.clkDiv_inst.next_cnt[0] ),
    .RESET_B(net101),
    .Q(\smpl_rt_clkdiv.clkDiv_inst.cnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12467_ (.CLK(clknet_leaf_33_clk),
    .D(\smpl_rt_clkdiv.clkDiv_inst.next_cnt[1] ),
    .RESET_B(net99),
    .Q(\smpl_rt_clkdiv.clkDiv_inst.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12468_ (.CLK(clknet_leaf_34_clk),
    .D(\smpl_rt_clkdiv.clkDiv_inst.next_cnt[2] ),
    .RESET_B(net99),
    .Q(\smpl_rt_clkdiv.clkDiv_inst.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12469_ (.CLK(clknet_leaf_33_clk),
    .D(\smpl_rt_clkdiv.clkDiv_inst.next_cnt[3] ),
    .RESET_B(net101),
    .Q(\smpl_rt_clkdiv.clkDiv_inst.cnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12470_ (.CLK(clknet_leaf_33_clk),
    .D(\smpl_rt_clkdiv.clkDiv_inst.next_cnt[4] ),
    .RESET_B(net100),
    .Q(\smpl_rt_clkdiv.clkDiv_inst.cnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12471_ (.CLK(clknet_leaf_31_clk),
    .D(\smpl_rt_clkdiv.clkDiv_inst.next_cnt[5] ),
    .RESET_B(net100),
    .Q(\smpl_rt_clkdiv.clkDiv_inst.cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12472_ (.CLK(clknet_leaf_32_clk),
    .D(\smpl_rt_clkdiv.clkDiv_inst.next_cnt[6] ),
    .RESET_B(net99),
    .Q(\smpl_rt_clkdiv.clkDiv_inst.cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12473_ (.CLK(clknet_leaf_32_clk),
    .D(\smpl_rt_clkdiv.clkDiv_inst.next_cnt[7] ),
    .RESET_B(net99),
    .Q(\smpl_rt_clkdiv.clkDiv_inst.cnt[7] ));
 sky130_fd_sc_hd__dfrtp_4 _12474_ (.CLK(clknet_leaf_116_clk),
    .D(\FSM.next_mode[0] ),
    .RESET_B(net150),
    .Q(net17));
 sky130_fd_sc_hd__dfrtp_4 _12475_ (.CLK(clknet_leaf_116_clk),
    .D(\FSM.next_mode[1] ),
    .RESET_B(net150),
    .Q(net18));
 sky130_fd_sc_hd__dfrtp_1 _12476_ (.CLK(clknet_leaf_106_clk),
    .D(_00038_),
    .RESET_B(net151),
    .Q(\sig_norm.acc[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12477_ (.CLK(clknet_leaf_107_clk),
    .D(_00039_),
    .RESET_B(net152),
    .Q(\sig_norm.acc[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12478_ (.CLK(clknet_leaf_108_clk),
    .D(_00040_),
    .RESET_B(net152),
    .Q(\sig_norm.acc[2] ));
 sky130_fd_sc_hd__dfrtp_2 _12479_ (.CLK(clknet_leaf_108_clk),
    .D(_00041_),
    .RESET_B(net152),
    .Q(\sig_norm.acc[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12480_ (.CLK(clknet_leaf_108_clk),
    .D(_00042_),
    .RESET_B(net152),
    .Q(\sig_norm.acc[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12481_ (.CLK(clknet_leaf_108_clk),
    .D(net1028),
    .RESET_B(net151),
    .Q(\sig_norm.acc[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12482_ (.CLK(clknet_leaf_108_clk),
    .D(_00044_),
    .RESET_B(net151),
    .Q(\sig_norm.acc[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12483_ (.CLK(clknet_leaf_108_clk),
    .D(_00045_),
    .RESET_B(net151),
    .Q(\sig_norm.acc[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12484_ (.CLK(clknet_leaf_107_clk),
    .D(_00046_),
    .RESET_B(net151),
    .Q(\sig_norm.acc[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12485_ (.CLK(clknet_leaf_106_clk),
    .D(_00047_),
    .RESET_B(net151),
    .Q(\sig_norm.acc[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12486_ (.CLK(clknet_leaf_107_clk),
    .D(_00048_),
    .RESET_B(net151),
    .Q(\sig_norm.acc[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12487_ (.CLK(clknet_leaf_108_clk),
    .D(_00049_),
    .RESET_B(net151),
    .Q(\sig_norm.acc[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12488_ (.CLK(clknet_leaf_107_clk),
    .D(_00050_),
    .RESET_B(net151),
    .Q(\sig_norm.acc[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12489_ (.CLK(clknet_leaf_107_clk),
    .D(_00051_),
    .RESET_B(net151),
    .Q(\sig_norm.quo[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12490_ (.CLK(clknet_leaf_109_clk),
    .D(_00052_),
    .RESET_B(net158),
    .Q(\sig_norm.quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12491_ (.CLK(clknet_leaf_107_clk),
    .D(_00053_),
    .RESET_B(net158),
    .Q(\sig_norm.quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12492_ (.CLK(clknet_leaf_107_clk),
    .D(_00054_),
    .RESET_B(net153),
    .Q(\sig_norm.quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12493_ (.CLK(clknet_leaf_107_clk),
    .D(_00055_),
    .RESET_B(net152),
    .Q(\sig_norm.quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12494_ (.CLK(clknet_leaf_106_clk),
    .D(_00056_),
    .RESET_B(net153),
    .Q(\sig_norm.quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12495_ (.CLK(clknet_leaf_104_clk),
    .D(_00057_),
    .RESET_B(net153),
    .Q(\sig_norm.quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12496_ (.CLK(clknet_leaf_102_clk),
    .D(_00058_),
    .RESET_B(net158),
    .Q(\sig_norm.quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12497_ (.CLK(clknet_leaf_102_clk),
    .D(_00059_),
    .RESET_B(net156),
    .Q(\sig_norm.quo[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12498_ (.CLK(clknet_leaf_103_clk),
    .D(_00060_),
    .RESET_B(net156),
    .Q(\sig_norm.quo[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12499_ (.CLK(clknet_leaf_103_clk),
    .D(_00061_),
    .RESET_B(net156),
    .Q(\sig_norm.quo[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12500_ (.CLK(clknet_leaf_102_clk),
    .D(net429),
    .RESET_B(net156),
    .Q(\sig_norm.acc_next[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12501_ (.CLK(clknet_leaf_106_clk),
    .D(_00063_),
    .RESET_B(net153),
    .Q(\PWM.final_in[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12502_ (.CLK(clknet_leaf_106_clk),
    .D(_00064_),
    .RESET_B(net154),
    .Q(\PWM.final_in[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12503_ (.CLK(clknet_leaf_106_clk),
    .D(_00065_),
    .RESET_B(net154),
    .Q(\PWM.final_in[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12504_ (.CLK(clknet_leaf_106_clk),
    .D(_00066_),
    .RESET_B(net154),
    .Q(\PWM.final_in[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12505_ (.CLK(clknet_leaf_104_clk),
    .D(_00067_),
    .RESET_B(net154),
    .Q(\PWM.final_in[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12506_ (.CLK(clknet_leaf_104_clk),
    .D(_00068_),
    .RESET_B(net154),
    .Q(\PWM.final_in[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12507_ (.CLK(clknet_leaf_103_clk),
    .D(_00069_),
    .RESET_B(net156),
    .Q(\PWM.final_in[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12508_ (.CLK(clknet_leaf_103_clk),
    .D(_00070_),
    .RESET_B(net156),
    .Q(\PWM.final_in[7] ));
 sky130_fd_sc_hd__dfrtp_4 _12509_ (.CLK(clknet_leaf_84_clk),
    .D(_00071_),
    .RESET_B(net202),
    .Q(\genblk2[9].wave_shpr.div.i[0] ));
 sky130_fd_sc_hd__dfrtp_2 _12510_ (.CLK(clknet_leaf_84_clk),
    .D(net1040),
    .RESET_B(net202),
    .Q(\genblk2[9].wave_shpr.div.i[1] ));
 sky130_fd_sc_hd__dfrtp_2 _12511_ (.CLK(clknet_leaf_84_clk),
    .D(_00073_),
    .RESET_B(net202),
    .Q(\genblk2[9].wave_shpr.div.i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12512_ (.CLK(clknet_leaf_84_clk),
    .D(_00074_),
    .RESET_B(net202),
    .Q(\genblk2[9].wave_shpr.div.i[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12513_ (.CLK(clknet_leaf_84_clk),
    .D(_00075_),
    .RESET_B(net202),
    .Q(\genblk2[9].wave_shpr.div.i[4] ));
 sky130_fd_sc_hd__dfrtp_4 _12514_ (.CLK(clknet_leaf_106_clk),
    .D(_00025_),
    .RESET_B(net153),
    .Q(\PWM.start ));
 sky130_fd_sc_hd__dfrtp_1 _12515_ (.CLK(clknet_leaf_106_clk),
    .D(_00024_),
    .RESET_B(net154),
    .Q(\sig_norm.busy ));
 sky130_fd_sc_hd__dfrtp_1 _12516_ (.CLK(clknet_leaf_105_clk),
    .D(\PWM.next_counter[0] ),
    .RESET_B(net155),
    .Q(\PWM.counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12517_ (.CLK(clknet_leaf_105_clk),
    .D(\PWM.next_counter[1] ),
    .RESET_B(net155),
    .Q(\PWM.counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12518_ (.CLK(clknet_leaf_105_clk),
    .D(\PWM.next_counter[2] ),
    .RESET_B(net155),
    .Q(\PWM.counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12519_ (.CLK(clknet_leaf_104_clk),
    .D(\PWM.next_counter[3] ),
    .RESET_B(net157),
    .Q(\PWM.counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12520_ (.CLK(clknet_leaf_104_clk),
    .D(\PWM.next_counter[4] ),
    .RESET_B(net157),
    .Q(\PWM.counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12521_ (.CLK(clknet_leaf_103_clk),
    .D(\PWM.next_counter[5] ),
    .RESET_B(net156),
    .Q(\PWM.counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12522_ (.CLK(clknet_leaf_103_clk),
    .D(\PWM.next_counter[6] ),
    .RESET_B(net156),
    .Q(\PWM.counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12523_ (.CLK(clknet_leaf_103_clk),
    .D(\PWM.next_counter[7] ),
    .RESET_B(net157),
    .Q(\PWM.counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12524_ (.CLK(clknet_leaf_59_clk),
    .D(_00076_),
    .RESET_B(net193),
    .Q(\genblk2[0].wave_shpr.div.b1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12525_ (.CLK(clknet_leaf_67_clk),
    .D(_00077_),
    .RESET_B(net194),
    .Q(\genblk2[0].wave_shpr.div.b1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12526_ (.CLK(clknet_leaf_66_clk),
    .D(_00078_),
    .RESET_B(net197),
    .Q(\genblk2[0].wave_shpr.div.b1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12527_ (.CLK(clknet_leaf_67_clk),
    .D(_00079_),
    .RESET_B(net193),
    .Q(\genblk2[0].wave_shpr.div.b1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12528_ (.CLK(clknet_leaf_43_clk),
    .D(_00080_),
    .RESET_B(net124),
    .Q(\genblk2[0].wave_shpr.div.b1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12529_ (.CLK(clknet_leaf_59_clk),
    .D(_00081_),
    .RESET_B(net187),
    .Q(\genblk2[0].wave_shpr.div.b1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12530_ (.CLK(clknet_leaf_61_clk),
    .D(_00082_),
    .RESET_B(net188),
    .Q(\genblk2[0].wave_shpr.div.b1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12531_ (.CLK(clknet_leaf_61_clk),
    .D(_00083_),
    .RESET_B(net186),
    .Q(\genblk2[0].wave_shpr.div.b1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12532_ (.CLK(clknet_leaf_61_clk),
    .D(_00084_),
    .RESET_B(net186),
    .Q(\genblk2[0].wave_shpr.div.b1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12533_ (.CLK(clknet_leaf_61_clk),
    .D(_00085_),
    .RESET_B(net186),
    .Q(\genblk2[0].wave_shpr.div.b1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12534_ (.CLK(clknet_leaf_45_clk),
    .D(_00086_),
    .RESET_B(net186),
    .Q(\genblk2[0].wave_shpr.div.b1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12535_ (.CLK(clknet_leaf_45_clk),
    .D(_00087_),
    .RESET_B(net186),
    .Q(\genblk2[0].wave_shpr.div.b1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12536_ (.CLK(clknet_leaf_44_clk),
    .D(_00088_),
    .RESET_B(net123),
    .Q(\genblk2[0].wave_shpr.div.b1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12537_ (.CLK(clknet_leaf_41_clk),
    .D(_00089_),
    .RESET_B(net123),
    .Q(\genblk2[0].wave_shpr.div.b1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12538_ (.CLK(clknet_leaf_63_clk),
    .D(_00090_),
    .RESET_B(net190),
    .Q(\genblk2[0].wave_shpr.div.b1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12539_ (.CLK(clknet_leaf_62_clk),
    .D(_00091_),
    .RESET_B(net189),
    .Q(\genblk2[0].wave_shpr.div.b1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12540_ (.CLK(clknet_leaf_62_clk),
    .D(_00092_),
    .RESET_B(net189),
    .Q(\genblk2[0].wave_shpr.div.b1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12541_ (.CLK(clknet_leaf_64_clk),
    .D(_00093_),
    .RESET_B(net189),
    .Q(\genblk2[0].wave_shpr.div.b1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12542_ (.CLK(clknet_leaf_100_clk),
    .D(net287),
    .RESET_B(net164),
    .Q(\PWM.pwm_out ));
 sky130_fd_sc_hd__dfrtp_4 _12543_ (.CLK(clknet_leaf_60_clk),
    .D(\genblk1[0].osc.clkdiv_C.next_cnt[0] ),
    .RESET_B(net187),
    .Q(\genblk1[0].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _12544_ (.CLK(clknet_leaf_60_clk),
    .D(\genblk1[0].osc.clkdiv_C.next_cnt[1] ),
    .RESET_B(net192),
    .Q(\genblk1[0].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _12545_ (.CLK(clknet_leaf_60_clk),
    .D(\genblk1[0].osc.clkdiv_C.next_cnt[2] ),
    .RESET_B(net187),
    .Q(\genblk1[0].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_4 _12546_ (.CLK(clknet_leaf_61_clk),
    .D(\genblk1[0].osc.clkdiv_C.next_cnt[3] ),
    .RESET_B(net188),
    .Q(\genblk1[0].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__dfrtp_4 _12547_ (.CLK(clknet_leaf_61_clk),
    .D(\genblk1[0].osc.clkdiv_C.next_cnt[4] ),
    .RESET_B(net186),
    .Q(\genblk1[0].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__dfrtp_4 _12548_ (.CLK(clknet_leaf_61_clk),
    .D(\genblk1[0].osc.clkdiv_C.next_cnt[5] ),
    .RESET_B(net186),
    .Q(\genblk1[0].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__dfrtp_2 _12549_ (.CLK(clknet_leaf_60_clk),
    .D(\genblk1[0].osc.clkdiv_C.next_cnt[6] ),
    .RESET_B(net186),
    .Q(\genblk1[0].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__dfrtp_4 _12550_ (.CLK(clknet_leaf_60_clk),
    .D(\genblk1[0].osc.clkdiv_C.next_cnt[7] ),
    .RESET_B(net186),
    .Q(\genblk1[0].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__dfrtp_4 _12551_ (.CLK(clknet_leaf_60_clk),
    .D(\genblk1[0].osc.clkdiv_C.next_cnt[8] ),
    .RESET_B(net187),
    .Q(\genblk1[0].osc.clkdiv_C.cnt[8] ));
 sky130_fd_sc_hd__dfrtp_4 _12552_ (.CLK(clknet_leaf_60_clk),
    .D(\genblk1[0].osc.clkdiv_C.next_cnt[9] ),
    .RESET_B(net186),
    .Q(\genblk1[0].osc.clkdiv_C.cnt[9] ));
 sky130_fd_sc_hd__dfrtp_4 _12553_ (.CLK(clknet_leaf_55_clk),
    .D(\genblk1[0].osc.clkdiv_C.next_cnt[10] ),
    .RESET_B(net176),
    .Q(\genblk1[0].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__dfrtp_4 _12554_ (.CLK(clknet_leaf_55_clk),
    .D(\genblk1[0].osc.clkdiv_C.next_cnt[11] ),
    .RESET_B(net175),
    .Q(\genblk1[0].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__dfrtp_4 _12555_ (.CLK(clknet_leaf_55_clk),
    .D(\genblk1[0].osc.clkdiv_C.next_cnt[12] ),
    .RESET_B(net175),
    .Q(\genblk1[0].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__dfrtp_4 _12556_ (.CLK(clknet_leaf_55_clk),
    .D(\genblk1[0].osc.clkdiv_C.next_cnt[13] ),
    .RESET_B(net175),
    .Q(\genblk1[0].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__dfrtp_4 _12557_ (.CLK(clknet_leaf_55_clk),
    .D(\genblk1[0].osc.clkdiv_C.next_cnt[14] ),
    .RESET_B(net175),
    .Q(\genblk1[0].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__dfrtp_4 _12558_ (.CLK(clknet_leaf_55_clk),
    .D(\genblk1[0].osc.clkdiv_C.next_cnt[15] ),
    .RESET_B(net176),
    .Q(\genblk1[0].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__dfrtp_4 _12559_ (.CLK(clknet_leaf_56_clk),
    .D(\genblk1[0].osc.clkdiv_C.next_cnt[16] ),
    .RESET_B(net181),
    .Q(\genblk1[0].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__dfrtp_4 _12560_ (.CLK(clknet_leaf_57_clk),
    .D(\genblk1[0].osc.clkdiv_C.next_cnt[17] ),
    .RESET_B(net181),
    .Q(\genblk1[0].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__dfrtp_4 _12561_ (.CLK(clknet_leaf_29_clk),
    .D(\genblk1[1].osc.clkdiv_C.next_cnt[0] ),
    .RESET_B(net96),
    .Q(\genblk1[1].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _12562_ (.CLK(clknet_leaf_30_clk),
    .D(\genblk1[1].osc.clkdiv_C.next_cnt[1] ),
    .RESET_B(net96),
    .Q(\genblk1[1].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_2 _12563_ (.CLK(clknet_leaf_30_clk),
    .D(\genblk1[1].osc.clkdiv_C.next_cnt[2] ),
    .RESET_B(net96),
    .Q(\genblk1[1].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_4 _12564_ (.CLK(clknet_leaf_29_clk),
    .D(\genblk1[1].osc.clkdiv_C.next_cnt[3] ),
    .RESET_B(net96),
    .Q(\genblk1[1].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__dfrtp_4 _12565_ (.CLK(clknet_leaf_28_clk),
    .D(\genblk1[1].osc.clkdiv_C.next_cnt[4] ),
    .RESET_B(net89),
    .Q(\genblk1[1].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__dfrtp_4 _12566_ (.CLK(clknet_leaf_28_clk),
    .D(\genblk1[1].osc.clkdiv_C.next_cnt[5] ),
    .RESET_B(net89),
    .Q(\genblk1[1].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__dfrtp_2 _12567_ (.CLK(clknet_leaf_27_clk),
    .D(\genblk1[1].osc.clkdiv_C.next_cnt[6] ),
    .RESET_B(net89),
    .Q(\genblk1[1].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__dfrtp_4 _12568_ (.CLK(clknet_leaf_27_clk),
    .D(\genblk1[1].osc.clkdiv_C.next_cnt[7] ),
    .RESET_B(net90),
    .Q(\genblk1[1].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__dfrtp_4 _12569_ (.CLK(clknet_leaf_27_clk),
    .D(\genblk1[1].osc.clkdiv_C.next_cnt[8] ),
    .RESET_B(net90),
    .Q(\genblk1[1].osc.clkdiv_C.cnt[8] ));
 sky130_fd_sc_hd__dfrtp_4 _12570_ (.CLK(clknet_leaf_28_clk),
    .D(\genblk1[1].osc.clkdiv_C.next_cnt[9] ),
    .RESET_B(net90),
    .Q(\genblk1[1].osc.clkdiv_C.cnt[9] ));
 sky130_fd_sc_hd__dfrtp_4 _12571_ (.CLK(clknet_leaf_28_clk),
    .D(\genblk1[1].osc.clkdiv_C.next_cnt[10] ),
    .RESET_B(net89),
    .Q(\genblk1[1].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__dfrtp_4 _12572_ (.CLK(clknet_leaf_28_clk),
    .D(\genblk1[1].osc.clkdiv_C.next_cnt[11] ),
    .RESET_B(net89),
    .Q(\genblk1[1].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__dfrtp_4 _12573_ (.CLK(clknet_leaf_29_clk),
    .D(\genblk1[1].osc.clkdiv_C.next_cnt[12] ),
    .RESET_B(net89),
    .Q(\genblk1[1].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__dfrtp_4 _12574_ (.CLK(clknet_leaf_29_clk),
    .D(\genblk1[1].osc.clkdiv_C.next_cnt[13] ),
    .RESET_B(net89),
    .Q(\genblk1[1].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__dfrtp_4 _12575_ (.CLK(clknet_leaf_29_clk),
    .D(\genblk1[1].osc.clkdiv_C.next_cnt[14] ),
    .RESET_B(net95),
    .Q(\genblk1[1].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__dfrtp_4 _12576_ (.CLK(clknet_leaf_29_clk),
    .D(\genblk1[1].osc.clkdiv_C.next_cnt[15] ),
    .RESET_B(net95),
    .Q(\genblk1[1].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__dfrtp_4 _12577_ (.CLK(clknet_leaf_21_clk),
    .D(\genblk1[1].osc.clkdiv_C.next_cnt[16] ),
    .RESET_B(net95),
    .Q(\genblk1[1].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__dfrtp_4 _12578_ (.CLK(clknet_leaf_29_clk),
    .D(\genblk1[1].osc.clkdiv_C.next_cnt[17] ),
    .RESET_B(net96),
    .Q(\genblk1[1].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__dfrtp_4 _12579_ (.CLK(clknet_leaf_14_clk),
    .D(\genblk1[2].osc.clkdiv_C.next_cnt[0] ),
    .RESET_B(net70),
    .Q(\genblk1[2].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _12580_ (.CLK(clknet_leaf_14_clk),
    .D(\genblk1[2].osc.clkdiv_C.next_cnt[1] ),
    .RESET_B(net70),
    .Q(\genblk1[2].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _12581_ (.CLK(clknet_leaf_14_clk),
    .D(\genblk1[2].osc.clkdiv_C.next_cnt[2] ),
    .RESET_B(net70),
    .Q(\genblk1[2].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_2 _12582_ (.CLK(clknet_leaf_14_clk),
    .D(\genblk1[2].osc.clkdiv_C.next_cnt[3] ),
    .RESET_B(net74),
    .Q(\genblk1[2].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__dfrtp_4 _12583_ (.CLK(clknet_leaf_124_clk),
    .D(\genblk1[2].osc.clkdiv_C.next_cnt[4] ),
    .RESET_B(net72),
    .Q(\genblk1[2].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__dfrtp_2 _12584_ (.CLK(clknet_leaf_124_clk),
    .D(\genblk1[2].osc.clkdiv_C.next_cnt[5] ),
    .RESET_B(net76),
    .Q(\genblk1[2].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__dfrtp_2 _12585_ (.CLK(clknet_leaf_124_clk),
    .D(\genblk1[2].osc.clkdiv_C.next_cnt[6] ),
    .RESET_B(net76),
    .Q(\genblk1[2].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__dfrtp_4 _12586_ (.CLK(clknet_leaf_14_clk),
    .D(\genblk1[2].osc.clkdiv_C.next_cnt[7] ),
    .RESET_B(net74),
    .Q(\genblk1[2].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12587_ (.CLK(clknet_leaf_14_clk),
    .D(\genblk1[2].osc.clkdiv_C.next_cnt[8] ),
    .RESET_B(net72),
    .Q(\genblk1[2].osc.clkdiv_C.cnt[8] ));
 sky130_fd_sc_hd__dfrtp_4 _12588_ (.CLK(clknet_leaf_14_clk),
    .D(\genblk1[2].osc.clkdiv_C.next_cnt[9] ),
    .RESET_B(net72),
    .Q(\genblk1[2].osc.clkdiv_C.cnt[9] ));
 sky130_fd_sc_hd__dfrtp_2 _12589_ (.CLK(clknet_leaf_14_clk),
    .D(\genblk1[2].osc.clkdiv_C.next_cnt[10] ),
    .RESET_B(net72),
    .Q(\genblk1[2].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__dfrtp_4 _12590_ (.CLK(clknet_leaf_13_clk),
    .D(\genblk1[2].osc.clkdiv_C.next_cnt[11] ),
    .RESET_B(net70),
    .Q(\genblk1[2].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__dfrtp_4 _12591_ (.CLK(clknet_leaf_13_clk),
    .D(\genblk1[2].osc.clkdiv_C.next_cnt[12] ),
    .RESET_B(net70),
    .Q(\genblk1[2].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__dfrtp_2 _12592_ (.CLK(clknet_leaf_13_clk),
    .D(\genblk1[2].osc.clkdiv_C.next_cnt[13] ),
    .RESET_B(net70),
    .Q(\genblk1[2].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__dfrtp_4 _12593_ (.CLK(clknet_leaf_13_clk),
    .D(\genblk1[2].osc.clkdiv_C.next_cnt[14] ),
    .RESET_B(net70),
    .Q(\genblk1[2].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__dfrtp_2 _12594_ (.CLK(clknet_leaf_12_clk),
    .D(\genblk1[2].osc.clkdiv_C.next_cnt[15] ),
    .RESET_B(net52),
    .Q(\genblk1[2].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__dfrtp_4 _12595_ (.CLK(clknet_leaf_11_clk),
    .D(\genblk1[2].osc.clkdiv_C.next_cnt[16] ),
    .RESET_B(net56),
    .Q(\genblk1[2].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__dfrtp_2 _12596_ (.CLK(clknet_leaf_15_clk),
    .D(\genblk1[2].osc.clkdiv_C.next_cnt[17] ),
    .RESET_B(net73),
    .Q(\genblk1[2].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__dfrtp_4 _12597_ (.CLK(clknet_leaf_21_clk),
    .D(\genblk1[3].osc.clkdiv_C.next_cnt[0] ),
    .RESET_B(net97),
    .Q(\genblk1[3].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _12598_ (.CLK(clknet_leaf_21_clk),
    .D(\genblk1[3].osc.clkdiv_C.next_cnt[1] ),
    .RESET_B(net97),
    .Q(\genblk1[3].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _12599_ (.CLK(clknet_leaf_21_clk),
    .D(\genblk1[3].osc.clkdiv_C.next_cnt[2] ),
    .RESET_B(net97),
    .Q(\genblk1[3].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_2 _12600_ (.CLK(clknet_leaf_21_clk),
    .D(\genblk1[3].osc.clkdiv_C.next_cnt[3] ),
    .RESET_B(net97),
    .Q(\genblk1[3].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__dfrtp_4 _12601_ (.CLK(clknet_leaf_21_clk),
    .D(\genblk1[3].osc.clkdiv_C.next_cnt[4] ),
    .RESET_B(net97),
    .Q(\genblk1[3].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__dfrtp_4 _12602_ (.CLK(clknet_leaf_21_clk),
    .D(\genblk1[3].osc.clkdiv_C.next_cnt[5] ),
    .RESET_B(net95),
    .Q(\genblk1[3].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__dfrtp_4 _12603_ (.CLK(clknet_leaf_21_clk),
    .D(\genblk1[3].osc.clkdiv_C.next_cnt[6] ),
    .RESET_B(net97),
    .Q(\genblk1[3].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__dfrtp_4 _12604_ (.CLK(clknet_leaf_21_clk),
    .D(\genblk1[3].osc.clkdiv_C.next_cnt[7] ),
    .RESET_B(net97),
    .Q(\genblk1[3].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__dfrtp_4 _12605_ (.CLK(clknet_leaf_22_clk),
    .D(\genblk1[3].osc.clkdiv_C.next_cnt[8] ),
    .RESET_B(net94),
    .Q(\genblk1[3].osc.clkdiv_C.cnt[8] ));
 sky130_fd_sc_hd__dfrtp_2 _12606_ (.CLK(clknet_leaf_22_clk),
    .D(\genblk1[3].osc.clkdiv_C.next_cnt[9] ),
    .RESET_B(net92),
    .Q(\genblk1[3].osc.clkdiv_C.cnt[9] ));
 sky130_fd_sc_hd__dfrtp_4 _12607_ (.CLK(clknet_leaf_22_clk),
    .D(\genblk1[3].osc.clkdiv_C.next_cnt[10] ),
    .RESET_B(net94),
    .Q(\genblk1[3].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12608_ (.CLK(clknet_leaf_23_clk),
    .D(\genblk1[3].osc.clkdiv_C.next_cnt[11] ),
    .RESET_B(net94),
    .Q(\genblk1[3].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__dfrtp_4 _12609_ (.CLK(clknet_leaf_22_clk),
    .D(\genblk1[3].osc.clkdiv_C.next_cnt[12] ),
    .RESET_B(net94),
    .Q(\genblk1[3].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__dfrtp_4 _12610_ (.CLK(clknet_leaf_22_clk),
    .D(\genblk1[3].osc.clkdiv_C.next_cnt[13] ),
    .RESET_B(net93),
    .Q(\genblk1[3].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__dfrtp_4 _12611_ (.CLK(clknet_leaf_23_clk),
    .D(\genblk1[3].osc.clkdiv_C.next_cnt[14] ),
    .RESET_B(net94),
    .Q(\genblk1[3].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__dfrtp_4 _12612_ (.CLK(clknet_leaf_23_clk),
    .D(\genblk1[3].osc.clkdiv_C.next_cnt[15] ),
    .RESET_B(net94),
    .Q(\genblk1[3].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__dfrtp_2 _12613_ (.CLK(clknet_leaf_23_clk),
    .D(\genblk1[3].osc.clkdiv_C.next_cnt[16] ),
    .RESET_B(net94),
    .Q(\genblk1[3].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12614_ (.CLK(clknet_leaf_23_clk),
    .D(\genblk1[3].osc.clkdiv_C.next_cnt[17] ),
    .RESET_B(net109),
    .Q(\genblk1[3].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__dfrtp_4 _12615_ (.CLK(clknet_leaf_121_clk),
    .D(\genblk1[4].osc.clkdiv_C.next_cnt[0] ),
    .RESET_B(net81),
    .Q(\genblk1[4].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _12616_ (.CLK(clknet_leaf_18_clk),
    .D(\genblk1[4].osc.clkdiv_C.next_cnt[1] ),
    .RESET_B(net80),
    .Q(\genblk1[4].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _12617_ (.CLK(clknet_leaf_18_clk),
    .D(\genblk1[4].osc.clkdiv_C.next_cnt[2] ),
    .RESET_B(net80),
    .Q(\genblk1[4].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_4 _12618_ (.CLK(clknet_leaf_17_clk),
    .D(\genblk1[4].osc.clkdiv_C.next_cnt[3] ),
    .RESET_B(net80),
    .Q(\genblk1[4].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__dfrtp_4 _12619_ (.CLK(clknet_leaf_17_clk),
    .D(\genblk1[4].osc.clkdiv_C.next_cnt[4] ),
    .RESET_B(net83),
    .Q(\genblk1[4].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__dfrtp_4 _12620_ (.CLK(clknet_leaf_17_clk),
    .D(\genblk1[4].osc.clkdiv_C.next_cnt[5] ),
    .RESET_B(net83),
    .Q(\genblk1[4].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__dfrtp_4 _12621_ (.CLK(clknet_leaf_17_clk),
    .D(\genblk1[4].osc.clkdiv_C.next_cnt[6] ),
    .RESET_B(net80),
    .Q(\genblk1[4].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__dfrtp_4 _12622_ (.CLK(clknet_leaf_17_clk),
    .D(\genblk1[4].osc.clkdiv_C.next_cnt[7] ),
    .RESET_B(net83),
    .Q(\genblk1[4].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__dfrtp_4 _12623_ (.CLK(clknet_leaf_16_clk),
    .D(\genblk1[4].osc.clkdiv_C.next_cnt[8] ),
    .RESET_B(net74),
    .Q(\genblk1[4].osc.clkdiv_C.cnt[8] ));
 sky130_fd_sc_hd__dfrtp_4 _12624_ (.CLK(clknet_leaf_19_clk),
    .D(\genblk1[4].osc.clkdiv_C.next_cnt[9] ),
    .RESET_B(net109),
    .Q(\genblk1[4].osc.clkdiv_C.cnt[9] ));
 sky130_fd_sc_hd__dfrtp_4 _12625_ (.CLK(clknet_leaf_16_clk),
    .D(\genblk1[4].osc.clkdiv_C.next_cnt[10] ),
    .RESET_B(net74),
    .Q(\genblk1[4].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__dfrtp_4 _12626_ (.CLK(clknet_leaf_16_clk),
    .D(\genblk1[4].osc.clkdiv_C.next_cnt[11] ),
    .RESET_B(net74),
    .Q(\genblk1[4].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__dfrtp_4 _12627_ (.CLK(clknet_leaf_120_clk),
    .D(\genblk1[4].osc.clkdiv_C.next_cnt[12] ),
    .RESET_B(net81),
    .Q(\genblk1[4].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__dfrtp_4 _12628_ (.CLK(clknet_leaf_18_clk),
    .D(\genblk1[4].osc.clkdiv_C.next_cnt[13] ),
    .RESET_B(net81),
    .Q(\genblk1[4].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__dfrtp_4 _12629_ (.CLK(clknet_leaf_120_clk),
    .D(\genblk1[4].osc.clkdiv_C.next_cnt[14] ),
    .RESET_B(net82),
    .Q(\genblk1[4].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__dfrtp_2 _12630_ (.CLK(clknet_leaf_18_clk),
    .D(\genblk1[4].osc.clkdiv_C.next_cnt[15] ),
    .RESET_B(net82),
    .Q(\genblk1[4].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__dfrtp_4 _12631_ (.CLK(clknet_leaf_18_clk),
    .D(\genblk1[4].osc.clkdiv_C.next_cnt[16] ),
    .RESET_B(net112),
    .Q(\genblk1[4].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__dfrtp_2 _12632_ (.CLK(clknet_leaf_18_clk),
    .D(\genblk1[4].osc.clkdiv_C.next_cnt[17] ),
    .RESET_B(net112),
    .Q(\genblk1[4].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__dfrtp_4 _12633_ (.CLK(clknet_leaf_16_clk),
    .D(\genblk1[5].osc.clkdiv_C.next_cnt[0] ),
    .RESET_B(net74),
    .Q(\genblk1[5].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _12634_ (.CLK(clknet_leaf_16_clk),
    .D(\genblk1[5].osc.clkdiv_C.next_cnt[1] ),
    .RESET_B(net74),
    .Q(\genblk1[5].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _12635_ (.CLK(clknet_leaf_16_clk),
    .D(\genblk1[5].osc.clkdiv_C.next_cnt[2] ),
    .RESET_B(net74),
    .Q(\genblk1[5].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_4 _12636_ (.CLK(clknet_leaf_19_clk),
    .D(\genblk1[5].osc.clkdiv_C.next_cnt[3] ),
    .RESET_B(net109),
    .Q(\genblk1[5].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__dfrtp_4 _12637_ (.CLK(clknet_leaf_16_clk),
    .D(\genblk1[5].osc.clkdiv_C.next_cnt[4] ),
    .RESET_B(net73),
    .Q(\genblk1[5].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__dfrtp_2 _12638_ (.CLK(clknet_leaf_19_clk),
    .D(\genblk1[5].osc.clkdiv_C.next_cnt[5] ),
    .RESET_B(net109),
    .Q(\genblk1[5].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__dfrtp_4 _12639_ (.CLK(clknet_leaf_16_clk),
    .D(\genblk1[5].osc.clkdiv_C.next_cnt[6] ),
    .RESET_B(net73),
    .Q(\genblk1[5].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__dfrtp_4 _12640_ (.CLK(clknet_leaf_15_clk),
    .D(\genblk1[5].osc.clkdiv_C.next_cnt[7] ),
    .RESET_B(net73),
    .Q(\genblk1[5].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__dfrtp_2 _12641_ (.CLK(clknet_leaf_10_clk),
    .D(\genblk1[5].osc.clkdiv_C.next_cnt[8] ),
    .RESET_B(net56),
    .Q(\genblk1[5].osc.clkdiv_C.cnt[8] ));
 sky130_fd_sc_hd__dfrtp_2 _12642_ (.CLK(clknet_leaf_10_clk),
    .D(\genblk1[5].osc.clkdiv_C.next_cnt[9] ),
    .RESET_B(net56),
    .Q(\genblk1[5].osc.clkdiv_C.cnt[9] ));
 sky130_fd_sc_hd__dfrtp_4 _12643_ (.CLK(clknet_leaf_10_clk),
    .D(\genblk1[5].osc.clkdiv_C.next_cnt[10] ),
    .RESET_B(net56),
    .Q(\genblk1[5].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__dfrtp_4 _12644_ (.CLK(clknet_leaf_10_clk),
    .D(\genblk1[5].osc.clkdiv_C.next_cnt[11] ),
    .RESET_B(net57),
    .Q(\genblk1[5].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__dfrtp_4 _12645_ (.CLK(clknet_leaf_24_clk),
    .D(\genblk1[5].osc.clkdiv_C.next_cnt[12] ),
    .RESET_B(net92),
    .Q(\genblk1[5].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__dfrtp_4 _12646_ (.CLK(clknet_leaf_24_clk),
    .D(\genblk1[5].osc.clkdiv_C.next_cnt[13] ),
    .RESET_B(net92),
    .Q(\genblk1[5].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__dfrtp_4 _12647_ (.CLK(clknet_leaf_9_clk),
    .D(\genblk1[5].osc.clkdiv_C.next_cnt[14] ),
    .RESET_B(net54),
    .Q(\genblk1[5].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__dfrtp_2 _12648_ (.CLK(clknet_leaf_9_clk),
    .D(\genblk1[5].osc.clkdiv_C.next_cnt[15] ),
    .RESET_B(net54),
    .Q(\genblk1[5].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__dfrtp_4 _12649_ (.CLK(clknet_leaf_10_clk),
    .D(\genblk1[5].osc.clkdiv_C.next_cnt[16] ),
    .RESET_B(net55),
    .Q(\genblk1[5].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12650_ (.CLK(clknet_leaf_10_clk),
    .D(\genblk1[5].osc.clkdiv_C.next_cnt[17] ),
    .RESET_B(net57),
    .Q(\genblk1[5].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__dfrtp_4 _12651_ (.CLK(clknet_leaf_28_clk),
    .D(\genblk1[6].osc.clkdiv_C.next_cnt[0] ),
    .RESET_B(net89),
    .Q(\genblk1[6].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _12652_ (.CLK(clknet_leaf_27_clk),
    .D(\genblk1[6].osc.clkdiv_C.next_cnt[1] ),
    .RESET_B(net89),
    .Q(\genblk1[6].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12653_ (.CLK(clknet_leaf_27_clk),
    .D(\genblk1[6].osc.clkdiv_C.next_cnt[2] ),
    .RESET_B(net89),
    .Q(\genblk1[6].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_4 _12654_ (.CLK(clknet_leaf_27_clk),
    .D(\genblk1[6].osc.clkdiv_C.next_cnt[3] ),
    .RESET_B(net90),
    .Q(\genblk1[6].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__dfrtp_4 _12655_ (.CLK(clknet_leaf_27_clk),
    .D(\genblk1[6].osc.clkdiv_C.next_cnt[4] ),
    .RESET_B(net90),
    .Q(\genblk1[6].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__dfrtp_4 _12656_ (.CLK(clknet_leaf_27_clk),
    .D(\genblk1[6].osc.clkdiv_C.next_cnt[5] ),
    .RESET_B(net90),
    .Q(\genblk1[6].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__dfrtp_2 _12657_ (.CLK(clknet_leaf_27_clk),
    .D(\genblk1[6].osc.clkdiv_C.next_cnt[6] ),
    .RESET_B(net90),
    .Q(\genblk1[6].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__dfrtp_4 _12658_ (.CLK(clknet_leaf_27_clk),
    .D(\genblk1[6].osc.clkdiv_C.next_cnt[7] ),
    .RESET_B(net90),
    .Q(\genblk1[6].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__dfrtp_4 _12659_ (.CLK(clknet_leaf_27_clk),
    .D(\genblk1[6].osc.clkdiv_C.next_cnt[8] ),
    .RESET_B(net90),
    .Q(\genblk1[6].osc.clkdiv_C.cnt[8] ));
 sky130_fd_sc_hd__dfrtp_4 _12660_ (.CLK(clknet_leaf_26_clk),
    .D(\genblk1[6].osc.clkdiv_C.next_cnt[9] ),
    .RESET_B(net87),
    .Q(\genblk1[6].osc.clkdiv_C.cnt[9] ));
 sky130_fd_sc_hd__dfrtp_4 _12661_ (.CLK(clknet_leaf_26_clk),
    .D(\genblk1[6].osc.clkdiv_C.next_cnt[10] ),
    .RESET_B(net88),
    .Q(\genblk1[6].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__dfrtp_4 _12662_ (.CLK(clknet_leaf_25_clk),
    .D(\genblk1[6].osc.clkdiv_C.next_cnt[11] ),
    .RESET_B(net87),
    .Q(\genblk1[6].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__dfrtp_4 _12663_ (.CLK(clknet_leaf_26_clk),
    .D(\genblk1[6].osc.clkdiv_C.next_cnt[12] ),
    .RESET_B(net88),
    .Q(\genblk1[6].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__dfrtp_4 _12664_ (.CLK(clknet_leaf_26_clk),
    .D(\genblk1[6].osc.clkdiv_C.next_cnt[13] ),
    .RESET_B(net88),
    .Q(\genblk1[6].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__dfrtp_4 _12665_ (.CLK(clknet_leaf_25_clk),
    .D(\genblk1[6].osc.clkdiv_C.next_cnt[14] ),
    .RESET_B(net86),
    .Q(\genblk1[6].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__dfrtp_4 _12666_ (.CLK(clknet_leaf_25_clk),
    .D(\genblk1[6].osc.clkdiv_C.next_cnt[15] ),
    .RESET_B(net88),
    .Q(\genblk1[6].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__dfrtp_2 _12667_ (.CLK(clknet_leaf_24_clk),
    .D(\genblk1[6].osc.clkdiv_C.next_cnt[16] ),
    .RESET_B(net88),
    .Q(\genblk1[6].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12668_ (.CLK(clknet_leaf_24_clk),
    .D(\genblk1[6].osc.clkdiv_C.next_cnt[17] ),
    .RESET_B(net92),
    .Q(\genblk1[6].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__dfrtp_2 _12669_ (.CLK(clknet_leaf_90_clk),
    .D(\genblk1[7].osc.clkdiv_C.next_cnt[0] ),
    .RESET_B(net173),
    .Q(\genblk1[7].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _12670_ (.CLK(clknet_leaf_90_clk),
    .D(\genblk1[7].osc.clkdiv_C.next_cnt[1] ),
    .RESET_B(net173),
    .Q(\genblk1[7].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _12671_ (.CLK(clknet_leaf_89_clk),
    .D(\genblk1[7].osc.clkdiv_C.next_cnt[2] ),
    .RESET_B(net173),
    .Q(\genblk1[7].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_2 _12672_ (.CLK(clknet_leaf_90_clk),
    .D(\genblk1[7].osc.clkdiv_C.next_cnt[3] ),
    .RESET_B(net173),
    .Q(\genblk1[7].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__dfrtp_4 _12673_ (.CLK(clknet_leaf_90_clk),
    .D(\genblk1[7].osc.clkdiv_C.next_cnt[4] ),
    .RESET_B(net173),
    .Q(\genblk1[7].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__dfrtp_2 _12674_ (.CLK(clknet_leaf_90_clk),
    .D(\genblk1[7].osc.clkdiv_C.next_cnt[5] ),
    .RESET_B(net174),
    .Q(\genblk1[7].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__dfrtp_4 _12675_ (.CLK(clknet_leaf_90_clk),
    .D(\genblk1[7].osc.clkdiv_C.next_cnt[6] ),
    .RESET_B(net141),
    .Q(\genblk1[7].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__dfrtp_4 _12676_ (.CLK(clknet_leaf_120_clk),
    .D(\genblk1[7].osc.clkdiv_C.next_cnt[7] ),
    .RESET_B(net82),
    .Q(\genblk1[7].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__dfrtp_4 _12677_ (.CLK(clknet_leaf_120_clk),
    .D(\genblk1[7].osc.clkdiv_C.next_cnt[8] ),
    .RESET_B(net142),
    .Q(\genblk1[7].osc.clkdiv_C.cnt[8] ));
 sky130_fd_sc_hd__dfrtp_4 _12678_ (.CLK(clknet_leaf_120_clk),
    .D(\genblk1[7].osc.clkdiv_C.next_cnt[9] ),
    .RESET_B(net142),
    .Q(\genblk1[7].osc.clkdiv_C.cnt[9] ));
 sky130_fd_sc_hd__dfrtp_4 _12679_ (.CLK(clknet_leaf_120_clk),
    .D(\genblk1[7].osc.clkdiv_C.next_cnt[10] ),
    .RESET_B(net82),
    .Q(\genblk1[7].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__dfrtp_4 _12680_ (.CLK(clknet_leaf_120_clk),
    .D(\genblk1[7].osc.clkdiv_C.next_cnt[11] ),
    .RESET_B(net82),
    .Q(\genblk1[7].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__dfrtp_2 _12681_ (.CLK(clknet_leaf_120_clk),
    .D(\genblk1[7].osc.clkdiv_C.next_cnt[12] ),
    .RESET_B(net82),
    .Q(\genblk1[7].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__dfrtp_4 _12682_ (.CLK(clknet_leaf_120_clk),
    .D(\genblk1[7].osc.clkdiv_C.next_cnt[13] ),
    .RESET_B(net81),
    .Q(\genblk1[7].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__dfrtp_2 _12683_ (.CLK(clknet_leaf_120_clk),
    .D(\genblk1[7].osc.clkdiv_C.next_cnt[14] ),
    .RESET_B(net81),
    .Q(\genblk1[7].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__dfrtp_4 _12684_ (.CLK(clknet_leaf_120_clk),
    .D(\genblk1[7].osc.clkdiv_C.next_cnt[15] ),
    .RESET_B(net141),
    .Q(\genblk1[7].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__dfrtp_2 _12685_ (.CLK(clknet_leaf_119_clk),
    .D(\genblk1[7].osc.clkdiv_C.next_cnt[16] ),
    .RESET_B(net141),
    .Q(\genblk1[7].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12686_ (.CLK(clknet_leaf_119_clk),
    .D(\genblk1[7].osc.clkdiv_C.next_cnt[17] ),
    .RESET_B(net141),
    .Q(\genblk1[7].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__dfrtp_4 _12687_ (.CLK(clknet_leaf_54_clk),
    .D(\genblk1[8].osc.clkdiv_C.next_cnt[0] ),
    .RESET_B(net174),
    .Q(\genblk1[8].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _12688_ (.CLK(clknet_leaf_53_clk),
    .D(\genblk1[8].osc.clkdiv_C.next_cnt[1] ),
    .RESET_B(net112),
    .Q(\genblk1[8].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12689_ (.CLK(clknet_leaf_53_clk),
    .D(\genblk1[8].osc.clkdiv_C.next_cnt[2] ),
    .RESET_B(net174),
    .Q(\genblk1[8].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_4 _12690_ (.CLK(clknet_leaf_53_clk),
    .D(\genblk1[8].osc.clkdiv_C.next_cnt[3] ),
    .RESET_B(net174),
    .Q(\genblk1[8].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__dfrtp_4 _12691_ (.CLK(clknet_leaf_54_clk),
    .D(\genblk1[8].osc.clkdiv_C.next_cnt[4] ),
    .RESET_B(net174),
    .Q(\genblk1[8].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__dfrtp_4 _12692_ (.CLK(clknet_leaf_53_clk),
    .D(\genblk1[8].osc.clkdiv_C.next_cnt[5] ),
    .RESET_B(net172),
    .Q(\genblk1[8].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__dfrtp_4 _12693_ (.CLK(clknet_leaf_54_clk),
    .D(\genblk1[8].osc.clkdiv_C.next_cnt[6] ),
    .RESET_B(net172),
    .Q(\genblk1[8].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__dfrtp_4 _12694_ (.CLK(clknet_leaf_54_clk),
    .D(\genblk1[8].osc.clkdiv_C.next_cnt[7] ),
    .RESET_B(net172),
    .Q(\genblk1[8].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__dfrtp_4 _12695_ (.CLK(clknet_leaf_54_clk),
    .D(\genblk1[8].osc.clkdiv_C.next_cnt[8] ),
    .RESET_B(net172),
    .Q(\genblk1[8].osc.clkdiv_C.cnt[8] ));
 sky130_fd_sc_hd__dfrtp_4 _12696_ (.CLK(clknet_leaf_54_clk),
    .D(\genblk1[8].osc.clkdiv_C.next_cnt[9] ),
    .RESET_B(net172),
    .Q(\genblk1[8].osc.clkdiv_C.cnt[9] ));
 sky130_fd_sc_hd__dfrtp_4 _12697_ (.CLK(clknet_leaf_54_clk),
    .D(\genblk1[8].osc.clkdiv_C.next_cnt[10] ),
    .RESET_B(net172),
    .Q(\genblk1[8].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__dfrtp_4 _12698_ (.CLK(clknet_leaf_54_clk),
    .D(\genblk1[8].osc.clkdiv_C.next_cnt[11] ),
    .RESET_B(net172),
    .Q(\genblk1[8].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__dfrtp_4 _12699_ (.CLK(clknet_leaf_54_clk),
    .D(\genblk1[8].osc.clkdiv_C.next_cnt[12] ),
    .RESET_B(net172),
    .Q(\genblk1[8].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__dfrtp_2 _12700_ (.CLK(clknet_leaf_89_clk),
    .D(\genblk1[8].osc.clkdiv_C.next_cnt[13] ),
    .RESET_B(net172),
    .Q(\genblk1[8].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__dfrtp_4 _12701_ (.CLK(clknet_leaf_89_clk),
    .D(\genblk1[8].osc.clkdiv_C.next_cnt[14] ),
    .RESET_B(net172),
    .Q(\genblk1[8].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__dfrtp_4 _12702_ (.CLK(clknet_leaf_89_clk),
    .D(\genblk1[8].osc.clkdiv_C.next_cnt[15] ),
    .RESET_B(net173),
    .Q(\genblk1[8].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__dfrtp_4 _12703_ (.CLK(clknet_leaf_89_clk),
    .D(\genblk1[8].osc.clkdiv_C.next_cnt[16] ),
    .RESET_B(net173),
    .Q(\genblk1[8].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12704_ (.CLK(clknet_leaf_89_clk),
    .D(\genblk1[8].osc.clkdiv_C.next_cnt[17] ),
    .RESET_B(net173),
    .Q(\genblk1[8].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__dfrtp_4 _12705_ (.CLK(clknet_leaf_86_clk),
    .D(\genblk1[9].osc.clkdiv_C.next_cnt[0] ),
    .RESET_B(net181),
    .Q(\genblk1[9].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _12706_ (.CLK(clknet_leaf_86_clk),
    .D(\genblk1[9].osc.clkdiv_C.next_cnt[1] ),
    .RESET_B(net183),
    .Q(\genblk1[9].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _12707_ (.CLK(clknet_leaf_56_clk),
    .D(\genblk1[9].osc.clkdiv_C.next_cnt[2] ),
    .RESET_B(net181),
    .Q(\genblk1[9].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_4 _12708_ (.CLK(clknet_leaf_56_clk),
    .D(\genblk1[9].osc.clkdiv_C.next_cnt[3] ),
    .RESET_B(net181),
    .Q(\genblk1[9].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__dfrtp_4 _12709_ (.CLK(clknet_leaf_56_clk),
    .D(\genblk1[9].osc.clkdiv_C.next_cnt[4] ),
    .RESET_B(net181),
    .Q(\genblk1[9].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__dfrtp_4 _12710_ (.CLK(clknet_leaf_56_clk),
    .D(\genblk1[9].osc.clkdiv_C.next_cnt[5] ),
    .RESET_B(net181),
    .Q(\genblk1[9].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__dfrtp_4 _12711_ (.CLK(clknet_leaf_56_clk),
    .D(\genblk1[9].osc.clkdiv_C.next_cnt[6] ),
    .RESET_B(net175),
    .Q(\genblk1[9].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__dfrtp_4 _12712_ (.CLK(clknet_leaf_55_clk),
    .D(\genblk1[9].osc.clkdiv_C.next_cnt[7] ),
    .RESET_B(net175),
    .Q(\genblk1[9].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12713_ (.CLK(clknet_leaf_55_clk),
    .D(\genblk1[9].osc.clkdiv_C.next_cnt[8] ),
    .RESET_B(net175),
    .Q(\genblk1[9].osc.clkdiv_C.cnt[8] ));
 sky130_fd_sc_hd__dfrtp_2 _12714_ (.CLK(clknet_leaf_54_clk),
    .D(\genblk1[9].osc.clkdiv_C.next_cnt[9] ),
    .RESET_B(net175),
    .Q(\genblk1[9].osc.clkdiv_C.cnt[9] ));
 sky130_fd_sc_hd__dfrtp_4 _12715_ (.CLK(clknet_leaf_54_clk),
    .D(\genblk1[9].osc.clkdiv_C.next_cnt[10] ),
    .RESET_B(net175),
    .Q(\genblk1[9].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__dfrtp_4 _12716_ (.CLK(clknet_leaf_56_clk),
    .D(\genblk1[9].osc.clkdiv_C.next_cnt[11] ),
    .RESET_B(net175),
    .Q(\genblk1[9].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__dfrtp_4 _12717_ (.CLK(clknet_leaf_86_clk),
    .D(\genblk1[9].osc.clkdiv_C.next_cnt[12] ),
    .RESET_B(net181),
    .Q(\genblk1[9].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__dfrtp_4 _12718_ (.CLK(clknet_leaf_86_clk),
    .D(\genblk1[9].osc.clkdiv_C.next_cnt[13] ),
    .RESET_B(net181),
    .Q(\genblk1[9].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__dfrtp_4 _12719_ (.CLK(clknet_leaf_86_clk),
    .D(\genblk1[9].osc.clkdiv_C.next_cnt[14] ),
    .RESET_B(net181),
    .Q(\genblk1[9].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__dfrtp_4 _12720_ (.CLK(clknet_leaf_86_clk),
    .D(\genblk1[9].osc.clkdiv_C.next_cnt[15] ),
    .RESET_B(net183),
    .Q(\genblk1[9].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__dfrtp_4 _12721_ (.CLK(clknet_leaf_86_clk),
    .D(\genblk1[9].osc.clkdiv_C.next_cnt[16] ),
    .RESET_B(net183),
    .Q(\genblk1[9].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__dfrtp_4 _12722_ (.CLK(clknet_leaf_86_clk),
    .D(\genblk1[9].osc.clkdiv_C.next_cnt[17] ),
    .RESET_B(net183),
    .Q(\genblk1[9].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__dfrtp_4 _12723_ (.CLK(clknet_leaf_37_clk),
    .D(\genblk1[10].osc.clkdiv_C.next_cnt[0] ),
    .RESET_B(net113),
    .Q(\genblk1[10].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _12724_ (.CLK(clknet_leaf_37_clk),
    .D(\genblk1[10].osc.clkdiv_C.next_cnt[1] ),
    .RESET_B(net113),
    .Q(\genblk1[10].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _12725_ (.CLK(clknet_leaf_37_clk),
    .D(\genblk1[10].osc.clkdiv_C.next_cnt[2] ),
    .RESET_B(net113),
    .Q(\genblk1[10].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_4 _12726_ (.CLK(clknet_leaf_37_clk),
    .D(\genblk1[10].osc.clkdiv_C.next_cnt[3] ),
    .RESET_B(net113),
    .Q(\genblk1[10].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__dfrtp_4 _12727_ (.CLK(clknet_leaf_38_clk),
    .D(\genblk1[10].osc.clkdiv_C.next_cnt[4] ),
    .RESET_B(net113),
    .Q(\genblk1[10].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__dfrtp_4 _12728_ (.CLK(clknet_leaf_38_clk),
    .D(\genblk1[10].osc.clkdiv_C.next_cnt[5] ),
    .RESET_B(net113),
    .Q(\genblk1[10].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__dfrtp_4 _12729_ (.CLK(clknet_leaf_38_clk),
    .D(\genblk1[10].osc.clkdiv_C.next_cnt[6] ),
    .RESET_B(net115),
    .Q(\genblk1[10].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__dfrtp_4 _12730_ (.CLK(clknet_leaf_39_clk),
    .D(\genblk1[10].osc.clkdiv_C.next_cnt[7] ),
    .RESET_B(net115),
    .Q(\genblk1[10].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12731_ (.CLK(clknet_leaf_38_clk),
    .D(\genblk1[10].osc.clkdiv_C.next_cnt[8] ),
    .RESET_B(net115),
    .Q(\genblk1[10].osc.clkdiv_C.cnt[8] ));
 sky130_fd_sc_hd__dfrtp_4 _12732_ (.CLK(clknet_leaf_38_clk),
    .D(\genblk1[10].osc.clkdiv_C.next_cnt[9] ),
    .RESET_B(net115),
    .Q(\genblk1[10].osc.clkdiv_C.cnt[9] ));
 sky130_fd_sc_hd__dfrtp_4 _12733_ (.CLK(clknet_leaf_38_clk),
    .D(\genblk1[10].osc.clkdiv_C.next_cnt[10] ),
    .RESET_B(net115),
    .Q(\genblk1[10].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__dfrtp_4 _12734_ (.CLK(clknet_leaf_38_clk),
    .D(\genblk1[10].osc.clkdiv_C.next_cnt[11] ),
    .RESET_B(net113),
    .Q(\genblk1[10].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__dfrtp_2 _12735_ (.CLK(clknet_leaf_38_clk),
    .D(\genblk1[10].osc.clkdiv_C.next_cnt[12] ),
    .RESET_B(net114),
    .Q(\genblk1[10].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__dfrtp_4 _12736_ (.CLK(clknet_leaf_37_clk),
    .D(\genblk1[10].osc.clkdiv_C.next_cnt[13] ),
    .RESET_B(net114),
    .Q(\genblk1[10].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__dfrtp_2 _12737_ (.CLK(clknet_leaf_37_clk),
    .D(\genblk1[10].osc.clkdiv_C.next_cnt[14] ),
    .RESET_B(net114),
    .Q(\genblk1[10].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__dfrtp_2 _12738_ (.CLK(clknet_leaf_38_clk),
    .D(\genblk1[10].osc.clkdiv_C.next_cnt[15] ),
    .RESET_B(net114),
    .Q(\genblk1[10].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__dfrtp_2 _12739_ (.CLK(clknet_leaf_48_clk),
    .D(\genblk1[10].osc.clkdiv_C.next_cnt[16] ),
    .RESET_B(net114),
    .Q(\genblk1[10].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12740_ (.CLK(clknet_leaf_48_clk),
    .D(\genblk1[10].osc.clkdiv_C.next_cnt[17] ),
    .RESET_B(net119),
    .Q(\genblk1[10].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__dfrtp_4 _12741_ (.CLK(clknet_leaf_49_clk),
    .D(\genblk1[11].osc.clkdiv_C.next_cnt[0] ),
    .RESET_B(net108),
    .Q(\genblk1[11].osc.clkdiv_C.cnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _12742_ (.CLK(clknet_leaf_50_clk),
    .D(\genblk1[11].osc.clkdiv_C.next_cnt[1] ),
    .RESET_B(net108),
    .Q(\genblk1[11].osc.clkdiv_C.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _12743_ (.CLK(clknet_leaf_49_clk),
    .D(\genblk1[11].osc.clkdiv_C.next_cnt[2] ),
    .RESET_B(net108),
    .Q(\genblk1[11].osc.clkdiv_C.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_4 _12744_ (.CLK(clknet_leaf_49_clk),
    .D(\genblk1[11].osc.clkdiv_C.next_cnt[3] ),
    .RESET_B(net108),
    .Q(\genblk1[11].osc.clkdiv_C.cnt[3] ));
 sky130_fd_sc_hd__dfrtp_4 _12745_ (.CLK(clknet_leaf_50_clk),
    .D(\genblk1[11].osc.clkdiv_C.next_cnt[4] ),
    .RESET_B(net108),
    .Q(\genblk1[11].osc.clkdiv_C.cnt[4] ));
 sky130_fd_sc_hd__dfrtp_4 _12746_ (.CLK(clknet_leaf_49_clk),
    .D(\genblk1[11].osc.clkdiv_C.next_cnt[5] ),
    .RESET_B(net108),
    .Q(\genblk1[11].osc.clkdiv_C.cnt[5] ));
 sky130_fd_sc_hd__dfrtp_4 _12747_ (.CLK(clknet_leaf_49_clk),
    .D(\genblk1[11].osc.clkdiv_C.next_cnt[6] ),
    .RESET_B(net108),
    .Q(\genblk1[11].osc.clkdiv_C.cnt[6] ));
 sky130_fd_sc_hd__dfrtp_4 _12748_ (.CLK(clknet_leaf_50_clk),
    .D(\genblk1[11].osc.clkdiv_C.next_cnt[7] ),
    .RESET_B(net111),
    .Q(\genblk1[11].osc.clkdiv_C.cnt[7] ));
 sky130_fd_sc_hd__dfrtp_2 _12749_ (.CLK(clknet_leaf_46_clk),
    .D(\genblk1[11].osc.clkdiv_C.next_cnt[8] ),
    .RESET_B(net119),
    .Q(\genblk1[11].osc.clkdiv_C.cnt[8] ));
 sky130_fd_sc_hd__dfrtp_2 _12750_ (.CLK(clknet_leaf_46_clk),
    .D(\genblk1[11].osc.clkdiv_C.next_cnt[9] ),
    .RESET_B(net119),
    .Q(\genblk1[11].osc.clkdiv_C.cnt[9] ));
 sky130_fd_sc_hd__dfrtp_2 _12751_ (.CLK(clknet_leaf_50_clk),
    .D(\genblk1[11].osc.clkdiv_C.next_cnt[10] ),
    .RESET_B(net111),
    .Q(\genblk1[11].osc.clkdiv_C.cnt[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12752_ (.CLK(clknet_leaf_50_clk),
    .D(\genblk1[11].osc.clkdiv_C.next_cnt[11] ),
    .RESET_B(net111),
    .Q(\genblk1[11].osc.clkdiv_C.cnt[11] ));
 sky130_fd_sc_hd__dfrtp_4 _12753_ (.CLK(clknet_leaf_51_clk),
    .D(\genblk1[11].osc.clkdiv_C.next_cnt[12] ),
    .RESET_B(net110),
    .Q(\genblk1[11].osc.clkdiv_C.cnt[12] ));
 sky130_fd_sc_hd__dfrtp_2 _12754_ (.CLK(clknet_leaf_51_clk),
    .D(\genblk1[11].osc.clkdiv_C.next_cnt[13] ),
    .RESET_B(net110),
    .Q(\genblk1[11].osc.clkdiv_C.cnt[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12755_ (.CLK(clknet_leaf_52_clk),
    .D(\genblk1[11].osc.clkdiv_C.next_cnt[14] ),
    .RESET_B(net110),
    .Q(\genblk1[11].osc.clkdiv_C.cnt[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12756_ (.CLK(clknet_leaf_50_clk),
    .D(\genblk1[11].osc.clkdiv_C.next_cnt[15] ),
    .RESET_B(net110),
    .Q(\genblk1[11].osc.clkdiv_C.cnt[15] ));
 sky130_fd_sc_hd__dfrtp_4 _12757_ (.CLK(clknet_leaf_52_clk),
    .D(\genblk1[11].osc.clkdiv_C.next_cnt[16] ),
    .RESET_B(net110),
    .Q(\genblk1[11].osc.clkdiv_C.cnt[16] ));
 sky130_fd_sc_hd__dfrtp_4 _12758_ (.CLK(clknet_leaf_52_clk),
    .D(\genblk1[11].osc.clkdiv_C.next_cnt[17] ),
    .RESET_B(net110),
    .Q(\genblk1[11].osc.clkdiv_C.cnt[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12759_ (.CLK(clknet_leaf_58_clk),
    .D(_00000_),
    .RESET_B(net192),
    .Q(\genblk2[0].wave_shpr.div.busy ));
 sky130_fd_sc_hd__dfrtp_1 _12760_ (.CLK(clknet_leaf_93_clk),
    .D(_00001_),
    .RESET_B(net146),
    .Q(\genblk2[0].wave_shpr.div.done ));
 sky130_fd_sc_hd__dfrtp_4 _12761_ (.CLK(clknet_leaf_20_clk),
    .D(_00094_),
    .RESET_B(net108),
    .Q(\freq_div.state[0] ));
 sky130_fd_sc_hd__dfstp_2 _12762_ (.CLK(clknet_leaf_20_clk),
    .D(_00095_),
    .SET_B(net109),
    .Q(\freq_div.state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _12763_ (.CLK(clknet_leaf_20_clk),
    .D(_00096_),
    .RESET_B(net108),
    .Q(\freq_div.state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _12764_ (.CLK(clknet_leaf_92_clk),
    .D(_00097_),
    .RESET_B(net148),
    .Q(\genblk2[0].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__dfrtp_2 _12765_ (.CLK(clknet_leaf_93_clk),
    .D(_00098_),
    .RESET_B(net146),
    .Q(\genblk2[0].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12766_ (.CLK(clknet_leaf_91_clk),
    .D(_00099_),
    .RESET_B(net146),
    .Q(\genblk2[0].wave_shpr.div.fin_quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12767_ (.CLK(clknet_leaf_93_clk),
    .D(_00100_),
    .RESET_B(net148),
    .Q(\genblk2[0].wave_shpr.div.fin_quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12768_ (.CLK(clknet_leaf_93_clk),
    .D(_00101_),
    .RESET_B(net148),
    .Q(\genblk2[0].wave_shpr.div.fin_quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12769_ (.CLK(clknet_leaf_93_clk),
    .D(_00102_),
    .RESET_B(net148),
    .Q(\genblk2[0].wave_shpr.div.fin_quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12770_ (.CLK(clknet_leaf_93_clk),
    .D(_00103_),
    .RESET_B(net148),
    .Q(\genblk2[0].wave_shpr.div.fin_quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12771_ (.CLK(clknet_leaf_93_clk),
    .D(_00104_),
    .RESET_B(net148),
    .Q(\genblk2[0].wave_shpr.div.fin_quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12772_ (.CLK(clknet_leaf_47_clk),
    .D(_00105_),
    .RESET_B(net121),
    .Q(\genblk2[10].wave_shpr.div.b1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12773_ (.CLK(clknet_leaf_47_clk),
    .D(_00106_),
    .RESET_B(net119),
    .Q(\genblk2[10].wave_shpr.div.b1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12774_ (.CLK(clknet_leaf_44_clk),
    .D(_00107_),
    .RESET_B(net120),
    .Q(\genblk2[10].wave_shpr.div.b1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12775_ (.CLK(clknet_leaf_41_clk),
    .D(_00108_),
    .RESET_B(net123),
    .Q(\genblk2[10].wave_shpr.div.b1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12776_ (.CLK(clknet_leaf_43_clk),
    .D(_00109_),
    .RESET_B(net124),
    .Q(\genblk2[10].wave_shpr.div.b1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12777_ (.CLK(clknet_leaf_43_clk),
    .D(_00110_),
    .RESET_B(net124),
    .Q(\genblk2[10].wave_shpr.div.b1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12778_ (.CLK(clknet_leaf_41_clk),
    .D(_00111_),
    .RESET_B(net123),
    .Q(\genblk2[10].wave_shpr.div.b1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12779_ (.CLK(clknet_leaf_41_clk),
    .D(_00112_),
    .RESET_B(net116),
    .Q(\genblk2[10].wave_shpr.div.b1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12780_ (.CLK(clknet_leaf_40_clk),
    .D(_00113_),
    .RESET_B(net116),
    .Q(\genblk2[10].wave_shpr.div.b1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12781_ (.CLK(clknet_leaf_40_clk),
    .D(_00114_),
    .RESET_B(net115),
    .Q(\genblk2[10].wave_shpr.div.b1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12782_ (.CLK(clknet_leaf_40_clk),
    .D(_00115_),
    .RESET_B(net117),
    .Q(\genblk2[10].wave_shpr.div.b1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12783_ (.CLK(clknet_leaf_40_clk),
    .D(_00116_),
    .RESET_B(net117),
    .Q(\genblk2[10].wave_shpr.div.b1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12784_ (.CLK(clknet_leaf_40_clk),
    .D(_00117_),
    .RESET_B(net123),
    .Q(\genblk2[10].wave_shpr.div.b1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12785_ (.CLK(clknet_leaf_41_clk),
    .D(_00118_),
    .RESET_B(net123),
    .Q(\genblk2[10].wave_shpr.div.b1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12786_ (.CLK(clknet_leaf_43_clk),
    .D(_00119_),
    .RESET_B(net124),
    .Q(\genblk2[10].wave_shpr.div.b1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12787_ (.CLK(clknet_leaf_43_clk),
    .D(_00120_),
    .RESET_B(net124),
    .Q(\genblk2[10].wave_shpr.div.b1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12788_ (.CLK(clknet_leaf_43_clk),
    .D(_00121_),
    .RESET_B(net124),
    .Q(\genblk2[10].wave_shpr.div.b1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12789_ (.CLK(clknet_leaf_43_clk),
    .D(_00122_),
    .RESET_B(net124),
    .Q(\genblk2[10].wave_shpr.div.b1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12790_ (.CLK(clknet_leaf_57_clk),
    .D(_00123_),
    .RESET_B(net182),
    .Q(\genblk2[0].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12791_ (.CLK(clknet_leaf_91_clk),
    .D(_00124_),
    .RESET_B(net146),
    .Q(\genblk2[0].wave_shpr.div.quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12792_ (.CLK(clknet_leaf_91_clk),
    .D(_00125_),
    .RESET_B(net148),
    .Q(\genblk2[0].wave_shpr.div.quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12793_ (.CLK(clknet_leaf_93_clk),
    .D(net559),
    .RESET_B(net148),
    .Q(\genblk2[0].wave_shpr.div.quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12794_ (.CLK(clknet_leaf_93_clk),
    .D(_00127_),
    .RESET_B(net148),
    .Q(\genblk2[0].wave_shpr.div.quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12795_ (.CLK(clknet_leaf_92_clk),
    .D(net601),
    .RESET_B(net148),
    .Q(\genblk2[0].wave_shpr.div.quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12796_ (.CLK(clknet_leaf_92_clk),
    .D(_00129_),
    .RESET_B(net149),
    .Q(\genblk2[0].wave_shpr.div.quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12797_ (.CLK(clknet_leaf_57_clk),
    .D(net270),
    .RESET_B(net183),
    .Q(\genblk2[0].wave_shpr.div.quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12798_ (.CLK(clknet_leaf_57_clk),
    .D(_00131_),
    .RESET_B(net183),
    .Q(\genblk2[0].wave_shpr.div.quo[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12799_ (.CLK(clknet_leaf_59_clk),
    .D(net278),
    .RESET_B(net192),
    .Q(\genblk2[0].wave_shpr.div.quo[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12800_ (.CLK(clknet_leaf_59_clk),
    .D(_00133_),
    .RESET_B(net192),
    .Q(\genblk2[0].wave_shpr.div.quo[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12801_ (.CLK(clknet_leaf_59_clk),
    .D(net570),
    .RESET_B(net193),
    .Q(\genblk2[0].wave_shpr.div.quo[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12802_ (.CLK(clknet_leaf_59_clk),
    .D(_00135_),
    .RESET_B(net193),
    .Q(\genblk2[0].wave_shpr.div.quo[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12803_ (.CLK(clknet_leaf_59_clk),
    .D(_00136_),
    .RESET_B(net188),
    .Q(\genblk2[0].wave_shpr.div.quo[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12804_ (.CLK(clknet_leaf_59_clk),
    .D(net496),
    .RESET_B(net188),
    .Q(\genblk2[0].wave_shpr.div.quo[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12805_ (.CLK(clknet_leaf_59_clk),
    .D(net544),
    .RESET_B(net187),
    .Q(\genblk2[0].wave_shpr.div.quo[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12806_ (.CLK(clknet_leaf_59_clk),
    .D(_00139_),
    .RESET_B(net187),
    .Q(\genblk2[0].wave_shpr.div.quo[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12807_ (.CLK(clknet_leaf_59_clk),
    .D(_00140_),
    .RESET_B(net187),
    .Q(\genblk2[0].wave_shpr.div.quo[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12808_ (.CLK(clknet_leaf_60_clk),
    .D(net411),
    .RESET_B(net187),
    .Q(\genblk2[0].wave_shpr.div.quo[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12809_ (.CLK(clknet_leaf_60_clk),
    .D(_00142_),
    .RESET_B(net187),
    .Q(\genblk2[0].wave_shpr.div.quo[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12810_ (.CLK(clknet_leaf_59_clk),
    .D(net299),
    .RESET_B(net187),
    .Q(\genblk2[0].wave_shpr.div.quo[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12811_ (.CLK(clknet_leaf_59_clk),
    .D(_00144_),
    .RESET_B(net192),
    .Q(\genblk2[0].wave_shpr.div.quo[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12812_ (.CLK(clknet_leaf_58_clk),
    .D(net266),
    .RESET_B(net192),
    .Q(\genblk2[0].wave_shpr.div.quo[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12813_ (.CLK(clknet_leaf_58_clk),
    .D(_00146_),
    .RESET_B(net192),
    .Q(\genblk2[0].wave_shpr.div.quo[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12814_ (.CLK(clknet_leaf_58_clk),
    .D(net455),
    .RESET_B(net192),
    .Q(\genblk2[0].wave_shpr.div.quo[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12815_ (.CLK(clknet_leaf_58_clk),
    .D(net579),
    .RESET_B(net192),
    .Q(\genblk2[0].wave_shpr.div.acc_next[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12816_ (.CLK(clknet_leaf_58_clk),
    .D(_00149_),
    .RESET_B(net192),
    .Q(\genblk2[0].wave_shpr.div.acc[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12817_ (.CLK(clknet_leaf_59_clk),
    .D(_00150_),
    .RESET_B(net193),
    .Q(\genblk2[0].wave_shpr.div.acc[1] ));
 sky130_fd_sc_hd__dfrtp_2 _12818_ (.CLK(clknet_leaf_67_clk),
    .D(_00151_),
    .RESET_B(net193),
    .Q(\genblk2[0].wave_shpr.div.acc[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12819_ (.CLK(clknet_leaf_66_clk),
    .D(_00152_),
    .RESET_B(net196),
    .Q(\genblk2[0].wave_shpr.div.acc[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12820_ (.CLK(clknet_leaf_66_clk),
    .D(_00153_),
    .RESET_B(net196),
    .Q(\genblk2[0].wave_shpr.div.acc[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12821_ (.CLK(clknet_leaf_67_clk),
    .D(net824),
    .RESET_B(net196),
    .Q(\genblk2[0].wave_shpr.div.acc[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12822_ (.CLK(clknet_leaf_62_clk),
    .D(_00155_),
    .RESET_B(net189),
    .Q(\genblk2[0].wave_shpr.div.acc[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12823_ (.CLK(clknet_leaf_62_clk),
    .D(_00156_),
    .RESET_B(net189),
    .Q(\genblk2[0].wave_shpr.div.acc[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12824_ (.CLK(clknet_leaf_62_clk),
    .D(_00157_),
    .RESET_B(net189),
    .Q(\genblk2[0].wave_shpr.div.acc[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12825_ (.CLK(clknet_leaf_62_clk),
    .D(_00158_),
    .RESET_B(net190),
    .Q(\genblk2[0].wave_shpr.div.acc[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12826_ (.CLK(clknet_leaf_62_clk),
    .D(_00159_),
    .RESET_B(net190),
    .Q(\genblk2[0].wave_shpr.div.acc[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12827_ (.CLK(clknet_leaf_62_clk),
    .D(_00160_),
    .RESET_B(net190),
    .Q(\genblk2[0].wave_shpr.div.acc[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12828_ (.CLK(clknet_leaf_62_clk),
    .D(_00161_),
    .RESET_B(net190),
    .Q(\genblk2[0].wave_shpr.div.acc[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12829_ (.CLK(clknet_leaf_64_clk),
    .D(_00162_),
    .RESET_B(net189),
    .Q(\genblk2[0].wave_shpr.div.acc[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12830_ (.CLK(clknet_leaf_62_clk),
    .D(_00163_),
    .RESET_B(net189),
    .Q(\genblk2[0].wave_shpr.div.acc[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12831_ (.CLK(clknet_leaf_64_clk),
    .D(_00164_),
    .RESET_B(net189),
    .Q(\genblk2[0].wave_shpr.div.acc[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12832_ (.CLK(clknet_leaf_64_clk),
    .D(_00165_),
    .RESET_B(net189),
    .Q(\genblk2[0].wave_shpr.div.acc[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12833_ (.CLK(clknet_leaf_64_clk),
    .D(_00166_),
    .RESET_B(net196),
    .Q(\genblk2[0].wave_shpr.div.acc[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12834_ (.CLK(clknet_leaf_64_clk),
    .D(_00167_),
    .RESET_B(net196),
    .Q(\genblk2[0].wave_shpr.div.acc[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12835_ (.CLK(clknet_leaf_64_clk),
    .D(net689),
    .RESET_B(net196),
    .Q(\genblk2[0].wave_shpr.div.acc[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12836_ (.CLK(clknet_leaf_64_clk),
    .D(_00169_),
    .RESET_B(net196),
    .Q(\genblk2[0].wave_shpr.div.acc[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12837_ (.CLK(clknet_leaf_65_clk),
    .D(_00170_),
    .RESET_B(net196),
    .Q(\genblk2[0].wave_shpr.div.acc[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12838_ (.CLK(clknet_leaf_65_clk),
    .D(_00171_),
    .RESET_B(net196),
    .Q(\genblk2[0].wave_shpr.div.acc[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12839_ (.CLK(clknet_leaf_65_clk),
    .D(_00172_),
    .RESET_B(net197),
    .Q(\genblk2[0].wave_shpr.div.acc[23] ));
 sky130_fd_sc_hd__dfrtp_2 _12840_ (.CLK(clknet_leaf_65_clk),
    .D(net1306),
    .RESET_B(net197),
    .Q(\genblk2[0].wave_shpr.div.acc[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12841_ (.CLK(clknet_leaf_64_clk),
    .D(_00174_),
    .RESET_B(net196),
    .Q(\genblk2[0].wave_shpr.div.acc[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12842_ (.CLK(clknet_leaf_65_clk),
    .D(_00175_),
    .RESET_B(net197),
    .Q(\genblk2[0].wave_shpr.div.acc[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12843_ (.CLK(clknet_leaf_30_clk),
    .D(_00006_),
    .RESET_B(net104),
    .Q(\genblk2[1].wave_shpr.div.busy ));
 sky130_fd_sc_hd__dfrtp_1 _12844_ (.CLK(clknet_leaf_116_clk),
    .D(_00007_),
    .RESET_B(net150),
    .Q(\genblk2[1].wave_shpr.div.done ));
 sky130_fd_sc_hd__dfrtp_2 _12845_ (.CLK(clknet_leaf_68_clk),
    .D(_00176_),
    .RESET_B(net194),
    .Q(\genblk2[11].wave_shpr.div.i[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12846_ (.CLK(clknet_leaf_68_clk),
    .D(_00177_),
    .RESET_B(net211),
    .Q(\genblk2[11].wave_shpr.div.i[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12847_ (.CLK(clknet_leaf_58_clk),
    .D(_00178_),
    .RESET_B(net211),
    .Q(\genblk2[11].wave_shpr.div.i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12848_ (.CLK(clknet_leaf_58_clk),
    .D(_00179_),
    .RESET_B(net194),
    .Q(\genblk2[11].wave_shpr.div.i[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12849_ (.CLK(clknet_leaf_58_clk),
    .D(_00180_),
    .RESET_B(net194),
    .Q(\genblk2[11].wave_shpr.div.i[4] ));
 sky130_fd_sc_hd__dfrtp_4 _12850_ (.CLK(clknet_leaf_118_clk),
    .D(_00181_),
    .RESET_B(net138),
    .Q(\genblk2[1].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__dfrtp_2 _12851_ (.CLK(clknet_leaf_118_clk),
    .D(_00182_),
    .RESET_B(net138),
    .Q(\genblk2[1].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__dfrtp_2 _12852_ (.CLK(clknet_leaf_118_clk),
    .D(_00183_),
    .RESET_B(net138),
    .Q(\genblk2[1].wave_shpr.div.fin_quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12853_ (.CLK(clknet_leaf_119_clk),
    .D(_00184_),
    .RESET_B(net139),
    .Q(\genblk2[1].wave_shpr.div.fin_quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12854_ (.CLK(clknet_leaf_119_clk),
    .D(_00185_),
    .RESET_B(net139),
    .Q(\genblk2[1].wave_shpr.div.fin_quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12855_ (.CLK(clknet_leaf_91_clk),
    .D(_00186_),
    .RESET_B(net146),
    .Q(\genblk2[1].wave_shpr.div.fin_quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12856_ (.CLK(clknet_leaf_91_clk),
    .D(_00187_),
    .RESET_B(net146),
    .Q(\genblk2[1].wave_shpr.div.fin_quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12857_ (.CLK(clknet_leaf_91_clk),
    .D(_00188_),
    .RESET_B(net146),
    .Q(\genblk2[1].wave_shpr.div.fin_quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12858_ (.CLK(clknet_leaf_134_clk),
    .D(_00189_),
    .RESET_B(net60),
    .Q(\genblk2[2].wave_shpr.div.b1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12859_ (.CLK(clknet_leaf_132_clk),
    .D(_00190_),
    .RESET_B(net64),
    .Q(\genblk2[2].wave_shpr.div.b1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12860_ (.CLK(clknet_leaf_129_clk),
    .D(_00191_),
    .RESET_B(net64),
    .Q(\genblk2[2].wave_shpr.div.b1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12861_ (.CLK(clknet_leaf_129_clk),
    .D(_00192_),
    .RESET_B(net64),
    .Q(\genblk2[2].wave_shpr.div.b1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12862_ (.CLK(clknet_leaf_126_clk),
    .D(_00193_),
    .RESET_B(net61),
    .Q(\genblk2[2].wave_shpr.div.b1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12863_ (.CLK(clknet_leaf_129_clk),
    .D(_00194_),
    .RESET_B(net66),
    .Q(\genblk2[2].wave_shpr.div.b1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12864_ (.CLK(clknet_leaf_129_clk),
    .D(_00195_),
    .RESET_B(net64),
    .Q(\genblk2[2].wave_shpr.div.b1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12865_ (.CLK(clknet_leaf_135_clk),
    .D(_00196_),
    .RESET_B(net61),
    .Q(\genblk2[2].wave_shpr.div.b1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12866_ (.CLK(clknet_leaf_135_clk),
    .D(_00197_),
    .RESET_B(net61),
    .Q(\genblk2[2].wave_shpr.div.b1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12867_ (.CLK(clknet_leaf_134_clk),
    .D(_00198_),
    .RESET_B(net60),
    .Q(\genblk2[2].wave_shpr.div.b1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12868_ (.CLK(clknet_leaf_134_clk),
    .D(_00199_),
    .RESET_B(net60),
    .Q(\genblk2[2].wave_shpr.div.b1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12869_ (.CLK(clknet_leaf_134_clk),
    .D(_00200_),
    .RESET_B(net60),
    .Q(\genblk2[2].wave_shpr.div.b1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12870_ (.CLK(clknet_leaf_134_clk),
    .D(_00201_),
    .RESET_B(net59),
    .Q(\genblk2[2].wave_shpr.div.b1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12871_ (.CLK(clknet_leaf_134_clk),
    .D(_00202_),
    .RESET_B(net59),
    .Q(\genblk2[2].wave_shpr.div.b1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12872_ (.CLK(clknet_leaf_134_clk),
    .D(_00203_),
    .RESET_B(net59),
    .Q(\genblk2[2].wave_shpr.div.b1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12873_ (.CLK(clknet_leaf_138_clk),
    .D(_00204_),
    .RESET_B(net39),
    .Q(\genblk2[2].wave_shpr.div.b1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12874_ (.CLK(clknet_leaf_136_clk),
    .D(_00205_),
    .RESET_B(net42),
    .Q(\genblk2[2].wave_shpr.div.b1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12875_ (.CLK(clknet_leaf_138_clk),
    .D(_00206_),
    .RESET_B(net39),
    .Q(\genblk2[2].wave_shpr.div.b1[17] ));
 sky130_fd_sc_hd__dfrtp_4 _12876_ (.CLK(clknet_leaf_49_clk),
    .D(_00207_),
    .RESET_B(net113),
    .Q(\genblk2[1].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12877_ (.CLK(clknet_leaf_119_clk),
    .D(_00208_),
    .RESET_B(net141),
    .Q(\genblk2[1].wave_shpr.div.quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12878_ (.CLK(clknet_leaf_119_clk),
    .D(net685),
    .RESET_B(net143),
    .Q(\genblk2[1].wave_shpr.div.quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12879_ (.CLK(clknet_leaf_119_clk),
    .D(_00210_),
    .RESET_B(net139),
    .Q(\genblk2[1].wave_shpr.div.quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12880_ (.CLK(clknet_leaf_119_clk),
    .D(_00211_),
    .RESET_B(net146),
    .Q(\genblk2[1].wave_shpr.div.quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12881_ (.CLK(clknet_leaf_91_clk),
    .D(net415),
    .RESET_B(net146),
    .Q(\genblk2[1].wave_shpr.div.quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12882_ (.CLK(clknet_leaf_91_clk),
    .D(_00213_),
    .RESET_B(net146),
    .Q(\genblk2[1].wave_shpr.div.quo[6] ));
 sky130_fd_sc_hd__dfrtp_2 _12883_ (.CLK(clknet_leaf_55_clk),
    .D(net293),
    .RESET_B(net176),
    .Q(\genblk2[1].wave_shpr.div.quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12884_ (.CLK(clknet_leaf_30_clk),
    .D(net461),
    .RESET_B(net97),
    .Q(\genblk2[1].wave_shpr.div.quo[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12885_ (.CLK(clknet_leaf_30_clk),
    .D(_00216_),
    .RESET_B(net97),
    .Q(\genblk2[1].wave_shpr.div.quo[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12886_ (.CLK(clknet_leaf_30_clk),
    .D(_00217_),
    .RESET_B(net98),
    .Q(\genblk2[1].wave_shpr.div.quo[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12887_ (.CLK(clknet_leaf_30_clk),
    .D(_00218_),
    .RESET_B(net96),
    .Q(\genblk2[1].wave_shpr.div.quo[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12888_ (.CLK(clknet_leaf_30_clk),
    .D(_00219_),
    .RESET_B(net96),
    .Q(\genblk2[1].wave_shpr.div.quo[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12889_ (.CLK(clknet_leaf_30_clk),
    .D(_00220_),
    .RESET_B(net96),
    .Q(\genblk2[1].wave_shpr.div.quo[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12890_ (.CLK(clknet_leaf_28_clk),
    .D(_00221_),
    .RESET_B(net91),
    .Q(\genblk2[1].wave_shpr.div.quo[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12891_ (.CLK(clknet_leaf_28_clk),
    .D(net512),
    .RESET_B(net91),
    .Q(\genblk2[1].wave_shpr.div.quo[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12892_ (.CLK(clknet_leaf_28_clk),
    .D(net463),
    .RESET_B(net91),
    .Q(\genblk2[1].wave_shpr.div.quo[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12893_ (.CLK(clknet_leaf_28_clk),
    .D(_00224_),
    .RESET_B(net91),
    .Q(\genblk2[1].wave_shpr.div.quo[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12894_ (.CLK(clknet_leaf_32_clk),
    .D(net427),
    .RESET_B(net99),
    .Q(\genblk2[1].wave_shpr.div.quo[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12895_ (.CLK(clknet_leaf_32_clk),
    .D(_00226_),
    .RESET_B(net99),
    .Q(\genblk2[1].wave_shpr.div.quo[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12896_ (.CLK(clknet_leaf_32_clk),
    .D(_00227_),
    .RESET_B(net99),
    .Q(\genblk2[1].wave_shpr.div.quo[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12897_ (.CLK(clknet_leaf_31_clk),
    .D(net258),
    .RESET_B(net99),
    .Q(\genblk2[1].wave_shpr.div.quo[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12898_ (.CLK(clknet_leaf_31_clk),
    .D(_00229_),
    .RESET_B(net102),
    .Q(\genblk2[1].wave_shpr.div.quo[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12899_ (.CLK(clknet_leaf_30_clk),
    .D(net341),
    .RESET_B(net102),
    .Q(\genblk2[1].wave_shpr.div.quo[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12900_ (.CLK(clknet_leaf_30_clk),
    .D(net633),
    .RESET_B(net102),
    .Q(\genblk2[1].wave_shpr.div.quo[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12901_ (.CLK(clknet_leaf_30_clk),
    .D(net589),
    .RESET_B(net102),
    .Q(\genblk2[1].wave_shpr.div.acc_next[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12902_ (.CLK(clknet_leaf_30_clk),
    .D(_00233_),
    .RESET_B(net104),
    .Q(\genblk2[1].wave_shpr.div.acc[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12903_ (.CLK(clknet_leaf_37_clk),
    .D(net753),
    .RESET_B(net104),
    .Q(\genblk2[1].wave_shpr.div.acc[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12904_ (.CLK(clknet_leaf_37_clk),
    .D(_00235_),
    .RESET_B(net104),
    .Q(\genblk2[1].wave_shpr.div.acc[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12905_ (.CLK(clknet_leaf_37_clk),
    .D(_00236_),
    .RESET_B(net104),
    .Q(\genblk2[1].wave_shpr.div.acc[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12906_ (.CLK(clknet_leaf_36_clk),
    .D(_00237_),
    .RESET_B(net104),
    .Q(\genblk2[1].wave_shpr.div.acc[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12907_ (.CLK(clknet_leaf_36_clk),
    .D(_00238_),
    .RESET_B(net102),
    .Q(\genblk2[1].wave_shpr.div.acc[5] ));
 sky130_fd_sc_hd__dfrtp_2 _12908_ (.CLK(clknet_leaf_36_clk),
    .D(_00239_),
    .RESET_B(net103),
    .Q(\genblk2[1].wave_shpr.div.acc[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12909_ (.CLK(clknet_leaf_31_clk),
    .D(_00240_),
    .RESET_B(net100),
    .Q(\genblk2[1].wave_shpr.div.acc[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12910_ (.CLK(clknet_leaf_33_clk),
    .D(_00241_),
    .RESET_B(net100),
    .Q(\genblk2[1].wave_shpr.div.acc[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12911_ (.CLK(clknet_leaf_34_clk),
    .D(_00242_),
    .RESET_B(net107),
    .Q(\genblk2[1].wave_shpr.div.acc[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12912_ (.CLK(clknet_leaf_34_clk),
    .D(_00243_),
    .RESET_B(net107),
    .Q(\genblk2[1].wave_shpr.div.acc[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12913_ (.CLK(clknet_leaf_34_clk),
    .D(_00244_),
    .RESET_B(net106),
    .Q(\genblk2[1].wave_shpr.div.acc[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12914_ (.CLK(clknet_leaf_36_clk),
    .D(net367),
    .RESET_B(net106),
    .Q(\genblk2[1].wave_shpr.div.acc[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12915_ (.CLK(clknet_leaf_36_clk),
    .D(_00246_),
    .RESET_B(net105),
    .Q(\genblk2[1].wave_shpr.div.acc[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12916_ (.CLK(clknet_leaf_35_clk),
    .D(_00247_),
    .RESET_B(net105),
    .Q(\genblk2[1].wave_shpr.div.acc[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12917_ (.CLK(clknet_leaf_35_clk),
    .D(_00248_),
    .RESET_B(net105),
    .Q(\genblk2[1].wave_shpr.div.acc[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12918_ (.CLK(clknet_leaf_39_clk),
    .D(_00249_),
    .RESET_B(net115),
    .Q(\genblk2[1].wave_shpr.div.acc[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12919_ (.CLK(clknet_leaf_39_clk),
    .D(_00250_),
    .RESET_B(net115),
    .Q(\genblk2[1].wave_shpr.div.acc[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12920_ (.CLK(clknet_leaf_35_clk),
    .D(_00251_),
    .RESET_B(net118),
    .Q(\genblk2[1].wave_shpr.div.acc[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12921_ (.CLK(clknet_leaf_35_clk),
    .D(_00252_),
    .RESET_B(net105),
    .Q(\genblk2[1].wave_shpr.div.acc[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12922_ (.CLK(clknet_leaf_35_clk),
    .D(_00253_),
    .RESET_B(net105),
    .Q(\genblk2[1].wave_shpr.div.acc[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12923_ (.CLK(clknet_leaf_35_clk),
    .D(_00254_),
    .RESET_B(net105),
    .Q(\genblk2[1].wave_shpr.div.acc[21] ));
 sky130_fd_sc_hd__dfrtp_2 _12924_ (.CLK(clknet_leaf_35_clk),
    .D(_00255_),
    .RESET_B(net105),
    .Q(\genblk2[1].wave_shpr.div.acc[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12925_ (.CLK(clknet_leaf_35_clk),
    .D(_00256_),
    .RESET_B(net106),
    .Q(\genblk2[1].wave_shpr.div.acc[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12926_ (.CLK(clknet_leaf_35_clk),
    .D(_00257_),
    .RESET_B(net106),
    .Q(\genblk2[1].wave_shpr.div.acc[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12927_ (.CLK(clknet_leaf_35_clk),
    .D(_00258_),
    .RESET_B(net106),
    .Q(\genblk2[1].wave_shpr.div.acc[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12928_ (.CLK(clknet_leaf_35_clk),
    .D(_00259_),
    .RESET_B(net118),
    .Q(\genblk2[1].wave_shpr.div.acc[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12929_ (.CLK(clknet_leaf_123_clk),
    .D(_00008_),
    .RESET_B(net76),
    .Q(\genblk2[2].wave_shpr.div.busy ));
 sky130_fd_sc_hd__dfrtp_1 _12930_ (.CLK(clknet_leaf_116_clk),
    .D(_00009_),
    .RESET_B(net150),
    .Q(\genblk2[2].wave_shpr.div.done ));
 sky130_fd_sc_hd__dfrtp_2 _12931_ (.CLK(clknet_leaf_31_clk),
    .D(_00260_),
    .RESET_B(net102),
    .Q(\genblk2[1].wave_shpr.div.i[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12932_ (.CLK(clknet_leaf_31_clk),
    .D(_00261_),
    .RESET_B(net103),
    .Q(\genblk2[1].wave_shpr.div.i[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12933_ (.CLK(clknet_leaf_31_clk),
    .D(_00262_),
    .RESET_B(net102),
    .Q(\genblk2[1].wave_shpr.div.i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12934_ (.CLK(clknet_leaf_30_clk),
    .D(_00263_),
    .RESET_B(net102),
    .Q(\genblk2[1].wave_shpr.div.i[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12935_ (.CLK(clknet_leaf_30_clk),
    .D(_00264_),
    .RESET_B(net102),
    .Q(\genblk2[1].wave_shpr.div.i[4] ));
 sky130_fd_sc_hd__dfrtp_4 _12936_ (.CLK(clknet_leaf_113_clk),
    .D(_00265_),
    .RESET_B(net130),
    .Q(\genblk2[2].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__dfrtp_2 _12937_ (.CLK(clknet_leaf_111_clk),
    .D(_00266_),
    .RESET_B(net130),
    .Q(\genblk2[2].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12938_ (.CLK(clknet_leaf_111_clk),
    .D(_00267_),
    .RESET_B(net136),
    .Q(\genblk2[2].wave_shpr.div.fin_quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12939_ (.CLK(clknet_leaf_110_clk),
    .D(_00268_),
    .RESET_B(net136),
    .Q(\genblk2[2].wave_shpr.div.fin_quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12940_ (.CLK(clknet_leaf_110_clk),
    .D(_00269_),
    .RESET_B(net136),
    .Q(\genblk2[2].wave_shpr.div.fin_quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12941_ (.CLK(clknet_leaf_111_clk),
    .D(_00270_),
    .RESET_B(net136),
    .Q(\genblk2[2].wave_shpr.div.fin_quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12942_ (.CLK(clknet_leaf_111_clk),
    .D(_00271_),
    .RESET_B(net130),
    .Q(\genblk2[2].wave_shpr.div.fin_quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12943_ (.CLK(clknet_leaf_111_clk),
    .D(_00272_),
    .RESET_B(net130),
    .Q(\genblk2[2].wave_shpr.div.fin_quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12944_ (.CLK(clknet_leaf_2_clk),
    .D(_00273_),
    .RESET_B(net42),
    .Q(\genblk2[3].wave_shpr.div.b1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12945_ (.CLK(clknet_leaf_13_clk),
    .D(_00274_),
    .RESET_B(net69),
    .Q(\genblk2[3].wave_shpr.div.b1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12946_ (.CLK(clknet_leaf_125_clk),
    .D(_00275_),
    .RESET_B(net69),
    .Q(\genblk2[3].wave_shpr.div.b1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12947_ (.CLK(clknet_leaf_125_clk),
    .D(_00276_),
    .RESET_B(net69),
    .Q(\genblk2[3].wave_shpr.div.b1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12948_ (.CLK(clknet_leaf_125_clk),
    .D(_00277_),
    .RESET_B(net71),
    .Q(\genblk2[3].wave_shpr.div.b1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12949_ (.CLK(clknet_leaf_121_clk),
    .D(_00278_),
    .RESET_B(net77),
    .Q(\genblk2[3].wave_shpr.div.b1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12950_ (.CLK(clknet_leaf_125_clk),
    .D(_00279_),
    .RESET_B(net71),
    .Q(\genblk2[3].wave_shpr.div.b1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12951_ (.CLK(clknet_leaf_125_clk),
    .D(_00280_),
    .RESET_B(net71),
    .Q(\genblk2[3].wave_shpr.div.b1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12952_ (.CLK(clknet_leaf_125_clk),
    .D(_00281_),
    .RESET_B(net61),
    .Q(\genblk2[3].wave_shpr.div.b1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12953_ (.CLK(clknet_leaf_136_clk),
    .D(_00282_),
    .RESET_B(net62),
    .Q(\genblk2[3].wave_shpr.div.b1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12954_ (.CLK(clknet_leaf_136_clk),
    .D(_00283_),
    .RESET_B(net62),
    .Q(\genblk2[3].wave_shpr.div.b1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12955_ (.CLK(clknet_leaf_136_clk),
    .D(_00284_),
    .RESET_B(net62),
    .Q(\genblk2[3].wave_shpr.div.b1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12956_ (.CLK(clknet_leaf_136_clk),
    .D(_00285_),
    .RESET_B(net42),
    .Q(\genblk2[3].wave_shpr.div.b1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12957_ (.CLK(clknet_leaf_114_clk),
    .D(_00286_),
    .RESET_B(net132),
    .Q(\genblk2[3].wave_shpr.div.b1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12958_ (.CLK(clknet_leaf_136_clk),
    .D(_00287_),
    .RESET_B(net42),
    .Q(\genblk2[3].wave_shpr.div.b1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12959_ (.CLK(clknet_leaf_136_clk),
    .D(_00288_),
    .RESET_B(net42),
    .Q(\genblk2[3].wave_shpr.div.b1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12960_ (.CLK(clknet_leaf_137_clk),
    .D(_00289_),
    .RESET_B(net39),
    .Q(\genblk2[3].wave_shpr.div.b1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12961_ (.CLK(clknet_leaf_139_clk),
    .D(_00290_),
    .RESET_B(net39),
    .Q(\genblk2[3].wave_shpr.div.b1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12962_ (.CLK(clknet_leaf_130_clk),
    .D(_00291_),
    .RESET_B(net65),
    .Q(\genblk2[2].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12963_ (.CLK(clknet_leaf_111_clk),
    .D(_00292_),
    .RESET_B(net130),
    .Q(\genblk2[2].wave_shpr.div.quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12964_ (.CLK(clknet_leaf_111_clk),
    .D(_00293_),
    .RESET_B(net130),
    .Q(\genblk2[2].wave_shpr.div.quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12965_ (.CLK(clknet_leaf_110_clk),
    .D(_00294_),
    .RESET_B(net130),
    .Q(\genblk2[2].wave_shpr.div.quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12966_ (.CLK(clknet_leaf_111_clk),
    .D(net337),
    .RESET_B(net130),
    .Q(\genblk2[2].wave_shpr.div.quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12967_ (.CLK(clknet_leaf_111_clk),
    .D(net697),
    .RESET_B(net130),
    .Q(\genblk2[2].wave_shpr.div.quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12968_ (.CLK(clknet_leaf_111_clk),
    .D(_00297_),
    .RESET_B(net130),
    .Q(\genblk2[2].wave_shpr.div.quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12969_ (.CLK(clknet_leaf_111_clk),
    .D(_00298_),
    .RESET_B(net128),
    .Q(\genblk2[2].wave_shpr.div.quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12970_ (.CLK(clknet_leaf_113_clk),
    .D(net276),
    .RESET_B(net128),
    .Q(\genblk2[2].wave_shpr.div.quo[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12971_ (.CLK(clknet_leaf_125_clk),
    .D(net301),
    .RESET_B(net71),
    .Q(\genblk2[2].wave_shpr.div.quo[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12972_ (.CLK(clknet_leaf_125_clk),
    .D(_00301_),
    .RESET_B(net71),
    .Q(\genblk2[2].wave_shpr.div.quo[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12973_ (.CLK(clknet_leaf_124_clk),
    .D(net442),
    .RESET_B(net71),
    .Q(\genblk2[2].wave_shpr.div.quo[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12974_ (.CLK(clknet_leaf_124_clk),
    .D(net554),
    .RESET_B(net71),
    .Q(\genblk2[2].wave_shpr.div.quo[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12975_ (.CLK(clknet_leaf_124_clk),
    .D(_00304_),
    .RESET_B(net71),
    .Q(\genblk2[2].wave_shpr.div.quo[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12976_ (.CLK(clknet_leaf_123_clk),
    .D(net458),
    .RESET_B(net71),
    .Q(\genblk2[2].wave_shpr.div.quo[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12977_ (.CLK(clknet_leaf_123_clk),
    .D(_00306_),
    .RESET_B(net72),
    .Q(\genblk2[2].wave_shpr.div.quo[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12978_ (.CLK(clknet_leaf_124_clk),
    .D(net316),
    .RESET_B(net72),
    .Q(\genblk2[2].wave_shpr.div.quo[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12979_ (.CLK(clknet_leaf_124_clk),
    .D(_00308_),
    .RESET_B(net72),
    .Q(\genblk2[2].wave_shpr.div.quo[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12980_ (.CLK(clknet_leaf_14_clk),
    .D(_00309_),
    .RESET_B(net72),
    .Q(\genblk2[2].wave_shpr.div.quo[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12981_ (.CLK(clknet_leaf_124_clk),
    .D(_00310_),
    .RESET_B(net75),
    .Q(\genblk2[2].wave_shpr.div.quo[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12982_ (.CLK(clknet_leaf_125_clk),
    .D(net323),
    .RESET_B(net70),
    .Q(\genblk2[2].wave_shpr.div.quo[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12983_ (.CLK(clknet_leaf_125_clk),
    .D(_00312_),
    .RESET_B(net69),
    .Q(\genblk2[2].wave_shpr.div.quo[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12984_ (.CLK(clknet_leaf_13_clk),
    .D(net262),
    .RESET_B(net69),
    .Q(\genblk2[2].wave_shpr.div.quo[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12985_ (.CLK(clknet_leaf_13_clk),
    .D(_00314_),
    .RESET_B(net69),
    .Q(\genblk2[2].wave_shpr.div.quo[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12986_ (.CLK(clknet_leaf_13_clk),
    .D(_00315_),
    .RESET_B(net69),
    .Q(\genblk2[2].wave_shpr.div.quo[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12987_ (.CLK(clknet_leaf_125_clk),
    .D(net260),
    .RESET_B(net69),
    .Q(\genblk2[2].wave_shpr.div.acc_next[0] ));
 sky130_fd_sc_hd__dfrtp_2 _12988_ (.CLK(clknet_leaf_124_clk),
    .D(net915),
    .RESET_B(net71),
    .Q(\genblk2[2].wave_shpr.div.acc[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12989_ (.CLK(clknet_leaf_132_clk),
    .D(_00318_),
    .RESET_B(net64),
    .Q(\genblk2[2].wave_shpr.div.acc[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12990_ (.CLK(clknet_leaf_131_clk),
    .D(_00319_),
    .RESET_B(net65),
    .Q(\genblk2[2].wave_shpr.div.acc[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12991_ (.CLK(clknet_leaf_130_clk),
    .D(_00320_),
    .RESET_B(net65),
    .Q(\genblk2[2].wave_shpr.div.acc[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12992_ (.CLK(clknet_leaf_131_clk),
    .D(_00321_),
    .RESET_B(net64),
    .Q(\genblk2[2].wave_shpr.div.acc[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12993_ (.CLK(clknet_leaf_131_clk),
    .D(_00322_),
    .RESET_B(net64),
    .Q(\genblk2[2].wave_shpr.div.acc[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12994_ (.CLK(clknet_leaf_131_clk),
    .D(_00323_),
    .RESET_B(net64),
    .Q(\genblk2[2].wave_shpr.div.acc[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12995_ (.CLK(clknet_leaf_131_clk),
    .D(_00324_),
    .RESET_B(net64),
    .Q(\genblk2[2].wave_shpr.div.acc[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12996_ (.CLK(clknet_leaf_132_clk),
    .D(_00325_),
    .RESET_B(net60),
    .Q(\genblk2[2].wave_shpr.div.acc[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12997_ (.CLK(clknet_leaf_132_clk),
    .D(_00326_),
    .RESET_B(net60),
    .Q(\genblk2[2].wave_shpr.div.acc[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12998_ (.CLK(clknet_leaf_131_clk),
    .D(_00327_),
    .RESET_B(net64),
    .Q(\genblk2[2].wave_shpr.div.acc[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12999_ (.CLK(clknet_leaf_132_clk),
    .D(_00328_),
    .RESET_B(net60),
    .Q(\genblk2[2].wave_shpr.div.acc[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13000_ (.CLK(clknet_leaf_132_clk),
    .D(_00329_),
    .RESET_B(net63),
    .Q(\genblk2[2].wave_shpr.div.acc[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13001_ (.CLK(clknet_leaf_133_clk),
    .D(_00330_),
    .RESET_B(net59),
    .Q(\genblk2[2].wave_shpr.div.acc[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13002_ (.CLK(clknet_leaf_133_clk),
    .D(_00331_),
    .RESET_B(net59),
    .Q(\genblk2[2].wave_shpr.div.acc[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13003_ (.CLK(clknet_leaf_133_clk),
    .D(_00332_),
    .RESET_B(net59),
    .Q(\genblk2[2].wave_shpr.div.acc[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13004_ (.CLK(clknet_leaf_138_clk),
    .D(_00333_),
    .RESET_B(net39),
    .Q(\genblk2[2].wave_shpr.div.acc[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13005_ (.CLK(clknet_leaf_138_clk),
    .D(_00334_),
    .RESET_B(net40),
    .Q(\genblk2[2].wave_shpr.div.acc[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13006_ (.CLK(clknet_leaf_133_clk),
    .D(net581),
    .RESET_B(net40),
    .Q(\genblk2[2].wave_shpr.div.acc[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13007_ (.CLK(clknet_leaf_138_clk),
    .D(net606),
    .RESET_B(net40),
    .Q(\genblk2[2].wave_shpr.div.acc[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13008_ (.CLK(clknet_leaf_133_clk),
    .D(_00337_),
    .RESET_B(net59),
    .Q(\genblk2[2].wave_shpr.div.acc[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13009_ (.CLK(clknet_leaf_133_clk),
    .D(_00338_),
    .RESET_B(net59),
    .Q(\genblk2[2].wave_shpr.div.acc[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13010_ (.CLK(clknet_leaf_133_clk),
    .D(_00339_),
    .RESET_B(net59),
    .Q(\genblk2[2].wave_shpr.div.acc[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13011_ (.CLK(clknet_leaf_133_clk),
    .D(_00340_),
    .RESET_B(net59),
    .Q(\genblk2[2].wave_shpr.div.acc[23] ));
 sky130_fd_sc_hd__dfrtp_2 _13012_ (.CLK(clknet_leaf_133_clk),
    .D(_00341_),
    .RESET_B(net60),
    .Q(\genblk2[2].wave_shpr.div.acc[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13013_ (.CLK(clknet_leaf_133_clk),
    .D(_00342_),
    .RESET_B(net60),
    .Q(\genblk2[2].wave_shpr.div.acc[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13014_ (.CLK(clknet_leaf_132_clk),
    .D(_00343_),
    .RESET_B(net60),
    .Q(\genblk2[2].wave_shpr.div.acc[26] ));
 sky130_fd_sc_hd__dfrtp_1 _13015_ (.CLK(clknet_leaf_12_clk),
    .D(_00010_),
    .RESET_B(net52),
    .Q(\genblk2[3].wave_shpr.div.busy ));
 sky130_fd_sc_hd__dfrtp_1 _13016_ (.CLK(clknet_leaf_121_clk),
    .D(_00011_),
    .RESET_B(net77),
    .Q(\genblk2[3].wave_shpr.div.done ));
 sky130_fd_sc_hd__dfrtp_2 _13017_ (.CLK(clknet_leaf_124_clk),
    .D(_00344_),
    .RESET_B(net76),
    .Q(\genblk2[2].wave_shpr.div.i[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13018_ (.CLK(clknet_leaf_123_clk),
    .D(_00345_),
    .RESET_B(net76),
    .Q(\genblk2[2].wave_shpr.div.i[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13019_ (.CLK(clknet_leaf_123_clk),
    .D(_00346_),
    .RESET_B(net76),
    .Q(\genblk2[2].wave_shpr.div.i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13020_ (.CLK(clknet_leaf_123_clk),
    .D(_00347_),
    .RESET_B(net77),
    .Q(\genblk2[2].wave_shpr.div.i[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13021_ (.CLK(clknet_leaf_122_clk),
    .D(_00348_),
    .RESET_B(net76),
    .Q(\genblk2[2].wave_shpr.div.i[4] ));
 sky130_fd_sc_hd__dfrtp_2 _13022_ (.CLK(clknet_leaf_128_clk),
    .D(_00349_),
    .RESET_B(net67),
    .Q(\genblk2[3].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__dfrtp_2 _13023_ (.CLK(clknet_leaf_113_clk),
    .D(_00350_),
    .RESET_B(net128),
    .Q(\genblk2[3].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__dfrtp_2 _13024_ (.CLK(clknet_leaf_114_clk),
    .D(_00351_),
    .RESET_B(net132),
    .Q(\genblk2[3].wave_shpr.div.fin_quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13025_ (.CLK(clknet_leaf_113_clk),
    .D(_00352_),
    .RESET_B(net134),
    .Q(\genblk2[3].wave_shpr.div.fin_quo[3] ));
 sky130_fd_sc_hd__dfrtp_2 _13026_ (.CLK(clknet_leaf_113_clk),
    .D(_00353_),
    .RESET_B(net134),
    .Q(\genblk2[3].wave_shpr.div.fin_quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13027_ (.CLK(clknet_leaf_113_clk),
    .D(_00354_),
    .RESET_B(net131),
    .Q(\genblk2[3].wave_shpr.div.fin_quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13028_ (.CLK(clknet_leaf_113_clk),
    .D(_00355_),
    .RESET_B(net131),
    .Q(\genblk2[3].wave_shpr.div.fin_quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13029_ (.CLK(clknet_leaf_113_clk),
    .D(_00356_),
    .RESET_B(net131),
    .Q(\genblk2[3].wave_shpr.div.fin_quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13030_ (.CLK(clknet_leaf_122_clk),
    .D(_00357_),
    .RESET_B(net79),
    .Q(\genblk2[4].wave_shpr.div.b1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13031_ (.CLK(clknet_leaf_122_clk),
    .D(_00358_),
    .RESET_B(net79),
    .Q(\genblk2[4].wave_shpr.div.b1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13032_ (.CLK(clknet_leaf_121_clk),
    .D(_00359_),
    .RESET_B(net78),
    .Q(\genblk2[4].wave_shpr.div.b1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13033_ (.CLK(clknet_leaf_123_clk),
    .D(_00360_),
    .RESET_B(net79),
    .Q(\genblk2[4].wave_shpr.div.b1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13034_ (.CLK(clknet_leaf_127_clk),
    .D(_00361_),
    .RESET_B(net66),
    .Q(\genblk2[4].wave_shpr.div.b1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13035_ (.CLK(clknet_leaf_122_clk),
    .D(_00362_),
    .RESET_B(net76),
    .Q(\genblk2[4].wave_shpr.div.b1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13036_ (.CLK(clknet_leaf_123_clk),
    .D(_00363_),
    .RESET_B(net76),
    .Q(\genblk2[4].wave_shpr.div.b1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13037_ (.CLK(clknet_leaf_125_clk),
    .D(_00364_),
    .RESET_B(net72),
    .Q(\genblk2[4].wave_shpr.div.b1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13038_ (.CLK(clknet_leaf_126_clk),
    .D(_00365_),
    .RESET_B(net66),
    .Q(\genblk2[4].wave_shpr.div.b1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13039_ (.CLK(clknet_leaf_126_clk),
    .D(_00366_),
    .RESET_B(net61),
    .Q(\genblk2[4].wave_shpr.div.b1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13040_ (.CLK(clknet_leaf_126_clk),
    .D(_00367_),
    .RESET_B(net61),
    .Q(\genblk2[4].wave_shpr.div.b1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13041_ (.CLK(clknet_leaf_126_clk),
    .D(_00368_),
    .RESET_B(net66),
    .Q(\genblk2[4].wave_shpr.div.b1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13042_ (.CLK(clknet_leaf_128_clk),
    .D(_00369_),
    .RESET_B(net67),
    .Q(\genblk2[4].wave_shpr.div.b1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13043_ (.CLK(clknet_leaf_128_clk),
    .D(_00370_),
    .RESET_B(net66),
    .Q(\genblk2[4].wave_shpr.div.b1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13044_ (.CLK(clknet_leaf_128_clk),
    .D(_00371_),
    .RESET_B(net67),
    .Q(\genblk2[4].wave_shpr.div.b1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13045_ (.CLK(clknet_leaf_128_clk),
    .D(_00372_),
    .RESET_B(net67),
    .Q(\genblk2[4].wave_shpr.div.b1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13046_ (.CLK(clknet_leaf_112_clk),
    .D(_00373_),
    .RESET_B(net128),
    .Q(\genblk2[4].wave_shpr.div.b1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13047_ (.CLK(clknet_leaf_129_clk),
    .D(_00374_),
    .RESET_B(net65),
    .Q(\genblk2[4].wave_shpr.div.b1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13048_ (.CLK(clknet_leaf_135_clk),
    .D(_00375_),
    .RESET_B(net62),
    .Q(\genblk2[3].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13049_ (.CLK(clknet_leaf_112_clk),
    .D(_00376_),
    .RESET_B(net132),
    .Q(\genblk2[3].wave_shpr.div.quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13050_ (.CLK(clknet_leaf_113_clk),
    .D(net327),
    .RESET_B(net128),
    .Q(\genblk2[3].wave_shpr.div.quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13051_ (.CLK(clknet_leaf_113_clk),
    .D(net738),
    .RESET_B(net128),
    .Q(\genblk2[3].wave_shpr.div.quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13052_ (.CLK(clknet_leaf_113_clk),
    .D(net780),
    .RESET_B(net131),
    .Q(\genblk2[3].wave_shpr.div.quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13053_ (.CLK(clknet_leaf_113_clk),
    .D(_00380_),
    .RESET_B(net128),
    .Q(\genblk2[3].wave_shpr.div.quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13054_ (.CLK(clknet_leaf_113_clk),
    .D(net815),
    .RESET_B(net128),
    .Q(\genblk2[3].wave_shpr.div.quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13055_ (.CLK(clknet_leaf_113_clk),
    .D(_00382_),
    .RESET_B(net128),
    .Q(\genblk2[3].wave_shpr.div.quo[7] ));
 sky130_fd_sc_hd__dfrtp_2 _13056_ (.CLK(clknet_leaf_134_clk),
    .D(_00383_),
    .RESET_B(net63),
    .Q(\genblk2[3].wave_shpr.div.quo[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13057_ (.CLK(clknet_leaf_24_clk),
    .D(net539),
    .RESET_B(net92),
    .Q(\genblk2[3].wave_shpr.div.quo[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13058_ (.CLK(clknet_leaf_24_clk),
    .D(_00385_),
    .RESET_B(net92),
    .Q(\genblk2[3].wave_shpr.div.quo[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13059_ (.CLK(clknet_leaf_24_clk),
    .D(_00386_),
    .RESET_B(net92),
    .Q(\genblk2[3].wave_shpr.div.quo[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13060_ (.CLK(clknet_leaf_21_clk),
    .D(_00387_),
    .RESET_B(net95),
    .Q(\genblk2[3].wave_shpr.div.quo[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13061_ (.CLK(clknet_leaf_29_clk),
    .D(net388),
    .RESET_B(net95),
    .Q(\genblk2[3].wave_shpr.div.quo[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13062_ (.CLK(clknet_leaf_29_clk),
    .D(net635),
    .RESET_B(net95),
    .Q(\genblk2[3].wave_shpr.div.quo[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13063_ (.CLK(clknet_leaf_29_clk),
    .D(_00390_),
    .RESET_B(net95),
    .Q(\genblk2[3].wave_shpr.div.quo[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13064_ (.CLK(clknet_leaf_29_clk),
    .D(_00391_),
    .RESET_B(net95),
    .Q(\genblk2[3].wave_shpr.div.quo[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13065_ (.CLK(clknet_leaf_22_clk),
    .D(net377),
    .RESET_B(net95),
    .Q(\genblk2[3].wave_shpr.div.quo[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13066_ (.CLK(clknet_leaf_22_clk),
    .D(net452),
    .RESET_B(net93),
    .Q(\genblk2[3].wave_shpr.div.quo[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13067_ (.CLK(clknet_leaf_22_clk),
    .D(_00394_),
    .RESET_B(net93),
    .Q(\genblk2[3].wave_shpr.div.quo[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13068_ (.CLK(clknet_leaf_24_clk),
    .D(net297),
    .RESET_B(net93),
    .Q(\genblk2[3].wave_shpr.div.quo[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13069_ (.CLK(clknet_leaf_24_clk),
    .D(net546),
    .RESET_B(net93),
    .Q(\genblk2[3].wave_shpr.div.quo[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13070_ (.CLK(clknet_leaf_24_clk),
    .D(_00397_),
    .RESET_B(net92),
    .Q(\genblk2[3].wave_shpr.div.quo[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13071_ (.CLK(clknet_leaf_24_clk),
    .D(_00398_),
    .RESET_B(net92),
    .Q(\genblk2[3].wave_shpr.div.quo[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13072_ (.CLK(clknet_leaf_23_clk),
    .D(net491),
    .RESET_B(net94),
    .Q(\genblk2[3].wave_shpr.div.quo[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13073_ (.CLK(clknet_leaf_23_clk),
    .D(net562),
    .RESET_B(net98),
    .Q(\genblk2[3].wave_shpr.div.acc_next[0] ));
 sky130_fd_sc_hd__dfrtp_2 _13074_ (.CLK(clknet_leaf_11_clk),
    .D(net437),
    .RESET_B(net56),
    .Q(\genblk2[3].wave_shpr.div.acc[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13075_ (.CLK(clknet_leaf_2_clk),
    .D(_00402_),
    .RESET_B(net42),
    .Q(\genblk2[3].wave_shpr.div.acc[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13076_ (.CLK(clknet_leaf_136_clk),
    .D(_00403_),
    .RESET_B(net62),
    .Q(\genblk2[3].wave_shpr.div.acc[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13077_ (.CLK(clknet_leaf_125_clk),
    .D(_00404_),
    .RESET_B(net62),
    .Q(\genblk2[3].wave_shpr.div.acc[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13078_ (.CLK(clknet_leaf_125_clk),
    .D(_00405_),
    .RESET_B(net61),
    .Q(\genblk2[3].wave_shpr.div.acc[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13079_ (.CLK(clknet_leaf_125_clk),
    .D(_00406_),
    .RESET_B(net61),
    .Q(\genblk2[3].wave_shpr.div.acc[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13080_ (.CLK(clknet_leaf_125_clk),
    .D(_00407_),
    .RESET_B(net63),
    .Q(\genblk2[3].wave_shpr.div.acc[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13081_ (.CLK(clknet_leaf_126_clk),
    .D(_00408_),
    .RESET_B(net63),
    .Q(\genblk2[3].wave_shpr.div.acc[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13082_ (.CLK(clknet_leaf_126_clk),
    .D(_00409_),
    .RESET_B(net61),
    .Q(\genblk2[3].wave_shpr.div.acc[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13083_ (.CLK(clknet_leaf_135_clk),
    .D(_00410_),
    .RESET_B(net61),
    .Q(\genblk2[3].wave_shpr.div.acc[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13084_ (.CLK(clknet_leaf_135_clk),
    .D(_00411_),
    .RESET_B(net62),
    .Q(\genblk2[3].wave_shpr.div.acc[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13085_ (.CLK(clknet_leaf_135_clk),
    .D(_00412_),
    .RESET_B(net62),
    .Q(\genblk2[3].wave_shpr.div.acc[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13086_ (.CLK(clknet_leaf_136_clk),
    .D(net943),
    .RESET_B(net42),
    .Q(\genblk2[3].wave_shpr.div.acc[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13087_ (.CLK(clknet_leaf_136_clk),
    .D(_00414_),
    .RESET_B(net42),
    .Q(\genblk2[3].wave_shpr.div.acc[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13088_ (.CLK(clknet_leaf_137_clk),
    .D(_00415_),
    .RESET_B(net40),
    .Q(\genblk2[3].wave_shpr.div.acc[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13089_ (.CLK(clknet_leaf_137_clk),
    .D(_00416_),
    .RESET_B(net40),
    .Q(\genblk2[3].wave_shpr.div.acc[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13090_ (.CLK(clknet_leaf_137_clk),
    .D(_00417_),
    .RESET_B(net39),
    .Q(\genblk2[3].wave_shpr.div.acc[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13091_ (.CLK(clknet_leaf_137_clk),
    .D(_00418_),
    .RESET_B(net39),
    .Q(\genblk2[3].wave_shpr.div.acc[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13092_ (.CLK(clknet_leaf_137_clk),
    .D(_00419_),
    .RESET_B(net39),
    .Q(\genblk2[3].wave_shpr.div.acc[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13093_ (.CLK(clknet_leaf_139_clk),
    .D(_00420_),
    .RESET_B(net39),
    .Q(\genblk2[3].wave_shpr.div.acc[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13094_ (.CLK(clknet_leaf_1_clk),
    .D(_00421_),
    .RESET_B(net38),
    .Q(\genblk2[3].wave_shpr.div.acc[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13095_ (.CLK(clknet_leaf_1_clk),
    .D(_00422_),
    .RESET_B(net41),
    .Q(\genblk2[3].wave_shpr.div.acc[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13096_ (.CLK(clknet_leaf_137_clk),
    .D(_00423_),
    .RESET_B(net41),
    .Q(\genblk2[3].wave_shpr.div.acc[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13097_ (.CLK(clknet_leaf_137_clk),
    .D(_00424_),
    .RESET_B(net41),
    .Q(\genblk2[3].wave_shpr.div.acc[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13098_ (.CLK(clknet_leaf_137_clk),
    .D(_00425_),
    .RESET_B(net39),
    .Q(\genblk2[3].wave_shpr.div.acc[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13099_ (.CLK(clknet_leaf_137_clk),
    .D(_00426_),
    .RESET_B(net42),
    .Q(\genblk2[3].wave_shpr.div.acc[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13100_ (.CLK(clknet_leaf_136_clk),
    .D(_00427_),
    .RESET_B(net42),
    .Q(\genblk2[3].wave_shpr.div.acc[26] ));
 sky130_fd_sc_hd__dfrtp_1 _13101_ (.CLK(clknet_leaf_122_clk),
    .D(_00012_),
    .RESET_B(net78),
    .Q(\genblk2[4].wave_shpr.div.busy ));
 sky130_fd_sc_hd__dfrtp_1 _13102_ (.CLK(clknet_leaf_118_clk),
    .D(_00013_),
    .RESET_B(net139),
    .Q(\genblk2[4].wave_shpr.div.done ));
 sky130_fd_sc_hd__dfrtp_2 _13103_ (.CLK(clknet_leaf_12_clk),
    .D(_00428_),
    .RESET_B(net51),
    .Q(\genblk2[3].wave_shpr.div.i[0] ));
 sky130_fd_sc_hd__dfrtp_2 _13104_ (.CLK(clknet_leaf_13_clk),
    .D(_00429_),
    .RESET_B(net52),
    .Q(\genblk2[3].wave_shpr.div.i[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13105_ (.CLK(clknet_leaf_12_clk),
    .D(_00430_),
    .RESET_B(net52),
    .Q(\genblk2[3].wave_shpr.div.i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13106_ (.CLK(clknet_leaf_12_clk),
    .D(_00431_),
    .RESET_B(net52),
    .Q(\genblk2[3].wave_shpr.div.i[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13107_ (.CLK(clknet_leaf_13_clk),
    .D(_00432_),
    .RESET_B(net53),
    .Q(\genblk2[3].wave_shpr.div.i[4] ));
 sky130_fd_sc_hd__dfrtp_4 _13108_ (.CLK(clknet_leaf_127_clk),
    .D(_00433_),
    .RESET_B(net133),
    .Q(\genblk2[4].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__dfrtp_2 _13109_ (.CLK(clknet_leaf_114_clk),
    .D(_00434_),
    .RESET_B(net133),
    .Q(\genblk2[4].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13110_ (.CLK(clknet_leaf_114_clk),
    .D(_00435_),
    .RESET_B(net133),
    .Q(\genblk2[4].wave_shpr.div.fin_quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13111_ (.CLK(clknet_leaf_115_clk),
    .D(_00436_),
    .RESET_B(net134),
    .Q(\genblk2[4].wave_shpr.div.fin_quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13112_ (.CLK(clknet_leaf_115_clk),
    .D(_00437_),
    .RESET_B(net134),
    .Q(\genblk2[4].wave_shpr.div.fin_quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13113_ (.CLK(clknet_leaf_115_clk),
    .D(_00438_),
    .RESET_B(net134),
    .Q(\genblk2[4].wave_shpr.div.fin_quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13114_ (.CLK(clknet_leaf_115_clk),
    .D(_00439_),
    .RESET_B(net135),
    .Q(\genblk2[4].wave_shpr.div.fin_quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13115_ (.CLK(clknet_leaf_115_clk),
    .D(_00440_),
    .RESET_B(net135),
    .Q(\genblk2[4].wave_shpr.div.fin_quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13116_ (.CLK(clknet_leaf_2_clk),
    .D(_00441_),
    .RESET_B(net52),
    .Q(\genblk2[5].wave_shpr.div.b1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13117_ (.CLK(clknet_leaf_13_clk),
    .D(_00442_),
    .RESET_B(net52),
    .Q(\genblk2[5].wave_shpr.div.b1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13118_ (.CLK(clknet_leaf_125_clk),
    .D(_00443_),
    .RESET_B(net69),
    .Q(\genblk2[5].wave_shpr.div.b1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13119_ (.CLK(clknet_leaf_2_clk),
    .D(_00444_),
    .RESET_B(net51),
    .Q(\genblk2[5].wave_shpr.div.b1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13120_ (.CLK(clknet_leaf_136_clk),
    .D(_00445_),
    .RESET_B(net43),
    .Q(\genblk2[5].wave_shpr.div.b1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13121_ (.CLK(clknet_leaf_136_clk),
    .D(_00446_),
    .RESET_B(net43),
    .Q(\genblk2[5].wave_shpr.div.b1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13122_ (.CLK(clknet_leaf_136_clk),
    .D(_00447_),
    .RESET_B(net43),
    .Q(\genblk2[5].wave_shpr.div.b1[6] ));
 sky130_fd_sc_hd__dfrtp_2 _13123_ (.CLK(clknet_leaf_124_clk),
    .D(_00448_),
    .RESET_B(net77),
    .Q(\genblk2[5].wave_shpr.div.b1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13124_ (.CLK(clknet_leaf_3_clk),
    .D(_00449_),
    .RESET_B(net51),
    .Q(\genblk2[5].wave_shpr.div.b1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13125_ (.CLK(clknet_leaf_3_clk),
    .D(_00450_),
    .RESET_B(net51),
    .Q(\genblk2[5].wave_shpr.div.b1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13126_ (.CLK(clknet_leaf_3_clk),
    .D(_00451_),
    .RESET_B(net51),
    .Q(\genblk2[5].wave_shpr.div.b1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13127_ (.CLK(clknet_leaf_3_clk),
    .D(_00452_),
    .RESET_B(net46),
    .Q(\genblk2[5].wave_shpr.div.b1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13128_ (.CLK(clknet_leaf_3_clk),
    .D(_00453_),
    .RESET_B(net46),
    .Q(\genblk2[5].wave_shpr.div.b1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13129_ (.CLK(clknet_leaf_3_clk),
    .D(_00454_),
    .RESET_B(net46),
    .Q(\genblk2[5].wave_shpr.div.b1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13130_ (.CLK(clknet_leaf_3_clk),
    .D(_00455_),
    .RESET_B(net46),
    .Q(\genblk2[5].wave_shpr.div.b1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13131_ (.CLK(clknet_leaf_4_clk),
    .D(_00456_),
    .RESET_B(net46),
    .Q(\genblk2[5].wave_shpr.div.b1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13132_ (.CLK(clknet_leaf_3_clk),
    .D(_00457_),
    .RESET_B(net46),
    .Q(\genblk2[5].wave_shpr.div.b1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13133_ (.CLK(clknet_leaf_0_clk),
    .D(_00458_),
    .RESET_B(net41),
    .Q(\genblk2[5].wave_shpr.div.b1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13134_ (.CLK(clknet_leaf_115_clk),
    .D(_00459_),
    .RESET_B(net133),
    .Q(\genblk2[4].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13135_ (.CLK(clknet_leaf_114_clk),
    .D(net419),
    .RESET_B(net133),
    .Q(\genblk2[4].wave_shpr.div.quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13136_ (.CLK(clknet_leaf_115_clk),
    .D(net465),
    .RESET_B(net133),
    .Q(\genblk2[4].wave_shpr.div.quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13137_ (.CLK(clknet_leaf_115_clk),
    .D(_00462_),
    .RESET_B(net135),
    .Q(\genblk2[4].wave_shpr.div.quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13138_ (.CLK(clknet_leaf_115_clk),
    .D(net733),
    .RESET_B(net135),
    .Q(\genblk2[4].wave_shpr.div.quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13139_ (.CLK(clknet_leaf_115_clk),
    .D(net750),
    .RESET_B(net133),
    .Q(\genblk2[4].wave_shpr.div.quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13140_ (.CLK(clknet_leaf_115_clk),
    .D(_00465_),
    .RESET_B(net133),
    .Q(\genblk2[4].wave_shpr.div.quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13141_ (.CLK(clknet_leaf_115_clk),
    .D(_00466_),
    .RESET_B(net135),
    .Q(\genblk2[4].wave_shpr.div.quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13142_ (.CLK(clknet_leaf_115_clk),
    .D(_00467_),
    .RESET_B(net135),
    .Q(\genblk2[4].wave_shpr.div.quo[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13143_ (.CLK(clknet_leaf_121_clk),
    .D(net252),
    .RESET_B(net81),
    .Q(\genblk2[4].wave_shpr.div.quo[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13144_ (.CLK(clknet_leaf_121_clk),
    .D(net673),
    .RESET_B(net81),
    .Q(\genblk2[4].wave_shpr.div.quo[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13145_ (.CLK(clknet_leaf_121_clk),
    .D(net603),
    .RESET_B(net81),
    .Q(\genblk2[4].wave_shpr.div.quo[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13146_ (.CLK(clknet_leaf_121_clk),
    .D(_00471_),
    .RESET_B(net81),
    .Q(\genblk2[4].wave_shpr.div.quo[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13147_ (.CLK(clknet_leaf_121_clk),
    .D(net638),
    .RESET_B(net80),
    .Q(\genblk2[4].wave_shpr.div.quo[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13148_ (.CLK(clknet_leaf_121_clk),
    .D(_00473_),
    .RESET_B(net81),
    .Q(\genblk2[4].wave_shpr.div.quo[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13149_ (.CLK(clknet_leaf_121_clk),
    .D(net597),
    .RESET_B(net80),
    .Q(\genblk2[4].wave_shpr.div.quo[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13150_ (.CLK(clknet_leaf_121_clk),
    .D(net681),
    .RESET_B(net80),
    .Q(\genblk2[4].wave_shpr.div.quo[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13151_ (.CLK(clknet_leaf_17_clk),
    .D(net532),
    .RESET_B(net80),
    .Q(\genblk2[4].wave_shpr.div.quo[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13152_ (.CLK(clknet_leaf_17_clk),
    .D(_00477_),
    .RESET_B(net80),
    .Q(\genblk2[4].wave_shpr.div.quo[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13153_ (.CLK(clknet_leaf_121_clk),
    .D(net256),
    .RESET_B(net77),
    .Q(\genblk2[4].wave_shpr.div.quo[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13154_ (.CLK(clknet_leaf_121_clk),
    .D(_00479_),
    .RESET_B(net77),
    .Q(\genblk2[4].wave_shpr.div.quo[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13155_ (.CLK(clknet_leaf_121_clk),
    .D(net627),
    .RESET_B(net80),
    .Q(\genblk2[4].wave_shpr.div.quo[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13156_ (.CLK(clknet_leaf_121_clk),
    .D(net666),
    .RESET_B(net78),
    .Q(\genblk2[4].wave_shpr.div.quo[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13157_ (.CLK(clknet_leaf_121_clk),
    .D(_00482_),
    .RESET_B(net78),
    .Q(\genblk2[4].wave_shpr.div.quo[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13158_ (.CLK(clknet_leaf_121_clk),
    .D(_00483_),
    .RESET_B(net78),
    .Q(\genblk2[4].wave_shpr.div.quo[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13159_ (.CLK(clknet_leaf_121_clk),
    .D(net644),
    .RESET_B(net78),
    .Q(\genblk2[4].wave_shpr.div.acc_next[0] ));
 sky130_fd_sc_hd__dfrtp_2 _13160_ (.CLK(clknet_leaf_122_clk),
    .D(_00485_),
    .RESET_B(net78),
    .Q(\genblk2[4].wave_shpr.div.acc[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13161_ (.CLK(clknet_leaf_122_clk),
    .D(_00486_),
    .RESET_B(net79),
    .Q(\genblk2[4].wave_shpr.div.acc[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13162_ (.CLK(clknet_leaf_115_clk),
    .D(_00487_),
    .RESET_B(net67),
    .Q(\genblk2[4].wave_shpr.div.acc[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13163_ (.CLK(clknet_leaf_114_clk),
    .D(_00488_),
    .RESET_B(net67),
    .Q(\genblk2[4].wave_shpr.div.acc[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13164_ (.CLK(clknet_leaf_127_clk),
    .D(net843),
    .RESET_B(net67),
    .Q(\genblk2[4].wave_shpr.div.acc[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13165_ (.CLK(clknet_leaf_127_clk),
    .D(_00490_),
    .RESET_B(net68),
    .Q(\genblk2[4].wave_shpr.div.acc[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13166_ (.CLK(clknet_leaf_127_clk),
    .D(_00491_),
    .RESET_B(net79),
    .Q(\genblk2[4].wave_shpr.div.acc[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13167_ (.CLK(clknet_leaf_123_clk),
    .D(net972),
    .RESET_B(net76),
    .Q(\genblk2[4].wave_shpr.div.acc[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13168_ (.CLK(clknet_leaf_127_clk),
    .D(_00493_),
    .RESET_B(net66),
    .Q(\genblk2[4].wave_shpr.div.acc[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13169_ (.CLK(clknet_leaf_127_clk),
    .D(_00494_),
    .RESET_B(net66),
    .Q(\genblk2[4].wave_shpr.div.acc[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13170_ (.CLK(clknet_leaf_126_clk),
    .D(_00495_),
    .RESET_B(net68),
    .Q(\genblk2[4].wave_shpr.div.acc[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13171_ (.CLK(clknet_leaf_126_clk),
    .D(_00496_),
    .RESET_B(net66),
    .Q(\genblk2[4].wave_shpr.div.acc[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13172_ (.CLK(clknet_leaf_128_clk),
    .D(_00497_),
    .RESET_B(net66),
    .Q(\genblk2[4].wave_shpr.div.acc[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13173_ (.CLK(clknet_leaf_128_clk),
    .D(_00498_),
    .RESET_B(net66),
    .Q(\genblk2[4].wave_shpr.div.acc[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13174_ (.CLK(clknet_leaf_129_clk),
    .D(_00499_),
    .RESET_B(net65),
    .Q(\genblk2[4].wave_shpr.div.acc[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13175_ (.CLK(clknet_leaf_129_clk),
    .D(_00500_),
    .RESET_B(net67),
    .Q(\genblk2[4].wave_shpr.div.acc[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13176_ (.CLK(clknet_leaf_130_clk),
    .D(_00501_),
    .RESET_B(net65),
    .Q(\genblk2[4].wave_shpr.div.acc[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13177_ (.CLK(clknet_leaf_130_clk),
    .D(_00502_),
    .RESET_B(net65),
    .Q(\genblk2[4].wave_shpr.div.acc[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13178_ (.CLK(clknet_leaf_131_clk),
    .D(_00503_),
    .RESET_B(net65),
    .Q(\genblk2[4].wave_shpr.div.acc[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13179_ (.CLK(clknet_leaf_131_clk),
    .D(_00504_),
    .RESET_B(net65),
    .Q(\genblk2[4].wave_shpr.div.acc[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13180_ (.CLK(clknet_leaf_130_clk),
    .D(_00505_),
    .RESET_B(net68),
    .Q(\genblk2[4].wave_shpr.div.acc[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13181_ (.CLK(clknet_leaf_112_clk),
    .D(_00506_),
    .RESET_B(net68),
    .Q(\genblk2[4].wave_shpr.div.acc[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13182_ (.CLK(clknet_leaf_130_clk),
    .D(net473),
    .RESET_B(net129),
    .Q(\genblk2[4].wave_shpr.div.acc[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13183_ (.CLK(clknet_leaf_112_clk),
    .D(_00508_),
    .RESET_B(net129),
    .Q(\genblk2[4].wave_shpr.div.acc[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13184_ (.CLK(clknet_leaf_112_clk),
    .D(_00509_),
    .RESET_B(net129),
    .Q(\genblk2[4].wave_shpr.div.acc[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13185_ (.CLK(clknet_leaf_112_clk),
    .D(_00510_),
    .RESET_B(net128),
    .Q(\genblk2[4].wave_shpr.div.acc[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13186_ (.CLK(clknet_leaf_112_clk),
    .D(_00511_),
    .RESET_B(net129),
    .Q(\genblk2[4].wave_shpr.div.acc[26] ));
 sky130_fd_sc_hd__dfrtp_1 _13187_ (.CLK(clknet_leaf_11_clk),
    .D(_00014_),
    .RESET_B(net56),
    .Q(\genblk2[5].wave_shpr.div.busy ));
 sky130_fd_sc_hd__dfrtp_1 _13188_ (.CLK(clknet_leaf_118_clk),
    .D(_00015_),
    .RESET_B(net139),
    .Q(\genblk2[5].wave_shpr.div.done ));
 sky130_fd_sc_hd__dfrtp_2 _13189_ (.CLK(clknet_leaf_122_clk),
    .D(_00512_),
    .RESET_B(net78),
    .Q(\genblk2[4].wave_shpr.div.i[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13190_ (.CLK(clknet_leaf_118_clk),
    .D(_00513_),
    .RESET_B(net138),
    .Q(\genblk2[4].wave_shpr.div.i[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13191_ (.CLK(clknet_leaf_122_clk),
    .D(net735),
    .RESET_B(net78),
    .Q(\genblk2[4].wave_shpr.div.i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13192_ (.CLK(clknet_leaf_122_clk),
    .D(_00515_),
    .RESET_B(net79),
    .Q(\genblk2[4].wave_shpr.div.i[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13193_ (.CLK(clknet_leaf_118_clk),
    .D(_00516_),
    .RESET_B(net138),
    .Q(\genblk2[4].wave_shpr.div.i[4] ));
 sky130_fd_sc_hd__dfrtp_4 _13194_ (.CLK(clknet_leaf_127_clk),
    .D(_00517_),
    .RESET_B(net67),
    .Q(\genblk2[5].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__dfrtp_2 _13195_ (.CLK(clknet_leaf_128_clk),
    .D(_00518_),
    .RESET_B(net132),
    .Q(\genblk2[5].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__dfrtp_2 _13196_ (.CLK(clknet_leaf_114_clk),
    .D(_00519_),
    .RESET_B(net134),
    .Q(\genblk2[5].wave_shpr.div.fin_quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13197_ (.CLK(clknet_leaf_113_clk),
    .D(_00520_),
    .RESET_B(net134),
    .Q(\genblk2[5].wave_shpr.div.fin_quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13198_ (.CLK(clknet_leaf_114_clk),
    .D(_00521_),
    .RESET_B(net134),
    .Q(\genblk2[5].wave_shpr.div.fin_quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13199_ (.CLK(clknet_leaf_114_clk),
    .D(_00522_),
    .RESET_B(net134),
    .Q(\genblk2[5].wave_shpr.div.fin_quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13200_ (.CLK(clknet_leaf_115_clk),
    .D(_00523_),
    .RESET_B(net134),
    .Q(\genblk2[5].wave_shpr.div.fin_quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13201_ (.CLK(clknet_leaf_114_clk),
    .D(_00524_),
    .RESET_B(net132),
    .Q(\genblk2[5].wave_shpr.div.fin_quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13202_ (.CLK(clknet_leaf_8_clk),
    .D(_00525_),
    .RESET_B(net55),
    .Q(\genblk2[6].wave_shpr.div.b1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13203_ (.CLK(clknet_leaf_8_clk),
    .D(_00526_),
    .RESET_B(net48),
    .Q(\genblk2[6].wave_shpr.div.b1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13204_ (.CLK(clknet_leaf_8_clk),
    .D(_00527_),
    .RESET_B(net48),
    .Q(\genblk2[6].wave_shpr.div.b1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13205_ (.CLK(clknet_leaf_8_clk),
    .D(_00528_),
    .RESET_B(net48),
    .Q(\genblk2[6].wave_shpr.div.b1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13206_ (.CLK(clknet_leaf_25_clk),
    .D(_00529_),
    .RESET_B(net88),
    .Q(\genblk2[6].wave_shpr.div.b1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13207_ (.CLK(clknet_leaf_25_clk),
    .D(_00530_),
    .RESET_B(net86),
    .Q(\genblk2[6].wave_shpr.div.b1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13208_ (.CLK(clknet_leaf_8_clk),
    .D(_00531_),
    .RESET_B(net88),
    .Q(\genblk2[6].wave_shpr.div.b1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13209_ (.CLK(clknet_leaf_25_clk),
    .D(_00532_),
    .RESET_B(net86),
    .Q(\genblk2[6].wave_shpr.div.b1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13210_ (.CLK(clknet_leaf_25_clk),
    .D(_00533_),
    .RESET_B(net86),
    .Q(\genblk2[6].wave_shpr.div.b1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13211_ (.CLK(clknet_leaf_25_clk),
    .D(_00534_),
    .RESET_B(net86),
    .Q(\genblk2[6].wave_shpr.div.b1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13212_ (.CLK(clknet_leaf_25_clk),
    .D(_00535_),
    .RESET_B(net86),
    .Q(\genblk2[6].wave_shpr.div.b1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13213_ (.CLK(clknet_leaf_7_clk),
    .D(_00536_),
    .RESET_B(net49),
    .Q(\genblk2[6].wave_shpr.div.b1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13214_ (.CLK(clknet_leaf_6_clk),
    .D(_00537_),
    .RESET_B(net48),
    .Q(\genblk2[6].wave_shpr.div.b1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13215_ (.CLK(clknet_leaf_6_clk),
    .D(_00538_),
    .RESET_B(net48),
    .Q(\genblk2[6].wave_shpr.div.b1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13216_ (.CLK(clknet_leaf_6_clk),
    .D(_00539_),
    .RESET_B(net46),
    .Q(\genblk2[6].wave_shpr.div.b1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13217_ (.CLK(clknet_leaf_6_clk),
    .D(_00540_),
    .RESET_B(net48),
    .Q(\genblk2[6].wave_shpr.div.b1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13218_ (.CLK(clknet_leaf_5_clk),
    .D(_00541_),
    .RESET_B(net46),
    .Q(\genblk2[6].wave_shpr.div.b1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13219_ (.CLK(clknet_leaf_3_clk),
    .D(_00542_),
    .RESET_B(net47),
    .Q(\genblk2[6].wave_shpr.div.b1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13220_ (.CLK(clknet_leaf_136_clk),
    .D(_00543_),
    .RESET_B(net62),
    .Q(\genblk2[5].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13221_ (.CLK(clknet_leaf_114_clk),
    .D(_00544_),
    .RESET_B(net132),
    .Q(\genblk2[5].wave_shpr.div.quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13222_ (.CLK(clknet_leaf_114_clk),
    .D(net880),
    .RESET_B(net132),
    .Q(\genblk2[5].wave_shpr.div.quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13223_ (.CLK(clknet_leaf_114_clk),
    .D(_00546_),
    .RESET_B(net132),
    .Q(\genblk2[5].wave_shpr.div.quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13224_ (.CLK(clknet_leaf_114_clk),
    .D(_00547_),
    .RESET_B(net132),
    .Q(\genblk2[5].wave_shpr.div.quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13225_ (.CLK(clknet_leaf_114_clk),
    .D(_00548_),
    .RESET_B(net133),
    .Q(\genblk2[5].wave_shpr.div.quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13226_ (.CLK(clknet_leaf_127_clk),
    .D(net254),
    .RESET_B(net132),
    .Q(\genblk2[5].wave_shpr.div.quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13227_ (.CLK(clknet_leaf_127_clk),
    .D(_00550_),
    .RESET_B(net67),
    .Q(\genblk2[5].wave_shpr.div.quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13228_ (.CLK(clknet_leaf_125_clk),
    .D(net309),
    .RESET_B(net69),
    .Q(\genblk2[5].wave_shpr.div.quo[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13229_ (.CLK(clknet_leaf_15_clk),
    .D(_00552_),
    .RESET_B(net56),
    .Q(\genblk2[5].wave_shpr.div.quo[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13230_ (.CLK(clknet_leaf_11_clk),
    .D(net311),
    .RESET_B(net73),
    .Q(\genblk2[5].wave_shpr.div.quo[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13231_ (.CLK(clknet_leaf_11_clk),
    .D(_00554_),
    .RESET_B(net73),
    .Q(\genblk2[5].wave_shpr.div.quo[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13232_ (.CLK(clknet_leaf_15_clk),
    .D(net501),
    .RESET_B(net73),
    .Q(\genblk2[5].wave_shpr.div.quo[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13233_ (.CLK(clknet_leaf_15_clk),
    .D(_00556_),
    .RESET_B(net73),
    .Q(\genblk2[5].wave_shpr.div.quo[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13234_ (.CLK(clknet_leaf_16_clk),
    .D(net295),
    .RESET_B(net73),
    .Q(\genblk2[5].wave_shpr.div.quo[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13235_ (.CLK(clknet_leaf_15_clk),
    .D(net250),
    .RESET_B(net73),
    .Q(\genblk2[5].wave_shpr.div.quo[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13236_ (.CLK(clknet_leaf_15_clk),
    .D(_00559_),
    .RESET_B(net74),
    .Q(\genblk2[5].wave_shpr.div.quo[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13237_ (.CLK(clknet_leaf_10_clk),
    .D(_00560_),
    .RESET_B(net57),
    .Q(\genblk2[5].wave_shpr.div.quo[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13238_ (.CLK(clknet_leaf_11_clk),
    .D(net236),
    .RESET_B(net57),
    .Q(\genblk2[5].wave_shpr.div.quo[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13239_ (.CLK(clknet_leaf_10_clk),
    .D(_00562_),
    .RESET_B(net57),
    .Q(\genblk2[5].wave_shpr.div.quo[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13240_ (.CLK(clknet_leaf_11_clk),
    .D(net234),
    .RESET_B(net57),
    .Q(\genblk2[5].wave_shpr.div.quo[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13241_ (.CLK(clknet_leaf_10_clk),
    .D(_00564_),
    .RESET_B(net55),
    .Q(\genblk2[5].wave_shpr.div.quo[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13242_ (.CLK(clknet_leaf_9_clk),
    .D(net246),
    .RESET_B(net55),
    .Q(\genblk2[5].wave_shpr.div.quo[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13243_ (.CLK(clknet_leaf_9_clk),
    .D(_00566_),
    .RESET_B(net55),
    .Q(\genblk2[5].wave_shpr.div.quo[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13244_ (.CLK(clknet_leaf_9_clk),
    .D(_00567_),
    .RESET_B(net54),
    .Q(\genblk2[5].wave_shpr.div.quo[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13245_ (.CLK(clknet_leaf_11_clk),
    .D(net325),
    .RESET_B(net54),
    .Q(\genblk2[5].wave_shpr.div.acc_next[0] ));
 sky130_fd_sc_hd__dfrtp_2 _13246_ (.CLK(clknet_leaf_11_clk),
    .D(net494),
    .RESET_B(net56),
    .Q(\genblk2[5].wave_shpr.div.acc[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13247_ (.CLK(clknet_leaf_2_clk),
    .D(_00570_),
    .RESET_B(net52),
    .Q(\genblk2[5].wave_shpr.div.acc[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13248_ (.CLK(clknet_leaf_13_clk),
    .D(net911),
    .RESET_B(net52),
    .Q(\genblk2[5].wave_shpr.div.acc[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13249_ (.CLK(clknet_leaf_2_clk),
    .D(_00572_),
    .RESET_B(net52),
    .Q(\genblk2[5].wave_shpr.div.acc[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13250_ (.CLK(clknet_leaf_2_clk),
    .D(_00573_),
    .RESET_B(net43),
    .Q(\genblk2[5].wave_shpr.div.acc[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13251_ (.CLK(clknet_leaf_2_clk),
    .D(_00574_),
    .RESET_B(net41),
    .Q(\genblk2[5].wave_shpr.div.acc[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13252_ (.CLK(clknet_leaf_1_clk),
    .D(_00575_),
    .RESET_B(net41),
    .Q(\genblk2[5].wave_shpr.div.acc[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13253_ (.CLK(clknet_leaf_1_clk),
    .D(_00576_),
    .RESET_B(net41),
    .Q(\genblk2[5].wave_shpr.div.acc[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13254_ (.CLK(clknet_leaf_2_clk),
    .D(_00577_),
    .RESET_B(net43),
    .Q(\genblk2[5].wave_shpr.div.acc[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13255_ (.CLK(clknet_leaf_2_clk),
    .D(_00578_),
    .RESET_B(net51),
    .Q(\genblk2[5].wave_shpr.div.acc[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13256_ (.CLK(clknet_leaf_3_clk),
    .D(net773),
    .RESET_B(net51),
    .Q(\genblk2[5].wave_shpr.div.acc[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13257_ (.CLK(clknet_leaf_3_clk),
    .D(_00580_),
    .RESET_B(net46),
    .Q(\genblk2[5].wave_shpr.div.acc[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13258_ (.CLK(clknet_leaf_2_clk),
    .D(_00581_),
    .RESET_B(net51),
    .Q(\genblk2[5].wave_shpr.div.acc[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13259_ (.CLK(clknet_leaf_2_clk),
    .D(_00582_),
    .RESET_B(net43),
    .Q(\genblk2[5].wave_shpr.div.acc[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13260_ (.CLK(clknet_leaf_0_clk),
    .D(_00583_),
    .RESET_B(net38),
    .Q(\genblk2[5].wave_shpr.div.acc[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13261_ (.CLK(clknet_leaf_0_clk),
    .D(_00584_),
    .RESET_B(net38),
    .Q(\genblk2[5].wave_shpr.div.acc[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13262_ (.CLK(clknet_leaf_0_clk),
    .D(_00585_),
    .RESET_B(net38),
    .Q(\genblk2[5].wave_shpr.div.acc[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13263_ (.CLK(clknet_leaf_0_clk),
    .D(_00586_),
    .RESET_B(net38),
    .Q(\genblk2[5].wave_shpr.div.acc[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13264_ (.CLK(clknet_leaf_1_clk),
    .D(_00587_),
    .RESET_B(net38),
    .Q(\genblk2[5].wave_shpr.div.acc[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13265_ (.CLK(clknet_leaf_0_clk),
    .D(_00588_),
    .RESET_B(net38),
    .Q(\genblk2[5].wave_shpr.div.acc[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13266_ (.CLK(clknet_leaf_0_clk),
    .D(_00589_),
    .RESET_B(net38),
    .Q(\genblk2[5].wave_shpr.div.acc[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13267_ (.CLK(clknet_leaf_1_clk),
    .D(_00590_),
    .RESET_B(net38),
    .Q(\genblk2[5].wave_shpr.div.acc[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13268_ (.CLK(clknet_leaf_1_clk),
    .D(_00591_),
    .RESET_B(net44),
    .Q(\genblk2[5].wave_shpr.div.acc[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13269_ (.CLK(clknet_leaf_1_clk),
    .D(_00592_),
    .RESET_B(net41),
    .Q(\genblk2[5].wave_shpr.div.acc[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13270_ (.CLK(clknet_leaf_1_clk),
    .D(_00593_),
    .RESET_B(net43),
    .Q(\genblk2[5].wave_shpr.div.acc[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13271_ (.CLK(clknet_leaf_137_clk),
    .D(_00594_),
    .RESET_B(net41),
    .Q(\genblk2[5].wave_shpr.div.acc[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13272_ (.CLK(clknet_leaf_136_clk),
    .D(_00595_),
    .RESET_B(net41),
    .Q(\genblk2[5].wave_shpr.div.acc[26] ));
 sky130_fd_sc_hd__dfrtp_1 _13273_ (.CLK(clknet_leaf_12_clk),
    .D(_00016_),
    .RESET_B(net51),
    .Q(\genblk2[6].wave_shpr.div.busy ));
 sky130_fd_sc_hd__dfrtp_1 _13274_ (.CLK(clknet_leaf_118_clk),
    .D(_00017_),
    .RESET_B(net138),
    .Q(\genblk2[6].wave_shpr.div.done ));
 sky130_fd_sc_hd__dfrtp_4 _13275_ (.CLK(clknet_leaf_12_clk),
    .D(_00596_),
    .RESET_B(net54),
    .Q(\genblk2[5].wave_shpr.div.i[0] ));
 sky130_fd_sc_hd__dfrtp_2 _13276_ (.CLK(clknet_leaf_12_clk),
    .D(_00597_),
    .RESET_B(net54),
    .Q(\genblk2[5].wave_shpr.div.i[1] ));
 sky130_fd_sc_hd__dfrtp_2 _13277_ (.CLK(clknet_leaf_12_clk),
    .D(_00598_),
    .RESET_B(net54),
    .Q(\genblk2[5].wave_shpr.div.i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13278_ (.CLK(clknet_leaf_11_clk),
    .D(_00599_),
    .RESET_B(net56),
    .Q(\genblk2[5].wave_shpr.div.i[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13279_ (.CLK(clknet_leaf_11_clk),
    .D(_00600_),
    .RESET_B(net56),
    .Q(\genblk2[5].wave_shpr.div.i[4] ));
 sky130_fd_sc_hd__dfrtp_4 _13280_ (.CLK(clknet_leaf_122_clk),
    .D(_00601_),
    .RESET_B(net79),
    .Q(\genblk2[6].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__dfrtp_2 _13281_ (.CLK(clknet_leaf_122_clk),
    .D(_00602_),
    .RESET_B(net79),
    .Q(\genblk2[6].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__dfrtp_2 _13282_ (.CLK(clknet_leaf_117_clk),
    .D(_00603_),
    .RESET_B(net137),
    .Q(\genblk2[6].wave_shpr.div.fin_quo[2] ));
 sky130_fd_sc_hd__dfrtp_2 _13283_ (.CLK(clknet_leaf_117_clk),
    .D(_00604_),
    .RESET_B(net137),
    .Q(\genblk2[6].wave_shpr.div.fin_quo[3] ));
 sky130_fd_sc_hd__dfrtp_2 _13284_ (.CLK(clknet_leaf_117_clk),
    .D(_00605_),
    .RESET_B(net137),
    .Q(\genblk2[6].wave_shpr.div.fin_quo[4] ));
 sky130_fd_sc_hd__dfrtp_2 _13285_ (.CLK(clknet_leaf_117_clk),
    .D(_00606_),
    .RESET_B(net137),
    .Q(\genblk2[6].wave_shpr.div.fin_quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13286_ (.CLK(clknet_leaf_118_clk),
    .D(_00607_),
    .RESET_B(net137),
    .Q(\genblk2[6].wave_shpr.div.fin_quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13287_ (.CLK(clknet_leaf_118_clk),
    .D(_00608_),
    .RESET_B(net138),
    .Q(\genblk2[6].wave_shpr.div.fin_quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13288_ (.CLK(clknet_leaf_90_clk),
    .D(_00609_),
    .RESET_B(net147),
    .Q(\genblk2[7].wave_shpr.div.b1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13289_ (.CLK(clknet_leaf_92_clk),
    .D(_00610_),
    .RESET_B(net147),
    .Q(\genblk2[7].wave_shpr.div.b1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13290_ (.CLK(clknet_leaf_88_clk),
    .D(_00611_),
    .RESET_B(net177),
    .Q(\genblk2[7].wave_shpr.div.b1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13291_ (.CLK(clknet_leaf_88_clk),
    .D(_00612_),
    .RESET_B(net177),
    .Q(\genblk2[7].wave_shpr.div.b1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13292_ (.CLK(clknet_leaf_88_clk),
    .D(_00613_),
    .RESET_B(net177),
    .Q(\genblk2[7].wave_shpr.div.b1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13293_ (.CLK(clknet_leaf_87_clk),
    .D(_00614_),
    .RESET_B(net179),
    .Q(\genblk2[7].wave_shpr.div.b1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13294_ (.CLK(clknet_leaf_87_clk),
    .D(_00615_),
    .RESET_B(net179),
    .Q(\genblk2[7].wave_shpr.div.b1[6] ));
 sky130_fd_sc_hd__dfrtp_2 _13295_ (.CLK(clknet_leaf_53_clk),
    .D(_00616_),
    .RESET_B(net112),
    .Q(\genblk2[7].wave_shpr.div.b1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13296_ (.CLK(clknet_leaf_87_clk),
    .D(_00617_),
    .RESET_B(net179),
    .Q(\genblk2[7].wave_shpr.div.b1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13297_ (.CLK(clknet_leaf_86_clk),
    .D(_00618_),
    .RESET_B(net179),
    .Q(\genblk2[7].wave_shpr.div.b1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13298_ (.CLK(clknet_leaf_84_clk),
    .D(_00619_),
    .RESET_B(net202),
    .Q(\genblk2[7].wave_shpr.div.b1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13299_ (.CLK(clknet_leaf_84_clk),
    .D(_00620_),
    .RESET_B(net202),
    .Q(\genblk2[7].wave_shpr.div.b1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13300_ (.CLK(clknet_leaf_83_clk),
    .D(_00621_),
    .RESET_B(net199),
    .Q(\genblk2[7].wave_shpr.div.b1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13301_ (.CLK(clknet_leaf_84_clk),
    .D(_00622_),
    .RESET_B(net202),
    .Q(\genblk2[7].wave_shpr.div.b1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13302_ (.CLK(clknet_leaf_87_clk),
    .D(_00623_),
    .RESET_B(net179),
    .Q(\genblk2[7].wave_shpr.div.b1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13303_ (.CLK(clknet_leaf_87_clk),
    .D(_00624_),
    .RESET_B(net201),
    .Q(\genblk2[7].wave_shpr.div.b1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13304_ (.CLK(clknet_leaf_96_clk),
    .D(_00625_),
    .RESET_B(net161),
    .Q(\genblk2[7].wave_shpr.div.b1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13305_ (.CLK(clknet_leaf_96_clk),
    .D(_00626_),
    .RESET_B(net161),
    .Q(\genblk2[7].wave_shpr.div.b1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13306_ (.CLK(clknet_leaf_3_clk),
    .D(_00627_),
    .RESET_B(net51),
    .Q(\genblk2[6].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13307_ (.CLK(clknet_leaf_122_clk),
    .D(_00628_),
    .RESET_B(net137),
    .Q(\genblk2[6].wave_shpr.div.quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13308_ (.CLK(clknet_leaf_117_clk),
    .D(_00629_),
    .RESET_B(net137),
    .Q(\genblk2[6].wave_shpr.div.quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13309_ (.CLK(clknet_leaf_117_clk),
    .D(_00630_),
    .RESET_B(net137),
    .Q(\genblk2[6].wave_shpr.div.quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13310_ (.CLK(clknet_leaf_118_clk),
    .D(net272),
    .RESET_B(net137),
    .Q(\genblk2[6].wave_shpr.div.quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13311_ (.CLK(clknet_leaf_118_clk),
    .D(net721),
    .RESET_B(net137),
    .Q(\genblk2[6].wave_shpr.div.quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13312_ (.CLK(clknet_leaf_118_clk),
    .D(_00633_),
    .RESET_B(net138),
    .Q(\genblk2[6].wave_shpr.div.quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13313_ (.CLK(clknet_leaf_121_clk),
    .D(net242),
    .RESET_B(net78),
    .Q(\genblk2[6].wave_shpr.div.quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13314_ (.CLK(clknet_leaf_12_clk),
    .D(_00635_),
    .RESET_B(net54),
    .Q(\genblk2[6].wave_shpr.div.quo[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13315_ (.CLK(clknet_leaf_9_clk),
    .D(net516),
    .RESET_B(net48),
    .Q(\genblk2[6].wave_shpr.div.quo[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13316_ (.CLK(clknet_leaf_9_clk),
    .D(_00637_),
    .RESET_B(net50),
    .Q(\genblk2[6].wave_shpr.div.quo[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13317_ (.CLK(clknet_leaf_24_clk),
    .D(net345),
    .RESET_B(net88),
    .Q(\genblk2[6].wave_shpr.div.quo[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13318_ (.CLK(clknet_leaf_25_clk),
    .D(net624),
    .RESET_B(net86),
    .Q(\genblk2[6].wave_shpr.div.quo[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13319_ (.CLK(clknet_leaf_26_clk),
    .D(net621),
    .RESET_B(net87),
    .Q(\genblk2[6].wave_shpr.div.quo[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13320_ (.CLK(clknet_leaf_26_clk),
    .D(net499),
    .RESET_B(net87),
    .Q(\genblk2[6].wave_shpr.div.quo[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13321_ (.CLK(clknet_leaf_26_clk),
    .D(_00642_),
    .RESET_B(net87),
    .Q(\genblk2[6].wave_shpr.div.quo[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13322_ (.CLK(clknet_leaf_26_clk),
    .D(_00643_),
    .RESET_B(net87),
    .Q(\genblk2[6].wave_shpr.div.quo[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13323_ (.CLK(clknet_leaf_26_clk),
    .D(_00644_),
    .RESET_B(net87),
    .Q(\genblk2[6].wave_shpr.div.quo[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13324_ (.CLK(clknet_leaf_26_clk),
    .D(_00645_),
    .RESET_B(net87),
    .Q(\genblk2[6].wave_shpr.div.quo[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13325_ (.CLK(clknet_leaf_26_clk),
    .D(_00646_),
    .RESET_B(net87),
    .Q(\genblk2[6].wave_shpr.div.quo[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13326_ (.CLK(clknet_leaf_25_clk),
    .D(net314),
    .RESET_B(net86),
    .Q(\genblk2[6].wave_shpr.div.quo[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13327_ (.CLK(clknet_leaf_25_clk),
    .D(net568),
    .RESET_B(net86),
    .Q(\genblk2[6].wave_shpr.div.quo[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13328_ (.CLK(clknet_leaf_25_clk),
    .D(_00649_),
    .RESET_B(net86),
    .Q(\genblk2[6].wave_shpr.div.quo[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13329_ (.CLK(clknet_leaf_25_clk),
    .D(_00650_),
    .RESET_B(net91),
    .Q(\genblk2[6].wave_shpr.div.quo[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13330_ (.CLK(clknet_leaf_24_clk),
    .D(net386),
    .RESET_B(net91),
    .Q(\genblk2[6].wave_shpr.div.quo[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13331_ (.CLK(clknet_leaf_24_clk),
    .D(_00652_),
    .RESET_B(net92),
    .Q(\genblk2[6].wave_shpr.div.acc_next[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13332_ (.CLK(clknet_leaf_9_clk),
    .D(net284),
    .RESET_B(net54),
    .Q(\genblk2[6].wave_shpr.div.acc[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13333_ (.CLK(clknet_leaf_9_clk),
    .D(_00654_),
    .RESET_B(net54),
    .Q(\genblk2[6].wave_shpr.div.acc[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13334_ (.CLK(clknet_leaf_6_clk),
    .D(_00655_),
    .RESET_B(net48),
    .Q(\genblk2[6].wave_shpr.div.acc[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13335_ (.CLK(clknet_leaf_6_clk),
    .D(_00656_),
    .RESET_B(net48),
    .Q(\genblk2[6].wave_shpr.div.acc[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13336_ (.CLK(clknet_leaf_6_clk),
    .D(_00657_),
    .RESET_B(net48),
    .Q(\genblk2[6].wave_shpr.div.acc[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13337_ (.CLK(clknet_leaf_8_clk),
    .D(_00658_),
    .RESET_B(net49),
    .Q(\genblk2[6].wave_shpr.div.acc[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13338_ (.CLK(clknet_leaf_8_clk),
    .D(_00659_),
    .RESET_B(net50),
    .Q(\genblk2[6].wave_shpr.div.acc[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13339_ (.CLK(clknet_leaf_7_clk),
    .D(_00660_),
    .RESET_B(net49),
    .Q(\genblk2[6].wave_shpr.div.acc[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13340_ (.CLK(clknet_leaf_7_clk),
    .D(_00661_),
    .RESET_B(net49),
    .Q(\genblk2[6].wave_shpr.div.acc[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13341_ (.CLK(clknet_leaf_7_clk),
    .D(_00662_),
    .RESET_B(net49),
    .Q(\genblk2[6].wave_shpr.div.acc[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13342_ (.CLK(clknet_leaf_7_clk),
    .D(_00663_),
    .RESET_B(net49),
    .Q(\genblk2[6].wave_shpr.div.acc[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13343_ (.CLK(clknet_leaf_7_clk),
    .D(_00664_),
    .RESET_B(net49),
    .Q(\genblk2[6].wave_shpr.div.acc[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13344_ (.CLK(clknet_leaf_7_clk),
    .D(_00665_),
    .RESET_B(net49),
    .Q(\genblk2[6].wave_shpr.div.acc[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13345_ (.CLK(clknet_leaf_6_clk),
    .D(_00666_),
    .RESET_B(net49),
    .Q(\genblk2[6].wave_shpr.div.acc[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13346_ (.CLK(clknet_leaf_6_clk),
    .D(_00667_),
    .RESET_B(net49),
    .Q(\genblk2[6].wave_shpr.div.acc[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13347_ (.CLK(clknet_leaf_5_clk),
    .D(_00668_),
    .RESET_B(net45),
    .Q(\genblk2[6].wave_shpr.div.acc[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13348_ (.CLK(clknet_leaf_5_clk),
    .D(_00669_),
    .RESET_B(net45),
    .Q(\genblk2[6].wave_shpr.div.acc[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13349_ (.CLK(clknet_leaf_4_clk),
    .D(_00670_),
    .RESET_B(net45),
    .Q(\genblk2[6].wave_shpr.div.acc[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13350_ (.CLK(clknet_leaf_5_clk),
    .D(_00671_),
    .RESET_B(net45),
    .Q(\genblk2[6].wave_shpr.div.acc[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13351_ (.CLK(clknet_leaf_5_clk),
    .D(_00672_),
    .RESET_B(net47),
    .Q(\genblk2[6].wave_shpr.div.acc[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13352_ (.CLK(clknet_leaf_4_clk),
    .D(_00673_),
    .RESET_B(net45),
    .Q(\genblk2[6].wave_shpr.div.acc[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13353_ (.CLK(clknet_leaf_4_clk),
    .D(_00674_),
    .RESET_B(net45),
    .Q(\genblk2[6].wave_shpr.div.acc[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13354_ (.CLK(clknet_leaf_4_clk),
    .D(_00675_),
    .RESET_B(net45),
    .Q(\genblk2[6].wave_shpr.div.acc[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13355_ (.CLK(clknet_leaf_4_clk),
    .D(_00676_),
    .RESET_B(net45),
    .Q(\genblk2[6].wave_shpr.div.acc[23] ));
 sky130_fd_sc_hd__dfrtp_2 _13356_ (.CLK(clknet_leaf_4_clk),
    .D(_00677_),
    .RESET_B(net45),
    .Q(\genblk2[6].wave_shpr.div.acc[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13357_ (.CLK(clknet_leaf_4_clk),
    .D(_00678_),
    .RESET_B(net45),
    .Q(\genblk2[6].wave_shpr.div.acc[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13358_ (.CLK(clknet_leaf_4_clk),
    .D(_00679_),
    .RESET_B(net46),
    .Q(\genblk2[6].wave_shpr.div.acc[26] ));
 sky130_fd_sc_hd__dfrtp_1 _13359_ (.CLK(clknet_leaf_91_clk),
    .D(_00018_),
    .RESET_B(net143),
    .Q(\genblk2[7].wave_shpr.div.busy ));
 sky130_fd_sc_hd__dfrtp_1 _13360_ (.CLK(clknet_leaf_116_clk),
    .D(_00019_),
    .RESET_B(net139),
    .Q(\genblk2[7].wave_shpr.div.done ));
 sky130_fd_sc_hd__dfrtp_2 _13361_ (.CLK(clknet_leaf_6_clk),
    .D(_00680_),
    .RESET_B(net47),
    .Q(\genblk2[6].wave_shpr.div.i[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13362_ (.CLK(clknet_leaf_6_clk),
    .D(_00681_),
    .RESET_B(net47),
    .Q(\genblk2[6].wave_shpr.div.i[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13363_ (.CLK(clknet_leaf_3_clk),
    .D(_00682_),
    .RESET_B(net53),
    .Q(\genblk2[6].wave_shpr.div.i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13364_ (.CLK(clknet_leaf_12_clk),
    .D(_00683_),
    .RESET_B(net53),
    .Q(\genblk2[6].wave_shpr.div.i[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13365_ (.CLK(clknet_leaf_12_clk),
    .D(_00684_),
    .RESET_B(net53),
    .Q(\genblk2[6].wave_shpr.div.i[4] ));
 sky130_fd_sc_hd__dfrtp_2 _13366_ (.CLK(clknet_leaf_91_clk),
    .D(_00685_),
    .RESET_B(net143),
    .Q(\genblk2[7].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__dfrtp_2 _13367_ (.CLK(clknet_leaf_116_clk),
    .D(_00686_),
    .RESET_B(net139),
    .Q(\genblk2[7].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13368_ (.CLK(clknet_leaf_116_clk),
    .D(_00687_),
    .RESET_B(net139),
    .Q(\genblk2[7].wave_shpr.div.fin_quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13369_ (.CLK(clknet_leaf_116_clk),
    .D(_00688_),
    .RESET_B(net140),
    .Q(\genblk2[7].wave_shpr.div.fin_quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13370_ (.CLK(clknet_leaf_116_clk),
    .D(_00689_),
    .RESET_B(net140),
    .Q(\genblk2[7].wave_shpr.div.fin_quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13371_ (.CLK(clknet_leaf_117_clk),
    .D(_00690_),
    .RESET_B(net140),
    .Q(\genblk2[7].wave_shpr.div.fin_quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13372_ (.CLK(clknet_leaf_115_clk),
    .D(_00691_),
    .RESET_B(net140),
    .Q(\genblk2[7].wave_shpr.div.fin_quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13373_ (.CLK(clknet_leaf_117_clk),
    .D(_00692_),
    .RESET_B(net140),
    .Q(\genblk2[7].wave_shpr.div.fin_quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13374_ (.CLK(clknet_leaf_96_clk),
    .D(_00693_),
    .RESET_B(net167),
    .Q(\genblk2[8].wave_shpr.div.b1[0] ));
 sky130_fd_sc_hd__dfrtp_2 _13375_ (.CLK(clknet_leaf_86_clk),
    .D(_00694_),
    .RESET_B(net179),
    .Q(\genblk2[8].wave_shpr.div.b1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13376_ (.CLK(clknet_leaf_96_clk),
    .D(_00695_),
    .RESET_B(net167),
    .Q(\genblk2[8].wave_shpr.div.b1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13377_ (.CLK(clknet_leaf_81_clk),
    .D(_00696_),
    .RESET_B(net199),
    .Q(\genblk2[8].wave_shpr.div.b1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13378_ (.CLK(clknet_leaf_81_clk),
    .D(_00697_),
    .RESET_B(net205),
    .Q(\genblk2[8].wave_shpr.div.b1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13379_ (.CLK(clknet_leaf_81_clk),
    .D(_00698_),
    .RESET_B(net199),
    .Q(\genblk2[8].wave_shpr.div.b1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13380_ (.CLK(clknet_leaf_80_clk),
    .D(_00699_),
    .RESET_B(net200),
    .Q(\genblk2[8].wave_shpr.div.b1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13381_ (.CLK(clknet_leaf_96_clk),
    .D(_00700_),
    .RESET_B(net167),
    .Q(\genblk2[8].wave_shpr.div.b1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13382_ (.CLK(clknet_leaf_83_clk),
    .D(_00701_),
    .RESET_B(net200),
    .Q(\genblk2[8].wave_shpr.div.b1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13383_ (.CLK(clknet_leaf_83_clk),
    .D(_00702_),
    .RESET_B(net200),
    .Q(\genblk2[8].wave_shpr.div.b1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13384_ (.CLK(clknet_leaf_83_clk),
    .D(_00703_),
    .RESET_B(net200),
    .Q(\genblk2[8].wave_shpr.div.b1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13385_ (.CLK(clknet_leaf_83_clk),
    .D(_00704_),
    .RESET_B(net200),
    .Q(\genblk2[8].wave_shpr.div.b1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13386_ (.CLK(clknet_leaf_86_clk),
    .D(_00705_),
    .RESET_B(net183),
    .Q(\genblk2[8].wave_shpr.div.b1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13387_ (.CLK(clknet_leaf_83_clk),
    .D(_00706_),
    .RESET_B(net200),
    .Q(\genblk2[8].wave_shpr.div.b1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13388_ (.CLK(clknet_leaf_78_clk),
    .D(_00707_),
    .RESET_B(net208),
    .Q(\genblk2[8].wave_shpr.div.b1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13389_ (.CLK(clknet_leaf_78_clk),
    .D(_00708_),
    .RESET_B(net205),
    .Q(\genblk2[8].wave_shpr.div.b1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13390_ (.CLK(clknet_leaf_79_clk),
    .D(_00709_),
    .RESET_B(net205),
    .Q(\genblk2[8].wave_shpr.div.b1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13391_ (.CLK(clknet_leaf_79_clk),
    .D(_00710_),
    .RESET_B(net206),
    .Q(\genblk2[8].wave_shpr.div.b1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13392_ (.CLK(clknet_leaf_91_clk),
    .D(_00711_),
    .RESET_B(net143),
    .Q(\genblk2[7].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13393_ (.CLK(clknet_leaf_118_clk),
    .D(_00712_),
    .RESET_B(net139),
    .Q(\genblk2[7].wave_shpr.div.quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13394_ (.CLK(clknet_leaf_116_clk),
    .D(net564),
    .RESET_B(net145),
    .Q(\genblk2[7].wave_shpr.div.quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13395_ (.CLK(clknet_leaf_116_clk),
    .D(_00714_),
    .RESET_B(net140),
    .Q(\genblk2[7].wave_shpr.div.quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13396_ (.CLK(clknet_leaf_117_clk),
    .D(net332),
    .RESET_B(net140),
    .Q(\genblk2[7].wave_shpr.div.quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13397_ (.CLK(clknet_leaf_117_clk),
    .D(net662),
    .RESET_B(net140),
    .Q(\genblk2[7].wave_shpr.div.quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13398_ (.CLK(clknet_leaf_117_clk),
    .D(_00717_),
    .RESET_B(net140),
    .Q(\genblk2[7].wave_shpr.div.quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13399_ (.CLK(clknet_leaf_119_clk),
    .D(net318),
    .RESET_B(net139),
    .Q(\genblk2[7].wave_shpr.div.quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13400_ (.CLK(clknet_leaf_119_clk),
    .D(net422),
    .RESET_B(net143),
    .Q(\genblk2[7].wave_shpr.div.quo[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13401_ (.CLK(clknet_leaf_92_clk),
    .D(_00720_),
    .RESET_B(net143),
    .Q(\genblk2[7].wave_shpr.div.quo[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13402_ (.CLK(clknet_leaf_90_clk),
    .D(net303),
    .RESET_B(net147),
    .Q(\genblk2[7].wave_shpr.div.quo[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13403_ (.CLK(clknet_leaf_92_clk),
    .D(_00722_),
    .RESET_B(net147),
    .Q(\genblk2[7].wave_shpr.div.quo[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13404_ (.CLK(clknet_leaf_90_clk),
    .D(net371),
    .RESET_B(net143),
    .Q(\genblk2[7].wave_shpr.div.quo[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13405_ (.CLK(clknet_leaf_90_clk),
    .D(_00724_),
    .RESET_B(net143),
    .Q(\genblk2[7].wave_shpr.div.quo[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13406_ (.CLK(clknet_leaf_90_clk),
    .D(_00725_),
    .RESET_B(net144),
    .Q(\genblk2[7].wave_shpr.div.quo[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13407_ (.CLK(clknet_leaf_90_clk),
    .D(_00726_),
    .RESET_B(net144),
    .Q(\genblk2[7].wave_shpr.div.quo[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13408_ (.CLK(clknet_leaf_90_clk),
    .D(_00727_),
    .RESET_B(net142),
    .Q(\genblk2[7].wave_shpr.div.quo[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13409_ (.CLK(clknet_leaf_90_clk),
    .D(net549),
    .RESET_B(net144),
    .Q(\genblk2[7].wave_shpr.div.quo[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13410_ (.CLK(clknet_leaf_90_clk),
    .D(_00729_),
    .RESET_B(net144),
    .Q(\genblk2[7].wave_shpr.div.quo[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13411_ (.CLK(clknet_leaf_91_clk),
    .D(_00730_),
    .RESET_B(net144),
    .Q(\genblk2[7].wave_shpr.div.quo[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13412_ (.CLK(clknet_leaf_120_clk),
    .D(net232),
    .RESET_B(net142),
    .Q(\genblk2[7].wave_shpr.div.quo[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13413_ (.CLK(clknet_leaf_120_clk),
    .D(net528),
    .RESET_B(net142),
    .Q(\genblk2[7].wave_shpr.div.quo[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13414_ (.CLK(clknet_leaf_120_clk),
    .D(_00733_),
    .RESET_B(net141),
    .Q(\genblk2[7].wave_shpr.div.quo[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13415_ (.CLK(clknet_leaf_120_clk),
    .D(net488),
    .RESET_B(net141),
    .Q(\genblk2[7].wave_shpr.div.quo[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13416_ (.CLK(clknet_leaf_119_clk),
    .D(net535),
    .RESET_B(net141),
    .Q(\genblk2[7].wave_shpr.div.quo[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13417_ (.CLK(clknet_leaf_119_clk),
    .D(_00736_),
    .RESET_B(net141),
    .Q(\genblk2[7].wave_shpr.div.acc_next[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13418_ (.CLK(clknet_leaf_119_clk),
    .D(_00737_),
    .RESET_B(net141),
    .Q(\genblk2[7].wave_shpr.div.acc[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13419_ (.CLK(clknet_leaf_91_clk),
    .D(_00738_),
    .RESET_B(net147),
    .Q(\genblk2[7].wave_shpr.div.acc[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13420_ (.CLK(clknet_leaf_91_clk),
    .D(_00739_),
    .RESET_B(net147),
    .Q(\genblk2[7].wave_shpr.div.acc[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13421_ (.CLK(clknet_leaf_92_clk),
    .D(_00740_),
    .RESET_B(net147),
    .Q(\genblk2[7].wave_shpr.div.acc[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13422_ (.CLK(clknet_leaf_92_clk),
    .D(_00741_),
    .RESET_B(net149),
    .Q(\genblk2[7].wave_shpr.div.acc[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13423_ (.CLK(clknet_leaf_87_clk),
    .D(_00742_),
    .RESET_B(net179),
    .Q(\genblk2[7].wave_shpr.div.acc[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13424_ (.CLK(clknet_leaf_87_clk),
    .D(_00743_),
    .RESET_B(net179),
    .Q(\genblk2[7].wave_shpr.div.acc[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13425_ (.CLK(clknet_leaf_87_clk),
    .D(_00744_),
    .RESET_B(net201),
    .Q(\genblk2[7].wave_shpr.div.acc[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13426_ (.CLK(clknet_leaf_82_clk),
    .D(_00745_),
    .RESET_B(net201),
    .Q(\genblk2[7].wave_shpr.div.acc[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13427_ (.CLK(clknet_leaf_87_clk),
    .D(_00746_),
    .RESET_B(net201),
    .Q(\genblk2[7].wave_shpr.div.acc[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13428_ (.CLK(clknet_leaf_82_clk),
    .D(net798),
    .RESET_B(net201),
    .Q(\genblk2[7].wave_shpr.div.acc[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13429_ (.CLK(clknet_leaf_83_clk),
    .D(_00748_),
    .RESET_B(net201),
    .Q(\genblk2[7].wave_shpr.div.acc[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13430_ (.CLK(clknet_leaf_82_clk),
    .D(net853),
    .RESET_B(net201),
    .Q(\genblk2[7].wave_shpr.div.acc[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13431_ (.CLK(clknet_leaf_82_clk),
    .D(_00750_),
    .RESET_B(net201),
    .Q(\genblk2[7].wave_shpr.div.acc[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13432_ (.CLK(clknet_leaf_82_clk),
    .D(_00751_),
    .RESET_B(net201),
    .Q(\genblk2[7].wave_shpr.div.acc[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13433_ (.CLK(clknet_leaf_82_clk),
    .D(_00752_),
    .RESET_B(net201),
    .Q(\genblk2[7].wave_shpr.div.acc[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13434_ (.CLK(clknet_leaf_81_clk),
    .D(net1011),
    .RESET_B(net199),
    .Q(\genblk2[7].wave_shpr.div.acc[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13435_ (.CLK(clknet_leaf_95_clk),
    .D(_00754_),
    .RESET_B(net161),
    .Q(\genblk2[7].wave_shpr.div.acc[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13436_ (.CLK(clknet_leaf_95_clk),
    .D(_00755_),
    .RESET_B(net159),
    .Q(\genblk2[7].wave_shpr.div.acc[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13437_ (.CLK(clknet_leaf_95_clk),
    .D(_00756_),
    .RESET_B(net161),
    .Q(\genblk2[7].wave_shpr.div.acc[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13438_ (.CLK(clknet_leaf_95_clk),
    .D(_00757_),
    .RESET_B(net159),
    .Q(\genblk2[7].wave_shpr.div.acc[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13439_ (.CLK(clknet_leaf_94_clk),
    .D(_00758_),
    .RESET_B(net162),
    .Q(\genblk2[7].wave_shpr.div.acc[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13440_ (.CLK(clknet_leaf_95_clk),
    .D(_00759_),
    .RESET_B(net162),
    .Q(\genblk2[7].wave_shpr.div.acc[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13441_ (.CLK(clknet_leaf_95_clk),
    .D(_00760_),
    .RESET_B(net162),
    .Q(\genblk2[7].wave_shpr.div.acc[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13442_ (.CLK(clknet_leaf_92_clk),
    .D(_00761_),
    .RESET_B(net149),
    .Q(\genblk2[7].wave_shpr.div.acc[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13443_ (.CLK(clknet_leaf_92_clk),
    .D(_00762_),
    .RESET_B(net149),
    .Q(\genblk2[7].wave_shpr.div.acc[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13444_ (.CLK(clknet_leaf_95_clk),
    .D(net382),
    .RESET_B(net149),
    .Q(\genblk2[7].wave_shpr.div.acc[26] ));
 sky130_fd_sc_hd__dfrtp_1 _13445_ (.CLK(clknet_leaf_81_clk),
    .D(_00020_),
    .RESET_B(net199),
    .Q(\genblk2[8].wave_shpr.div.busy ));
 sky130_fd_sc_hd__dfrtp_1 _13446_ (.CLK(clknet_leaf_99_clk),
    .D(_00021_),
    .RESET_B(net166),
    .Q(\genblk2[8].wave_shpr.div.done ));
 sky130_fd_sc_hd__dfrtp_2 _13447_ (.CLK(clknet_leaf_90_clk),
    .D(_00764_),
    .RESET_B(net144),
    .Q(\genblk2[7].wave_shpr.div.i[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13448_ (.CLK(clknet_leaf_91_clk),
    .D(_00765_),
    .RESET_B(net147),
    .Q(\genblk2[7].wave_shpr.div.i[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13449_ (.CLK(clknet_leaf_91_clk),
    .D(_00766_),
    .RESET_B(net144),
    .Q(\genblk2[7].wave_shpr.div.i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13450_ (.CLK(clknet_leaf_119_clk),
    .D(_00767_),
    .RESET_B(net143),
    .Q(\genblk2[7].wave_shpr.div.i[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13451_ (.CLK(clknet_leaf_119_clk),
    .D(_00768_),
    .RESET_B(net143),
    .Q(\genblk2[7].wave_shpr.div.i[4] ));
 sky130_fd_sc_hd__dfrtp_4 _13452_ (.CLK(clknet_leaf_99_clk),
    .D(_00769_),
    .RESET_B(net166),
    .Q(\genblk2[8].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__dfrtp_4 _13453_ (.CLK(clknet_leaf_99_clk),
    .D(_00770_),
    .RESET_B(net168),
    .Q(\genblk2[8].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__dfrtp_4 _13454_ (.CLK(clknet_leaf_99_clk),
    .D(_00771_),
    .RESET_B(net164),
    .Q(\genblk2[8].wave_shpr.div.fin_quo[2] ));
 sky130_fd_sc_hd__dfrtp_2 _13455_ (.CLK(clknet_leaf_99_clk),
    .D(_00772_),
    .RESET_B(net168),
    .Q(\genblk2[8].wave_shpr.div.fin_quo[3] ));
 sky130_fd_sc_hd__dfrtp_2 _13456_ (.CLK(clknet_leaf_100_clk),
    .D(_00773_),
    .RESET_B(net164),
    .Q(\genblk2[8].wave_shpr.div.fin_quo[4] ));
 sky130_fd_sc_hd__dfrtp_4 _13457_ (.CLK(clknet_leaf_99_clk),
    .D(_00774_),
    .RESET_B(net165),
    .Q(\genblk2[8].wave_shpr.div.fin_quo[5] ));
 sky130_fd_sc_hd__dfrtp_2 _13458_ (.CLK(clknet_leaf_99_clk),
    .D(_00775_),
    .RESET_B(net165),
    .Q(\genblk2[8].wave_shpr.div.fin_quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13459_ (.CLK(clknet_leaf_99_clk),
    .D(_00776_),
    .RESET_B(net166),
    .Q(\genblk2[8].wave_shpr.div.fin_quo[7] ));
 sky130_fd_sc_hd__dfrtp_2 _13460_ (.CLK(clknet_leaf_84_clk),
    .D(_00777_),
    .RESET_B(net203),
    .Q(\genblk2[9].wave_shpr.div.b1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13461_ (.CLK(clknet_leaf_84_clk),
    .D(_00778_),
    .RESET_B(net203),
    .Q(\genblk2[9].wave_shpr.div.b1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13462_ (.CLK(clknet_leaf_83_clk),
    .D(_00779_),
    .RESET_B(net203),
    .Q(\genblk2[9].wave_shpr.div.b1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13463_ (.CLK(clknet_leaf_83_clk),
    .D(_00780_),
    .RESET_B(net203),
    .Q(\genblk2[9].wave_shpr.div.b1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13464_ (.CLK(clknet_leaf_83_clk),
    .D(_00781_),
    .RESET_B(net203),
    .Q(\genblk2[9].wave_shpr.div.b1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13465_ (.CLK(clknet_leaf_75_clk),
    .D(_00782_),
    .RESET_B(net203),
    .Q(\genblk2[9].wave_shpr.div.b1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13466_ (.CLK(clknet_leaf_75_clk),
    .D(_00783_),
    .RESET_B(net203),
    .Q(\genblk2[9].wave_shpr.div.b1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13467_ (.CLK(clknet_leaf_75_clk),
    .D(_00784_),
    .RESET_B(net203),
    .Q(\genblk2[9].wave_shpr.div.b1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13468_ (.CLK(clknet_leaf_75_clk),
    .D(_00785_),
    .RESET_B(net203),
    .Q(\genblk2[9].wave_shpr.div.b1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13469_ (.CLK(clknet_leaf_85_clk),
    .D(_00786_),
    .RESET_B(net204),
    .Q(\genblk2[9].wave_shpr.div.b1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13470_ (.CLK(clknet_leaf_74_clk),
    .D(_00787_),
    .RESET_B(net203),
    .Q(\genblk2[9].wave_shpr.div.b1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13471_ (.CLK(clknet_leaf_75_clk),
    .D(_00788_),
    .RESET_B(net204),
    .Q(\genblk2[9].wave_shpr.div.b1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13472_ (.CLK(clknet_leaf_74_clk),
    .D(_00789_),
    .RESET_B(net212),
    .Q(\genblk2[9].wave_shpr.div.b1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13473_ (.CLK(clknet_leaf_74_clk),
    .D(_00790_),
    .RESET_B(net215),
    .Q(\genblk2[9].wave_shpr.div.b1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13474_ (.CLK(clknet_leaf_71_clk),
    .D(_00791_),
    .RESET_B(net215),
    .Q(\genblk2[9].wave_shpr.div.b1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13475_ (.CLK(clknet_leaf_71_clk),
    .D(_00792_),
    .RESET_B(net216),
    .Q(\genblk2[9].wave_shpr.div.b1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13476_ (.CLK(clknet_leaf_72_clk),
    .D(_00793_),
    .RESET_B(net216),
    .Q(\genblk2[9].wave_shpr.div.b1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13477_ (.CLK(clknet_leaf_72_clk),
    .D(_00794_),
    .RESET_B(net216),
    .Q(\genblk2[9].wave_shpr.div.b1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13478_ (.CLK(clknet_leaf_99_clk),
    .D(_00795_),
    .RESET_B(net168),
    .Q(\genblk2[8].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13479_ (.CLK(clknet_leaf_99_clk),
    .D(net744),
    .RESET_B(net168),
    .Q(\genblk2[8].wave_shpr.div.quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13480_ (.CLK(clknet_leaf_99_clk),
    .D(_00797_),
    .RESET_B(net168),
    .Q(\genblk2[8].wave_shpr.div.quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13481_ (.CLK(clknet_leaf_100_clk),
    .D(_00798_),
    .RESET_B(net168),
    .Q(\genblk2[8].wave_shpr.div.quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13482_ (.CLK(clknet_leaf_99_clk),
    .D(net347),
    .RESET_B(net168),
    .Q(\genblk2[8].wave_shpr.div.quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13483_ (.CLK(clknet_leaf_99_clk),
    .D(_00800_),
    .RESET_B(net168),
    .Q(\genblk2[8].wave_shpr.div.quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13484_ (.CLK(clknet_leaf_99_clk),
    .D(_00801_),
    .RESET_B(net168),
    .Q(\genblk2[8].wave_shpr.div.quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13485_ (.CLK(clknet_leaf_97_clk),
    .D(_00802_),
    .RESET_B(net167),
    .Q(\genblk2[8].wave_shpr.div.quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13486_ (.CLK(clknet_leaf_79_clk),
    .D(net405),
    .RESET_B(net206),
    .Q(\genblk2[8].wave_shpr.div.quo[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13487_ (.CLK(clknet_leaf_89_clk),
    .D(_00804_),
    .RESET_B(net177),
    .Q(\genblk2[8].wave_shpr.div.quo[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13488_ (.CLK(clknet_leaf_88_clk),
    .D(net330),
    .RESET_B(net177),
    .Q(\genblk2[8].wave_shpr.div.quo[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13489_ (.CLK(clknet_leaf_88_clk),
    .D(net470),
    .RESET_B(net177),
    .Q(\genblk2[8].wave_shpr.div.quo[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13490_ (.CLK(clknet_leaf_88_clk),
    .D(_00807_),
    .RESET_B(net177),
    .Q(\genblk2[8].wave_shpr.div.quo[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13491_ (.CLK(clknet_leaf_88_clk),
    .D(_00808_),
    .RESET_B(net177),
    .Q(\genblk2[8].wave_shpr.div.quo[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13492_ (.CLK(clknet_leaf_87_clk),
    .D(_00809_),
    .RESET_B(net177),
    .Q(\genblk2[8].wave_shpr.div.quo[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13493_ (.CLK(clknet_leaf_86_clk),
    .D(net238),
    .RESET_B(net177),
    .Q(\genblk2[8].wave_shpr.div.quo[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13494_ (.CLK(clknet_leaf_86_clk),
    .D(_00811_),
    .RESET_B(net178),
    .Q(\genblk2[8].wave_shpr.div.quo[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13495_ (.CLK(clknet_leaf_88_clk),
    .D(_00812_),
    .RESET_B(net178),
    .Q(\genblk2[8].wave_shpr.div.quo[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13496_ (.CLK(clknet_leaf_86_clk),
    .D(net264),
    .RESET_B(net178),
    .Q(\genblk2[8].wave_shpr.div.quo[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13497_ (.CLK(clknet_leaf_86_clk),
    .D(net618),
    .RESET_B(net178),
    .Q(\genblk2[8].wave_shpr.div.quo[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13498_ (.CLK(clknet_leaf_86_clk),
    .D(_00815_),
    .RESET_B(net178),
    .Q(\genblk2[8].wave_shpr.div.quo[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13499_ (.CLK(clknet_leaf_86_clk),
    .D(_00816_),
    .RESET_B(net179),
    .Q(\genblk2[8].wave_shpr.div.quo[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13500_ (.CLK(clknet_leaf_87_clk),
    .D(_00817_),
    .RESET_B(net179),
    .Q(\genblk2[8].wave_shpr.div.quo[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13501_ (.CLK(clknet_leaf_86_clk),
    .D(net230),
    .RESET_B(net180),
    .Q(\genblk2[8].wave_shpr.div.quo[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13502_ (.CLK(clknet_leaf_87_clk),
    .D(_00819_),
    .RESET_B(net180),
    .Q(\genblk2[8].wave_shpr.div.quo[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13503_ (.CLK(clknet_leaf_87_clk),
    .D(_00820_),
    .RESET_B(net180),
    .Q(\genblk2[8].wave_shpr.div.acc_next[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13504_ (.CLK(clknet_leaf_81_clk),
    .D(_00821_),
    .RESET_B(net199),
    .Q(\genblk2[8].wave_shpr.div.acc[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13505_ (.CLK(clknet_leaf_98_clk),
    .D(_00822_),
    .RESET_B(net167),
    .Q(\genblk2[8].wave_shpr.div.acc[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13506_ (.CLK(clknet_leaf_98_clk),
    .D(_00823_),
    .RESET_B(net167),
    .Q(\genblk2[8].wave_shpr.div.acc[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13507_ (.CLK(clknet_leaf_80_clk),
    .D(_00824_),
    .RESET_B(net205),
    .Q(\genblk2[8].wave_shpr.div.acc[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13508_ (.CLK(clknet_leaf_79_clk),
    .D(_00825_),
    .RESET_B(net205),
    .Q(\genblk2[8].wave_shpr.div.acc[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13509_ (.CLK(clknet_leaf_80_clk),
    .D(_00826_),
    .RESET_B(net205),
    .Q(\genblk2[8].wave_shpr.div.acc[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13510_ (.CLK(clknet_leaf_80_clk),
    .D(_00827_),
    .RESET_B(net205),
    .Q(\genblk2[8].wave_shpr.div.acc[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13511_ (.CLK(clknet_leaf_78_clk),
    .D(_00828_),
    .RESET_B(net205),
    .Q(\genblk2[8].wave_shpr.div.acc[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13512_ (.CLK(clknet_leaf_78_clk),
    .D(_00829_),
    .RESET_B(net205),
    .Q(\genblk2[8].wave_shpr.div.acc[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13513_ (.CLK(clknet_leaf_78_clk),
    .D(_00830_),
    .RESET_B(net205),
    .Q(\genblk2[8].wave_shpr.div.acc[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13514_ (.CLK(clknet_leaf_78_clk),
    .D(_00831_),
    .RESET_B(net207),
    .Q(\genblk2[8].wave_shpr.div.acc[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13515_ (.CLK(clknet_leaf_78_clk),
    .D(_00832_),
    .RESET_B(net206),
    .Q(\genblk2[8].wave_shpr.div.acc[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13516_ (.CLK(clknet_leaf_78_clk),
    .D(_00833_),
    .RESET_B(net208),
    .Q(\genblk2[8].wave_shpr.div.acc[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13517_ (.CLK(clknet_leaf_77_clk),
    .D(_00834_),
    .RESET_B(net208),
    .Q(\genblk2[8].wave_shpr.div.acc[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13518_ (.CLK(clknet_leaf_78_clk),
    .D(_00835_),
    .RESET_B(net206),
    .Q(\genblk2[8].wave_shpr.div.acc[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13519_ (.CLK(clknet_leaf_79_clk),
    .D(_00836_),
    .RESET_B(net206),
    .Q(\genblk2[8].wave_shpr.div.acc[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13520_ (.CLK(clknet_leaf_79_clk),
    .D(_00837_),
    .RESET_B(net206),
    .Q(\genblk2[8].wave_shpr.div.acc[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13521_ (.CLK(clknet_leaf_79_clk),
    .D(_00838_),
    .RESET_B(net206),
    .Q(\genblk2[8].wave_shpr.div.acc[17] ));
 sky130_fd_sc_hd__dfrtp_2 _13522_ (.CLK(clknet_leaf_79_clk),
    .D(_00839_),
    .RESET_B(net206),
    .Q(\genblk2[8].wave_shpr.div.acc[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13523_ (.CLK(clknet_leaf_98_clk),
    .D(_00840_),
    .RESET_B(net169),
    .Q(\genblk2[8].wave_shpr.div.acc[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13524_ (.CLK(clknet_leaf_98_clk),
    .D(_00841_),
    .RESET_B(net169),
    .Q(\genblk2[8].wave_shpr.div.acc[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13525_ (.CLK(clknet_leaf_98_clk),
    .D(_00842_),
    .RESET_B(net169),
    .Q(\genblk2[8].wave_shpr.div.acc[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13526_ (.CLK(clknet_leaf_98_clk),
    .D(_00843_),
    .RESET_B(net169),
    .Q(\genblk2[8].wave_shpr.div.acc[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13527_ (.CLK(clknet_leaf_98_clk),
    .D(_00844_),
    .RESET_B(net169),
    .Q(\genblk2[8].wave_shpr.div.acc[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13528_ (.CLK(clknet_leaf_98_clk),
    .D(_00845_),
    .RESET_B(net169),
    .Q(\genblk2[8].wave_shpr.div.acc[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13529_ (.CLK(clknet_leaf_98_clk),
    .D(_00846_),
    .RESET_B(net169),
    .Q(\genblk2[8].wave_shpr.div.acc[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13530_ (.CLK(clknet_leaf_98_clk),
    .D(_00847_),
    .RESET_B(net169),
    .Q(\genblk2[8].wave_shpr.div.acc[26] ));
 sky130_fd_sc_hd__dfrtp_1 _13531_ (.CLK(clknet_leaf_84_clk),
    .D(_00022_),
    .RESET_B(net202),
    .Q(\genblk2[9].wave_shpr.div.busy ));
 sky130_fd_sc_hd__dfrtp_1 _13532_ (.CLK(clknet_leaf_97_clk),
    .D(_00023_),
    .RESET_B(net166),
    .Q(\genblk2[9].wave_shpr.div.done ));
 sky130_fd_sc_hd__dfrtp_2 _13533_ (.CLK(clknet_leaf_81_clk),
    .D(_00848_),
    .RESET_B(net199),
    .Q(\genblk2[8].wave_shpr.div.i[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13534_ (.CLK(clknet_leaf_81_clk),
    .D(_00849_),
    .RESET_B(net199),
    .Q(\genblk2[8].wave_shpr.div.i[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13535_ (.CLK(clknet_leaf_81_clk),
    .D(_00850_),
    .RESET_B(net199),
    .Q(\genblk2[8].wave_shpr.div.i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13536_ (.CLK(clknet_leaf_81_clk),
    .D(_00851_),
    .RESET_B(net199),
    .Q(\genblk2[8].wave_shpr.div.i[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13537_ (.CLK(clknet_leaf_81_clk),
    .D(_00852_),
    .RESET_B(net200),
    .Q(\genblk2[8].wave_shpr.div.i[4] ));
 sky130_fd_sc_hd__dfrtp_2 _13538_ (.CLK(clknet_leaf_100_clk),
    .D(_00853_),
    .RESET_B(net165),
    .Q(\genblk2[9].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__dfrtp_2 _13539_ (.CLK(clknet_leaf_100_clk),
    .D(_00854_),
    .RESET_B(net165),
    .Q(\genblk2[9].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13540_ (.CLK(clknet_leaf_101_clk),
    .D(_00855_),
    .RESET_B(net164),
    .Q(\genblk2[9].wave_shpr.div.fin_quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13541_ (.CLK(clknet_leaf_101_clk),
    .D(_00856_),
    .RESET_B(net165),
    .Q(\genblk2[9].wave_shpr.div.fin_quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13542_ (.CLK(clknet_leaf_101_clk),
    .D(_00857_),
    .RESET_B(net165),
    .Q(\genblk2[9].wave_shpr.div.fin_quo[4] ));
 sky130_fd_sc_hd__dfrtp_2 _13543_ (.CLK(clknet_leaf_101_clk),
    .D(_00858_),
    .RESET_B(net164),
    .Q(\genblk2[9].wave_shpr.div.fin_quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13544_ (.CLK(clknet_leaf_101_clk),
    .D(_00859_),
    .RESET_B(net164),
    .Q(\genblk2[9].wave_shpr.div.fin_quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13545_ (.CLK(clknet_leaf_101_clk),
    .D(_00860_),
    .RESET_B(net165),
    .Q(\genblk2[9].wave_shpr.div.fin_quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13546_ (.CLK(clknet_leaf_109_clk),
    .D(_00861_),
    .RESET_B(net152),
    .Q(\sig_norm.b1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13547_ (.CLK(clknet_leaf_109_clk),
    .D(_00862_),
    .RESET_B(net152),
    .Q(\sig_norm.b1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13548_ (.CLK(clknet_leaf_110_clk),
    .D(_00863_),
    .RESET_B(net152),
    .Q(\sig_norm.b1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13549_ (.CLK(clknet_leaf_110_clk),
    .D(_00864_),
    .RESET_B(net152),
    .Q(\sig_norm.b1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13550_ (.CLK(clknet_leaf_100_clk),
    .D(_00865_),
    .RESET_B(net170),
    .Q(\genblk2[9].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13551_ (.CLK(clknet_leaf_100_clk),
    .D(_00866_),
    .RESET_B(net165),
    .Q(\genblk2[9].wave_shpr.div.quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13552_ (.CLK(clknet_leaf_100_clk),
    .D(net650),
    .RESET_B(net165),
    .Q(\genblk2[9].wave_shpr.div.quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13553_ (.CLK(clknet_leaf_100_clk),
    .D(net687),
    .RESET_B(net164),
    .Q(\genblk2[9].wave_shpr.div.quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13554_ (.CLK(clknet_leaf_100_clk),
    .D(_00869_),
    .RESET_B(net164),
    .Q(\genblk2[9].wave_shpr.div.quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13555_ (.CLK(clknet_leaf_101_clk),
    .D(net587),
    .RESET_B(net164),
    .Q(\genblk2[9].wave_shpr.div.quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13556_ (.CLK(clknet_leaf_101_clk),
    .D(_00871_),
    .RESET_B(net164),
    .Q(\genblk2[9].wave_shpr.div.quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13557_ (.CLK(clknet_leaf_97_clk),
    .D(net268),
    .RESET_B(net169),
    .Q(\genblk2[9].wave_shpr.div.quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13558_ (.CLK(clknet_leaf_78_clk),
    .D(_00873_),
    .RESET_B(net208),
    .Q(\genblk2[9].wave_shpr.div.quo[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13559_ (.CLK(clknet_leaf_85_clk),
    .D(_00874_),
    .RESET_B(net184),
    .Q(\genblk2[9].wave_shpr.div.quo[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13560_ (.CLK(clknet_leaf_84_clk),
    .D(net291),
    .RESET_B(net184),
    .Q(\genblk2[9].wave_shpr.div.quo[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13561_ (.CLK(clknet_leaf_85_clk),
    .D(_00876_),
    .RESET_B(net184),
    .Q(\genblk2[9].wave_shpr.div.quo[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13562_ (.CLK(clknet_leaf_85_clk),
    .D(_00877_),
    .RESET_B(net184),
    .Q(\genblk2[9].wave_shpr.div.quo[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13563_ (.CLK(clknet_leaf_57_clk),
    .D(net244),
    .RESET_B(net184),
    .Q(\genblk2[9].wave_shpr.div.quo[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13564_ (.CLK(clknet_leaf_57_clk),
    .D(_00879_),
    .RESET_B(net182),
    .Q(\genblk2[9].wave_shpr.div.quo[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13565_ (.CLK(clknet_leaf_57_clk),
    .D(_00880_),
    .RESET_B(net182),
    .Q(\genblk2[9].wave_shpr.div.quo[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13566_ (.CLK(clknet_leaf_56_clk),
    .D(net305),
    .RESET_B(net182),
    .Q(\genblk2[9].wave_shpr.div.quo[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13567_ (.CLK(clknet_leaf_55_clk),
    .D(net350),
    .RESET_B(net176),
    .Q(\genblk2[9].wave_shpr.div.quo[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13568_ (.CLK(clknet_leaf_55_clk),
    .D(_00883_),
    .RESET_B(net176),
    .Q(\genblk2[9].wave_shpr.div.quo[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13569_ (.CLK(clknet_leaf_55_clk),
    .D(_00884_),
    .RESET_B(net182),
    .Q(\genblk2[9].wave_shpr.div.quo[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13570_ (.CLK(clknet_leaf_56_clk),
    .D(net363),
    .RESET_B(net182),
    .Q(\genblk2[9].wave_shpr.div.quo[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13571_ (.CLK(clknet_leaf_56_clk),
    .D(_00886_),
    .RESET_B(net182),
    .Q(\genblk2[9].wave_shpr.div.quo[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13572_ (.CLK(clknet_leaf_85_clk),
    .D(_00887_),
    .RESET_B(net184),
    .Q(\genblk2[9].wave_shpr.div.quo[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13573_ (.CLK(clknet_leaf_86_clk),
    .D(net227),
    .RESET_B(net183),
    .Q(\genblk2[9].wave_shpr.div.quo[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13574_ (.CLK(clknet_leaf_85_clk),
    .D(_00889_),
    .RESET_B(net183),
    .Q(\genblk2[9].wave_shpr.div.quo[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13575_ (.CLK(clknet_leaf_84_clk),
    .D(net307),
    .RESET_B(net183),
    .Q(\genblk2[9].wave_shpr.div.acc_next[0] ));
 sky130_fd_sc_hd__dfrtp_2 _13576_ (.CLK(clknet_leaf_84_clk),
    .D(net1210),
    .RESET_B(net202),
    .Q(\genblk2[9].wave_shpr.div.acc[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13577_ (.CLK(clknet_leaf_76_clk),
    .D(_00892_),
    .RESET_B(net207),
    .Q(\genblk2[9].wave_shpr.div.acc[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13578_ (.CLK(clknet_leaf_78_clk),
    .D(_00893_),
    .RESET_B(net207),
    .Q(\genblk2[9].wave_shpr.div.acc[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13579_ (.CLK(clknet_leaf_76_clk),
    .D(_00894_),
    .RESET_B(net207),
    .Q(\genblk2[9].wave_shpr.div.acc[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13580_ (.CLK(clknet_leaf_76_clk),
    .D(_00895_),
    .RESET_B(net207),
    .Q(\genblk2[9].wave_shpr.div.acc[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13581_ (.CLK(clknet_leaf_76_clk),
    .D(_00896_),
    .RESET_B(net207),
    .Q(\genblk2[9].wave_shpr.div.acc[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13582_ (.CLK(clknet_leaf_76_clk),
    .D(_00897_),
    .RESET_B(net207),
    .Q(\genblk2[9].wave_shpr.div.acc[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13583_ (.CLK(clknet_leaf_76_clk),
    .D(_00898_),
    .RESET_B(net207),
    .Q(\genblk2[9].wave_shpr.div.acc[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13584_ (.CLK(clknet_leaf_75_clk),
    .D(_00899_),
    .RESET_B(net207),
    .Q(\genblk2[9].wave_shpr.div.acc[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13585_ (.CLK(clknet_leaf_76_clk),
    .D(_00900_),
    .RESET_B(net207),
    .Q(\genblk2[9].wave_shpr.div.acc[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13586_ (.CLK(clknet_leaf_72_clk),
    .D(_00901_),
    .RESET_B(net215),
    .Q(\genblk2[9].wave_shpr.div.acc[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13587_ (.CLK(clknet_leaf_73_clk),
    .D(_00902_),
    .RESET_B(net215),
    .Q(\genblk2[9].wave_shpr.div.acc[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13588_ (.CLK(clknet_leaf_72_clk),
    .D(_00903_),
    .RESET_B(net215),
    .Q(\genblk2[9].wave_shpr.div.acc[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13589_ (.CLK(clknet_leaf_72_clk),
    .D(_00904_),
    .RESET_B(net215),
    .Q(\genblk2[9].wave_shpr.div.acc[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13590_ (.CLK(clknet_leaf_73_clk),
    .D(_00905_),
    .RESET_B(net215),
    .Q(\genblk2[9].wave_shpr.div.acc[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13591_ (.CLK(clknet_leaf_72_clk),
    .D(_00906_),
    .RESET_B(net216),
    .Q(\genblk2[9].wave_shpr.div.acc[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13592_ (.CLK(clknet_leaf_72_clk),
    .D(_00907_),
    .RESET_B(net216),
    .Q(\genblk2[9].wave_shpr.div.acc[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13593_ (.CLK(clknet_leaf_72_clk),
    .D(_00908_),
    .RESET_B(net216),
    .Q(\genblk2[9].wave_shpr.div.acc[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13594_ (.CLK(clknet_leaf_72_clk),
    .D(_00909_),
    .RESET_B(net216),
    .Q(\genblk2[9].wave_shpr.div.acc[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13595_ (.CLK(clknet_leaf_72_clk),
    .D(_00910_),
    .RESET_B(net216),
    .Q(\genblk2[9].wave_shpr.div.acc[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13596_ (.CLK(clknet_leaf_77_clk),
    .D(net936),
    .RESET_B(net208),
    .Q(\genblk2[9].wave_shpr.div.acc[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13597_ (.CLK(clknet_leaf_77_clk),
    .D(_00912_),
    .RESET_B(net208),
    .Q(\genblk2[9].wave_shpr.div.acc[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13598_ (.CLK(clknet_leaf_76_clk),
    .D(net647),
    .RESET_B(net208),
    .Q(\genblk2[9].wave_shpr.div.acc[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13599_ (.CLK(clknet_leaf_77_clk),
    .D(_00914_),
    .RESET_B(net208),
    .Q(\genblk2[9].wave_shpr.div.acc[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13600_ (.CLK(clknet_leaf_76_clk),
    .D(_00915_),
    .RESET_B(net208),
    .Q(\genblk2[9].wave_shpr.div.acc[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13601_ (.CLK(clknet_leaf_77_clk),
    .D(_00916_),
    .RESET_B(net209),
    .Q(\genblk2[9].wave_shpr.div.acc[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13602_ (.CLK(clknet_leaf_77_clk),
    .D(_00917_),
    .RESET_B(net209),
    .Q(\genblk2[9].wave_shpr.div.acc[26] ));
 sky130_fd_sc_hd__dfrtp_1 _13603_ (.CLK(clknet_leaf_45_clk),
    .D(_00002_),
    .RESET_B(net121),
    .Q(\genblk2[10].wave_shpr.div.busy ));
 sky130_fd_sc_hd__dfrtp_1 _13604_ (.CLK(clknet_leaf_97_clk),
    .D(_00003_),
    .RESET_B(net166),
    .Q(\genblk2[10].wave_shpr.div.done ));
 sky130_fd_sc_hd__dfrtp_2 _13605_ (.CLK(clknet_leaf_59_clk),
    .D(_00918_),
    .RESET_B(net193),
    .Q(\genblk2[0].wave_shpr.div.i[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13606_ (.CLK(clknet_leaf_67_clk),
    .D(_00919_),
    .RESET_B(net194),
    .Q(\genblk2[0].wave_shpr.div.i[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13607_ (.CLK(clknet_leaf_68_clk),
    .D(_00920_),
    .RESET_B(net194),
    .Q(\genblk2[0].wave_shpr.div.i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13608_ (.CLK(clknet_leaf_58_clk),
    .D(_00921_),
    .RESET_B(net194),
    .Q(\genblk2[0].wave_shpr.div.i[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13609_ (.CLK(clknet_leaf_58_clk),
    .D(_00922_),
    .RESET_B(net194),
    .Q(\genblk2[0].wave_shpr.div.i[4] ));
 sky130_fd_sc_hd__dfrtp_2 _13610_ (.CLK(clknet_leaf_93_clk),
    .D(_00923_),
    .RESET_B(net159),
    .Q(\genblk2[10].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__dfrtp_2 _13611_ (.CLK(clknet_leaf_93_clk),
    .D(_00924_),
    .RESET_B(net159),
    .Q(\genblk2[10].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13612_ (.CLK(clknet_leaf_94_clk),
    .D(_00925_),
    .RESET_B(net159),
    .Q(\genblk2[10].wave_shpr.div.fin_quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13613_ (.CLK(clknet_leaf_94_clk),
    .D(_00926_),
    .RESET_B(net159),
    .Q(\genblk2[10].wave_shpr.div.fin_quo[3] ));
 sky130_fd_sc_hd__dfrtp_2 _13614_ (.CLK(clknet_leaf_94_clk),
    .D(_00927_),
    .RESET_B(net159),
    .Q(\genblk2[10].wave_shpr.div.fin_quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13615_ (.CLK(clknet_leaf_94_clk),
    .D(_00928_),
    .RESET_B(net160),
    .Q(\genblk2[10].wave_shpr.div.fin_quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13616_ (.CLK(clknet_leaf_94_clk),
    .D(_00929_),
    .RESET_B(net160),
    .Q(\genblk2[10].wave_shpr.div.fin_quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13617_ (.CLK(clknet_leaf_94_clk),
    .D(_00930_),
    .RESET_B(net160),
    .Q(\genblk2[10].wave_shpr.div.fin_quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13618_ (.CLK(clknet_leaf_84_clk),
    .D(_00931_),
    .RESET_B(net204),
    .Q(\genblk2[11].wave_shpr.div.b1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13619_ (.CLK(clknet_leaf_68_clk),
    .D(_00932_),
    .RESET_B(net211),
    .Q(\genblk2[11].wave_shpr.div.b1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13620_ (.CLK(clknet_leaf_75_clk),
    .D(_00933_),
    .RESET_B(net204),
    .Q(\genblk2[11].wave_shpr.div.b1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13621_ (.CLK(clknet_leaf_74_clk),
    .D(_00934_),
    .RESET_B(net212),
    .Q(\genblk2[11].wave_shpr.div.b1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13622_ (.CLK(clknet_leaf_75_clk),
    .D(_00935_),
    .RESET_B(net204),
    .Q(\genblk2[11].wave_shpr.div.b1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13623_ (.CLK(clknet_leaf_85_clk),
    .D(_00936_),
    .RESET_B(net204),
    .Q(\genblk2[11].wave_shpr.div.b1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13624_ (.CLK(clknet_leaf_68_clk),
    .D(_00937_),
    .RESET_B(net194),
    .Q(\genblk2[11].wave_shpr.div.b1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13625_ (.CLK(clknet_leaf_68_clk),
    .D(_00938_),
    .RESET_B(net194),
    .Q(\genblk2[11].wave_shpr.div.b1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13626_ (.CLK(clknet_leaf_67_clk),
    .D(_00939_),
    .RESET_B(net195),
    .Q(\genblk2[11].wave_shpr.div.b1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13627_ (.CLK(clknet_leaf_66_clk),
    .D(_00940_),
    .RESET_B(net197),
    .Q(\genblk2[11].wave_shpr.div.b1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13628_ (.CLK(clknet_leaf_65_clk),
    .D(_00941_),
    .RESET_B(net197),
    .Q(\genblk2[11].wave_shpr.div.b1[10] ));
 sky130_fd_sc_hd__dfrtp_4 _13629_ (.CLK(clknet_leaf_38_clk),
    .D(_00942_),
    .RESET_B(net116),
    .Q(\genblk2[11].wave_shpr.div.b1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13630_ (.CLK(clknet_leaf_67_clk),
    .D(_00943_),
    .RESET_B(net195),
    .Q(\genblk2[11].wave_shpr.div.b1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13631_ (.CLK(clknet_leaf_66_clk),
    .D(_00944_),
    .RESET_B(net197),
    .Q(\genblk2[11].wave_shpr.div.b1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13632_ (.CLK(clknet_leaf_69_clk),
    .D(_00945_),
    .RESET_B(net213),
    .Q(\genblk2[11].wave_shpr.div.b1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13633_ (.CLK(clknet_leaf_69_clk),
    .D(_00946_),
    .RESET_B(net213),
    .Q(\genblk2[11].wave_shpr.div.b1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13634_ (.CLK(clknet_leaf_69_clk),
    .D(_00947_),
    .RESET_B(net211),
    .Q(\genblk2[11].wave_shpr.div.b1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13635_ (.CLK(clknet_leaf_69_clk),
    .D(_00948_),
    .RESET_B(net212),
    .Q(\genblk2[11].wave_shpr.div.b1[17] ));
 sky130_fd_sc_hd__dfrtp_4 _13636_ (.CLK(clknet_leaf_68_clk),
    .D(_00949_),
    .RESET_B(net195),
    .Q(\genblk2[10].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13637_ (.CLK(clknet_leaf_93_clk),
    .D(_00950_),
    .RESET_B(net159),
    .Q(\genblk2[10].wave_shpr.div.quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13638_ (.CLK(clknet_leaf_94_clk),
    .D(net221),
    .RESET_B(net159),
    .Q(\genblk2[10].wave_shpr.div.quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13639_ (.CLK(clknet_leaf_94_clk),
    .D(_00952_),
    .RESET_B(net159),
    .Q(\genblk2[10].wave_shpr.div.quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13640_ (.CLK(clknet_leaf_94_clk),
    .D(net683),
    .RESET_B(net160),
    .Q(\genblk2[10].wave_shpr.div.quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13641_ (.CLK(clknet_leaf_94_clk),
    .D(_00954_),
    .RESET_B(net160),
    .Q(\genblk2[10].wave_shpr.div.quo[5] ));
 sky130_fd_sc_hd__dfrtp_4 _13642_ (.CLK(clknet_leaf_95_clk),
    .D(_00955_),
    .RESET_B(net161),
    .Q(\genblk2[10].wave_shpr.div.quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13643_ (.CLK(clknet_leaf_68_clk),
    .D(_00956_),
    .RESET_B(net211),
    .Q(\genblk2[10].wave_shpr.div.quo[7] ));
 sky130_fd_sc_hd__dfrtp_4 _13644_ (.CLK(clknet_leaf_69_clk),
    .D(net321),
    .RESET_B(net211),
    .Q(\genblk2[10].wave_shpr.div.quo[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13645_ (.CLK(clknet_leaf_48_clk),
    .D(net433),
    .RESET_B(net114),
    .Q(\genblk2[10].wave_shpr.div.quo[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13646_ (.CLK(clknet_leaf_48_clk),
    .D(_00959_),
    .RESET_B(net114),
    .Q(\genblk2[10].wave_shpr.div.quo[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13647_ (.CLK(clknet_leaf_47_clk),
    .D(_00960_),
    .RESET_B(net114),
    .Q(\genblk2[10].wave_shpr.div.quo[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13648_ (.CLK(clknet_leaf_38_clk),
    .D(net224),
    .RESET_B(net126),
    .Q(\genblk2[10].wave_shpr.div.quo[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13649_ (.CLK(clknet_leaf_38_clk),
    .D(_00962_),
    .RESET_B(net126),
    .Q(\genblk2[10].wave_shpr.div.quo[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13650_ (.CLK(clknet_leaf_38_clk),
    .D(_00963_),
    .RESET_B(net116),
    .Q(\genblk2[10].wave_shpr.div.quo[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13651_ (.CLK(clknet_leaf_41_clk),
    .D(_00964_),
    .RESET_B(net116),
    .Q(\genblk2[10].wave_shpr.div.quo[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13652_ (.CLK(clknet_leaf_40_clk),
    .D(_00965_),
    .RESET_B(net116),
    .Q(\genblk2[10].wave_shpr.div.quo[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13653_ (.CLK(clknet_leaf_41_clk),
    .D(net354),
    .RESET_B(net116),
    .Q(\genblk2[10].wave_shpr.div.quo[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13654_ (.CLK(clknet_leaf_41_clk),
    .D(_00967_),
    .RESET_B(net116),
    .Q(\genblk2[10].wave_shpr.div.quo[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13655_ (.CLK(clknet_leaf_41_clk),
    .D(_00968_),
    .RESET_B(net116),
    .Q(\genblk2[10].wave_shpr.div.quo[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13656_ (.CLK(clknet_leaf_44_clk),
    .D(_00969_),
    .RESET_B(net116),
    .Q(\genblk2[10].wave_shpr.div.quo[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13657_ (.CLK(clknet_leaf_48_clk),
    .D(_00970_),
    .RESET_B(net120),
    .Q(\genblk2[10].wave_shpr.div.quo[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13658_ (.CLK(clknet_leaf_44_clk),
    .D(net335),
    .RESET_B(net120),
    .Q(\genblk2[10].wave_shpr.div.quo[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13659_ (.CLK(clknet_leaf_47_clk),
    .D(net475),
    .RESET_B(net120),
    .Q(\genblk2[10].wave_shpr.div.quo[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13660_ (.CLK(clknet_leaf_47_clk),
    .D(net447),
    .RESET_B(net120),
    .Q(\genblk2[10].wave_shpr.div.quo[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13661_ (.CLK(clknet_leaf_47_clk),
    .D(_00974_),
    .RESET_B(net120),
    .Q(\genblk2[10].wave_shpr.div.acc_next[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13662_ (.CLK(clknet_leaf_45_clk),
    .D(net248),
    .RESET_B(net121),
    .Q(\genblk2[10].wave_shpr.div.acc[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13663_ (.CLK(clknet_leaf_44_clk),
    .D(_00976_),
    .RESET_B(net121),
    .Q(\genblk2[10].wave_shpr.div.acc[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13664_ (.CLK(clknet_leaf_43_clk),
    .D(_00977_),
    .RESET_B(net124),
    .Q(\genblk2[10].wave_shpr.div.acc[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13665_ (.CLK(clknet_leaf_43_clk),
    .D(_00978_),
    .RESET_B(net123),
    .Q(\genblk2[10].wave_shpr.div.acc[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13666_ (.CLK(clknet_leaf_41_clk),
    .D(net869),
    .RESET_B(net123),
    .Q(\genblk2[10].wave_shpr.div.acc[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13667_ (.CLK(clknet_leaf_42_clk),
    .D(_00980_),
    .RESET_B(net124),
    .Q(\genblk2[10].wave_shpr.div.acc[5] ));
 sky130_fd_sc_hd__dfrtp_2 _13668_ (.CLK(clknet_leaf_42_clk),
    .D(_00981_),
    .RESET_B(net123),
    .Q(\genblk2[10].wave_shpr.div.acc[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13669_ (.CLK(clknet_leaf_41_clk),
    .D(_00982_),
    .RESET_B(net125),
    .Q(\genblk2[10].wave_shpr.div.acc[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13670_ (.CLK(clknet_leaf_40_clk),
    .D(_00983_),
    .RESET_B(net117),
    .Q(\genblk2[10].wave_shpr.div.acc[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13671_ (.CLK(clknet_leaf_40_clk),
    .D(_00984_),
    .RESET_B(net118),
    .Q(\genblk2[10].wave_shpr.div.acc[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13672_ (.CLK(clknet_leaf_40_clk),
    .D(_00985_),
    .RESET_B(net117),
    .Q(\genblk2[10].wave_shpr.div.acc[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13673_ (.CLK(clknet_leaf_40_clk),
    .D(_00986_),
    .RESET_B(net117),
    .Q(\genblk2[10].wave_shpr.div.acc[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13674_ (.CLK(clknet_leaf_41_clk),
    .D(_00987_),
    .RESET_B(net125),
    .Q(\genblk2[10].wave_shpr.div.acc[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13675_ (.CLK(clknet_leaf_42_clk),
    .D(_00988_),
    .RESET_B(net125),
    .Q(\genblk2[10].wave_shpr.div.acc[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13676_ (.CLK(clknet_leaf_42_clk),
    .D(_00989_),
    .RESET_B(net124),
    .Q(\genblk2[10].wave_shpr.div.acc[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13677_ (.CLK(clknet_leaf_42_clk),
    .D(_00990_),
    .RESET_B(net125),
    .Q(\genblk2[10].wave_shpr.div.acc[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13678_ (.CLK(clknet_leaf_42_clk),
    .D(_00991_),
    .RESET_B(net125),
    .Q(\genblk2[10].wave_shpr.div.acc[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13679_ (.CLK(clknet_leaf_43_clk),
    .D(net860),
    .RESET_B(net190),
    .Q(\genblk2[10].wave_shpr.div.acc[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13680_ (.CLK(clknet_leaf_63_clk),
    .D(_00993_),
    .RESET_B(net190),
    .Q(\genblk2[10].wave_shpr.div.acc[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13681_ (.CLK(clknet_leaf_63_clk),
    .D(_00994_),
    .RESET_B(net125),
    .Q(\genblk2[10].wave_shpr.div.acc[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13682_ (.CLK(clknet_leaf_42_clk),
    .D(_00995_),
    .RESET_B(net190),
    .Q(\genblk2[10].wave_shpr.div.acc[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13683_ (.CLK(clknet_leaf_63_clk),
    .D(_00996_),
    .RESET_B(net190),
    .Q(\genblk2[10].wave_shpr.div.acc[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13684_ (.CLK(clknet_leaf_63_clk),
    .D(_00997_),
    .RESET_B(net191),
    .Q(\genblk2[10].wave_shpr.div.acc[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13685_ (.CLK(clknet_leaf_63_clk),
    .D(_00998_),
    .RESET_B(net191),
    .Q(\genblk2[10].wave_shpr.div.acc[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13686_ (.CLK(clknet_leaf_63_clk),
    .D(_00999_),
    .RESET_B(net191),
    .Q(\genblk2[10].wave_shpr.div.acc[24] ));
 sky130_fd_sc_hd__dfrtp_2 _13687_ (.CLK(clknet_leaf_63_clk),
    .D(_01000_),
    .RESET_B(net191),
    .Q(\genblk2[10].wave_shpr.div.acc[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13688_ (.CLK(clknet_leaf_63_clk),
    .D(_01001_),
    .RESET_B(net190),
    .Q(\genblk2[10].wave_shpr.div.acc[26] ));
 sky130_fd_sc_hd__dfrtp_1 _13689_ (.CLK(clknet_leaf_57_clk),
    .D(_00004_),
    .RESET_B(net184),
    .Q(\genblk2[11].wave_shpr.div.busy ));
 sky130_fd_sc_hd__dfrtp_1 _13690_ (.CLK(clknet_leaf_97_clk),
    .D(_00005_),
    .RESET_B(net166),
    .Q(\genblk2[11].wave_shpr.div.done ));
 sky130_fd_sc_hd__dfrtp_2 _13691_ (.CLK(clknet_leaf_44_clk),
    .D(_01002_),
    .RESET_B(net122),
    .Q(\genblk2[10].wave_shpr.div.i[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13692_ (.CLK(clknet_leaf_44_clk),
    .D(_01003_),
    .RESET_B(net122),
    .Q(\genblk2[10].wave_shpr.div.i[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13693_ (.CLK(clknet_leaf_45_clk),
    .D(_01004_),
    .RESET_B(net122),
    .Q(\genblk2[10].wave_shpr.div.i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13694_ (.CLK(clknet_leaf_45_clk),
    .D(_01005_),
    .RESET_B(net122),
    .Q(\genblk2[10].wave_shpr.div.i[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13695_ (.CLK(clknet_leaf_45_clk),
    .D(_01006_),
    .RESET_B(net188),
    .Q(\genblk2[10].wave_shpr.div.i[4] ));
 sky130_fd_sc_hd__dfrtp_4 _13696_ (.CLK(clknet_leaf_96_clk),
    .D(_01007_),
    .RESET_B(net161),
    .Q(\genblk2[11].wave_shpr.div.fin_quo[0] ));
 sky130_fd_sc_hd__dfrtp_2 _13697_ (.CLK(clknet_leaf_96_clk),
    .D(_01008_),
    .RESET_B(net160),
    .Q(\genblk2[11].wave_shpr.div.fin_quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13698_ (.CLK(clknet_leaf_94_clk),
    .D(_01009_),
    .RESET_B(net160),
    .Q(\genblk2[11].wave_shpr.div.fin_quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13699_ (.CLK(clknet_leaf_94_clk),
    .D(_01010_),
    .RESET_B(net160),
    .Q(\genblk2[11].wave_shpr.div.fin_quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13700_ (.CLK(clknet_leaf_97_clk),
    .D(_01011_),
    .RESET_B(net166),
    .Q(\genblk2[11].wave_shpr.div.fin_quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13701_ (.CLK(clknet_leaf_99_clk),
    .D(_01012_),
    .RESET_B(net166),
    .Q(\genblk2[11].wave_shpr.div.fin_quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13702_ (.CLK(clknet_leaf_97_clk),
    .D(_01013_),
    .RESET_B(net167),
    .Q(\genblk2[11].wave_shpr.div.fin_quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13703_ (.CLK(clknet_leaf_96_clk),
    .D(_01014_),
    .RESET_B(net161),
    .Q(\genblk2[11].wave_shpr.div.fin_quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13704_ (.CLK(clknet_leaf_37_clk),
    .D(_01015_),
    .RESET_B(net113),
    .Q(\genblk2[1].wave_shpr.div.b1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13705_ (.CLK(clknet_leaf_37_clk),
    .D(_01016_),
    .RESET_B(net113),
    .Q(\genblk2[1].wave_shpr.div.b1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13706_ (.CLK(clknet_leaf_37_clk),
    .D(_01017_),
    .RESET_B(net114),
    .Q(\genblk2[1].wave_shpr.div.b1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13707_ (.CLK(clknet_leaf_37_clk),
    .D(_01018_),
    .RESET_B(net104),
    .Q(\genblk2[1].wave_shpr.div.b1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13708_ (.CLK(clknet_leaf_36_clk),
    .D(_01019_),
    .RESET_B(net104),
    .Q(\genblk2[1].wave_shpr.div.b1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13709_ (.CLK(clknet_leaf_31_clk),
    .D(_01020_),
    .RESET_B(net103),
    .Q(\genblk2[1].wave_shpr.div.b1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13710_ (.CLK(clknet_leaf_31_clk),
    .D(_01021_),
    .RESET_B(net103),
    .Q(\genblk2[1].wave_shpr.div.b1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13711_ (.CLK(clknet_leaf_31_clk),
    .D(_01022_),
    .RESET_B(net100),
    .Q(\genblk2[1].wave_shpr.div.b1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13712_ (.CLK(clknet_leaf_31_clk),
    .D(_01023_),
    .RESET_B(net100),
    .Q(\genblk2[1].wave_shpr.div.b1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13713_ (.CLK(clknet_leaf_31_clk),
    .D(_01024_),
    .RESET_B(net99),
    .Q(\genblk2[1].wave_shpr.div.b1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13714_ (.CLK(clknet_leaf_31_clk),
    .D(_01025_),
    .RESET_B(net102),
    .Q(\genblk2[1].wave_shpr.div.b1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13715_ (.CLK(clknet_leaf_21_clk),
    .D(_01026_),
    .RESET_B(net97),
    .Q(\genblk2[1].wave_shpr.div.b1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13716_ (.CLK(clknet_leaf_36_clk),
    .D(_01027_),
    .RESET_B(net103),
    .Q(\genblk2[1].wave_shpr.div.b1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13717_ (.CLK(clknet_leaf_36_clk),
    .D(_01028_),
    .RESET_B(net105),
    .Q(\genblk2[1].wave_shpr.div.b1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13718_ (.CLK(clknet_leaf_36_clk),
    .D(_01029_),
    .RESET_B(net105),
    .Q(\genblk2[1].wave_shpr.div.b1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13719_ (.CLK(clknet_leaf_36_clk),
    .D(_01030_),
    .RESET_B(net105),
    .Q(\genblk2[1].wave_shpr.div.b1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13720_ (.CLK(clknet_leaf_39_clk),
    .D(_01031_),
    .RESET_B(net115),
    .Q(\genblk2[1].wave_shpr.div.b1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13721_ (.CLK(clknet_leaf_40_clk),
    .D(_01032_),
    .RESET_B(net118),
    .Q(\genblk2[1].wave_shpr.div.b1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13722_ (.CLK(clknet_leaf_97_clk),
    .D(_01033_),
    .RESET_B(net161),
    .Q(\genblk2[11].wave_shpr.div.quo[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13723_ (.CLK(clknet_leaf_96_clk),
    .D(net431),
    .RESET_B(net160),
    .Q(\genblk2[11].wave_shpr.div.quo[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13724_ (.CLK(clknet_leaf_96_clk),
    .D(_01035_),
    .RESET_B(net160),
    .Q(\genblk2[11].wave_shpr.div.quo[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13725_ (.CLK(clknet_leaf_97_clk),
    .D(net403),
    .RESET_B(net166),
    .Q(\genblk2[11].wave_shpr.div.quo[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13726_ (.CLK(clknet_leaf_97_clk),
    .D(_01037_),
    .RESET_B(net166),
    .Q(\genblk2[11].wave_shpr.div.quo[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13727_ (.CLK(clknet_leaf_97_clk),
    .D(_01038_),
    .RESET_B(net167),
    .Q(\genblk2[11].wave_shpr.div.quo[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13728_ (.CLK(clknet_leaf_97_clk),
    .D(_01039_),
    .RESET_B(net167),
    .Q(\genblk2[11].wave_shpr.div.quo[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13729_ (.CLK(clknet_leaf_74_clk),
    .D(_01040_),
    .RESET_B(net212),
    .Q(\genblk2[11].wave_shpr.div.quo[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13730_ (.CLK(clknet_leaf_74_clk),
    .D(_01041_),
    .RESET_B(net212),
    .Q(\genblk2[11].wave_shpr.div.quo[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13731_ (.CLK(clknet_leaf_45_clk),
    .D(net356),
    .RESET_B(net121),
    .Q(\genblk2[11].wave_shpr.div.quo[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13732_ (.CLK(clknet_leaf_45_clk),
    .D(_01043_),
    .RESET_B(net121),
    .Q(\genblk2[11].wave_shpr.div.quo[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13733_ (.CLK(clknet_leaf_45_clk),
    .D(net468),
    .RESET_B(net121),
    .Q(\genblk2[11].wave_shpr.div.quo[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13734_ (.CLK(clknet_leaf_46_clk),
    .D(net444),
    .RESET_B(net119),
    .Q(\genblk2[11].wave_shpr.div.quo[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13735_ (.CLK(clknet_leaf_46_clk),
    .D(_01046_),
    .RESET_B(net119),
    .Q(\genblk2[11].wave_shpr.div.quo[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13736_ (.CLK(clknet_leaf_47_clk),
    .D(net343),
    .RESET_B(net119),
    .Q(\genblk2[11].wave_shpr.div.quo[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13737_ (.CLK(clknet_leaf_47_clk),
    .D(_01048_),
    .RESET_B(net119),
    .Q(\genblk2[11].wave_shpr.div.quo[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13738_ (.CLK(clknet_leaf_46_clk),
    .D(net352),
    .RESET_B(net119),
    .Q(\genblk2[11].wave_shpr.div.quo[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13739_ (.CLK(clknet_leaf_46_clk),
    .D(_01050_),
    .RESET_B(net119),
    .Q(\genblk2[11].wave_shpr.div.quo[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13740_ (.CLK(clknet_leaf_46_clk),
    .D(_01051_),
    .RESET_B(net121),
    .Q(\genblk2[11].wave_shpr.div.quo[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13741_ (.CLK(clknet_leaf_46_clk),
    .D(_01052_),
    .RESET_B(net121),
    .Q(\genblk2[11].wave_shpr.div.quo[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13742_ (.CLK(clknet_leaf_46_clk),
    .D(_01053_),
    .RESET_B(net121),
    .Q(\genblk2[11].wave_shpr.div.quo[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13743_ (.CLK(clknet_leaf_51_clk),
    .D(net240),
    .RESET_B(net110),
    .Q(\genblk2[11].wave_shpr.div.quo[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13744_ (.CLK(clknet_leaf_51_clk),
    .D(_01055_),
    .RESET_B(net110),
    .Q(\genblk2[11].wave_shpr.div.quo[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13745_ (.CLK(clknet_leaf_51_clk),
    .D(net439),
    .RESET_B(net110),
    .Q(\genblk2[11].wave_shpr.div.quo[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13746_ (.CLK(clknet_leaf_51_clk),
    .D(net435),
    .RESET_B(net110),
    .Q(\genblk2[11].wave_shpr.div.quo[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13747_ (.CLK(clknet_leaf_51_clk),
    .D(net413),
    .RESET_B(net111),
    .Q(\genblk2[11].wave_shpr.div.acc_next[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13748_ (.CLK(clknet_leaf_85_clk),
    .D(net1221),
    .RESET_B(net184),
    .Q(\genblk2[11].wave_shpr.div.acc[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13749_ (.CLK(clknet_leaf_75_clk),
    .D(_01060_),
    .RESET_B(net211),
    .Q(\genblk2[11].wave_shpr.div.acc[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13750_ (.CLK(clknet_leaf_75_clk),
    .D(_01061_),
    .RESET_B(net211),
    .Q(\genblk2[11].wave_shpr.div.acc[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13751_ (.CLK(clknet_leaf_74_clk),
    .D(_01062_),
    .RESET_B(net212),
    .Q(\genblk2[11].wave_shpr.div.acc[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13752_ (.CLK(clknet_leaf_68_clk),
    .D(_01063_),
    .RESET_B(net211),
    .Q(\genblk2[11].wave_shpr.div.acc[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13753_ (.CLK(clknet_leaf_68_clk),
    .D(_01064_),
    .RESET_B(net211),
    .Q(\genblk2[11].wave_shpr.div.acc[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13754_ (.CLK(clknet_leaf_68_clk),
    .D(_01065_),
    .RESET_B(net212),
    .Q(\genblk2[11].wave_shpr.div.acc[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13755_ (.CLK(clknet_leaf_68_clk),
    .D(_01066_),
    .RESET_B(net212),
    .Q(\genblk2[11].wave_shpr.div.acc[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13756_ (.CLK(clknet_leaf_69_clk),
    .D(_01067_),
    .RESET_B(net212),
    .Q(\genblk2[11].wave_shpr.div.acc[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13757_ (.CLK(clknet_leaf_70_clk),
    .D(_01068_),
    .RESET_B(net213),
    .Q(\genblk2[11].wave_shpr.div.acc[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13758_ (.CLK(clknet_leaf_66_clk),
    .D(_01069_),
    .RESET_B(net197),
    .Q(\genblk2[11].wave_shpr.div.acc[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13759_ (.CLK(clknet_leaf_66_clk),
    .D(_01070_),
    .RESET_B(net213),
    .Q(\genblk2[11].wave_shpr.div.acc[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13760_ (.CLK(clknet_leaf_70_clk),
    .D(_01071_),
    .RESET_B(net213),
    .Q(\genblk2[11].wave_shpr.div.acc[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13761_ (.CLK(clknet_leaf_70_clk),
    .D(_01072_),
    .RESET_B(net214),
    .Q(\genblk2[11].wave_shpr.div.acc[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13762_ (.CLK(clknet_leaf_69_clk),
    .D(net994),
    .RESET_B(net214),
    .Q(\genblk2[11].wave_shpr.div.acc[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13763_ (.CLK(clknet_leaf_69_clk),
    .D(_01074_),
    .RESET_B(net214),
    .Q(\genblk2[11].wave_shpr.div.acc[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13764_ (.CLK(clknet_leaf_69_clk),
    .D(_01075_),
    .RESET_B(net214),
    .Q(\genblk2[11].wave_shpr.div.acc[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13765_ (.CLK(clknet_leaf_69_clk),
    .D(_01076_),
    .RESET_B(net213),
    .Q(\genblk2[11].wave_shpr.div.acc[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13766_ (.CLK(clknet_leaf_69_clk),
    .D(_01077_),
    .RESET_B(net213),
    .Q(\genblk2[11].wave_shpr.div.acc[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13767_ (.CLK(clknet_leaf_71_clk),
    .D(_01078_),
    .RESET_B(net214),
    .Q(\genblk2[11].wave_shpr.div.acc[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13768_ (.CLK(clknet_leaf_71_clk),
    .D(_01079_),
    .RESET_B(net217),
    .Q(\genblk2[11].wave_shpr.div.acc[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13769_ (.CLK(clknet_leaf_71_clk),
    .D(_01080_),
    .RESET_B(net217),
    .Q(\genblk2[11].wave_shpr.div.acc[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13770_ (.CLK(clknet_leaf_71_clk),
    .D(_01081_),
    .RESET_B(net215),
    .Q(\genblk2[11].wave_shpr.div.acc[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13771_ (.CLK(clknet_leaf_73_clk),
    .D(_01082_),
    .RESET_B(net215),
    .Q(\genblk2[11].wave_shpr.div.acc[23] ));
 sky130_fd_sc_hd__dfrtp_2 _13772_ (.CLK(clknet_leaf_73_clk),
    .D(_01083_),
    .RESET_B(net215),
    .Q(\genblk2[11].wave_shpr.div.acc[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13773_ (.CLK(clknet_leaf_74_clk),
    .D(_01084_),
    .RESET_B(net213),
    .Q(\genblk2[11].wave_shpr.div.acc[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13774_ (.CLK(clknet_leaf_73_clk),
    .D(_01085_),
    .RESET_B(net213),
    .Q(\genblk2[11].wave_shpr.div.acc[26] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_2 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 fanout101 (.A(net107),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_4 fanout102 (.A(net104),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 fanout103 (.A(net104),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_4 fanout104 (.A(net107),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_4 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__buf_2 fanout106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__buf_2 fanout107 (.A(net127),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__buf_2 fanout109 (.A(net127),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_4 fanout110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__buf_2 fanout112 (.A(net127),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_4 fanout113 (.A(net114),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 fanout114 (.A(net126),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 fanout115 (.A(net118),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_4 fanout116 (.A(net118),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 fanout117 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__buf_2 fanout118 (.A(net126),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 fanout119 (.A(net122),
    .X(net119));
 sky130_fd_sc_hd__buf_2 fanout120 (.A(net122),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_4 fanout121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__buf_2 fanout122 (.A(net126),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_4 fanout123 (.A(net125),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_4 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__buf_2 fanout125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__buf_2 fanout126 (.A(net127),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_4 fanout127 (.A(net16),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_4 fanout128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 fanout129 (.A(net131),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_4 fanout130 (.A(net131),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 fanout131 (.A(net136),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(net133),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_4 fanout133 (.A(net135),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_4 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__buf_2 fanout135 (.A(net136),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_4 fanout136 (.A(net171),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_4 fanout137 (.A(net145),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_4 fanout138 (.A(net145),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_4 fanout139 (.A(net140),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_4 fanout140 (.A(net145),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_4 fanout141 (.A(net145),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 fanout142 (.A(net145),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_4 fanout143 (.A(net145),
    .X(net143));
 sky130_fd_sc_hd__buf_2 fanout144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_4 fanout145 (.A(net171),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_4 fanout146 (.A(net150),
    .X(net146));
 sky130_fd_sc_hd__buf_2 fanout147 (.A(net171),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 fanout148 (.A(net150),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 fanout149 (.A(net150),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_4 fanout150 (.A(net171),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_4 fanout151 (.A(net152),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_4 fanout152 (.A(net158),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_4 fanout153 (.A(net155),
    .X(net153));
 sky130_fd_sc_hd__buf_2 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_4 fanout155 (.A(net157),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 fanout157 (.A(net158),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_2 fanout158 (.A(net171),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_4 fanout159 (.A(net162),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_4 fanout160 (.A(net162),
    .X(net160));
 sky130_fd_sc_hd__buf_2 fanout161 (.A(net162),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 fanout162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 fanout163 (.A(net171),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_4 fanout164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_4 fanout165 (.A(net170),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_4 fanout166 (.A(net170),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_4 fanout167 (.A(net170),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_4 fanout168 (.A(net170),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_4 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__buf_2 fanout170 (.A(net171),
    .X(net170));
 sky130_fd_sc_hd__buf_4 fanout171 (.A(net16),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_4 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 fanout173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__buf_2 fanout174 (.A(net218),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_4 fanout175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_2 fanout176 (.A(net218),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_4 fanout177 (.A(net180),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_2 fanout178 (.A(net180),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_4 fanout179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__buf_2 fanout180 (.A(net185),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_4 fanout181 (.A(net185),
    .X(net181));
 sky130_fd_sc_hd__buf_2 fanout182 (.A(net185),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_4 fanout183 (.A(net185),
    .X(net183));
 sky130_fd_sc_hd__buf_2 fanout184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 fanout185 (.A(net218),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_4 fanout186 (.A(net188),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_4 fanout187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__buf_2 fanout188 (.A(net198),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_4 fanout189 (.A(net191),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_4 fanout190 (.A(net198),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_2 fanout191 (.A(net198),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(net193),
    .X(net192));
 sky130_fd_sc_hd__buf_2 fanout193 (.A(net195),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_4 fanout194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 fanout195 (.A(net198),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_4 fanout196 (.A(net198),
    .X(net196));
 sky130_fd_sc_hd__buf_2 fanout197 (.A(net198),
    .X(net197));
 sky130_fd_sc_hd__buf_2 fanout198 (.A(net218),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_4 fanout199 (.A(net210),
    .X(net199));
 sky130_fd_sc_hd__buf_2 fanout200 (.A(net210),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_4 fanout201 (.A(net210),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_4 fanout202 (.A(net204),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_4 fanout203 (.A(net204),
    .X(net203));
 sky130_fd_sc_hd__buf_2 fanout204 (.A(net210),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_4 fanout205 (.A(net209),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_4 fanout206 (.A(net209),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_4 fanout207 (.A(net208),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_4 fanout208 (.A(net209),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 fanout209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__buf_2 fanout210 (.A(net218),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_4 fanout211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_4 fanout212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_4 fanout213 (.A(net217),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 fanout214 (.A(net217),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_4 fanout215 (.A(net217),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_4 fanout216 (.A(net217),
    .X(net216));
 sky130_fd_sc_hd__buf_2 fanout217 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_4 fanout218 (.A(net16),
    .X(net218));
 sky130_fd_sc_hd__buf_4 fanout38 (.A(net44),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 fanout39 (.A(net44),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 fanout40 (.A(net44),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 fanout41 (.A(net43),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(net43),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 fanout43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 fanout44 (.A(net85),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 fanout45 (.A(net47),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__buf_2 fanout47 (.A(net50),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 fanout48 (.A(net50),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 fanout49 (.A(net50),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 fanout50 (.A(net85),
    .X(net50));
 sky130_fd_sc_hd__buf_4 fanout51 (.A(net53),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 fanout52 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__buf_2 fanout53 (.A(net58),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 fanout54 (.A(net58),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 fanout55 (.A(net58),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_4 fanout56 (.A(net58),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 fanout57 (.A(net58),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 fanout58 (.A(net85),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 fanout59 (.A(net63),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 fanout60 (.A(net63),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 fanout61 (.A(net62),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 fanout62 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__buf_2 fanout63 (.A(net85),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_4 fanout64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 fanout65 (.A(net68),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 fanout66 (.A(net68),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 fanout67 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 fanout68 (.A(net85),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_4 fanout69 (.A(net75),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 fanout70 (.A(net75),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_4 fanout71 (.A(net72),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_4 fanout72 (.A(net75),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_4 fanout73 (.A(net74),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_4 fanout74 (.A(net75),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 fanout75 (.A(net84),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 fanout76 (.A(net84),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 fanout77 (.A(net84),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_4 fanout78 (.A(net79),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_4 fanout79 (.A(net84),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_4 fanout80 (.A(net83),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_4 fanout81 (.A(net83),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 fanout82 (.A(net83),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 fanout83 (.A(net84),
    .X(net83));
 sky130_fd_sc_hd__buf_2 fanout84 (.A(net85),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 fanout85 (.A(net16),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_4 fanout86 (.A(net88),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_4 fanout87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_4 fanout88 (.A(net91),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_4 fanout89 (.A(net90),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 fanout90 (.A(net91),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_4 fanout91 (.A(net127),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_4 fanout92 (.A(net94),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 fanout93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_4 fanout94 (.A(net98),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_4 fanout95 (.A(net98),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_4 fanout96 (.A(net98),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_4 fanout97 (.A(net98),
    .X(net97));
 sky130_fd_sc_hd__buf_2 fanout98 (.A(net127),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_4 fanout99 (.A(net101),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\PWM.pwm_out ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\modein.delay_octave_up_in[0] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_00718_),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(\genblk2[0].wave_shpr.div.fin_quo[7] ),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(_03812_),
    .X(net1219));
 sky130_fd_sc_hd__clkbuf_2 hold1002 (.A(\genblk1[11].osc.clkdiv_C.cnt[17] ),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(_01059_),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(\genblk2[8].wave_shpr.div.acc[18] ),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(\genblk2[5].wave_shpr.div.b1[17] ),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(\genblk2[10].wave_shpr.div.b1[10] ),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(\genblk2[4].wave_shpr.div.b1[7] ),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(\genblk2[10].wave_shpr.div.acc[25] ),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(\genblk2[4].wave_shpr.div.b1[17] ),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\genblk2[8].wave_shpr.div.i[4] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(\genblk2[1].wave_shpr.div.acc[25] ),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(\genblk1[5].osc.clkdiv_C.cnt[13] ),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(\genblk2[9].wave_shpr.div.b1[3] ),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(\genblk2[9].wave_shpr.div.b1[10] ),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(\genblk2[4].wave_shpr.div.b1[10] ),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(\genblk2[6].wave_shpr.div.b1[11] ),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(\genblk2[7].wave_shpr.div.b1[17] ),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(\genblk2[1].wave_shpr.div.b1[3] ),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(\genblk2[9].wave_shpr.div.b1[8] ),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(\genblk1[3].osc.clkdiv_C.cnt[15] ),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\genblk2[10].wave_shpr.div.quo[7] ),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(\genblk2[0].wave_shpr.div.b1[3] ),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(\genblk2[9].wave_shpr.div.b1[17] ),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(\sig_norm.acc[4] ),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(\genblk2[10].wave_shpr.div.acc[6] ),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(\genblk2[11].wave_shpr.div.b1[6] ),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(\genblk2[0].wave_shpr.div.b1[1] ),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(\genblk2[10].wave_shpr.div.b1[8] ),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(\genblk2[3].wave_shpr.div.b1[4] ),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(\genblk2[8].wave_shpr.div.b1[9] ),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(\genblk2[2].wave_shpr.div.b1[1] ),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_00957_),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(\genblk2[6].wave_shpr.div.b1[12] ),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(\genblk2[10].wave_shpr.div.b1[3] ),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(\genblk2[7].wave_shpr.div.b1[3] ),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(\genblk2[10].wave_shpr.div.b1[13] ),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(\genblk1[7].osc.clkdiv_C.cnt[1] ),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(\genblk2[7].wave_shpr.div.b1[10] ),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(\genblk2[10].wave_shpr.div.b1[7] ),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(\genblk1[7].osc.clkdiv_C.cnt[17] ),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(\genblk1[2].osc.clkdiv_C.cnt[12] ),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(\genblk2[10].wave_shpr.div.acc[22] ),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\genblk2[2].wave_shpr.div.quo[19] ),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(\genblk2[6].wave_shpr.div.b1[6] ),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(\genblk2[9].wave_shpr.div.fin_quo[7] ),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(\genblk2[1].wave_shpr.div.acc[6] ),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(\sig_norm.quo[10] ),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(\genblk2[4].wave_shpr.div.b1[14] ),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(\genblk2[4].wave_shpr.div.quo[6] ),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(_04631_),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(\genblk2[11].wave_shpr.div.b1[3] ),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(\genblk2[5].wave_shpr.div.b1[11] ),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(\genblk2[1].wave_shpr.div.b1[4] ),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_00311_),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(\genblk2[9].wave_shpr.div.b1[4] ),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(\genblk1[11].osc.clkdiv_C.cnt[10] ),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(\genblk2[1].wave_shpr.div.b1[14] ),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(\genblk2[2].wave_shpr.div.b1[13] ),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(\genblk2[1].wave_shpr.div.b1[5] ),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(\genblk2[10].wave_shpr.div.b1[4] ),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(\genblk2[1].wave_shpr.div.b1[7] ),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(\genblk2[11].wave_shpr.div.b1[7] ),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(\genblk2[0].wave_shpr.div.b1[9] ),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(\genblk2[2].wave_shpr.div.b1[12] ),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\genblk2[5].wave_shpr.div.quo[24] ),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(\genblk2[11].wave_shpr.div.b1[17] ),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(\genblk2[5].wave_shpr.div.b1[12] ),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(\genblk2[8].wave_shpr.div.b1[8] ),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(\genblk2[4].wave_shpr.div.b1[13] ),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(\genblk2[2].wave_shpr.div.b1[14] ),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(\genblk2[5].wave_shpr.div.b1[10] ),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(\genblk2[10].wave_shpr.div.b1[9] ),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(\genblk2[3].wave_shpr.div.b1[12] ),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(\genblk2[7].wave_shpr.div.b1[9] ),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(\genblk2[5].wave_shpr.div.b1[4] ),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_00568_),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(\genblk2[7].wave_shpr.div.b1[2] ),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(\genblk2[0].wave_shpr.div.b1[7] ),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(\genblk2[3].wave_shpr.div.b1[3] ),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(\genblk2[0].wave_shpr.div.b1[14] ),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(\genblk2[10].wave_shpr.div.b1[11] ),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(\genblk2[7].wave_shpr.div.b1[5] ),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(\genblk2[9].wave_shpr.div.b1[2] ),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(\genblk2[1].wave_shpr.div.b1[2] ),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(\genblk1[9].osc.clkdiv_C.cnt[12] ),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(\genblk2[3].wave_shpr.div.b1[11] ),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\genblk2[3].wave_shpr.div.quo[1] ),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(\genblk2[3].wave_shpr.div.b1[8] ),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(\genblk2[1].wave_shpr.div.b1[13] ),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(\sig_norm.quo[7] ),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(\genblk2[7].wave_shpr.div.b1[12] ),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(\genblk2[10].wave_shpr.div.b1[17] ),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(\genblk2[5].wave_shpr.div.b1[9] ),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(\genblk2[2].wave_shpr.div.b1[10] ),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(\genblk2[0].wave_shpr.div.acc[24] ),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(_00173_),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(\PWM.counter[4] ),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_00377_),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(\genblk2[6].wave_shpr.div.b1[8] ),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(\genblk2[4].wave_shpr.div.quo[0] ),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(\genblk2[11].wave_shpr.div.quo[0] ),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(\genblk2[7].wave_shpr.div.quo[1] ),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(\genblk2[1].wave_shpr.div.quo[1] ),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(\genblk2[9].wave_shpr.div.quo[1] ),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(\genblk2[0].wave_shpr.div.quo[2] ),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(\genblk2[5].wave_shpr.div.quo[5] ),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(\genblk2[1].wave_shpr.div.quo[3] ),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(\genblk2[9].wave_shpr.div.quo[4] ),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\genblk2[8].wave_shpr.div.quo[22] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\genblk2[7].wave_shpr.div.i[4] ),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(\genblk2[7].wave_shpr.div.quo[3] ),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(\genblk2[6].wave_shpr.div.quo[3] ),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(\genblk2[6].wave_shpr.div.quo[2] ),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(\genblk2[8].wave_shpr.div.quo[3] ),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(\genblk2[0].wave_shpr.div.quo[1] ),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(\genblk2[10].wave_shpr.div.quo[3] ),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(\genblk2[10].wave_shpr.div.quo[5] ),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(\genblk2[8].wave_shpr.div.quo[5] ),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(\genblk2[5].wave_shpr.div.quo[3] ),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(\genblk2[2].wave_shpr.div.quo[3] ),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\genblk2[8].wave_shpr.div.quo[9] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(\genblk2[9].wave_shpr.div.quo[0] ),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(\genblk2[2].wave_shpr.div.quo[2] ),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(\genblk2[5].wave_shpr.div.quo[4] ),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\genblk2[8].wave_shpr.div.quo[0] ),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(\genblk2[11].wave_shpr.div.quo[5] ),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(\genblk2[4].wave_shpr.div.quo[3] ),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(\genblk2[0].wave_shpr.div.quo[4] ),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(\genblk2[8].wave_shpr.div.quo[6] ),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(\genblk2[5].wave_shpr.div.quo[1] ),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(\genblk2[8].wave_shpr.div.quo[2] ),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_00805_),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(\genblk2[6].wave_shpr.div.quo[1] ),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(\sig_norm.quo[4] ),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(\genblk2[4].wave_shpr.div.acc[7] ),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(\genblk2[11].wave_shpr.div.quo[6] ),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(\genblk2[5].wave_shpr.div.quo[0] ),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(\genblk2[2].wave_shpr.div.quo[1] ),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(\genblk2[5].wave_shpr.div.quo[6] ),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(\genblk2[5].wave_shpr.div.acc[20] ),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(\genblk2[3].wave_shpr.div.quo[5] ),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(\genblk2[7].wave_shpr.div.quo[0] ),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\genblk2[7].wave_shpr.div.quo[3] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(\genblk2[2].wave_shpr.div.quo[0] ),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1131 (.A(\genblk2[6].wave_shpr.div.quo[6] ),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_00715_),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\genblk2[3].wave_shpr.div.i[4] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\genblk2[10].wave_shpr.div.quo[21] ),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_00971_),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\genblk2[2].wave_shpr.div.quo[3] ),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_00295_),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_00818_),
    .X(net230));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold120 (.A(\smpl_rt_clkdiv.clkDiv_inst.cnt[0] ),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\genblk2[2].wave_shpr.div.quo[18] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\genblk2[1].wave_shpr.div.quo[22] ),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_00230_),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\genblk2[11].wave_shpr.div.quo[13] ),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_01047_),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\genblk2[6].wave_shpr.div.quo[10] ),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_00638_),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\genblk2[8].wave_shpr.div.quo[3] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_00799_),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\genblk2[7].wave_shpr.div.quo[19] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\genblk2[9].wave_shpr.div.acc[26] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\genblk2[9].wave_shpr.div.quo[16] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_00882_),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\genblk2[11].wave_shpr.div.quo[15] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_01049_),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\genblk2[10].wave_shpr.div.quo[16] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_00966_),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_2 hold137 (.A(\genblk2[11].wave_shpr.div.quo[8] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_01042_),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\genblk2[10].wave_shpr.div.quo[15] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_00731_),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\genblk2[11].wave_shpr.div.quo[7] ),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\smpl_rt_clkdiv.clkDiv_inst.cnt[2] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_01090_),
    .X(net360));
 sky130_fd_sc_hd__buf_1 hold143 (.A(\PWM.counter[0] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\genblk2[9].wave_shpr.div.quo[19] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_00885_),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\smpl_rt_clkdiv.clkDiv_inst.cnt[1] ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\smpl_rt_clkdiv.clkDiv_inst.cnt[6] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\genblk2[1].wave_shpr.div.acc[11] ),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_00245_),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\genblk2[5].wave_shpr.div.quo[19] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\smpl_rt_clkdiv.clkDiv_inst.cnt[3] ),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\genblk2[2].wave_shpr.div.b1[15] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\genblk2[7].wave_shpr.div.quo[11] ),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_00723_),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\sig_norm.quo[8] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\genblk2[10].wave_shpr.div.quo[14] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\genblk2[9].wave_shpr.div.b1[14] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\genblk2[3].wave_shpr.div.acc[26] ),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\genblk2[3].wave_shpr.div.quo[16] ),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_00392_),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_00563_),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\genblk2[5].wave_shpr.div.quo[16] ),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\genblk2[0].wave_shpr.div.quo[7] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\smpl_rt_clkdiv.clkDiv_inst.cnt[4] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\genblk2[7].wave_shpr.div.acc[26] ),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_00763_),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\genblk2[10].wave_shpr.div.quo[20] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\genblk2[11].wave_shpr.div.b1[14] ),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\genblk2[6].wave_shpr.div.quo[23] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_00651_),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\genblk2[3].wave_shpr.div.quo[12] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\genblk2[5].wave_shpr.div.quo[17] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_00388_),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\genblk2[8].wave_shpr.div.b1[2] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\genblk2[9].wave_shpr.div.b1[15] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\genblk2[8].wave_shpr.div.b1[15] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\genblk2[5].wave_shpr.div.acc[26] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\genblk2[2].wave_shpr.div.quo[17] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\genblk2[0].wave_shpr.div.b1[6] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\smpl_rt_clkdiv.clkDiv_inst.cnt[7] ),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\genblk2[0].wave_shpr.div.b1[16] ),
    .X(net396));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold179 (.A(\genblk2[11].wave_shpr.div.quo[6] ),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_00561_),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\genblk2[10].wave_shpr.div.quo[10] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\PWM.counter[7] ),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\genblk2[7].wave_shpr.div.quo[18] ),
    .X(net400));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold183 (.A(\genblk2[3].wave_shpr.div.quo[7] ),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\genblk2[11].wave_shpr.div.quo[2] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_01036_),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\genblk2[8].wave_shpr.div.quo[7] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_00803_),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\genblk2[1].wave_shpr.div.b1[15] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\smpl_rt_clkdiv.clkDiv_inst.cnt[5] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\genblk2[8].wave_shpr.div.quo[14] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\genblk2[4].wave_shpr.div.quo[7] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\genblk2[1].wave_shpr.div.b1[17] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\genblk2[0].wave_shpr.div.quo[17] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(_00141_),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\genblk2[11].wave_shpr.div.quo[24] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(_01058_),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\genblk2[1].wave_shpr.div.quo[4] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(_00212_),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\genblk2[9].wave_shpr.div.quo[21] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\genblk2[1].wave_shpr.div.quo[19] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\genblk2[10].wave_shpr.div.quo[1] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_00810_),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\genblk2[4].wave_shpr.div.quo[0] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_00460_),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\genblk2[11].wave_shpr.div.b1[8] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\genblk2[7].wave_shpr.div.quo[7] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_00719_),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\genblk2[5].wave_shpr.div.quo[8] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\genblk2[11].wave_shpr.div.b1[15] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\genblk2[1].wave_shpr.div.b1[16] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\genblk2[1].wave_shpr.div.quo[18] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(_00225_),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\genblk2[11].wave_shpr.div.quo[20] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\sig_norm.acc_next[0] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(_00062_),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\genblk2[11].wave_shpr.div.quo[0] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_01034_),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\genblk2[10].wave_shpr.div.quo[9] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_00958_),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\genblk2[11].wave_shpr.div.quo[23] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_01057_),
    .X(net435));
 sky130_fd_sc_hd__buf_1 hold218 (.A(\genblk1[3].osc.clkdiv_C.cnt[17] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_00401_),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_01054_),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\genblk2[11].wave_shpr.div.quo[22] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_01056_),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\genblk2[10].wave_shpr.div.quo[19] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\genblk2[2].wave_shpr.div.quo[10] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_00302_),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\genblk2[11].wave_shpr.div.quo[12] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_01045_),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\genblk2[8].wave_shpr.div.quo[24] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\genblk2[10].wave_shpr.div.quo[24] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_00973_),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\genblk2[6].wave_shpr.div.quo[6] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\genblk2[1].wave_shpr.div.acc[24] ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\genblk2[2].wave_shpr.div.quo[6] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\genblk2[8].wave_shpr.div.quo[8] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\genblk2[3].wave_shpr.div.quo[18] ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_00393_),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\genblk2[5].wave_shpr.div.quo[12] ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\genblk2[0].wave_shpr.div.quo[23] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_00147_),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\genblk2[8].wave_shpr.div.acc[22] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\genblk2[2].wave_shpr.div.quo[13] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_00634_),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_00305_),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\genblk2[5].wave_shpr.div.quo[23] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\genblk2[1].wave_shpr.div.quo[8] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(_00215_),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\genblk2[1].wave_shpr.div.quo[16] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_00223_),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\genblk2[4].wave_shpr.div.quo[1] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(_00461_),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\genblk2[0].wave_shpr.div.quo[18] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\genblk2[11].wave_shpr.div.quo[10] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\genblk2[9].wave_shpr.div.quo[12] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_01044_),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\genblk2[8].wave_shpr.div.quo[10] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_00806_),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\genblk2[5].wave_shpr.div.quo[22] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\genblk2[4].wave_shpr.div.acc[21] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_00507_),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\genblk2[10].wave_shpr.div.quo[22] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_00972_),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\genblk2[0].wave_shpr.div.quo[22] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\genblk2[6].wave_shpr.div.quo[9] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_00878_),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\genblk2[9].wave_shpr.div.b1[13] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\genblk2[11].wave_shpr.div.quo[9] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\genblk2[2].wave_shpr.div.quo[14] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\genblk2[9].wave_shpr.div.quo[11] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\genblk2[8].wave_shpr.div.quo[12] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\genblk2[11].wave_shpr.div.quo[19] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\genblk2[7].wave_shpr.div.b1[14] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\genblk2[9].wave_shpr.div.quo[14] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\genblk2[6].wave_shpr.div.quo[18] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\genblk2[7].wave_shpr.div.quo[22] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\genblk2[5].wave_shpr.div.quo[21] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_00734_),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\genblk2[11].wave_shpr.div.quo[14] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\genblk2[3].wave_shpr.div.quo[23] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_00399_),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\genblk2[7].wave_shpr.div.quo[8] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\genblk1[5].osc.clkdiv_C.cnt[17] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_00569_),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\genblk2[0].wave_shpr.div.quo[13] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_00137_),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\sig_norm.b1[1] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_00565_),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\genblk2[6].wave_shpr.div.quo[14] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(_00641_),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\genblk2[5].wave_shpr.div.quo[11] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(_00555_),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\genblk2[8].wave_shpr.div.quo[16] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\genblk2[5].wave_shpr.div.quo[20] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\genblk2[11].wave_shpr.div.quo[21] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\genblk2[8].wave_shpr.div.quo[23] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\genblk2[8].wave_shpr.div.quo[11] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\genblk2[5].wave_shpr.div.quo[18] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\genblk2[10].wave_shpr.div.acc_next[0] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\genblk2[4].wave_shpr.div.quo[6] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\genblk2[11].wave_shpr.div.quo[18] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\genblk2[11].wave_shpr.div.quo[17] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\genblk2[1].wave_shpr.div.quo[14] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(_00222_),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\genblk2[9].wave_shpr.div.quo[18] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\genblk2[3].wave_shpr.div.quo[15] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\genblk2[6].wave_shpr.div.quo[8] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(_00636_),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\genblk2[1].wave_shpr.div.quo[9] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_00951_),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_00975_),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\genblk2[10].wave_shpr.div.quo[18] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\genblk2[1].wave_shpr.div.quo[13] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\genblk2[2].wave_shpr.div.quo[23] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\genblk2[10].wave_shpr.div.quo[13] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\genblk2[0].wave_shpr.div.quo[16] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\genblk2[6].wave_shpr.div.quo[7] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\genblk2[3].wave_shpr.div.acc[21] ),
    .X(net524));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold307 (.A(\genblk2[3].wave_shpr.div.quo[11] ),
    .X(net525));
 sky130_fd_sc_hd__buf_1 hold308 (.A(\genblk2[9].wave_shpr.div.quo[8] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\genblk2[7].wave_shpr.div.quo[20] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\genblk2[5].wave_shpr.div.quo[14] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(_00732_),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\genblk2[3].wave_shpr.div.quo[22] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\genblk2[9].wave_shpr.div.quo[17] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\genblk2[4].wave_shpr.div.quo[17] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_00476_),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\genblk2[9].wave_shpr.div.quo[20] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\genblk2[7].wave_shpr.div.quo[24] ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(_00735_),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\genblk2[10].wave_shpr.div.acc[24] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\genblk2[1].wave_shpr.div.quo[12] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_00558_),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\genblk2[3].wave_shpr.div.quo[9] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(_00384_),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\genblk2[7].wave_shpr.div.acc_next[0] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\genblk2[9].wave_shpr.div.quo[13] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\genblk2[7].wave_shpr.div.quo[21] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\genblk2[0].wave_shpr.div.quo[15] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(_00138_),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\genblk2[3].wave_shpr.div.quo[20] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(_00396_),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\genblk2[10].wave_shpr.div.quo[17] ),
    .X(net547));
 sky130_fd_sc_hd__buf_1 hold33 (.A(\genblk2[4].wave_shpr.div.quo[8] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\genblk2[7].wave_shpr.div.quo[16] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(_00728_),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\genblk2[7].wave_shpr.div.quo[15] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\genblk2[5].wave_shpr.div.quo[15] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\genblk2[1].wave_shpr.div.quo[17] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\genblk2[2].wave_shpr.div.quo[12] ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(_00303_),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\genblk2[10].wave_shpr.div.quo[5] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\genblk2[9].wave_shpr.div.acc[21] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\genblk2[9].wave_shpr.div.quo[10] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_00468_),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\genblk2[0].wave_shpr.div.quo[2] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(_00126_),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\genblk2[6].wave_shpr.div.acc[18] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\genblk2[3].wave_shpr.div.quo[24] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(_00400_),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\genblk2[7].wave_shpr.div.quo[1] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(_00713_),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\genblk2[9].wave_shpr.div.quo[23] ),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\genblk2[5].wave_shpr.div.acc[21] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\genblk2[6].wave_shpr.div.quo[20] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\genblk2[5].wave_shpr.div.quo[5] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_00648_),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\genblk2[0].wave_shpr.div.quo[10] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_00134_),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\genblk2[11].wave_shpr.div.quo[16] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\genblk2[5].wave_shpr.div.quo[10] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\genblk2[2].wave_shpr.div.quo[16] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\genblk2[2].wave_shpr.div.quo[9] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\genblk2[8].wave_shpr.div.quo[21] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\genblk2[11].wave_shpr.div.acc[18] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\genblk2[0].wave_shpr.div.b1[15] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_00549_),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\genblk2[0].wave_shpr.div.acc_next[0] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(_00148_),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\genblk2[2].wave_shpr.div.acc[18] ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(_00335_),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\genblk2[6].wave_shpr.div.quo[17] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\genblk2[10].wave_shpr.div.quo[12] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\genblk2[0].wave_shpr.div.quo[12] ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\genblk2[7].wave_shpr.div.quo[17] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\genblk2[9].wave_shpr.div.quo[4] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(_00870_),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\genblk2[4].wave_shpr.div.quo[18] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\genblk2[1].wave_shpr.div.acc_next[0] ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(_00232_),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\genblk2[10].wave_shpr.div.acc[18] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\genblk2[4].wave_shpr.div.acc[19] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\genblk1[0].osc.clkdiv_C.cnt[7] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\genblk2[8].wave_shpr.div.b1[4] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\genblk2[6].wave_shpr.div.quo[15] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\genblk2[6].wave_shpr.div.quo[16] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\genblk2[4].wave_shpr.div.quo[14] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(_00474_),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_00478_),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\genblk2[0].wave_shpr.div.quo[9] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\genblk2[0].wave_shpr.div.quo[11] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\genblk2[0].wave_shpr.div.quo[4] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(_00128_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\genblk2[4].wave_shpr.div.quo[11] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(_00470_),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\genblk2[0].wave_shpr.div.acc[18] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\genblk2[2].wave_shpr.div.acc[19] ),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(_00336_),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\genblk2[3].wave_shpr.div.quo[21] ),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\genblk2[1].wave_shpr.div.quo[20] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\genblk2[1].wave_shpr.div.quo[21] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\genblk2[6].wave_shpr.div.quo[22] ),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\genblk2[1].wave_shpr.div.quo[10] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\genblk2[8].wave_shpr.div.quo[15] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\sig_norm.acc[7] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\genblk2[7].wave_shpr.div.quo[14] ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\genblk2[3].wave_shpr.div.b1[9] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\genblk2[8].wave_shpr.div.acc[26] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\genblk2[6].wave_shpr.div.quo[21] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\genblk2[8].wave_shpr.div.quo[18] ),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_2 hold4 (.A(\modein.delay_in[0] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_00228_),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_00814_),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\genblk2[11].wave_shpr.div.acc[23] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\genblk2[6].wave_shpr.div.quo[13] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(_00640_),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\genblk2[6].wave_shpr.div.acc[19] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\genblk2[6].wave_shpr.div.quo[11] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(_00639_),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\genblk2[5].wave_shpr.div.b1[5] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\genblk2[4].wave_shpr.div.quo[20] ),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(_00480_),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\genblk2[2].wave_shpr.div.quo[24] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\genblk2[7].wave_shpr.div.acc[18] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\sig_norm.acc[1] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\genblk2[5].wave_shpr.div.acc[18] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\genblk2[3].wave_shpr.div.quo[10] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\genblk2[1].wave_shpr.div.quo[24] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(_00231_),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\genblk2[3].wave_shpr.div.quo[14] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(_00389_),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\genblk2[0].wave_shpr.div.quo[20] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\genblk2[4].wave_shpr.div.quo[13] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_00316_),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(_00472_),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\genblk2[2].wave_shpr.div.quo[22] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\genblk2[7].wave_shpr.div.quo[13] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\genblk2[11].wave_shpr.div.acc[19] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\PWM.counter[1] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\genblk2[4].wave_shpr.div.acc_next[0] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(_00484_),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\genblk2[1].wave_shpr.div.quo[11] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\genblk2[9].wave_shpr.div.acc[22] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(_00913_),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\genblk2[2].wave_shpr.div.quo[21] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\genblk2[2].wave_shpr.div.acc[20] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\genblk2[9].wave_shpr.div.quo[1] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_00867_),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\genblk2[10].wave_shpr.div.b1[5] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\genblk2[0].wave_shpr.div.quo[5] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\genblk2[0].wave_shpr.div.acc[23] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\genblk2[5].wave_shpr.div.acc[22] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\genblk2[0].wave_shpr.div.quo[1] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\genblk2[2].wave_shpr.div.quo[20] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\genblk2[3].wave_shpr.div.acc[18] ),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_00313_),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\genblk2[4].wave_shpr.div.quo[19] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\genblk2[6].wave_shpr.div.acc[23] ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\genblk2[8].wave_shpr.div.quo[20] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\genblk2[7].wave_shpr.div.quo[4] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(_00716_),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\sig_norm.acc[10] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\genblk2[1].wave_shpr.div.acc[18] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\genblk2[4].wave_shpr.div.quo[22] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(_00481_),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\genblk2[4].wave_shpr.div.b1[16] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\genblk2[8].wave_shpr.div.quo[17] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\genblk2[6].wave_shpr.div.quo[24] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\genblk2[9].wave_shpr.div.acc[18] ),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\genblk2[7].wave_shpr.div.quo[12] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\genblk2[6].wave_shpr.div.quo[2] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\genblk2[4].wave_shpr.div.quo[10] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(_00469_),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\genblk2[10].wave_shpr.div.b1[15] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\genblk2[4].wave_shpr.div.quo[12] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\genblk2[8].wave_shpr.div.quo[6] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\genblk2[8].wave_shpr.div.quo[19] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_00813_),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\sig_norm.acc[8] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\genblk2[7].wave_shpr.div.acc[21] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\genblk2[4].wave_shpr.div.quo[16] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(_00475_),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\genblk2[10].wave_shpr.div.quo[3] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(_00953_),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\genblk2[1].wave_shpr.div.quo[1] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(_00209_),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\genblk2[9].wave_shpr.div.quo[2] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(_00868_),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\genblk2[0].wave_shpr.div.quo[21] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\genblk2[0].wave_shpr.div.acc[19] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(_00168_),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\genblk2[8].wave_shpr.div.acc[20] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\genblk1[8].osc.clkdiv_C.cnt[17] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\genblk2[5].wave_shpr.div.b1[2] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\genblk2[7].wave_shpr.div.quo[2] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\genblk2[4].wave_shpr.div.acc[20] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\genblk1[10].osc.clkdiv_C.cnt[17] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\genblk2[2].wave_shpr.div.quo[4] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(_00296_),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_00145_),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\genblk2[4].wave_shpr.div.quo[23] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\genblk2[8].wave_shpr.div.acc[2] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\genblk2[9].wave_shpr.div.quo[3] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\genblk2[1].wave_shpr.div.quo[3] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\genblk2[0].wave_shpr.div.b1[17] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\genblk2[8].wave_shpr.div.b1[16] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\genblk2[8].wave_shpr.div.acc[23] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\genblk2[10].wave_shpr.div.acc[20] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\genblk2[7].wave_shpr.div.acc[22] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\genblk2[2].wave_shpr.div.acc[23] ),
    .X(net707));
 sky130_fd_sc_hd__buf_1 hold49 (.A(\genblk2[9].wave_shpr.div.quo[6] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\genblk2[5].wave_shpr.div.b1[6] ),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\genblk2[8].wave_shpr.div.quo[2] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\genblk2[3].wave_shpr.div.acc[22] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\genblk2[2].wave_shpr.div.i[2] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\genblk2[9].wave_shpr.div.quo[5] ),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\genblk2[9].wave_shpr.div.b1[16] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\genblk2[4].wave_shpr.div.quo[24] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\genblk2[0].wave_shpr.div.acc[0] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\genblk2[2].wave_shpr.div.quo[5] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\sig_norm.acc[9] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\genblk2[10].wave_shpr.div.quo[11] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_00872_),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(\genblk1[1].osc.clkdiv_C.cnt[0] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\genblk2[2].wave_shpr.div.quo[2] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\genblk2[6].wave_shpr.div.quo[4] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(_00632_),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\genblk2[8].wave_shpr.div.b1[14] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\genblk2[10].wave_shpr.div.quo[4] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\genblk2[10].wave_shpr.div.quo[2] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\genblk2[3].wave_shpr.div.i[2] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\genblk2[8].wave_shpr.div.i[2] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\genblk2[0].wave_shpr.div.b1[5] ),
    .X(net727));
 sky130_fd_sc_hd__buf_1 hold51 (.A(\genblk2[0].wave_shpr.div.quo[6] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\genblk2[0].wave_shpr.div.quo[3] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\genblk2[5].wave_shpr.div.quo[4] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\genblk2[3].wave_shpr.div.b1[16] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\genblk2[11].wave_shpr.div.quo[5] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\genblk2[4].wave_shpr.div.quo[3] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(_00463_),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(\genblk2[4].wave_shpr.div.i[2] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(_00514_),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\genblk2[7].wave_shpr.div.quo[10] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\genblk2[3].wave_shpr.div.quo[2] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_00130_),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(_00378_),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\genblk2[6].wave_shpr.div.i[2] ),
    .X(net739));
 sky130_fd_sc_hd__buf_1 hold522 (.A(\genblk2[10].wave_shpr.div.quo[0] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\genblk2[11].wave_shpr.div.i[2] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\genblk2[6].wave_shpr.div.quo[5] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\genblk2[8].wave_shpr.div.quo[0] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(_00796_),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\genblk2[5].wave_shpr.div.quo[3] ),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(\genblk2[9].wave_shpr.div.quo[0] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\genblk2[6].wave_shpr.div.b1[14] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\genblk2[6].wave_shpr.div.quo[3] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\genblk2[10].wave_shpr.div.i[2] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\genblk2[4].wave_shpr.div.quo[4] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(_00464_),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\genblk2[8].wave_shpr.div.quo[5] ),
    .X(net751));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold534 (.A(\genblk2[1].wave_shpr.div.acc[0] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(_00234_),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\genblk2[7].wave_shpr.div.quo[5] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\genblk2[1].wave_shpr.div.quo[2] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\genblk2[6].wave_shpr.div.quo[1] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\genblk2[1].wave_shpr.div.i[2] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_00631_),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(\genblk2[7].wave_shpr.div.b1[16] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\genblk2[10].wave_shpr.div.b1[14] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\modein.delay_in[1] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\genblk2[2].wave_shpr.div.b1[17] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(\genblk2[11].wave_shpr.div.acc[9] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\genblk2[4].wave_shpr.div.acc[26] ),
    .X(net763));
 sky130_fd_sc_hd__buf_1 hold546 (.A(\genblk2[1].wave_shpr.div.quo[0] ),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\sig_norm.i[2] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(_00028_),
    .X(net766));
 sky130_fd_sc_hd__buf_1 hold549 (.A(\genblk2[11].wave_shpr.div.quo[4] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\genblk2[0].wave_shpr.div.i[4] ),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(\genblk2[8].wave_shpr.div.b1[7] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\genblk2[11].wave_shpr.div.quo[1] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(\genblk2[5].wave_shpr.div.quo[6] ),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\genblk2[1].wave_shpr.div.quo[5] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\genblk2[5].wave_shpr.div.acc[9] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(_00579_),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(\genblk2[1].wave_shpr.div.acc[16] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\genblk2[0].wave_shpr.div.i[2] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(\genblk2[11].wave_shpr.div.quo[3] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\genblk2[4].wave_shpr.div.acc[25] ),
    .X(net777));
 sky130_fd_sc_hd__buf_1 hold56 (.A(\genblk2[8].wave_shpr.div.acc_next[0] ),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(\genblk2[4].wave_shpr.div.acc[12] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\genblk2[3].wave_shpr.div.quo[3] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(_00379_),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\genblk2[4].wave_shpr.div.quo[5] ),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\genblk2[2].wave_shpr.div.acc[1] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\genblk2[5].wave_shpr.div.i[3] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(\genblk2[4].wave_shpr.div.acc[15] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\genblk2[11].wave_shpr.div.acc[11] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(\genblk2[0].wave_shpr.div.acc[17] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\genblk2[4].wave_shpr.div.acc[23] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\genblk2[2].wave_shpr.div.quo[7] ),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(\genblk2[2].wave_shpr.div.acc[17] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\genblk2[9].wave_shpr.div.i[3] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(\genblk2[3].wave_shpr.div.acc[10] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\genblk2[3].wave_shpr.div.acc[11] ),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_2 hold574 (.A(\genblk2[6].wave_shpr.div.quo[0] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\genblk2[4].wave_shpr.div.quo[2] ),
    .X(net793));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold576 (.A(\genblk2[3].wave_shpr.div.quo[0] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\genblk2[8].wave_shpr.div.quo[4] ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(\genblk2[3].wave_shpr.div.acc[9] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\genblk2[7].wave_shpr.div.acc[10] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_00299_),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_00747_),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\genblk2[9].wave_shpr.div.acc[14] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(\genblk2[5].wave_shpr.div.b1[14] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\genblk2[7].wave_shpr.div.i[2] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(\genblk2[8].wave_shpr.div.acc[16] ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\genblk2[1].wave_shpr.div.acc[23] ),
    .X(net803));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold586 (.A(\genblk2[0].wave_shpr.div.quo[0] ),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\genblk2[7].wave_shpr.div.acc[14] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(\genblk2[6].wave_shpr.div.acc[9] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\genblk2[9].wave_shpr.div.acc[11] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\genblk2[0].wave_shpr.div.quo[8] ),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(\genblk2[7].wave_shpr.div.acc[13] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\genblk2[7].wave_shpr.div.acc[15] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\PWM.counter[5] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(_01165_),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\genblk2[2].wave_shpr.div.quo[1] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\genblk2[1].wave_shpr.div.acc[10] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(\genblk2[3].wave_shpr.div.quo[5] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(_00381_),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(\genblk2[11].wave_shpr.div.acc[10] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\genblk2[9].wave_shpr.div.i[4] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_00961_),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_00132_),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(\genblk2[6].wave_shpr.div.acc[15] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\genblk2[6].wave_shpr.div.acc[6] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(\genblk2[3].wave_shpr.div.quo[6] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\genblk2[0].wave_shpr.div.acc[26] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(\genblk2[7].wave_shpr.div.quo[0] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\genblk2[0].wave_shpr.div.acc[5] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(_00154_),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\genblk2[1].wave_shpr.div.acc[5] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(\genblk2[6].wave_shpr.div.acc[7] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\genblk2[1].wave_shpr.div.acc[8] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\sig_norm.i[3] ),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(\genblk2[5].wave_shpr.div.acc[17] ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\genblk2[1].wave_shpr.div.acc[4] ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(\genblk2[2].wave_shpr.div.acc[11] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\PWM.counter[2] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(_01160_),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\genblk2[8].wave_shpr.div.acc[13] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(\genblk2[5].wave_shpr.div.b1[16] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\genblk2[5].wave_shpr.div.acc[15] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(\genblk2[2].wave_shpr.div.acc[7] ),
    .X(net836));
 sky130_fd_sc_hd__buf_1 hold619 (.A(\genblk1[6].osc.clkdiv_C.cnt[0] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\genblk2[6].wave_shpr.div.i[4] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(\genblk2[6].wave_shpr.div.acc[12] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\genblk2[9].wave_shpr.div.acc[8] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(\genblk2[0].wave_shpr.div.acc[15] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\genblk2[11].wave_shpr.div.acc[6] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(\genblk2[4].wave_shpr.div.acc[4] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(_00489_),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\genblk2[10].wave_shpr.div.acc[11] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\genblk2[2].wave_shpr.div.acc[16] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(\genblk2[8].wave_shpr.div.acc[14] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\genblk2[1].wave_shpr.div.acc[9] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\genblk2[4].wave_shpr.div.i[4] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\genblk1[7].osc.clkdiv_C.cnt[17] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\genblk2[3].wave_shpr.div.quo[4] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\genblk2[4].wave_shpr.div.acc[14] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\genblk1[4].osc.clkdiv_C.cnt[17] ),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(\genblk2[7].wave_shpr.div.acc[12] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(_00749_),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(\genblk2[0].wave_shpr.div.acc[3] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\genblk2[5].wave_shpr.div.i[4] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(_04964_),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\genblk2[2].wave_shpr.div.acc[12] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\genblk2[2].wave_shpr.div.i[4] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\genblk2[10].wave_shpr.div.acc[13] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\genblk2[10].wave_shpr.div.acc[17] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(_00992_),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\genblk2[0].wave_shpr.div.b1[0] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(\genblk2[3].wave_shpr.div.acc[14] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\genblk2[5].wave_shpr.div.acc[6] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(\genblk2[8].wave_shpr.div.b1[0] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\genblk2[1].wave_shpr.div.acc[13] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(\genblk2[0].wave_shpr.div.acc[6] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\genblk2[6].wave_shpr.div.acc[8] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\genblk2[6].wave_shpr.div.acc_next[0] ),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(\genblk2[10].wave_shpr.div.acc[4] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(_00979_),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(\genblk2[10].wave_shpr.div.acc[16] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\genblk2[8].wave_shpr.div.quo[1] ),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(\genblk2[8].wave_shpr.div.acc[3] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\genblk2[7].wave_shpr.div.acc[23] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\genblk2[1].wave_shpr.div.acc[20] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\genblk2[11].wave_shpr.div.acc[12] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(\genblk2[11].wave_shpr.div.acc[8] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\genblk2[7].wave_shpr.div.acc[4] ),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_00653_),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(\genblk2[11].wave_shpr.div.acc[17] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\genblk2[5].wave_shpr.div.quo[1] ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(_00545_),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\genblk2[4].wave_shpr.div.acc[16] ),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(\genblk2[5].wave_shpr.div.quo[2] ),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\genblk2[6].wave_shpr.div.acc[13] ),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(\genblk2[9].wave_shpr.div.acc[10] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\genblk2[5].wave_shpr.div.acc[5] ),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(\genblk2[9].wave_shpr.div.acc[4] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\genblk2[2].wave_shpr.div.acc[6] ),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\genblk2[1].wave_shpr.div.i[4] ),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(\genblk2[5].wave_shpr.div.acc[4] ),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\genblk2[0].wave_shpr.div.acc[12] ),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(\genblk2[3].wave_shpr.div.acc[7] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\genblk2[4].wave_shpr.div.acc[8] ),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(\genblk2[9].wave_shpr.div.acc[23] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\genblk2[7].wave_shpr.div.acc[7] ),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(\genblk2[7].wave_shpr.div.acc[11] ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\genblk2[2].wave_shpr.div.acc[9] ),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(\genblk2[5].wave_shpr.div.acc[19] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\genblk2[11].wave_shpr.div.acc[15] ),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\PWM.final_sample_in[7] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\genblk2[8].wave_shpr.div.acc[5] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\genblk2[6].wave_shpr.div.acc[17] ),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\genblk2[6].wave_shpr.div.acc[11] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\genblk2[4].wave_shpr.div.acc[13] ),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(\genblk2[5].wave_shpr.div.acc[14] ),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\genblk2[2].wave_shpr.div.acc[8] ),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(\genblk2[3].wave_shpr.div.acc[19] ),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(\genblk2[1].wave_shpr.div.acc[15] ),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(\genblk2[10].wave_shpr.div.acc[23] ),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(\genblk2[6].wave_shpr.div.acc[5] ),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\PWM.next_pwm_out ),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(\genblk2[8].wave_shpr.div.acc[10] ),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\genblk2[8].wave_shpr.div.acc[12] ),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(\genblk2[5].wave_shpr.div.acc[2] ),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(_00571_),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\genblk2[9].wave_shpr.div.acc[15] ),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\genblk2[0].wave_shpr.div.acc[14] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(\genblk2[2].wave_shpr.div.acc_next[0] ),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(_00317_),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(\genblk2[7].wave_shpr.div.acc[9] ),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(\genblk2[8].wave_shpr.div.acc[11] ),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\modein.delay_octave_down_in[0] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\genblk2[11].wave_shpr.div.i[4] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(\genblk2[2].wave_shpr.div.acc[3] ),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\genblk2[2].wave_shpr.div.acc[5] ),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(\genblk2[0].wave_shpr.div.acc[13] ),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\genblk2[6].wave_shpr.div.acc[14] ),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(\genblk2[8].wave_shpr.div.acc[9] ),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(\genblk2[7].wave_shpr.div.acc[20] ),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(\genblk2[7].wave_shpr.div.acc[17] ),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\genblk2[5].wave_shpr.div.acc[16] ),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(\genblk2[4].wave_shpr.div.acc[17] ),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\genblk2[5].wave_shpr.div.acc[8] ),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\genblk2[10].wave_shpr.div.i[4] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(\genblk2[4].wave_shpr.div.acc[9] ),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\genblk2[10].wave_shpr.div.acc[7] ),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(\genblk2[3].wave_shpr.div.acc[15] ),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\genblk2[11].wave_shpr.div.acc[21] ),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(\genblk2[8].wave_shpr.div.acc[6] ),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\genblk2[0].wave_shpr.div.acc[22] ),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(\genblk2[0].wave_shpr.div.acc[10] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\genblk2[9].wave_shpr.div.acc[20] ),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(_00911_),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\genblk2[4].wave_shpr.div.acc[2] ),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\genblk2[9].wave_shpr.div.quo[9] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(\genblk2[9].wave_shpr.div.acc[6] ),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\sig_norm.i[0] ),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(_00026_),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\genblk2[3].wave_shpr.div.acc[6] ),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(\genblk2[3].wave_shpr.div.acc[12] ),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(_00413_),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(\genblk2[10].wave_shpr.div.acc[15] ),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\genblk2[10].wave_shpr.div.acc[14] ),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(\genblk2[8].wave_shpr.div.acc[24] ),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\genblk2[8].wave_shpr.div.acc[15] ),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_00875_),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(\genblk2[3].wave_shpr.div.acc[17] ),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\genblk2[11].wave_shpr.div.acc[13] ),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(\genblk2[8].wave_shpr.div.acc[7] ),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\genblk2[10].wave_shpr.div.acc[10] ),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(\genblk2[2].wave_shpr.div.acc[10] ),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\genblk2[2].wave_shpr.div.acc[13] ),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(\genblk2[10].wave_shpr.div.acc[8] ),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\genblk2[11].wave_shpr.div.acc[22] ),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(\genblk2[0].wave_shpr.div.acc[9] ),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\genblk2[10].wave_shpr.div.acc[12] ),
    .X(net957));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold74 (.A(\genblk2[1].wave_shpr.div.quo[6] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(\genblk2[11].wave_shpr.div.acc[5] ),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\genblk2[10].wave_shpr.div.b1[16] ),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(\genblk2[11].wave_shpr.div.acc[26] ),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\genblk2[5].wave_shpr.div.acc[3] ),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(\genblk2[2].wave_shpr.div.acc[26] ),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\genblk2[3].wave_shpr.div.acc[5] ),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(\genblk2[0].wave_shpr.div.acc[7] ),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\genblk2[1].wave_shpr.div.acc[3] ),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(\genblk2[3].wave_shpr.div.acc[8] ),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\genblk2[9].wave_shpr.div.acc[13] ),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_00214_),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(\genblk2[2].wave_shpr.div.acc[22] ),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\genblk2[10].wave_shpr.div.acc[3] ),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(\genblk2[4].wave_shpr.div.acc[5] ),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\genblk2[4].wave_shpr.div.acc[7] ),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(_00492_),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(\genblk2[1].wave_shpr.div.acc[17] ),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(\genblk2[9].wave_shpr.div.acc[9] ),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\genblk2[2].wave_shpr.div.acc[4] ),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(\genblk2[3].wave_shpr.div.acc[2] ),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\genblk2[10].wave_shpr.div.acc[5] ),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\genblk2[5].wave_shpr.div.quo[13] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(\genblk2[8].wave_shpr.div.acc[8] ),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\genblk2[3].wave_shpr.div.acc[4] ),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(\genblk2[8].wave_shpr.div.acc[4] ),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\genblk2[5].wave_shpr.div.acc[13] ),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(\genblk2[5].wave_shpr.div.acc[20] ),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\genblk2[1].wave_shpr.div.acc[19] ),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(\genblk2[9].wave_shpr.div.acc[7] ),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(\genblk2[11].wave_shpr.div.acc[4] ),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(\genblk2[6].wave_shpr.div.acc[4] ),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\genblk2[9].wave_shpr.div.acc[17] ),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_00557_),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(\genblk2[7].wave_shpr.div.acc[6] ),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\genblk2[10].wave_shpr.div.acc[2] ),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(\genblk2[1].wave_shpr.div.acc[2] ),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\genblk2[8].wave_shpr.div.acc[17] ),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(\genblk2[7].wave_shpr.div.acc[3] ),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\genblk2[11].wave_shpr.div.acc[14] ),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(_01073_),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\genblk2[1].wave_shpr.div.acc[7] ),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(\PWM.counter[3] ),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\genblk2[11].wave_shpr.div.acc[7] ),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\genblk2[3].wave_shpr.div.quo[19] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(\genblk2[4].wave_shpr.div.acc[6] ),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\genblk2[9].wave_shpr.div.acc[5] ),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(\genblk2[3].wave_shpr.div.acc[23] ),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\genblk2[6].wave_shpr.div.acc[21] ),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(\genblk2[2].wave_shpr.div.acc[14] ),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\genblk2[6].wave_shpr.div.acc[10] ),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(\genblk2[0].wave_shpr.div.acc[11] ),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\genblk2[8].wave_shpr.div.b1[13] ),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(\genblk2[9].wave_shpr.div.acc[3] ),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\genblk2[11].wave_shpr.div.b1[0] ),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_00395_),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(\genblk2[4].wave_shpr.div.acc[11] ),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\genblk2[7].wave_shpr.div.acc[8] ),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(\genblk2[7].wave_shpr.div.acc[16] ),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(_00753_),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(\genblk2[5].wave_shpr.div.acc[23] ),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\genblk2[7].wave_shpr.div.acc[2] ),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(\genblk2[5].wave_shpr.div.acc[12] ),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\genblk2[6].wave_shpr.div.acc[3] ),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(\genblk2[3].wave_shpr.div.acc[16] ),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(\genblk2[3].wave_shpr.div.acc[13] ),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\genblk2[9].wave_shpr.div.quo[22] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\genblk2[0].wave_shpr.div.quo[19] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(\genblk2[8].wave_shpr.div.acc[21] ),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(\genblk2[1].wave_shpr.div.acc[14] ),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(\genblk2[11].wave_shpr.div.acc[3] ),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\genblk2[3].wave_shpr.div.acc[25] ),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(\genblk2[9].wave_shpr.div.acc[2] ),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\genblk2[9].wave_shpr.div.acc[19] ),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(\genblk2[4].wave_shpr.div.acc[10] ),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\genblk2[2].wave_shpr.div.b1[16] ),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(\genblk2[9].wave_shpr.div.acc[24] ),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\sig_norm.acc[5] ),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_00143_),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(_00043_),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\genblk2[7].wave_shpr.div.acc[24] ),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(\genblk2[7].wave_shpr.div.acc[5] ),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\genblk2[6].wave_shpr.div.acc[22] ),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(\genblk2[0].wave_shpr.div.acc[21] ),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\genblk2[0].wave_shpr.div.acc[4] ),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(\genblk2[2].wave_shpr.div.acc[21] ),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\genblk2[10].wave_shpr.div.acc[9] ),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(\genblk2[2].wave_shpr.div.acc[15] ),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\genblk2[5].wave_shpr.div.acc[7] ),
    .X(net1037));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold82 (.A(\genblk2[2].wave_shpr.div.quo[8] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(\genblk2[5].wave_shpr.div.acc[24] ),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\genblk2[9].wave_shpr.div.i[1] ),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(_00072_),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\genblk2[5].wave_shpr.div.acc[25] ),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(\genblk2[9].wave_shpr.div.b1[9] ),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\genblk2[6].wave_shpr.div.acc[26] ),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(\genblk2[11].wave_shpr.div.acc[1] ),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\genblk2[9].wave_shpr.div.acc[25] ),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(\genblk2[9].wave_shpr.div.acc[12] ),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(\genblk2[2].wave_shpr.div.b1[2] ),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_00300_),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(\genblk2[7].wave_shpr.div.acc[19] ),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(\genblk2[0].wave_shpr.div.acc[8] ),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(\genblk2[0].wave_shpr.div.acc[16] ),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\genblk1[2].osc.clkdiv_C.cnt[0] ),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(\genblk2[8].wave_shpr.div.acc[25] ),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\genblk2[7].wave_shpr.div.acc[25] ),
    .X(net1053));
 sky130_fd_sc_hd__buf_1 hold836 (.A(\genblk2[2].wave_shpr.div.quo[0] ),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(\genblk2[3].wave_shpr.div.acc[20] ),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(\genblk2[5].wave_shpr.div.quo[0] ),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(\genblk2[3].wave_shpr.div.acc[3] ),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\genblk2[7].wave_shpr.div.quo[9] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(\genblk1[7].osc.clkdiv_C.cnt[0] ),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(\genblk2[9].wave_shpr.div.acc[1] ),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(\genblk2[9].wave_shpr.div.acc[16] ),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\genblk2[5].wave_shpr.div.acc[11] ),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(\genblk2[5].wave_shpr.div.acc[1] ),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(\genblk1[6].osc.clkdiv_C.cnt[17] ),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(\genblk2[3].wave_shpr.div.acc[24] ),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(\sig_norm.acc[3] ),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(\genblk2[0].wave_shpr.div.acc[1] ),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(\genblk2[3].wave_shpr.div.acc[1] ),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(_00721_),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(\genblk2[4].wave_shpr.div.acc[3] ),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(\sig_norm.acc[2] ),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(\genblk2[7].wave_shpr.div.acc[1] ),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\genblk2[4].wave_shpr.div.b1[0] ),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(\genblk1[5].osc.clkdiv_C.cnt[7] ),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(\sig_norm.b1[2] ),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(\genblk2[4].wave_shpr.div.acc[18] ),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(\genblk2[4].wave_shpr.div.b1[2] ),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(\genblk2[6].wave_shpr.div.acc[25] ),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(\genblk1[3].osc.clkdiv_C.cnt[4] ),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\genblk2[9].wave_shpr.div.quo[15] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(\genblk2[11].wave_shpr.div.acc[25] ),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(\genblk2[3].wave_shpr.div.i[1] ),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(\genblk1[10].osc.clkdiv_C.cnt[0] ),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(\genblk2[10].wave_shpr.div.acc[26] ),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(\genblk2[0].wave_shpr.div.acc[25] ),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(\sig_norm.quo[0] ),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(\genblk2[0].wave_shpr.div.b1[11] ),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(\genblk2[9].wave_shpr.div.quo[7] ),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(\genblk2[11].wave_shpr.div.b1[16] ),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(\genblk2[10].wave_shpr.div.acc[21] ),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_00881_),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(\sig_norm.b1[3] ),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(\genblk1[0].osc.clkdiv_C.cnt[0] ),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(\genblk2[10].wave_shpr.div.i[1] ),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(\genblk2[1].wave_shpr.div.i[1] ),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(\genblk1[8].osc.clkdiv_C.cnt[0] ),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(\genblk2[6].wave_shpr.div.acc[16] ),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(\genblk2[2].wave_shpr.div.acc[25] ),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(\genblk1[3].osc.clkdiv_C.cnt[7] ),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(\genblk2[6].wave_shpr.div.b1[16] ),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(\genblk2[5].wave_shpr.div.b1[7] ),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\genblk2[9].wave_shpr.div.quo[24] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(\genblk2[8].wave_shpr.div.i[1] ),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(\genblk2[3].wave_shpr.div.b1[5] ),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(\genblk2[4].wave_shpr.div.b1[1] ),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\genblk1[3].osc.clkdiv_C.cnt[0] ),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(\PWM.final_in[2] ),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\PWM.final_in[1] ),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(\genblk1[6].osc.clkdiv_C.cnt[14] ),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(\genblk1[5].osc.clkdiv_C.cnt[4] ),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(\genblk2[0].wave_shpr.div.i[1] ),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(\genblk2[1].wave_shpr.div.acc[26] ),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_00890_),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(\genblk2[4].wave_shpr.div.i[1] ),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(\genblk2[1].wave_shpr.div.acc[21] ),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(\genblk2[2].wave_shpr.div.i[1] ),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(\PWM.final_sample_in[0] ),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(_02252_),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(\genblk2[7].wave_shpr.div.i[1] ),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(\genblk2[8].wave_shpr.div.acc[19] ),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(\genblk1[5].osc.clkdiv_C.cnt[15] ),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(\genblk2[8].wave_shpr.div.acc[1] ),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(\genblk2[5].wave_shpr.div.i[1] ),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_00888_),
    .X(net227));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold90 (.A(\genblk2[5].wave_shpr.div.quo[7] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(\genblk2[10].wave_shpr.div.acc[1] ),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(\genblk1[10].osc.clkdiv_C.cnt[12] ),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(\genblk1[5].osc.clkdiv_C.cnt[0] ),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(\genblk2[1].wave_shpr.div.b1[11] ),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(\genblk2[6].wave_shpr.div.acc[1] ),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(\genblk2[2].wave_shpr.div.i[3] ),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(\genblk2[11].wave_shpr.div.i[1] ),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(\genblk2[11].wave_shpr.div.acc[16] ),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(\sig_norm.quo[1] ),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(\genblk2[11].wave_shpr.div.acc[2] ),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_00551_),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(\PWM.final_in[7] ),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(\genblk2[4].wave_shpr.div.acc[1] ),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(\genblk2[6].wave_shpr.div.i[1] ),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(\sig_norm.acc[0] ),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(\PWM.final_in[6] ),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(\genblk1[0].osc.clkdiv_C.cnt[4] ),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(\PWM.final_in[0] ),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(\genblk2[10].wave_shpr.div.acc[19] ),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(\genblk1[9].osc.clkdiv_C.cnt[0] ),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(\genblk2[2].wave_shpr.div.acc[2] ),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\genblk2[5].wave_shpr.div.quo[9] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(\genblk2[6].wave_shpr.div.acc[20] ),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\genblk2[0].wave_shpr.div.acc[2] ),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(\genblk2[7].wave_shpr.div.b1[1] ),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(\sig_norm.acc[11] ),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(\PWM.final_sample_in[7] ),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\genblk1[10].osc.clkdiv_C.cnt[15] ),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(\genblk2[4].wave_shpr.div.acc[24] ),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\genblk1[3].osc.clkdiv_C.cnt[9] ),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(\genblk1[6].osc.clkdiv_C.cnt[13] ),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\genblk2[8].wave_shpr.div.b1[12] ),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_00553_),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(\genblk2[3].wave_shpr.div.i[3] ),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\genblk2[9].wave_shpr.div.i[2] ),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(\PWM.final_in[4] ),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(_03682_),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(\genblk2[3].wave_shpr.div.b1[13] ),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\genblk2[10].wave_shpr.div.i[3] ),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(\genblk2[5].wave_shpr.div.i[2] ),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(\sig_norm.acc[6] ),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(\sig_norm.quo[9] ),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(\PWM.final_sample_in[6] ),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\genblk2[8].wave_shpr.div.quo[13] ),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(\genblk2[0].wave_shpr.div.i[3] ),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(\genblk1[2].osc.clkdiv_C.cnt[10] ),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(\genblk2[4].wave_shpr.div.i[3] ),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(\sig_norm.b1[0] ),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(\genblk1[8].osc.clkdiv_C.cnt[4] ),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(\genblk2[11].wave_shpr.div.i[3] ),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(\genblk2[8].wave_shpr.div.i[3] ),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(\genblk2[6].wave_shpr.div.acc[2] ),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(\genblk1[2].osc.clkdiv_C.cnt[13] ),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(\genblk1[2].osc.clkdiv_C.cnt[15] ),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\genblk2[6].wave_shpr.div.quo[19] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(\PWM.final_in[5] ),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(_02257_),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(\sig_norm.quo[4] ),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(\genblk2[10].wave_shpr.div.b1[2] ),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(\PWM.final_in[3] ),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(\genblk2[10].wave_shpr.div.b1[6] ),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(\genblk2[1].wave_shpr.div.i[3] ),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(\genblk2[0].wave_shpr.div.acc[20] ),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(\sig_norm.quo[2] ),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(\genblk2[6].wave_shpr.div.i[3] ),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_00647_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(\genblk2[4].wave_shpr.div.b1[6] ),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(\smpl_rt_clkdiv.clkDiv_inst.cnt[6] ),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(\genblk1[6].osc.clkdiv_C.cnt[10] ),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(\genblk2[7].wave_shpr.div.i[3] ),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(\genblk1[8].osc.clkdiv_C.cnt[13] ),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(\genblk1[10].osc.clkdiv_C.cnt[8] ),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(\genblk2[0].wave_shpr.div.b1[10] ),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(\genblk1[8].osc.clkdiv_C.cnt[7] ),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(\genblk2[4].wave_shpr.div.b1[9] ),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(\genblk2[9].wave_shpr.div.b1[6] ),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\genblk2[2].wave_shpr.div.quo[15] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(\genblk2[4].wave_shpr.div.b1[4] ),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(\genblk1[7].osc.clkdiv_C.cnt[12] ),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(\genblk2[3].wave_shpr.div.b1[17] ),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(\genblk2[8].wave_shpr.div.b1[17] ),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(\genblk2[4].wave_shpr.div.b1[11] ),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(\genblk1[3].osc.clkdiv_C.cnt[12] ),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(\genblk1[9].osc.clkdiv_C.cnt[17] ),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(\genblk1[3].osc.clkdiv_C.cnt[14] ),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(\genblk1[0].osc.clkdiv_C.cnt[16] ),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(\genblk2[2].wave_shpr.div.quo[6] ),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_00307_),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(_04222_),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(\genblk2[10].wave_shpr.div.b1[12] ),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(\genblk2[7].wave_shpr.div.b1[4] ),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(\genblk2[7].wave_shpr.div.b1[8] ),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(\genblk2[7].wave_shpr.div.b1[6] ),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(\genblk2[11].wave_shpr.div.acc[20] ),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(\genblk2[11].wave_shpr.div.b1[10] ),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(\genblk2[4].wave_shpr.div.b1[12] ),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(\genblk2[4].wave_shpr.div.b1[8] ),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(\genblk1[2].osc.clkdiv_C.cnt[14] ),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\genblk2[7].wave_shpr.div.quo[6] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(\genblk2[9].wave_shpr.div.b1[5] ),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(\genblk2[9].wave_shpr.div.acc[0] ),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(_00891_),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(\genblk2[6].wave_shpr.div.b1[7] ),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(\genblk2[5].wave_shpr.div.b1[3] ),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(\genblk1[2].osc.clkdiv_C.cnt[11] ),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(\genblk2[8].wave_shpr.div.b1[3] ),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(\genblk2[7].wave_shpr.div.fin_quo[7] ),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(_05230_),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(\genblk2[11].wave_shpr.div.b1[9] ),
    .X(net1217));
 sky130_fd_sc_hd__buf_2 input1 (.A(pb[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(pb[4]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(pb[5]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(pb[6]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(pb[7]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(pb[8]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(pb[9]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_8 input16 (.A(reset),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(pb[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(pb[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(pb[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(pb[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(pb[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(pb[1]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(pb[2]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(pb[3]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 max_cap1 (.A(_05138_),
    .X(net1350));
 sky130_fd_sc_hd__buf_1 max_cap2 (.A(_04335_),
    .X(net1351));
 sky130_fd_sc_hd__buf_1 max_cap21 (.A(net1350),
    .X(net21));
 sky130_fd_sc_hd__buf_1 max_cap22 (.A(net1351),
    .X(net22));
 sky130_fd_sc_hd__buf_1 max_cap23 (.A(net1352),
    .X(net23));
 sky130_fd_sc_hd__buf_1 max_cap24 (.A(net1353),
    .X(net24));
 sky130_fd_sc_hd__buf_1 max_cap26 (.A(_03602_),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap29 (.A(_01372_),
    .X(net29));
 sky130_fd_sc_hd__buf_1 max_cap3 (.A(_03923_),
    .X(net1352));
 sky130_fd_sc_hd__buf_4 max_cap34 (.A(_01794_),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 max_cap36 (.A(_01423_),
    .X(net36));
 sky130_fd_sc_hd__buf_4 max_cap37 (.A(_01320_),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 max_cap4 (.A(net1354),
    .X(net1353));
 sky130_fd_sc_hd__clkbuf_1 max_cap6 (.A(_01692_),
    .X(net1355));
 sky130_fd_sc_hd__buf_1 max_cap7 (.A(_01760_),
    .X(net1356));
 sky130_fd_sc_hd__clkbuf_4 output17 (.A(net17),
    .X(mode_out[0]));
 sky130_fd_sc_hd__clkbuf_4 output18 (.A(net18),
    .X(mode_out[1]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(sigout));
 sky130_fd_sc_hd__buf_1 wire20 (.A(_06088_),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 wire25 (.A(_03112_),
    .X(net25));
 sky130_fd_sc_hd__buf_1 wire27 (.A(_01692_),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire28 (.A(net1356),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 wire30 (.A(_02635_),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 wire31 (.A(_02508_),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 wire32 (.A(_02302_),
    .X(net32));
 sky130_fd_sc_hd__buf_2 wire33 (.A(_02348_),
    .X(net33));
 sky130_fd_sc_hd__buf_2 wire35 (.A(_01239_),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 wire5 (.A(_02589_),
    .X(net1354));
endmodule

