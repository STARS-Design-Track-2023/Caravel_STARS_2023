// This is the unpowered netlist.
module calculator (blue,
    clk,
    nrst,
    red,
    pb,
    ss);
 output blue;
 input clk;
 input nrst;
 output red;
 input [9:0] pb;
 output [13:0] ss;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \u1.keycode[0] ;
 wire \u1.keycode[1] ;
 wire \u1.keycode[2] ;
 wire \u1.keycode[3] ;
 wire \u1.keycode[4] ;
 wire \u1.keycode[5] ;
 wire \u1.keycode[6] ;
 wire \u1.keycode[7] ;
 wire \u1.keycode[8] ;
 wire \u1.keypad_async[0] ;
 wire \u1.keypad_async[1] ;
 wire \u1.keypad_i[0] ;
 wire \u1.keypad_i[1] ;
 wire \u1.keypad_sync[0] ;
 wire \u1.keypad_sync[1] ;
 wire \u1.s_e_detect_w.i_signal ;
 wire \u1.s_e_detect_w.p_signal ;
 wire \u1.s_e_detect_w.s_signal ;
 wire \u1.state[0] ;
 wire \u1.state[10] ;
 wire \u1.state[11] ;
 wire \u1.state[12] ;
 wire \u1.state[13] ;
 wire \u1.state[14] ;
 wire \u1.state[1] ;
 wire \u1.state[2] ;
 wire \u1.state[3] ;
 wire \u1.state[4] ;
 wire \u1.state[6] ;
 wire \u1.state[7] ;
 wire \u1.state[8] ;
 wire \u1.state[9] ;
 wire \u1.store_dig ;
 wire \u3.keypad_13[0] ;
 wire \u3.keypad_13[1] ;
 wire \u3.keypad_async[0] ;
 wire \u3.keypad_async[1] ;
 wire \u3.keypad_sync[0] ;
 wire \u3.keypad_sync[1] ;
 wire \u3.out[1] ;
 wire \u4.op1[0] ;
 wire \u4.op1[1] ;
 wire \u4.op1[2] ;
 wire \u4.op1[3] ;
 wire \u4.op1[4] ;
 wire \u4.op1[5] ;
 wire \u4.op1[6] ;
 wire \u4.op1[7] ;
 wire \u4.op1[8] ;
 wire \u4.result_ready ;
 wire \u4.ssdec[0] ;
 wire \u4.ssdec[1] ;
 wire \u4.ssdec[2] ;
 wire \u4.ssdec[3] ;
 wire \u4.ssdec[4] ;
 wire \u4.ssdec[5] ;
 wire \u4.ssdec[6] ;
 wire \u4.ssdec[7] ;
 wire \u5.reg1[0] ;
 wire \u5.reg1[1] ;
 wire \u5.reg1[2] ;
 wire \u5.reg1[3] ;
 wire \u5.reg1[4] ;
 wire \u5.reg1[5] ;
 wire \u5.reg1[6] ;
 wire \u5.reg1[7] ;
 wire \u5.reg1[8] ;
 wire \u5.reg2[0] ;
 wire \u5.reg2[1] ;
 wire \u5.reg2[2] ;
 wire \u5.reg2[3] ;
 wire \u5.reg2[4] ;
 wire \u5.reg2[5] ;
 wire \u5.reg2[6] ;
 wire \u5.reg2[7] ;
 wire \u5.reg2[8] ;
 wire \u5.reg3[0] ;
 wire \u5.reg3[1] ;
 wire \u5.reg3[2] ;
 wire \u5.reg3[3] ;
 wire \u5.reg3[4] ;
 wire \u5.reg3[5] ;
 wire \u5.reg3[6] ;
 wire \u5.reg3[7] ;
 wire \u5.reg3[8] ;
 wire \u5.reg4[0] ;
 wire \u5.reg4[1] ;
 wire \u5.reg4[2] ;
 wire \u5.reg4[3] ;
 wire \u5.reg4[4] ;
 wire \u5.reg4[5] ;
 wire \u5.reg4[6] ;
 wire \u5.reg4[7] ;
 wire \u5.reg4[8] ;
 wire \u5.reg_num[0] ;
 wire \u5.reg_num[1] ;
 wire \u5.reg_num[2] ;
 wire \u5.reg_val[0] ;
 wire \u5.reg_val[1] ;
 wire \u5.reg_val[2] ;
 wire \u5.reg_val[3] ;
 wire \u5.reg_val[4] ;
 wire \u5.reg_val[5] ;
 wire \u5.reg_val[6] ;
 wire \u5.reg_val[7] ;
 wire \u5.reg_val[8] ;
 wire \u6.next_reg_num[0] ;
 wire \u6.next_reg_num[1] ;
 wire \u6.next_reg_num[2] ;
 wire \u6.reg_async[0] ;
 wire \u6.reg_async[1] ;
 wire \u6.reg_async[2] ;
 wire \u6.reg_async[3] ;
 wire \u6.reg_i[0] ;
 wire \u6.reg_i[1] ;
 wire \u6.reg_i[2] ;
 wire \u6.reg_i[3] ;
 wire \u6.reg_sync[0] ;
 wire \u6.reg_sync[1] ;
 wire \u6.reg_sync[2] ;
 wire \u6.reg_sync[3] ;
 wire \u7.assign_op1 ;
 wire \u7.assign_op2 ;
 wire \u7.s_e_detect.i_signal ;
 wire \u7.s_e_detect.p_signal ;
 wire \u7.s_e_detect.s_signal ;
 wire \u7.state[0] ;
 wire \u7.state[4] ;
 wire \u7.state[5] ;
 wire \u7.state[6] ;
 wire \u8.b_assign_op1 ;
 wire \u8.b_assign_op2 ;
 wire \u8.buff_opcode[1] ;
 wire \u8.new_op1[0] ;
 wire \u8.new_op1[1] ;
 wire \u8.new_op1[2] ;
 wire \u8.new_op1[3] ;
 wire \u8.new_op1[8] ;
 wire \u8.op1[4] ;
 wire \u8.op1[5] ;
 wire \u8.op1[6] ;
 wire \u8.op1[7] ;
 wire \u8.op2[0] ;
 wire \u8.op2[1] ;
 wire \u8.op2[2] ;
 wire \u8.op2[3] ;
 wire \u8.op2[4] ;
 wire \u8.op2[5] ;
 wire \u8.op2[6] ;
 wire \u8.op2[7] ;
 wire \u8.op2[8] ;

 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_92 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__or2b_1 _0469_ (.A(\u7.s_e_detect.p_signal ),
    .B_N(\u7.s_e_detect.s_signal ),
    .X(_0113_));
 sky130_fd_sc_hd__a21o_1 _0470_ (.A1(net67),
    .A2(_0113_),
    .B1(\u4.result_ready ),
    .X(_0011_));
 sky130_fd_sc_hd__or2b_1 _0471_ (.A(\u3.keypad_sync[1] ),
    .B_N(\u3.keypad_sync[0] ),
    .X(_0114_));
 sky130_fd_sc_hd__or2b_1 _0472_ (.A(\u3.keypad_sync[0] ),
    .B_N(\u3.keypad_sync[1] ),
    .X(_0115_));
 sky130_fd_sc_hd__a211o_1 _0473_ (.A1(_0114_),
    .A2(_0115_),
    .B1(\u3.keypad_13[1] ),
    .C1(\u3.keypad_13[0] ),
    .X(_0116_));
 sky130_fd_sc_hd__or3_1 _0474_ (.A(\u6.reg_i[1] ),
    .B(\u6.reg_i[0] ),
    .C(\u6.reg_i[3] ),
    .X(_0117_));
 sky130_fd_sc_hd__or4_1 _0475_ (.A(\u6.reg_sync[1] ),
    .B(\u6.reg_sync[0] ),
    .C(\u6.reg_sync[3] ),
    .D(\u6.reg_sync[2] ),
    .X(_0118_));
 sky130_fd_sc_hd__or3b_1 _0476_ (.A(\u6.reg_i[2] ),
    .B(_0117_),
    .C_N(_0118_),
    .X(_0119_));
 sky130_fd_sc_hd__clkbuf_2 _0477_ (.A(_0119_),
    .X(_0120_));
 sky130_fd_sc_hd__buf_6 _0478_ (.A(\u1.store_dig ),
    .X(_0121_));
 sky130_fd_sc_hd__a31o_1 _0479_ (.A1(net71),
    .A2(_0116_),
    .A3(_0120_),
    .B1(_0121_),
    .X(_0007_));
 sky130_fd_sc_hd__or2b_1 _0480_ (.A(\u1.s_e_detect_w.p_signal ),
    .B_N(\u1.s_e_detect_w.s_signal ),
    .X(_0122_));
 sky130_fd_sc_hd__a22o_1 _0481_ (.A1(net5),
    .A2(\u1.state[7] ),
    .B1(net69),
    .B2(_0122_),
    .X(_0006_));
 sky130_fd_sc_hd__or3_1 _0482_ (.A(\u5.reg_num[0] ),
    .B(\u5.reg_num[1] ),
    .C(\u5.reg_num[2] ),
    .X(_0123_));
 sky130_fd_sc_hd__and2_1 _0483_ (.A(\u7.state[6] ),
    .B(_0123_),
    .X(_0124_));
 sky130_fd_sc_hd__clkbuf_1 _0484_ (.A(_0124_),
    .X(_0003_));
 sky130_fd_sc_hd__inv_2 _0485_ (.A(\u1.state[0] ),
    .Y(_0125_));
 sky130_fd_sc_hd__nor2_1 _0486_ (.A(\u1.keypad_sync[0] ),
    .B(\u1.keypad_sync[1] ),
    .Y(_0126_));
 sky130_fd_sc_hd__or3_1 _0487_ (.A(\u1.keypad_i[1] ),
    .B(\u1.keypad_i[0] ),
    .C(_0126_),
    .X(_0127_));
 sky130_fd_sc_hd__clkbuf_4 _0488_ (.A(_0127_),
    .X(_0128_));
 sky130_fd_sc_hd__a2bb2o_1 _0489_ (.A1_N(_0125_),
    .A2_N(_0122_),
    .B1(_0128_),
    .B2(net66),
    .X(_0010_));
 sky130_fd_sc_hd__or3_1 _0490_ (.A(\u3.keypad_13[1] ),
    .B(net75),
    .C(_0115_),
    .X(_0129_));
 sky130_fd_sc_hd__inv_2 _0491_ (.A(net76),
    .Y(\u3.out[1] ));
 sky130_fd_sc_hd__and2_1 _0492_ (.A(\u7.state[4] ),
    .B(_0123_),
    .X(_0130_));
 sky130_fd_sc_hd__buf_1 _0493_ (.A(_0130_),
    .X(_0004_));
 sky130_fd_sc_hd__a211oi_1 _0494_ (.A1(_0114_),
    .A2(_0115_),
    .B1(\u3.keypad_13[1] ),
    .C1(\u3.keypad_13[0] ),
    .Y(_0131_));
 sky130_fd_sc_hd__and2_1 _0495_ (.A(net59),
    .B(_0131_),
    .X(_0132_));
 sky130_fd_sc_hd__clkbuf_1 _0496_ (.A(_0132_),
    .X(_0005_));
 sky130_fd_sc_hd__a21o_1 _0497_ (.A1(net59),
    .A2(_0116_),
    .B1(net47),
    .X(_0013_));
 sky130_fd_sc_hd__nor2_1 _0498_ (.A(\u5.reg_num[0] ),
    .B(\u5.reg_num[1] ),
    .Y(_0133_));
 sky130_fd_sc_hd__and2b_1 _0499_ (.A_N(\u5.reg_num[2] ),
    .B(_0133_),
    .X(_0134_));
 sky130_fd_sc_hd__and3b_1 _0500_ (.A_N(\u7.s_e_detect.p_signal ),
    .B(\u7.s_e_detect.s_signal ),
    .C(\u7.state[0] ),
    .X(_0135_));
 sky130_fd_sc_hd__a21o_1 _0501_ (.A1(net64),
    .A2(_0134_),
    .B1(_0135_),
    .X(_0012_));
 sky130_fd_sc_hd__a21o_1 _0502_ (.A1(net60),
    .A2(_0134_),
    .B1(net48),
    .X(_0014_));
 sky130_fd_sc_hd__inv_2 _0503_ (.A(net5),
    .Y(_0136_));
 sky130_fd_sc_hd__a21o_1 _0504_ (.A1(_0136_),
    .A2(\u1.state[7] ),
    .B1(\u1.state[8] ),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _0505_ (.A0(_0137_),
    .A1(\u1.state[4] ),
    .S(_0128_),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_1 _0506_ (.A(_0138_),
    .X(_0008_));
 sky130_fd_sc_hd__a311o_1 _0507_ (.A1(_0136_),
    .A2(\u1.state[7] ),
    .A3(_0128_),
    .B1(net61),
    .C1(\u1.state[3] ),
    .X(_0009_));
 sky130_fd_sc_hd__or2_1 _0508_ (.A(\u4.ssdec[1] ),
    .B(\u4.ssdec[0] ),
    .X(_0139_));
 sky130_fd_sc_hd__inv_2 _0509_ (.A(\u4.ssdec[1] ),
    .Y(_0140_));
 sky130_fd_sc_hd__a21oi_1 _0510_ (.A1(_0140_),
    .A2(\u4.ssdec[0] ),
    .B1(\u4.ssdec[2] ),
    .Y(_0141_));
 sky130_fd_sc_hd__a21oi_1 _0511_ (.A1(\u4.ssdec[2] ),
    .A2(_0139_),
    .B1(_0141_),
    .Y(_0142_));
 sky130_fd_sc_hd__nor2_1 _0512_ (.A(\u4.ssdec[2] ),
    .B(\u4.ssdec[1] ),
    .Y(_0143_));
 sky130_fd_sc_hd__nand2_2 _0513_ (.A(\u4.ssdec[3] ),
    .B(_0143_),
    .Y(_0144_));
 sky130_fd_sc_hd__o21ai_1 _0514_ (.A1(\u4.ssdec[3] ),
    .A2(_0142_),
    .B1(_0144_),
    .Y(net14));
 sky130_fd_sc_hd__and2_1 _0515_ (.A(\u4.ssdec[1] ),
    .B(\u4.ssdec[0] ),
    .X(_0145_));
 sky130_fd_sc_hd__and3b_1 _0516_ (.A_N(_0145_),
    .B(\u4.ssdec[2] ),
    .C(_0139_),
    .X(_0146_));
 sky130_fd_sc_hd__o21ai_1 _0517_ (.A1(\u4.ssdec[3] ),
    .A2(_0146_),
    .B1(_0144_),
    .Y(net19));
 sky130_fd_sc_hd__o21ba_1 _0518_ (.A1(\u4.ssdec[2] ),
    .A2(\u4.ssdec[0] ),
    .B1_N(\u4.ssdec[3] ),
    .X(_0147_));
 sky130_fd_sc_hd__or2_1 _0519_ (.A(_0143_),
    .B(_0147_),
    .X(_0148_));
 sky130_fd_sc_hd__clkbuf_1 _0520_ (.A(_0148_),
    .X(net20));
 sky130_fd_sc_hd__nor2_1 _0521_ (.A(_0141_),
    .B(_0146_),
    .Y(_0149_));
 sky130_fd_sc_hd__o21ai_2 _0522_ (.A1(\u4.ssdec[3] ),
    .A2(_0149_),
    .B1(_0144_),
    .Y(net21));
 sky130_fd_sc_hd__o21ba_1 _0523_ (.A1(_0140_),
    .A2(\u4.ssdec[3] ),
    .B1_N(_0143_),
    .X(_0150_));
 sky130_fd_sc_hd__nor2_1 _0524_ (.A(\u4.ssdec[0] ),
    .B(_0150_),
    .Y(net22));
 sky130_fd_sc_hd__and2b_1 _0525_ (.A_N(\u4.ssdec[2] ),
    .B(_0139_),
    .X(_0151_));
 sky130_fd_sc_hd__o31ai_2 _0526_ (.A1(\u4.ssdec[3] ),
    .A2(_0145_),
    .A3(_0151_),
    .B1(_0144_),
    .Y(net23));
 sky130_fd_sc_hd__a211o_1 _0527_ (.A1(\u4.ssdec[2] ),
    .A2(_0145_),
    .B1(_0143_),
    .C1(\u4.ssdec[3] ),
    .X(_0152_));
 sky130_fd_sc_hd__nand2_1 _0528_ (.A(_0144_),
    .B(_0152_),
    .Y(net24));
 sky130_fd_sc_hd__or4b_1 _0529_ (.A(\u6.reg_sync[1] ),
    .B(\u6.reg_sync[0] ),
    .C(\u6.reg_sync[3] ),
    .D_N(\u6.reg_sync[2] ),
    .X(_0153_));
 sky130_fd_sc_hd__or4b_1 _0530_ (.A(\u6.reg_sync[1] ),
    .B(\u6.reg_sync[3] ),
    .C(\u6.reg_sync[2] ),
    .D_N(\u6.reg_sync[0] ),
    .X(_0154_));
 sky130_fd_sc_hd__a21oi_1 _0531_ (.A1(_0153_),
    .A2(_0154_),
    .B1(_0120_),
    .Y(\u6.next_reg_num[0] ));
 sky130_fd_sc_hd__or4b_1 _0532_ (.A(\u6.reg_sync[0] ),
    .B(\u6.reg_sync[3] ),
    .C(\u6.reg_sync[2] ),
    .D_N(\u6.reg_sync[1] ),
    .X(_0155_));
 sky130_fd_sc_hd__a21oi_1 _0533_ (.A1(_0153_),
    .A2(_0155_),
    .B1(_0120_),
    .Y(\u6.next_reg_num[1] ));
 sky130_fd_sc_hd__or4b_1 _0534_ (.A(\u6.reg_sync[1] ),
    .B(\u6.reg_sync[0] ),
    .C(\u6.reg_sync[2] ),
    .D_N(\u6.reg_sync[3] ),
    .X(_0156_));
 sky130_fd_sc_hd__nor2_1 _0535_ (.A(_0120_),
    .B(_0156_),
    .Y(\u6.next_reg_num[2] ));
 sky130_fd_sc_hd__or2_1 _0536_ (.A(\u4.ssdec[5] ),
    .B(\u4.ssdec[4] ),
    .X(_0157_));
 sky130_fd_sc_hd__inv_2 _0537_ (.A(\u4.ssdec[5] ),
    .Y(_0158_));
 sky130_fd_sc_hd__a21oi_1 _0538_ (.A1(_0158_),
    .A2(\u4.ssdec[4] ),
    .B1(\u4.ssdec[6] ),
    .Y(_0159_));
 sky130_fd_sc_hd__a21oi_1 _0539_ (.A1(\u4.ssdec[6] ),
    .A2(_0157_),
    .B1(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__nor2_1 _0540_ (.A(\u4.ssdec[6] ),
    .B(\u4.ssdec[5] ),
    .Y(_0161_));
 sky130_fd_sc_hd__nand2_2 _0541_ (.A(\u4.ssdec[7] ),
    .B(_0161_),
    .Y(_0162_));
 sky130_fd_sc_hd__o21ai_1 _0542_ (.A1(\u4.ssdec[7] ),
    .A2(_0160_),
    .B1(_0162_),
    .Y(net25));
 sky130_fd_sc_hd__and2_1 _0543_ (.A(\u4.ssdec[5] ),
    .B(\u4.ssdec[4] ),
    .X(_0163_));
 sky130_fd_sc_hd__and3b_1 _0544_ (.A_N(_0163_),
    .B(\u4.ssdec[6] ),
    .C(_0157_),
    .X(_0164_));
 sky130_fd_sc_hd__o21ai_1 _0545_ (.A1(\u4.ssdec[7] ),
    .A2(_0164_),
    .B1(_0162_),
    .Y(net26));
 sky130_fd_sc_hd__o21ba_1 _0546_ (.A1(\u4.ssdec[6] ),
    .A2(\u4.ssdec[4] ),
    .B1_N(\u4.ssdec[7] ),
    .X(_0165_));
 sky130_fd_sc_hd__or2_1 _0547_ (.A(_0161_),
    .B(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__clkbuf_1 _0548_ (.A(_0166_),
    .X(net27));
 sky130_fd_sc_hd__nor2_1 _0549_ (.A(_0159_),
    .B(_0164_),
    .Y(_0167_));
 sky130_fd_sc_hd__o21ai_1 _0550_ (.A1(\u4.ssdec[7] ),
    .A2(_0167_),
    .B1(_0162_),
    .Y(net15));
 sky130_fd_sc_hd__o21ba_1 _0551_ (.A1(_0158_),
    .A2(\u4.ssdec[7] ),
    .B1_N(_0161_),
    .X(_0168_));
 sky130_fd_sc_hd__nor2_1 _0552_ (.A(\u4.ssdec[4] ),
    .B(_0168_),
    .Y(net16));
 sky130_fd_sc_hd__and2b_1 _0553_ (.A_N(\u4.ssdec[6] ),
    .B(_0157_),
    .X(_0169_));
 sky130_fd_sc_hd__o31ai_2 _0554_ (.A1(\u4.ssdec[7] ),
    .A2(_0163_),
    .A3(_0169_),
    .B1(_0162_),
    .Y(net17));
 sky130_fd_sc_hd__a211o_1 _0555_ (.A1(\u4.ssdec[6] ),
    .A2(_0163_),
    .B1(_0161_),
    .C1(\u4.ssdec[7] ),
    .X(_0170_));
 sky130_fd_sc_hd__nand2_1 _0556_ (.A(_0162_),
    .B(_0170_),
    .Y(net18));
 sky130_fd_sc_hd__inv_2 _0557_ (.A(net71),
    .Y(_0171_));
 sky130_fd_sc_hd__nor2_1 _0558_ (.A(_0171_),
    .B(_0120_),
    .Y(_0000_));
 sky130_fd_sc_hd__and3_1 _0559_ (.A(\u1.state[13] ),
    .B(_0131_),
    .C(_0120_),
    .X(_0172_));
 sky130_fd_sc_hd__clkbuf_1 _0560_ (.A(_0172_),
    .X(_0002_));
 sky130_fd_sc_hd__inv_2 _0561_ (.A(net65),
    .Y(_0173_));
 sky130_fd_sc_hd__nor2_1 _0562_ (.A(_0173_),
    .B(_0128_),
    .Y(_0001_));
 sky130_fd_sc_hd__nor2_8 _0563_ (.A(_0121_),
    .B(\u1.state[3] ),
    .Y(_0174_));
 sky130_fd_sc_hd__a22o_1 _0564_ (.A1(_0121_),
    .A2(\u1.keycode[0] ),
    .B1(net73),
    .B2(_0174_),
    .X(_0015_));
 sky130_fd_sc_hd__and2_1 _0565_ (.A(\u1.keycode[1] ),
    .B(\u1.keycode[0] ),
    .X(_0175_));
 sky130_fd_sc_hd__nor2_1 _0566_ (.A(\u1.keycode[1] ),
    .B(\u1.keycode[0] ),
    .Y(_0176_));
 sky130_fd_sc_hd__nor2_1 _0567_ (.A(_0175_),
    .B(_0176_),
    .Y(_0177_));
 sky130_fd_sc_hd__or2_1 _0568_ (.A(\u1.keycode[2] ),
    .B(_0175_),
    .X(_0178_));
 sky130_fd_sc_hd__xnor2_2 _0569_ (.A(\u1.keycode[3] ),
    .B(_0178_),
    .Y(_0179_));
 sky130_fd_sc_hd__o21ai_1 _0570_ (.A1(_0177_),
    .A2(_0179_),
    .B1(\u1.keycode[8] ),
    .Y(_0180_));
 sky130_fd_sc_hd__a31o_1 _0571_ (.A1(\u1.keycode[3] ),
    .A2(\u1.keycode[2] ),
    .A3(_0177_),
    .B1(_0180_),
    .X(_0181_));
 sky130_fd_sc_hd__or2_1 _0572_ (.A(\u1.keycode[1] ),
    .B(\u1.keycode[8] ),
    .X(_0182_));
 sky130_fd_sc_hd__a32o_1 _0573_ (.A1(_0121_),
    .A2(_0181_),
    .A3(_0182_),
    .B1(net96),
    .B2(_0174_),
    .X(_0016_));
 sky130_fd_sc_hd__or2_1 _0574_ (.A(\u1.keycode[1] ),
    .B(\u1.keycode[0] ),
    .X(_0183_));
 sky130_fd_sc_hd__o2111ai_1 _0575_ (.A1(\u1.keycode[3] ),
    .A2(_0175_),
    .B1(_0183_),
    .C1(\u1.keycode[2] ),
    .D1(\u1.keycode[8] ),
    .Y(_0184_));
 sky130_fd_sc_hd__a31o_1 _0576_ (.A1(\u1.keycode[1] ),
    .A2(\u1.keycode[0] ),
    .A3(\u1.keycode[8] ),
    .B1(\u1.keycode[2] ),
    .X(_0185_));
 sky130_fd_sc_hd__a32o_1 _0577_ (.A1(_0121_),
    .A2(_0184_),
    .A3(_0185_),
    .B1(net81),
    .B2(_0174_),
    .X(_0017_));
 sky130_fd_sc_hd__o31ai_4 _0578_ (.A1(\u1.keycode[2] ),
    .A2(_0175_),
    .A3(_0176_),
    .B1(_0179_),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _0579_ (.A(\u1.keycode[8] ),
    .Y(_0187_));
 sky130_fd_sc_hd__and2_1 _0580_ (.A(\u1.keycode[3] ),
    .B(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__a31o_1 _0581_ (.A1(\u1.keycode[8] ),
    .A2(_0179_),
    .A3(_0186_),
    .B1(_0188_),
    .X(_0189_));
 sky130_fd_sc_hd__a22o_1 _0582_ (.A1(net91),
    .A2(_0174_),
    .B1(_0189_),
    .B2(_0121_),
    .X(_0018_));
 sky130_fd_sc_hd__a21oi_1 _0583_ (.A1(\u1.keycode[8] ),
    .A2(_0186_),
    .B1(\u1.keycode[4] ),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_2 _0584_ (.A(_0121_),
    .Y(_0191_));
 sky130_fd_sc_hd__a31o_1 _0585_ (.A1(\u1.keycode[4] ),
    .A2(\u1.keycode[8] ),
    .A3(_0186_),
    .B1(_0191_),
    .X(_0192_));
 sky130_fd_sc_hd__a2bb2o_1 _0586_ (.A1_N(_0190_),
    .A2_N(_0192_),
    .B1(net84),
    .B2(_0174_),
    .X(_0019_));
 sky130_fd_sc_hd__or4_1 _0587_ (.A(\u1.keycode[3] ),
    .B(\u1.keycode[2] ),
    .C(\u1.keycode[7] ),
    .D(\u1.keycode[6] ),
    .X(_0193_));
 sky130_fd_sc_hd__o41a_1 _0588_ (.A1(\u1.keycode[5] ),
    .A2(\u1.keycode[4] ),
    .A3(_0183_),
    .A4(_0193_),
    .B1(\u1.keycode[8] ),
    .X(_0194_));
 sky130_fd_sc_hd__a21o_1 _0589_ (.A1(\u1.keycode[5] ),
    .A2(_0187_),
    .B1(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__o21a_1 _0590_ (.A1(\u1.keycode[4] ),
    .A2(_0186_),
    .B1(\u1.keycode[5] ),
    .X(_0196_));
 sky130_fd_sc_hd__nor3_1 _0591_ (.A(\u1.keycode[5] ),
    .B(\u1.keycode[4] ),
    .C(_0186_),
    .Y(_0197_));
 sky130_fd_sc_hd__or2_1 _0592_ (.A(_0196_),
    .B(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__nor2_1 _0593_ (.A(\u1.keycode[6] ),
    .B(_0196_),
    .Y(_0199_));
 sky130_fd_sc_hd__xnor2_1 _0594_ (.A(\u1.keycode[7] ),
    .B(_0199_),
    .Y(_0200_));
 sky130_fd_sc_hd__nor2_1 _0595_ (.A(_0198_),
    .B(_0200_),
    .Y(_0201_));
 sky130_fd_sc_hd__a21o_1 _0596_ (.A1(_0198_),
    .A2(_0200_),
    .B1(_0187_),
    .X(_0202_));
 sky130_fd_sc_hd__a21o_1 _0597_ (.A1(\u1.keycode[6] ),
    .A2(_0201_),
    .B1(_0202_),
    .X(_0203_));
 sky130_fd_sc_hd__a32o_1 _0598_ (.A1(_0121_),
    .A2(_0195_),
    .A3(_0203_),
    .B1(net77),
    .B2(_0174_),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _0599_ (.A(\u1.keycode[6] ),
    .B(_0196_),
    .X(_0204_));
 sky130_fd_sc_hd__or2_1 _0600_ (.A(_0199_),
    .B(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__o21ai_1 _0601_ (.A1(_0201_),
    .A2(_0205_),
    .B1(\u1.keycode[8] ),
    .Y(_0206_));
 sky130_fd_sc_hd__or2_1 _0602_ (.A(\u1.keycode[6] ),
    .B(\u1.keycode[8] ),
    .X(_0207_));
 sky130_fd_sc_hd__a32o_1 _0603_ (.A1(_0121_),
    .A2(_0206_),
    .A3(_0207_),
    .B1(net74),
    .B2(_0174_),
    .X(_0021_));
 sky130_fd_sc_hd__a32o_1 _0604_ (.A1(_0194_),
    .A2(_0201_),
    .A3(_0205_),
    .B1(_0187_),
    .B2(\u1.keycode[7] ),
    .X(_0208_));
 sky130_fd_sc_hd__a22o_1 _0605_ (.A1(net87),
    .A2(_0174_),
    .B1(_0208_),
    .B2(_0121_),
    .X(_0022_));
 sky130_fd_sc_hd__a22o_1 _0606_ (.A1(net132),
    .A2(_0174_),
    .B1(_0194_),
    .B2(_0121_),
    .X(_0023_));
 sky130_fd_sc_hd__o21ai_4 _0607_ (.A1(\u4.result_ready ),
    .A2(\u1.state[3] ),
    .B1(_0191_),
    .Y(_0209_));
 sky130_fd_sc_hd__and2_2 _0608_ (.A(_0191_),
    .B(\u1.state[3] ),
    .X(_0210_));
 sky130_fd_sc_hd__nor2_1 _0609_ (.A(_0209_),
    .B(_0210_),
    .Y(_0211_));
 sky130_fd_sc_hd__nand3_1 _0610_ (.A(\u8.op2[0] ),
    .B(\u8.op2[1] ),
    .C(\u8.buff_opcode[1] ),
    .Y(_0212_));
 sky130_fd_sc_hd__and4b_1 _0611_ (.A_N(\u8.op2[2] ),
    .B(\u8.buff_opcode[1] ),
    .C(\u8.op2[1] ),
    .D(\u8.op2[0] ),
    .X(_0213_));
 sky130_fd_sc_hd__a21o_1 _0612_ (.A1(\u8.op2[2] ),
    .A2(_0212_),
    .B1(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__or2_2 _0613_ (.A(\u8.new_op1[2] ),
    .B(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__nand2_1 _0614_ (.A(\u8.op2[1] ),
    .B(\u8.buff_opcode[1] ),
    .Y(_0216_));
 sky130_fd_sc_hd__and2b_1 _0615_ (.A_N(\u8.op2[0] ),
    .B(\u8.buff_opcode[1] ),
    .X(_0217_));
 sky130_fd_sc_hd__o22a_1 _0616_ (.A1(\u8.op2[0] ),
    .A2(_0216_),
    .B1(_0217_),
    .B2(\u8.op2[1] ),
    .X(_0218_));
 sky130_fd_sc_hd__xor2_2 _0617_ (.A(\u8.new_op1[1] ),
    .B(_0218_),
    .X(_0219_));
 sky130_fd_sc_hd__and2_1 _0618_ (.A(\u8.new_op1[1] ),
    .B(_0218_),
    .X(_0220_));
 sky130_fd_sc_hd__a31o_1 _0619_ (.A1(\u8.new_op1[0] ),
    .A2(\u8.op2[0] ),
    .A3(_0219_),
    .B1(_0220_),
    .X(_0221_));
 sky130_fd_sc_hd__nand2_1 _0620_ (.A(\u8.new_op1[2] ),
    .B(_0214_),
    .Y(_0222_));
 sky130_fd_sc_hd__a21boi_4 _0621_ (.A1(_0215_),
    .A2(_0221_),
    .B1_N(_0222_),
    .Y(_0223_));
 sky130_fd_sc_hd__inv_2 _0622_ (.A(\u8.buff_opcode[1] ),
    .Y(_0224_));
 sky130_fd_sc_hd__a211o_1 _0623_ (.A1(\u8.op2[0] ),
    .A2(\u8.op2[1] ),
    .B1(_0224_),
    .C1(\u8.op2[2] ),
    .X(_0225_));
 sky130_fd_sc_hd__xnor2_1 _0624_ (.A(\u8.op2[3] ),
    .B(_0225_),
    .Y(_0226_));
 sky130_fd_sc_hd__and2_1 _0625_ (.A(\u8.new_op1[3] ),
    .B(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__nor2_1 _0626_ (.A(\u8.new_op1[3] ),
    .B(_0226_),
    .Y(_0228_));
 sky130_fd_sc_hd__nor2_1 _0627_ (.A(_0227_),
    .B(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__xnor2_2 _0628_ (.A(_0223_),
    .B(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__nand2_1 _0629_ (.A(\u8.new_op1[0] ),
    .B(\u8.op2[0] ),
    .Y(_0231_));
 sky130_fd_sc_hd__xnor2_2 _0630_ (.A(_0231_),
    .B(_0219_),
    .Y(_0232_));
 sky130_fd_sc_hd__nand2_1 _0631_ (.A(_0222_),
    .B(_0215_),
    .Y(_0233_));
 sky130_fd_sc_hd__xnor2_1 _0632_ (.A(_0221_),
    .B(_0233_),
    .Y(_0234_));
 sky130_fd_sc_hd__or2_2 _0633_ (.A(_0232_),
    .B(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__o21bai_4 _0634_ (.A1(_0228_),
    .A2(_0223_),
    .B1_N(_0227_),
    .Y(_0236_));
 sky130_fd_sc_hd__a21oi_4 _0635_ (.A1(_0230_),
    .A2(_0235_),
    .B1(_0236_),
    .Y(_0237_));
 sky130_fd_sc_hd__xnor2_1 _0636_ (.A(\u8.op1[4] ),
    .B(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__xor2_1 _0637_ (.A(\u8.buff_opcode[1] ),
    .B(\u8.op2[4] ),
    .X(_0239_));
 sky130_fd_sc_hd__and2_2 _0638_ (.A(_0238_),
    .B(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__inv_2 _0639_ (.A(\u8.op1[4] ),
    .Y(_0241_));
 sky130_fd_sc_hd__or3b_1 _0640_ (.A(_0241_),
    .B(_0237_),
    .C_N(\u8.op1[5] ),
    .X(_0242_));
 sky130_fd_sc_hd__o21bai_1 _0641_ (.A1(_0241_),
    .A2(_0237_),
    .B1_N(\u8.op1[5] ),
    .Y(_0243_));
 sky130_fd_sc_hd__and3_1 _0642_ (.A(\u8.op2[5] ),
    .B(_0242_),
    .C(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__a21o_1 _0643_ (.A1(_0242_),
    .A2(_0243_),
    .B1(\u8.op2[5] ),
    .X(_0245_));
 sky130_fd_sc_hd__or2b_2 _0644_ (.A(_0244_),
    .B_N(_0245_),
    .X(_0246_));
 sky130_fd_sc_hd__xnor2_4 _0645_ (.A(_0240_),
    .B(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__a21o_1 _0646_ (.A1(_0240_),
    .A2(_0245_),
    .B1(_0244_),
    .X(_0248_));
 sky130_fd_sc_hd__nand2_1 _0647_ (.A(\u8.buff_opcode[1] ),
    .B(\u8.op2[5] ),
    .Y(_0249_));
 sky130_fd_sc_hd__xor2_2 _0648_ (.A(\u8.op2[6] ),
    .B(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__and3b_1 _0649_ (.A_N(_0237_),
    .B(\u8.op1[5] ),
    .C(\u8.op1[4] ),
    .X(_0251_));
 sky130_fd_sc_hd__xnor2_2 _0650_ (.A(\u8.op1[6] ),
    .B(_0251_),
    .Y(_0252_));
 sky130_fd_sc_hd__xnor2_1 _0651_ (.A(_0250_),
    .B(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__xnor2_2 _0652_ (.A(_0248_),
    .B(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__nor2_2 _0653_ (.A(_0247_),
    .B(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hd__nand2_1 _0654_ (.A(_0250_),
    .B(_0252_),
    .Y(_0256_));
 sky130_fd_sc_hd__nor2_1 _0655_ (.A(_0250_),
    .B(_0252_),
    .Y(_0257_));
 sky130_fd_sc_hd__a21o_1 _0656_ (.A1(_0248_),
    .A2(_0256_),
    .B1(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__or3_1 _0657_ (.A(_0224_),
    .B(\u8.op2[5] ),
    .C(\u8.op2[6] ),
    .X(_0259_));
 sky130_fd_sc_hd__xor2_2 _0658_ (.A(\u8.op2[7] ),
    .B(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__nand2_1 _0659_ (.A(\u8.op1[6] ),
    .B(_0251_),
    .Y(_0261_));
 sky130_fd_sc_hd__xor2_2 _0660_ (.A(\u8.op1[7] ),
    .B(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__xor2_1 _0661_ (.A(_0260_),
    .B(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__xnor2_2 _0662_ (.A(_0258_),
    .B(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__xor2_4 _0663_ (.A(\u8.buff_opcode[1] ),
    .B(\u8.op2[8] ),
    .X(_0265_));
 sky130_fd_sc_hd__nand2_1 _0664_ (.A(_0260_),
    .B(_0262_),
    .Y(_0266_));
 sky130_fd_sc_hd__nor2_1 _0665_ (.A(_0260_),
    .B(_0262_),
    .Y(_0267_));
 sky130_fd_sc_hd__a21oi_2 _0666_ (.A1(_0266_),
    .A2(_0258_),
    .B1(_0267_),
    .Y(_0268_));
 sky130_fd_sc_hd__o2111ai_4 _0667_ (.A1(_0255_),
    .A2(_0264_),
    .B1(_0265_),
    .C1(_0268_),
    .D1(\u8.new_op1[8] ),
    .Y(_0269_));
 sky130_fd_sc_hd__o21a_2 _0668_ (.A1(_0255_),
    .A2(_0264_),
    .B1(_0268_),
    .X(_0270_));
 sky130_fd_sc_hd__or3_1 _0669_ (.A(\u8.new_op1[8] ),
    .B(_0270_),
    .C(_0265_),
    .X(_0271_));
 sky130_fd_sc_hd__nand2_1 _0670_ (.A(_0269_),
    .B(_0271_),
    .Y(_0272_));
 sky130_fd_sc_hd__a22o_1 _0671_ (.A1(net72),
    .A2(_0209_),
    .B1(_0211_),
    .B2(_0272_),
    .X(_0024_));
 sky130_fd_sc_hd__or3_1 _0672_ (.A(\u4.result_ready ),
    .B(_0121_),
    .C(\u1.state[3] ),
    .X(_0273_));
 sky130_fd_sc_hd__clkbuf_4 _0673_ (.A(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__nand2_1 _0674_ (.A(_0121_),
    .B(_0187_),
    .Y(_0275_));
 sky130_fd_sc_hd__a21oi_2 _0675_ (.A1(\u8.new_op1[8] ),
    .A2(_0270_),
    .B1(_0265_),
    .Y(_0276_));
 sky130_fd_sc_hd__o21ai_2 _0676_ (.A1(\u8.new_op1[8] ),
    .A2(_0270_),
    .B1(_0269_),
    .Y(_0277_));
 sky130_fd_sc_hd__nor2_2 _0677_ (.A(_0276_),
    .B(_0277_),
    .Y(_0278_));
 sky130_fd_sc_hd__a22o_1 _0678_ (.A1(_0275_),
    .A2(_0209_),
    .B1(_0278_),
    .B2(_0174_),
    .X(_0279_));
 sky130_fd_sc_hd__o21a_1 _0679_ (.A1(net63),
    .A2(_0274_),
    .B1(_0279_),
    .X(_0025_));
 sky130_fd_sc_hd__or4_1 _0680_ (.A(\u1.state[0] ),
    .B(\u1.state[8] ),
    .C(\u1.state[4] ),
    .D(\u1.state[11] ),
    .X(_0280_));
 sky130_fd_sc_hd__or4b_2 _0681_ (.A(\u1.state[13] ),
    .B(_0280_),
    .C(\u1.state[7] ),
    .D_N(_0174_),
    .X(_0281_));
 sky130_fd_sc_hd__or4_1 _0682_ (.A(\u1.state[1] ),
    .B(\u1.state[2] ),
    .C(\u1.state[6] ),
    .D(\u1.state[9] ),
    .X(_0282_));
 sky130_fd_sc_hd__or4_2 _0683_ (.A(\u1.state[10] ),
    .B(\u1.state[14] ),
    .C(\u1.state[12] ),
    .D(_0282_),
    .X(_0283_));
 sky130_fd_sc_hd__o21bai_4 _0684_ (.A1(_0281_),
    .A2(_0283_),
    .B1_N(_0128_),
    .Y(_0284_));
 sky130_fd_sc_hd__a21oi_4 _0685_ (.A1(\u1.keypad_sync[0] ),
    .A2(\u1.keypad_sync[1] ),
    .B1(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__inv_2 _0686_ (.A(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__a2bb2o_1 _0687_ (.A1_N(\u1.keypad_sync[0] ),
    .A2_N(_0284_),
    .B1(_0286_),
    .B2(\u1.keycode[0] ),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _0688_ (.A0(\u1.keycode[1] ),
    .A1(\u1.keycode[0] ),
    .S(_0285_),
    .X(_0287_));
 sky130_fd_sc_hd__clkbuf_1 _0689_ (.A(_0287_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _0690_ (.A0(\u1.keycode[2] ),
    .A1(\u1.keycode[1] ),
    .S(_0285_),
    .X(_0288_));
 sky130_fd_sc_hd__clkbuf_1 _0691_ (.A(_0288_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _0692_ (.A0(\u1.keycode[3] ),
    .A1(\u1.keycode[2] ),
    .S(_0285_),
    .X(_0289_));
 sky130_fd_sc_hd__clkbuf_1 _0693_ (.A(_0289_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _0694_ (.A0(\u1.keycode[4] ),
    .A1(\u1.keycode[3] ),
    .S(_0285_),
    .X(_0290_));
 sky130_fd_sc_hd__clkbuf_1 _0695_ (.A(_0290_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _0696_ (.A0(\u1.keycode[5] ),
    .A1(\u1.keycode[4] ),
    .S(_0285_),
    .X(_0291_));
 sky130_fd_sc_hd__clkbuf_1 _0697_ (.A(_0291_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _0698_ (.A0(\u1.keycode[6] ),
    .A1(\u1.keycode[5] ),
    .S(_0285_),
    .X(_0292_));
 sky130_fd_sc_hd__clkbuf_1 _0699_ (.A(_0292_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _0700_ (.A0(\u1.keycode[7] ),
    .A1(\u1.keycode[6] ),
    .S(_0285_),
    .X(_0293_));
 sky130_fd_sc_hd__clkbuf_1 _0701_ (.A(_0293_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _0702_ (.A0(\u1.keycode[8] ),
    .A1(\u1.keycode[7] ),
    .S(_0285_),
    .X(_0294_));
 sky130_fd_sc_hd__clkbuf_1 _0703_ (.A(_0294_),
    .X(_0034_));
 sky130_fd_sc_hd__and2b_2 _0704_ (.A_N(\u5.reg_num[2] ),
    .B(\u5.reg_num[0] ),
    .X(_0295_));
 sky130_fd_sc_hd__nand3_4 _0705_ (.A(\u5.reg_num[1] ),
    .B(_0210_),
    .C(_0295_),
    .Y(_0296_));
 sky130_fd_sc_hd__mux2_1 _0706_ (.A0(\u4.op1[0] ),
    .A1(net89),
    .S(_0296_),
    .X(_0297_));
 sky130_fd_sc_hd__clkbuf_1 _0707_ (.A(_0297_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _0708_ (.A0(\u4.op1[1] ),
    .A1(net107),
    .S(_0296_),
    .X(_0298_));
 sky130_fd_sc_hd__clkbuf_1 _0709_ (.A(_0298_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _0710_ (.A0(\u4.op1[2] ),
    .A1(net112),
    .S(_0296_),
    .X(_0299_));
 sky130_fd_sc_hd__clkbuf_1 _0711_ (.A(_0299_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _0712_ (.A0(\u4.op1[3] ),
    .A1(net94),
    .S(_0296_),
    .X(_0300_));
 sky130_fd_sc_hd__clkbuf_1 _0713_ (.A(_0300_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _0714_ (.A0(\u4.op1[4] ),
    .A1(net115),
    .S(_0296_),
    .X(_0301_));
 sky130_fd_sc_hd__clkbuf_1 _0715_ (.A(_0301_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _0716_ (.A0(\u4.op1[5] ),
    .A1(net105),
    .S(_0296_),
    .X(_0302_));
 sky130_fd_sc_hd__clkbuf_1 _0717_ (.A(_0302_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _0718_ (.A0(\u4.op1[6] ),
    .A1(net99),
    .S(_0296_),
    .X(_0303_));
 sky130_fd_sc_hd__clkbuf_1 _0719_ (.A(_0303_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _0720_ (.A0(\u4.op1[7] ),
    .A1(net110),
    .S(_0296_),
    .X(_0304_));
 sky130_fd_sc_hd__clkbuf_1 _0721_ (.A(_0304_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _0722_ (.A0(\u4.op1[8] ),
    .A1(net93),
    .S(_0296_),
    .X(_0305_));
 sky130_fd_sc_hd__clkbuf_1 _0723_ (.A(_0305_),
    .X(_0043_));
 sky130_fd_sc_hd__and4bb_1 _0724_ (.A_N(\u5.reg_num[0] ),
    .B_N(\u5.reg_num[2] ),
    .C(_0210_),
    .D(\u5.reg_num[1] ),
    .X(_0306_));
 sky130_fd_sc_hd__clkbuf_4 _0725_ (.A(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _0726_ (.A0(net122),
    .A1(\u4.op1[0] ),
    .S(_0307_),
    .X(_0308_));
 sky130_fd_sc_hd__clkbuf_1 _0727_ (.A(_0308_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _0728_ (.A0(net80),
    .A1(\u4.op1[1] ),
    .S(_0307_),
    .X(_0309_));
 sky130_fd_sc_hd__clkbuf_1 _0729_ (.A(_0309_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _0730_ (.A0(net97),
    .A1(\u4.op1[2] ),
    .S(_0307_),
    .X(_0310_));
 sky130_fd_sc_hd__clkbuf_1 _0731_ (.A(_0310_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _0732_ (.A0(net104),
    .A1(\u4.op1[3] ),
    .S(_0307_),
    .X(_0311_));
 sky130_fd_sc_hd__clkbuf_1 _0733_ (.A(_0311_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _0734_ (.A0(net82),
    .A1(\u4.op1[4] ),
    .S(_0307_),
    .X(_0312_));
 sky130_fd_sc_hd__clkbuf_1 _0735_ (.A(_0312_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _0736_ (.A0(net103),
    .A1(\u4.op1[5] ),
    .S(_0307_),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_1 _0737_ (.A(_0313_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _0738_ (.A0(net85),
    .A1(\u4.op1[6] ),
    .S(_0307_),
    .X(_0314_));
 sky130_fd_sc_hd__clkbuf_1 _0739_ (.A(_0314_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _0740_ (.A0(net88),
    .A1(\u4.op1[7] ),
    .S(_0307_),
    .X(_0315_));
 sky130_fd_sc_hd__clkbuf_1 _0741_ (.A(_0315_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _0742_ (.A0(net101),
    .A1(\u4.op1[8] ),
    .S(_0307_),
    .X(_0316_));
 sky130_fd_sc_hd__clkbuf_1 _0743_ (.A(_0316_),
    .X(_0052_));
 sky130_fd_sc_hd__and3b_1 _0744_ (.A_N(\u5.reg_num[1] ),
    .B(_0210_),
    .C(_0295_),
    .X(_0317_));
 sky130_fd_sc_hd__clkbuf_4 _0745_ (.A(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _0746_ (.A0(net83),
    .A1(\u4.op1[0] ),
    .S(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__clkbuf_1 _0747_ (.A(_0319_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _0748_ (.A0(net109),
    .A1(\u4.op1[1] ),
    .S(_0318_),
    .X(_0320_));
 sky130_fd_sc_hd__clkbuf_1 _0749_ (.A(_0320_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _0750_ (.A0(net102),
    .A1(\u4.op1[2] ),
    .S(_0318_),
    .X(_0321_));
 sky130_fd_sc_hd__clkbuf_1 _0751_ (.A(_0321_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _0752_ (.A0(net86),
    .A1(\u4.op1[3] ),
    .S(_0318_),
    .X(_0322_));
 sky130_fd_sc_hd__clkbuf_1 _0753_ (.A(_0322_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _0754_ (.A0(net98),
    .A1(\u4.op1[4] ),
    .S(_0318_),
    .X(_0323_));
 sky130_fd_sc_hd__clkbuf_1 _0755_ (.A(_0323_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _0756_ (.A0(net113),
    .A1(\u4.op1[5] ),
    .S(_0318_),
    .X(_0324_));
 sky130_fd_sc_hd__clkbuf_1 _0757_ (.A(_0324_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _0758_ (.A0(net92),
    .A1(\u4.op1[6] ),
    .S(_0318_),
    .X(_0325_));
 sky130_fd_sc_hd__clkbuf_1 _0759_ (.A(_0325_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _0760_ (.A0(net79),
    .A1(\u4.op1[7] ),
    .S(_0318_),
    .X(_0326_));
 sky130_fd_sc_hd__clkbuf_1 _0761_ (.A(_0326_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _0762_ (.A0(net106),
    .A1(\u4.op1[8] ),
    .S(_0318_),
    .X(_0327_));
 sky130_fd_sc_hd__clkbuf_1 _0763_ (.A(_0327_),
    .X(_0061_));
 sky130_fd_sc_hd__or4_1 _0764_ (.A(\u7.assign_op1 ),
    .B(\u7.assign_op2 ),
    .C(\u7.state[5] ),
    .D(_0135_),
    .X(_0328_));
 sky130_fd_sc_hd__nor2_1 _0765_ (.A(\u7.state[4] ),
    .B(_0003_),
    .Y(_0329_));
 sky130_fd_sc_hd__a211oi_2 _0766_ (.A1(\u7.state[6] ),
    .A2(_0004_),
    .B1(_0328_),
    .C1(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__and4bb_1 _0767_ (.A_N(\u5.reg_num[0] ),
    .B_N(\u5.reg_num[2] ),
    .C(_0330_),
    .D(\u5.reg_num[1] ),
    .X(_0331_));
 sky130_fd_sc_hd__buf_4 _0768_ (.A(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__and3_1 _0769_ (.A(\u5.reg_num[1] ),
    .B(_0295_),
    .C(_0330_),
    .X(_0333_));
 sky130_fd_sc_hd__clkbuf_4 _0770_ (.A(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__and3_1 _0771_ (.A(\u5.reg_num[2] ),
    .B(_0133_),
    .C(_0330_),
    .X(_0335_));
 sky130_fd_sc_hd__buf_4 _0772_ (.A(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__nor3_2 _0773_ (.A(_0334_),
    .B(_0332_),
    .C(_0336_),
    .Y(_0337_));
 sky130_fd_sc_hd__a22o_1 _0774_ (.A1(\u5.reg3[0] ),
    .A2(_0334_),
    .B1(_0336_),
    .B2(\u5.reg4[0] ),
    .X(_0338_));
 sky130_fd_sc_hd__a221o_1 _0775_ (.A1(\u5.reg2[0] ),
    .A2(_0332_),
    .B1(_0337_),
    .B2(\u5.reg1[0] ),
    .C1(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__a211o_4 _0776_ (.A1(_0295_),
    .A2(_0330_),
    .B1(_0332_),
    .C1(_0336_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _0777_ (.A0(\u5.reg_val[0] ),
    .A1(_0339_),
    .S(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__clkbuf_1 _0778_ (.A(_0341_),
    .X(_0062_));
 sky130_fd_sc_hd__a22o_1 _0779_ (.A1(\u5.reg3[1] ),
    .A2(_0334_),
    .B1(_0336_),
    .B2(\u5.reg4[1] ),
    .X(_0342_));
 sky130_fd_sc_hd__a221o_1 _0780_ (.A1(\u5.reg2[1] ),
    .A2(_0332_),
    .B1(_0337_),
    .B2(\u5.reg1[1] ),
    .C1(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _0781_ (.A0(net136),
    .A1(_0343_),
    .S(_0340_),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_1 _0782_ (.A(_0344_),
    .X(_0063_));
 sky130_fd_sc_hd__a22o_1 _0783_ (.A1(\u5.reg3[2] ),
    .A2(_0334_),
    .B1(_0336_),
    .B2(\u5.reg4[2] ),
    .X(_0345_));
 sky130_fd_sc_hd__a221o_1 _0784_ (.A1(\u5.reg2[2] ),
    .A2(_0332_),
    .B1(net28),
    .B2(\u5.reg1[2] ),
    .C1(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _0785_ (.A0(\u5.reg_val[2] ),
    .A1(_0346_),
    .S(_0340_),
    .X(_0347_));
 sky130_fd_sc_hd__clkbuf_1 _0786_ (.A(_0347_),
    .X(_0064_));
 sky130_fd_sc_hd__a22o_1 _0787_ (.A1(\u5.reg3[3] ),
    .A2(_0334_),
    .B1(_0336_),
    .B2(\u5.reg4[3] ),
    .X(_0348_));
 sky130_fd_sc_hd__a221o_1 _0788_ (.A1(\u5.reg2[3] ),
    .A2(_0332_),
    .B1(_0337_),
    .B2(\u5.reg1[3] ),
    .C1(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _0789_ (.A0(net134),
    .A1(_0349_),
    .S(_0340_),
    .X(_0350_));
 sky130_fd_sc_hd__clkbuf_1 _0790_ (.A(_0350_),
    .X(_0065_));
 sky130_fd_sc_hd__a22o_1 _0791_ (.A1(\u5.reg3[4] ),
    .A2(_0334_),
    .B1(_0336_),
    .B2(\u5.reg4[4] ),
    .X(_0351_));
 sky130_fd_sc_hd__a221o_1 _0792_ (.A1(\u5.reg2[4] ),
    .A2(_0332_),
    .B1(net28),
    .B2(\u5.reg1[4] ),
    .C1(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _0793_ (.A0(\u5.reg_val[4] ),
    .A1(_0352_),
    .S(_0340_),
    .X(_0353_));
 sky130_fd_sc_hd__clkbuf_1 _0794_ (.A(_0353_),
    .X(_0066_));
 sky130_fd_sc_hd__a22o_1 _0795_ (.A1(\u5.reg3[5] ),
    .A2(_0334_),
    .B1(_0336_),
    .B2(\u5.reg4[5] ),
    .X(_0354_));
 sky130_fd_sc_hd__a221o_1 _0796_ (.A1(\u5.reg2[5] ),
    .A2(_0332_),
    .B1(net28),
    .B2(\u5.reg1[5] ),
    .C1(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _0797_ (.A0(\u5.reg_val[5] ),
    .A1(_0355_),
    .S(_0340_),
    .X(_0356_));
 sky130_fd_sc_hd__clkbuf_1 _0798_ (.A(_0356_),
    .X(_0067_));
 sky130_fd_sc_hd__a22o_1 _0799_ (.A1(\u5.reg3[6] ),
    .A2(_0334_),
    .B1(_0336_),
    .B2(\u5.reg4[6] ),
    .X(_0357_));
 sky130_fd_sc_hd__a221o_1 _0800_ (.A1(\u5.reg2[6] ),
    .A2(_0332_),
    .B1(net28),
    .B2(\u5.reg1[6] ),
    .C1(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _0801_ (.A0(\u5.reg_val[6] ),
    .A1(_0358_),
    .S(_0340_),
    .X(_0359_));
 sky130_fd_sc_hd__clkbuf_1 _0802_ (.A(_0359_),
    .X(_0068_));
 sky130_fd_sc_hd__a22o_1 _0803_ (.A1(\u5.reg3[7] ),
    .A2(_0334_),
    .B1(_0336_),
    .B2(\u5.reg4[7] ),
    .X(_0360_));
 sky130_fd_sc_hd__a221o_1 _0804_ (.A1(\u5.reg2[7] ),
    .A2(_0332_),
    .B1(net28),
    .B2(\u5.reg1[7] ),
    .C1(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _0805_ (.A0(\u5.reg_val[7] ),
    .A1(_0361_),
    .S(_0340_),
    .X(_0362_));
 sky130_fd_sc_hd__clkbuf_1 _0806_ (.A(_0362_),
    .X(_0069_));
 sky130_fd_sc_hd__a22o_1 _0807_ (.A1(\u5.reg3[8] ),
    .A2(_0334_),
    .B1(_0336_),
    .B2(\u5.reg4[8] ),
    .X(_0363_));
 sky130_fd_sc_hd__a221o_1 _0808_ (.A1(\u5.reg2[8] ),
    .A2(_0332_),
    .B1(_0337_),
    .B2(\u5.reg1[8] ),
    .C1(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _0809_ (.A0(\u5.reg_val[8] ),
    .A1(_0364_),
    .S(_0340_),
    .X(_0365_));
 sky130_fd_sc_hd__clkbuf_1 _0810_ (.A(_0365_),
    .X(_0070_));
 sky130_fd_sc_hd__or2_1 _0811_ (.A(\u8.new_op1[0] ),
    .B(\u8.op2[0] ),
    .X(_0366_));
 sky130_fd_sc_hd__and2_1 _0812_ (.A(_0231_),
    .B(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__a22o_1 _0813_ (.A1(_0121_),
    .A2(\u1.keycode[0] ),
    .B1(_0174_),
    .B2(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _0814_ (.A0(\u4.ssdec[0] ),
    .A1(_0368_),
    .S(_0274_),
    .X(_0369_));
 sky130_fd_sc_hd__clkbuf_1 _0815_ (.A(_0369_),
    .X(_0071_));
 sky130_fd_sc_hd__o21ai_1 _0816_ (.A1(_0191_),
    .A2(\u1.keycode[1] ),
    .B1(_0209_),
    .Y(_0370_));
 sky130_fd_sc_hd__xnor2_1 _0817_ (.A(_0232_),
    .B(_0237_),
    .Y(_0371_));
 sky130_fd_sc_hd__nand2_1 _0818_ (.A(_0367_),
    .B(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__nor2_1 _0819_ (.A(_0367_),
    .B(_0371_),
    .Y(_0373_));
 sky130_fd_sc_hd__inv_2 _0820_ (.A(_0373_),
    .Y(_0374_));
 sky130_fd_sc_hd__nand2_1 _0821_ (.A(_0372_),
    .B(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__nand2_1 _0822_ (.A(_0236_),
    .B(_0235_),
    .Y(_0376_));
 sky130_fd_sc_hd__mux2_1 _0823_ (.A0(_0376_),
    .A1(_0235_),
    .S(_0230_),
    .X(_0377_));
 sky130_fd_sc_hd__inv_2 _0824_ (.A(_0236_),
    .Y(_0378_));
 sky130_fd_sc_hd__o21ai_1 _0825_ (.A1(_0232_),
    .A2(_0237_),
    .B1(_0234_),
    .Y(_0379_));
 sky130_fd_sc_hd__o21a_1 _0826_ (.A1(_0378_),
    .A2(_0235_),
    .B1(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__and2_1 _0827_ (.A(_0372_),
    .B(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__nand2_1 _0828_ (.A(_0377_),
    .B(_0380_),
    .Y(_0382_));
 sky130_fd_sc_hd__o22a_1 _0829_ (.A1(_0377_),
    .A2(_0381_),
    .B1(_0382_),
    .B2(_0374_),
    .X(_0383_));
 sky130_fd_sc_hd__or3b_2 _0830_ (.A(_0276_),
    .B(_0277_),
    .C_N(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__o21ai_1 _0831_ (.A1(_0276_),
    .A2(_0277_),
    .B1(_0367_),
    .Y(_0385_));
 sky130_fd_sc_hd__a21oi_1 _0832_ (.A1(_0384_),
    .A2(_0385_),
    .B1(_0375_),
    .Y(_0386_));
 sky130_fd_sc_hd__or4b_1 _0833_ (.A(\u8.new_op1[1] ),
    .B(\u8.op2[5] ),
    .C(\u8.new_op1[8] ),
    .D_N(\u8.new_op1[3] ),
    .X(_0387_));
 sky130_fd_sc_hd__or4bb_1 _0834_ (.A(\u8.op2[0] ),
    .B(_0265_),
    .C_N(_0239_),
    .D_N(\u8.new_op1[0] ),
    .X(_0388_));
 sky130_fd_sc_hd__or4b_1 _0835_ (.A(_0218_),
    .B(_0387_),
    .C(_0388_),
    .D_N(_0250_),
    .X(_0389_));
 sky130_fd_sc_hd__or3b_1 _0836_ (.A(_0389_),
    .B(_0226_),
    .C_N(_0260_),
    .X(_0390_));
 sky130_fd_sc_hd__or3_1 _0837_ (.A(_0215_),
    .B(_0238_),
    .C(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__nand2_1 _0838_ (.A(_0242_),
    .B(_0243_),
    .Y(_0392_));
 sky130_fd_sc_hd__and4b_1 _0839_ (.A_N(_0391_),
    .B(_0392_),
    .C(_0252_),
    .D(_0262_),
    .X(_0393_));
 sky130_fd_sc_hd__and2b_2 _0840_ (.A_N(_0393_),
    .B(_0174_),
    .X(_0394_));
 sky130_fd_sc_hd__inv_2 _0841_ (.A(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__a311o_1 _0842_ (.A1(_0375_),
    .A2(_0384_),
    .A3(_0385_),
    .B1(_0386_),
    .C1(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__o2bb2a_1 _0843_ (.A1_N(_0370_),
    .A2_N(_0396_),
    .B1(\u4.ssdec[1] ),
    .B2(_0274_),
    .X(_0072_));
 sky130_fd_sc_hd__o21a_1 _0844_ (.A1(_0191_),
    .A2(\u1.keycode[2] ),
    .B1(_0209_),
    .X(_0397_));
 sky130_fd_sc_hd__or2_1 _0845_ (.A(_0276_),
    .B(_0277_),
    .X(_0398_));
 sky130_fd_sc_hd__a211o_1 _0846_ (.A1(_0372_),
    .A2(_0377_),
    .B1(_0380_),
    .C1(_0373_),
    .X(_0399_));
 sky130_fd_sc_hd__o21ai_1 _0847_ (.A1(_0398_),
    .A2(_0372_),
    .B1(_0380_),
    .Y(_0400_));
 sky130_fd_sc_hd__o211a_1 _0848_ (.A1(_0398_),
    .A2(_0399_),
    .B1(_0400_),
    .C1(_0394_),
    .X(_0401_));
 sky130_fd_sc_hd__o22a_1 _0849_ (.A1(net121),
    .A2(_0274_),
    .B1(_0397_),
    .B2(_0401_),
    .X(_0073_));
 sky130_fd_sc_hd__o21a_1 _0850_ (.A1(_0191_),
    .A2(\u1.keycode[3] ),
    .B1(_0209_),
    .X(_0402_));
 sky130_fd_sc_hd__nand3_1 _0851_ (.A(_0374_),
    .B(_0377_),
    .C(_0381_),
    .Y(_0403_));
 sky130_fd_sc_hd__mux2_1 _0852_ (.A0(_0377_),
    .A1(_0403_),
    .S(_0278_),
    .X(_0404_));
 sky130_fd_sc_hd__nor2_1 _0853_ (.A(_0395_),
    .B(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__o22a_1 _0854_ (.A1(\u4.ssdec[3] ),
    .A2(_0274_),
    .B1(_0402_),
    .B2(_0405_),
    .X(_0074_));
 sky130_fd_sc_hd__nor2_1 _0855_ (.A(_0238_),
    .B(_0239_),
    .Y(_0406_));
 sky130_fd_sc_hd__nor2_1 _0856_ (.A(_0240_),
    .B(_0406_),
    .Y(_0407_));
 sky130_fd_sc_hd__xnor2_1 _0857_ (.A(_0384_),
    .B(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__a22o_1 _0858_ (.A1(_0121_),
    .A2(\u1.keycode[4] ),
    .B1(_0394_),
    .B2(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _0859_ (.A0(\u4.ssdec[4] ),
    .A1(_0409_),
    .S(_0274_),
    .X(_0410_));
 sky130_fd_sc_hd__clkbuf_1 _0860_ (.A(_0410_),
    .X(_0075_));
 sky130_fd_sc_hd__o21a_1 _0861_ (.A1(_0191_),
    .A2(\u1.keycode[5] ),
    .B1(_0209_),
    .X(_0411_));
 sky130_fd_sc_hd__xor2_2 _0862_ (.A(_0247_),
    .B(_0270_),
    .X(_0412_));
 sky130_fd_sc_hd__nor2_1 _0863_ (.A(_0383_),
    .B(_0407_),
    .Y(_0413_));
 sky130_fd_sc_hd__and3_1 _0864_ (.A(_0278_),
    .B(_0412_),
    .C(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__a21oi_1 _0865_ (.A1(_0278_),
    .A2(_0413_),
    .B1(_0412_),
    .Y(_0415_));
 sky130_fd_sc_hd__o31a_1 _0866_ (.A1(_0393_),
    .A2(_0414_),
    .A3(_0415_),
    .B1(_0174_),
    .X(_0416_));
 sky130_fd_sc_hd__o22a_1 _0867_ (.A1(net124),
    .A2(_0274_),
    .B1(_0411_),
    .B2(_0416_),
    .X(_0076_));
 sky130_fd_sc_hd__nor2_1 _0868_ (.A(_0412_),
    .B(_0413_),
    .Y(_0417_));
 sky130_fd_sc_hd__inv_2 _0869_ (.A(_0268_),
    .Y(_0418_));
 sky130_fd_sc_hd__or2_1 _0870_ (.A(_0247_),
    .B(_0270_),
    .X(_0419_));
 sky130_fd_sc_hd__a22o_1 _0871_ (.A1(_0418_),
    .A2(_0255_),
    .B1(_0419_),
    .B2(_0254_),
    .X(_0420_));
 sky130_fd_sc_hd__a21o_1 _0872_ (.A1(_0278_),
    .A2(_0417_),
    .B1(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__a22oi_1 _0873_ (.A1(_0418_),
    .A2(_0255_),
    .B1(_0419_),
    .B2(_0254_),
    .Y(_0422_));
 sky130_fd_sc_hd__or2_1 _0874_ (.A(_0412_),
    .B(_0413_),
    .X(_0423_));
 sky130_fd_sc_hd__or3_1 _0875_ (.A(_0398_),
    .B(_0422_),
    .C(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__o21a_1 _0876_ (.A1(_0191_),
    .A2(\u1.keycode[6] ),
    .B1(_0209_),
    .X(_0425_));
 sky130_fd_sc_hd__a31o_1 _0877_ (.A1(_0394_),
    .A2(_0421_),
    .A3(_0424_),
    .B1(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__o21a_1 _0878_ (.A1(net114),
    .A2(_0274_),
    .B1(_0426_),
    .X(_0077_));
 sky130_fd_sc_hd__o21a_1 _0879_ (.A1(_0247_),
    .A2(_0254_),
    .B1(_0266_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _0880_ (.A0(_0255_),
    .A1(_0427_),
    .S(_0264_),
    .X(_0428_));
 sky130_fd_sc_hd__or4b_1 _0881_ (.A(_0398_),
    .B(_0420_),
    .C(_0417_),
    .D_N(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__a31o_1 _0882_ (.A1(_0278_),
    .A2(_0422_),
    .A3(_0423_),
    .B1(_0428_),
    .X(_0430_));
 sky130_fd_sc_hd__o21a_1 _0883_ (.A1(_0191_),
    .A2(\u1.keycode[7] ),
    .B1(_0209_),
    .X(_0431_));
 sky130_fd_sc_hd__a31o_1 _0884_ (.A1(_0394_),
    .A2(_0429_),
    .A3(_0430_),
    .B1(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__o21a_1 _0885_ (.A1(\u4.ssdec[7] ),
    .A2(_0274_),
    .B1(_0432_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _0886_ (.A0(\u8.op2[0] ),
    .A1(\u5.reg_val[0] ),
    .S(\u8.b_assign_op2 ),
    .X(_0433_));
 sky130_fd_sc_hd__clkbuf_1 _0887_ (.A(_0433_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _0888_ (.A0(\u8.op2[1] ),
    .A1(net130),
    .S(\u8.b_assign_op2 ),
    .X(_0434_));
 sky130_fd_sc_hd__clkbuf_1 _0889_ (.A(_0434_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _0890_ (.A0(\u8.op2[2] ),
    .A1(\u5.reg_val[2] ),
    .S(\u8.b_assign_op2 ),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_1 _0891_ (.A(_0435_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _0892_ (.A0(\u8.op2[3] ),
    .A1(net127),
    .S(\u8.b_assign_op2 ),
    .X(_0436_));
 sky130_fd_sc_hd__clkbuf_1 _0893_ (.A(_0436_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _0894_ (.A0(\u8.op2[4] ),
    .A1(\u5.reg_val[4] ),
    .S(\u8.b_assign_op2 ),
    .X(_0437_));
 sky130_fd_sc_hd__clkbuf_1 _0895_ (.A(_0437_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _0896_ (.A0(\u8.op2[5] ),
    .A1(\u5.reg_val[5] ),
    .S(\u8.b_assign_op2 ),
    .X(_0438_));
 sky130_fd_sc_hd__clkbuf_1 _0897_ (.A(_0438_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _0898_ (.A0(\u8.op2[6] ),
    .A1(\u5.reg_val[6] ),
    .S(\u8.b_assign_op2 ),
    .X(_0439_));
 sky130_fd_sc_hd__clkbuf_1 _0899_ (.A(_0439_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _0900_ (.A0(\u8.op2[7] ),
    .A1(\u5.reg_val[7] ),
    .S(\u8.b_assign_op2 ),
    .X(_0440_));
 sky130_fd_sc_hd__clkbuf_1 _0901_ (.A(_0440_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _0902_ (.A0(\u8.op2[8] ),
    .A1(\u5.reg_val[8] ),
    .S(\u8.b_assign_op2 ),
    .X(_0441_));
 sky130_fd_sc_hd__clkbuf_1 _0903_ (.A(_0441_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _0904_ (.A0(\u8.new_op1[0] ),
    .A1(net95),
    .S(\u8.b_assign_op1 ),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_1 _0905_ (.A(_0442_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _0906_ (.A0(\u8.new_op1[1] ),
    .A1(net135),
    .S(\u8.b_assign_op1 ),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_1 _0907_ (.A(_0443_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _0908_ (.A0(\u8.new_op1[2] ),
    .A1(\u5.reg_val[2] ),
    .S(\u8.b_assign_op1 ),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_1 _0909_ (.A(_0444_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _0910_ (.A0(\u8.new_op1[3] ),
    .A1(net127),
    .S(\u8.b_assign_op1 ),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_1 _0911_ (.A(_0445_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _0912_ (.A0(\u8.op1[4] ),
    .A1(\u5.reg_val[4] ),
    .S(\u8.b_assign_op1 ),
    .X(_0446_));
 sky130_fd_sc_hd__clkbuf_1 _0913_ (.A(_0446_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _0914_ (.A0(\u8.op1[5] ),
    .A1(\u5.reg_val[5] ),
    .S(\u8.b_assign_op1 ),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_1 _0915_ (.A(_0447_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _0916_ (.A0(\u8.op1[6] ),
    .A1(\u5.reg_val[6] ),
    .S(\u8.b_assign_op1 ),
    .X(_0448_));
 sky130_fd_sc_hd__clkbuf_1 _0917_ (.A(_0448_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _0918_ (.A0(\u8.op1[7] ),
    .A1(\u5.reg_val[7] ),
    .S(\u8.b_assign_op1 ),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_1 _0919_ (.A(_0449_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _0920_ (.A0(\u8.new_op1[8] ),
    .A1(\u5.reg_val[8] ),
    .S(\u8.b_assign_op1 ),
    .X(_0450_));
 sky130_fd_sc_hd__clkbuf_1 _0921_ (.A(_0450_),
    .X(_0096_));
 sky130_fd_sc_hd__and3_1 _0922_ (.A(\u5.reg_num[2] ),
    .B(_0133_),
    .C(_0210_),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_4 _0923_ (.A(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _0924_ (.A0(net90),
    .A1(\u4.op1[0] ),
    .S(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__clkbuf_1 _0925_ (.A(_0453_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _0926_ (.A0(net78),
    .A1(\u4.op1[1] ),
    .S(_0452_),
    .X(_0454_));
 sky130_fd_sc_hd__clkbuf_1 _0927_ (.A(_0454_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _0928_ (.A0(net108),
    .A1(\u4.op1[2] ),
    .S(_0452_),
    .X(_0455_));
 sky130_fd_sc_hd__clkbuf_1 _0929_ (.A(_0455_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _0930_ (.A0(net117),
    .A1(\u4.op1[3] ),
    .S(_0452_),
    .X(_0456_));
 sky130_fd_sc_hd__clkbuf_1 _0931_ (.A(_0456_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _0932_ (.A0(net120),
    .A1(\u4.op1[4] ),
    .S(_0452_),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_1 _0933_ (.A(_0457_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _0934_ (.A0(net100),
    .A1(\u4.op1[5] ),
    .S(_0452_),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_1 _0935_ (.A(_0458_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _0936_ (.A0(net125),
    .A1(\u4.op1[6] ),
    .S(_0452_),
    .X(_0459_));
 sky130_fd_sc_hd__clkbuf_1 _0937_ (.A(_0459_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _0938_ (.A0(net116),
    .A1(\u4.op1[7] ),
    .S(_0452_),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_1 _0939_ (.A(_0460_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _0940_ (.A0(net111),
    .A1(\u4.op1[8] ),
    .S(_0452_),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_1 _0941_ (.A(_0461_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _0942_ (.A0(\u1.state[6] ),
    .A1(\u1.state[14] ),
    .S(_0128_),
    .X(_0462_));
 sky130_fd_sc_hd__clkbuf_1 _0943_ (.A(_0462_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _0944_ (.A0(net126),
    .A1(\u1.state[12] ),
    .S(_0128_),
    .X(_0463_));
 sky130_fd_sc_hd__clkbuf_1 _0945_ (.A(_0463_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _0946_ (.A0(net133),
    .A1(\u1.state[10] ),
    .S(_0128_),
    .X(_0464_));
 sky130_fd_sc_hd__clkbuf_1 _0947_ (.A(_0464_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _0948_ (.A0(net118),
    .A1(\u1.state[9] ),
    .S(_0128_),
    .X(_0465_));
 sky130_fd_sc_hd__clkbuf_1 _0949_ (.A(net119),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _0950_ (.A0(\u1.state[10] ),
    .A1(net128),
    .S(_0128_),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_1 _0951_ (.A(net129),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _0952_ (.A0(net131),
    .A1(\u1.state[2] ),
    .S(_0128_),
    .X(_0467_));
 sky130_fd_sc_hd__clkbuf_1 _0953_ (.A(_0467_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _0954_ (.A0(net123),
    .A1(net118),
    .S(_0128_),
    .X(_0468_));
 sky130_fd_sc_hd__clkbuf_1 _0955_ (.A(_0468_),
    .X(_0112_));
 sky130_fd_sc_hd__dfstp_1 _0956_ (.CLK(clknet_4_10_0_clk),
    .D(net68),
    .SET_B(net32),
    .Q(\u7.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0957_ (.CLK(clknet_4_11_0_clk),
    .D(_0003_),
    .RESET_B(net32),
    .Q(\u7.assign_op2 ));
 sky130_fd_sc_hd__dfrtp_1 _0958_ (.CLK(clknet_4_11_0_clk),
    .D(_0004_),
    .RESET_B(net32),
    .Q(\u7.assign_op1 ));
 sky130_fd_sc_hd__dfrtp_4 _0959_ (.CLK(clknet_4_11_0_clk),
    .D(_0005_),
    .RESET_B(net32),
    .Q(\u4.result_ready ));
 sky130_fd_sc_hd__dfrtp_1 _0960_ (.CLK(clknet_4_9_0_clk),
    .D(_0012_),
    .RESET_B(net32),
    .Q(\u7.state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _0961_ (.CLK(clknet_4_8_0_clk),
    .D(_0013_),
    .RESET_B(net32),
    .Q(\u7.state[5] ));
 sky130_fd_sc_hd__dfrtp_1 _0962_ (.CLK(clknet_4_9_0_clk),
    .D(_0014_),
    .RESET_B(net33),
    .Q(\u7.state[6] ));
 sky130_fd_sc_hd__dfstp_1 _0963_ (.CLK(clknet_4_14_0_clk),
    .D(net70),
    .SET_B(net35),
    .Q(\u1.state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _0964_ (.CLK(clknet_4_14_0_clk),
    .D(_0000_),
    .RESET_B(net35),
    .Q(\u1.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _0965_ (.CLK(clknet_4_14_0_clk),
    .D(_0008_),
    .RESET_B(net35),
    .Q(\u1.state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _0966_ (.CLK(clknet_4_13_0_clk),
    .D(_0001_),
    .RESET_B(net35),
    .Q(\u1.store_dig ));
 sky130_fd_sc_hd__dfrtp_1 _0967_ (.CLK(clknet_4_14_0_clk),
    .D(net62),
    .RESET_B(net35),
    .Q(\u1.state[7] ));
 sky130_fd_sc_hd__dfrtp_1 _0968_ (.CLK(clknet_4_14_0_clk),
    .D(_0010_),
    .RESET_B(net35),
    .Q(\u1.state[8] ));
 sky130_fd_sc_hd__dfrtp_1 _0969_ (.CLK(clknet_4_14_0_clk),
    .D(_0002_),
    .RESET_B(net35),
    .Q(\u1.state[11] ));
 sky130_fd_sc_hd__dfrtp_1 _0970_ (.CLK(clknet_4_14_0_clk),
    .D(_0007_),
    .RESET_B(net35),
    .Q(\u1.state[13] ));
 sky130_fd_sc_hd__dfrtp_1 _0971_ (.CLK(clknet_4_7_0_clk),
    .D(net4),
    .RESET_B(net34),
    .Q(\u1.s_e_detect_w.i_signal ));
 sky130_fd_sc_hd__dfrtp_1 _0972_ (.CLK(clknet_4_13_0_clk),
    .D(net40),
    .RESET_B(net34),
    .Q(\u1.s_e_detect_w.s_signal ));
 sky130_fd_sc_hd__dfrtp_1 _0973_ (.CLK(clknet_4_12_0_clk),
    .D(net46),
    .RESET_B(net35),
    .Q(\u1.s_e_detect_w.p_signal ));
 sky130_fd_sc_hd__dfrtp_1 _0974_ (.CLK(clknet_4_5_0_clk),
    .D(net53),
    .RESET_B(net31),
    .Q(\u1.keypad_i[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0975_ (.CLK(clknet_4_5_0_clk),
    .D(net56),
    .RESET_B(net31),
    .Q(\u1.keypad_i[1] ));
 sky130_fd_sc_hd__dfrtp_2 _0976_ (.CLK(clknet_4_4_0_clk),
    .D(net43),
    .RESET_B(net31),
    .Q(\u1.keypad_sync[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0977_ (.CLK(clknet_4_5_0_clk),
    .D(net44),
    .RESET_B(net31),
    .Q(\u1.keypad_sync[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0978_ (.CLK(clknet_4_1_0_clk),
    .D(net2),
    .RESET_B(net29),
    .Q(\u1.keypad_async[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0979_ (.CLK(clknet_4_5_0_clk),
    .D(net3),
    .RESET_B(net31),
    .Q(\u1.keypad_async[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0980_ (.CLK(clknet_4_10_0_clk),
    .D(net52),
    .RESET_B(net32),
    .Q(\u3.keypad_13[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0981_ (.CLK(clknet_4_10_0_clk),
    .D(net51),
    .RESET_B(net32),
    .Q(\u3.keypad_13[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0982_ (.CLK(clknet_4_15_0_clk),
    .D(net39),
    .RESET_B(net35),
    .Q(\u3.keypad_sync[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0983_ (.CLK(clknet_4_10_0_clk),
    .D(net37),
    .RESET_B(net32),
    .Q(\u3.keypad_sync[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0984_ (.CLK(clknet_4_15_0_clk),
    .D(net6),
    .RESET_B(net35),
    .Q(\u3.keypad_async[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0985_ (.CLK(clknet_4_8_0_clk),
    .D(net7),
    .RESET_B(net32),
    .Q(\u3.keypad_async[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0986_ (.CLK(clknet_4_13_0_clk),
    .D(_0015_),
    .RESET_B(net34),
    .Q(\u4.op1[0] ));
 sky130_fd_sc_hd__dfrtp_2 _0987_ (.CLK(clknet_4_4_0_clk),
    .D(_0016_),
    .RESET_B(net30),
    .Q(\u4.op1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0988_ (.CLK(clknet_4_1_0_clk),
    .D(_0017_),
    .RESET_B(net31),
    .Q(\u4.op1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _0989_ (.CLK(clknet_4_6_0_clk),
    .D(_0018_),
    .RESET_B(net34),
    .Q(\u4.op1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _0990_ (.CLK(clknet_4_1_0_clk),
    .D(_0019_),
    .RESET_B(net30),
    .Q(\u4.op1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _0991_ (.CLK(clknet_4_4_0_clk),
    .D(_0020_),
    .RESET_B(net31),
    .Q(\u4.op1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _0992_ (.CLK(clknet_4_4_0_clk),
    .D(_0021_),
    .RESET_B(net31),
    .Q(\u4.op1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _0993_ (.CLK(clknet_4_5_0_clk),
    .D(_0022_),
    .RESET_B(net31),
    .Q(\u4.op1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _0994_ (.CLK(clknet_4_5_0_clk),
    .D(_0023_),
    .RESET_B(net31),
    .Q(\u4.op1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _0995_ (.CLK(clknet_4_0_0_clk),
    .D(_0024_),
    .RESET_B(net29),
    .Q(net13));
 sky130_fd_sc_hd__dfrtp_1 _0996_ (.CLK(clknet_4_0_0_clk),
    .D(_0025_),
    .RESET_B(net29),
    .Q(net12));
 sky130_fd_sc_hd__dfrtp_4 _0997_ (.CLK(clknet_4_5_0_clk),
    .D(_0026_),
    .RESET_B(net31),
    .Q(\u1.keycode[0] ));
 sky130_fd_sc_hd__dfrtp_4 _0998_ (.CLK(clknet_4_1_0_clk),
    .D(_0027_),
    .RESET_B(net29),
    .Q(\u1.keycode[1] ));
 sky130_fd_sc_hd__dfrtp_4 _0999_ (.CLK(clknet_4_1_0_clk),
    .D(_0028_),
    .RESET_B(net31),
    .Q(\u1.keycode[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1000_ (.CLK(clknet_4_1_0_clk),
    .D(_0029_),
    .RESET_B(net31),
    .Q(\u1.keycode[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1001_ (.CLK(clknet_4_1_0_clk),
    .D(_0030_),
    .RESET_B(net31),
    .Q(\u1.keycode[4] ));
 sky130_fd_sc_hd__dfrtp_4 _1002_ (.CLK(clknet_4_4_0_clk),
    .D(_0031_),
    .RESET_B(net31),
    .Q(\u1.keycode[5] ));
 sky130_fd_sc_hd__dfrtp_4 _1003_ (.CLK(clknet_4_4_0_clk),
    .D(_0032_),
    .RESET_B(net31),
    .Q(\u1.keycode[6] ));
 sky130_fd_sc_hd__dfrtp_4 _1004_ (.CLK(clknet_4_4_0_clk),
    .D(_0033_),
    .RESET_B(net31),
    .Q(\u1.keycode[7] ));
 sky130_fd_sc_hd__dfrtp_4 _1005_ (.CLK(clknet_4_4_0_clk),
    .D(_0034_),
    .RESET_B(net31),
    .Q(\u1.keycode[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1006_ (.CLK(clknet_4_11_0_clk),
    .D(net55),
    .RESET_B(net32),
    .Q(\u6.reg_i[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1007_ (.CLK(clknet_4_11_0_clk),
    .D(net58),
    .RESET_B(net32),
    .Q(\u6.reg_i[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1008_ (.CLK(clknet_4_11_0_clk),
    .D(net54),
    .RESET_B(net32),
    .Q(\u6.reg_i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1009_ (.CLK(clknet_4_11_0_clk),
    .D(net57),
    .RESET_B(net32),
    .Q(\u6.reg_i[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1010_ (.CLK(clknet_4_14_0_clk),
    .D(net41),
    .RESET_B(net35),
    .Q(\u6.reg_sync[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1011_ (.CLK(clknet_4_15_0_clk),
    .D(net38),
    .RESET_B(net35),
    .Q(\u6.reg_sync[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1012_ (.CLK(clknet_4_10_0_clk),
    .D(net45),
    .RESET_B(net32),
    .Q(\u6.reg_sync[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1013_ (.CLK(clknet_4_11_0_clk),
    .D(net49),
    .RESET_B(net36),
    .Q(\u6.reg_sync[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1014_ (.CLK(clknet_4_14_0_clk),
    .D(net8),
    .RESET_B(net35),
    .Q(\u6.reg_async[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1015_ (.CLK(clknet_4_13_0_clk),
    .D(net9),
    .RESET_B(net35),
    .Q(\u6.reg_async[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1016_ (.CLK(clknet_4_10_0_clk),
    .D(net10),
    .RESET_B(net32),
    .Q(\u6.reg_async[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1017_ (.CLK(clknet_4_1_0_clk),
    .D(net11),
    .RESET_B(net29),
    .Q(\u6.reg_async[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1018_ (.CLK(clknet_4_11_0_clk),
    .D(\u6.next_reg_num[0] ),
    .RESET_B(net33),
    .Q(\u5.reg_num[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1019_ (.CLK(clknet_4_11_0_clk),
    .D(\u6.next_reg_num[1] ),
    .RESET_B(net33),
    .Q(\u5.reg_num[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1020_ (.CLK(clknet_4_14_0_clk),
    .D(\u6.next_reg_num[2] ),
    .RESET_B(net33),
    .Q(\u5.reg_num[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1021_ (.CLK(clknet_4_12_0_clk),
    .D(_0035_),
    .RESET_B(net34),
    .Q(\u5.reg3[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1022_ (.CLK(clknet_4_12_0_clk),
    .D(_0036_),
    .RESET_B(net34),
    .Q(\u5.reg3[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1023_ (.CLK(clknet_4_6_0_clk),
    .D(_0037_),
    .RESET_B(net34),
    .Q(\u5.reg3[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1024_ (.CLK(clknet_4_7_0_clk),
    .D(_0038_),
    .RESET_B(net34),
    .Q(\u5.reg3[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1025_ (.CLK(clknet_4_3_0_clk),
    .D(_0039_),
    .RESET_B(net30),
    .Q(\u5.reg3[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1026_ (.CLK(clknet_4_4_0_clk),
    .D(_0040_),
    .RESET_B(net30),
    .Q(\u5.reg3[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1027_ (.CLK(clknet_4_4_0_clk),
    .D(_0041_),
    .RESET_B(net30),
    .Q(\u5.reg3[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1028_ (.CLK(clknet_4_5_0_clk),
    .D(_0042_),
    .RESET_B(net30),
    .Q(\u5.reg3[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1029_ (.CLK(clknet_4_7_0_clk),
    .D(_0043_),
    .RESET_B(net30),
    .Q(\u5.reg3[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1030_ (.CLK(clknet_4_13_0_clk),
    .D(_0044_),
    .RESET_B(net34),
    .Q(\u5.reg2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1031_ (.CLK(clknet_4_14_0_clk),
    .D(_0045_),
    .RESET_B(net34),
    .Q(\u5.reg2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1032_ (.CLK(clknet_4_6_0_clk),
    .D(_0046_),
    .RESET_B(net34),
    .Q(\u5.reg2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1033_ (.CLK(clknet_4_12_0_clk),
    .D(_0047_),
    .RESET_B(net34),
    .Q(\u5.reg2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1034_ (.CLK(clknet_4_6_0_clk),
    .D(_0048_),
    .RESET_B(net30),
    .Q(\u5.reg2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1035_ (.CLK(clknet_4_6_0_clk),
    .D(_0049_),
    .RESET_B(net30),
    .Q(\u5.reg2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1036_ (.CLK(clknet_4_7_0_clk),
    .D(_0050_),
    .RESET_B(net30),
    .Q(\u5.reg2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1037_ (.CLK(clknet_4_7_0_clk),
    .D(_0051_),
    .RESET_B(net30),
    .Q(\u5.reg2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1038_ (.CLK(clknet_4_7_0_clk),
    .D(_0052_),
    .RESET_B(net34),
    .Q(\u5.reg2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1039_ (.CLK(clknet_4_13_0_clk),
    .D(_0053_),
    .RESET_B(net34),
    .Q(\u5.reg1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1040_ (.CLK(clknet_4_12_0_clk),
    .D(_0054_),
    .RESET_B(net34),
    .Q(\u5.reg1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1041_ (.CLK(clknet_4_3_0_clk),
    .D(_0055_),
    .RESET_B(net34),
    .Q(\u5.reg1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1042_ (.CLK(clknet_4_12_0_clk),
    .D(_0056_),
    .RESET_B(net34),
    .Q(\u5.reg1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1043_ (.CLK(clknet_4_6_0_clk),
    .D(_0057_),
    .RESET_B(net30),
    .Q(\u5.reg1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1044_ (.CLK(clknet_4_6_0_clk),
    .D(_0058_),
    .RESET_B(net30),
    .Q(\u5.reg1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1045_ (.CLK(clknet_4_7_0_clk),
    .D(_0059_),
    .RESET_B(net30),
    .Q(\u5.reg1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1046_ (.CLK(clknet_4_5_0_clk),
    .D(_0060_),
    .RESET_B(net30),
    .Q(\u5.reg1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1047_ (.CLK(clknet_4_7_0_clk),
    .D(_0061_),
    .RESET_B(net36),
    .Q(\u5.reg1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1048_ (.CLK(clknet_4_9_0_clk),
    .D(_0062_),
    .RESET_B(net33),
    .Q(\u5.reg_val[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1049_ (.CLK(clknet_4_9_0_clk),
    .D(_0063_),
    .RESET_B(net33),
    .Q(\u5.reg_val[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1050_ (.CLK(clknet_4_9_0_clk),
    .D(_0064_),
    .RESET_B(net33),
    .Q(\u5.reg_val[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1051_ (.CLK(clknet_4_9_0_clk),
    .D(_0065_),
    .RESET_B(net33),
    .Q(\u5.reg_val[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1052_ (.CLK(clknet_4_3_0_clk),
    .D(_0066_),
    .RESET_B(net30),
    .Q(\u5.reg_val[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1053_ (.CLK(clknet_4_3_0_clk),
    .D(_0067_),
    .RESET_B(net30),
    .Q(\u5.reg_val[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1054_ (.CLK(clknet_4_3_0_clk),
    .D(_0068_),
    .RESET_B(net29),
    .Q(\u5.reg_val[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1055_ (.CLK(clknet_4_3_0_clk),
    .D(_0069_),
    .RESET_B(net29),
    .Q(\u5.reg_val[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1056_ (.CLK(clknet_4_3_0_clk),
    .D(_0070_),
    .RESET_B(net34),
    .Q(\u5.reg_val[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1057_ (.CLK(clknet_4_3_0_clk),
    .D(_0071_),
    .RESET_B(net29),
    .Q(\u4.ssdec[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1058_ (.CLK(clknet_4_1_0_clk),
    .D(_0072_),
    .RESET_B(net29),
    .Q(\u4.ssdec[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1059_ (.CLK(clknet_4_3_0_clk),
    .D(_0073_),
    .RESET_B(net29),
    .Q(\u4.ssdec[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1060_ (.CLK(clknet_4_3_0_clk),
    .D(_0074_),
    .RESET_B(net29),
    .Q(\u4.ssdec[3] ));
 sky130_fd_sc_hd__dfrtp_2 _1061_ (.CLK(clknet_4_0_0_clk),
    .D(_0075_),
    .RESET_B(net29),
    .Q(\u4.ssdec[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1062_ (.CLK(clknet_4_0_0_clk),
    .D(_0076_),
    .RESET_B(net29),
    .Q(\u4.ssdec[5] ));
 sky130_fd_sc_hd__dfrtp_4 _1063_ (.CLK(clknet_4_0_0_clk),
    .D(_0077_),
    .RESET_B(net29),
    .Q(\u4.ssdec[6] ));
 sky130_fd_sc_hd__dfrtp_4 _1064_ (.CLK(clknet_4_0_0_clk),
    .D(_0078_),
    .RESET_B(net29),
    .Q(\u4.ssdec[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1065_ (.CLK(clknet_4_10_0_clk),
    .D(net5),
    .RESET_B(net32),
    .Q(\u7.s_e_detect.i_signal ));
 sky130_fd_sc_hd__dfrtp_1 _1066_ (.CLK(clknet_4_10_0_clk),
    .D(net42),
    .RESET_B(net33),
    .Q(\u7.s_e_detect.s_signal ));
 sky130_fd_sc_hd__dfrtp_1 _1067_ (.CLK(clknet_4_10_0_clk),
    .D(net50),
    .RESET_B(net33),
    .Q(\u7.s_e_detect.p_signal ));
 sky130_fd_sc_hd__dfrtp_4 _1068_ (.CLK(clknet_4_10_0_clk),
    .D(\u3.out[1] ),
    .RESET_B(net32),
    .Q(\u8.buff_opcode[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1069_ (.CLK(clknet_4_9_0_clk),
    .D(_0079_),
    .RESET_B(net33),
    .Q(\u8.op2[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1070_ (.CLK(clknet_4_8_0_clk),
    .D(_0080_),
    .RESET_B(net32),
    .Q(\u8.op2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1071_ (.CLK(clknet_4_8_0_clk),
    .D(_0081_),
    .RESET_B(net33),
    .Q(\u8.op2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1072_ (.CLK(clknet_4_8_0_clk),
    .D(_0082_),
    .RESET_B(net33),
    .Q(\u8.op2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1073_ (.CLK(clknet_4_2_0_clk),
    .D(_0083_),
    .RESET_B(net29),
    .Q(\u8.op2[4] ));
 sky130_fd_sc_hd__dfrtp_2 _1074_ (.CLK(clknet_4_2_0_clk),
    .D(_0084_),
    .RESET_B(net29),
    .Q(\u8.op2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1075_ (.CLK(clknet_4_2_0_clk),
    .D(_0085_),
    .RESET_B(net29),
    .Q(\u8.op2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1076_ (.CLK(clknet_4_2_0_clk),
    .D(_0086_),
    .RESET_B(net29),
    .Q(\u8.op2[7] ));
 sky130_fd_sc_hd__dfrtp_2 _1077_ (.CLK(clknet_4_9_0_clk),
    .D(_0087_),
    .RESET_B(net33),
    .Q(\u8.op2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1078_ (.CLK(clknet_4_8_0_clk),
    .D(_0088_),
    .RESET_B(net33),
    .Q(\u8.new_op1[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1079_ (.CLK(clknet_4_8_0_clk),
    .D(_0089_),
    .RESET_B(net33),
    .Q(\u8.new_op1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1080_ (.CLK(clknet_4_8_0_clk),
    .D(_0090_),
    .RESET_B(net33),
    .Q(\u8.new_op1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1081_ (.CLK(clknet_4_8_0_clk),
    .D(_0091_),
    .RESET_B(net33),
    .Q(\u8.new_op1[3] ));
 sky130_fd_sc_hd__dfrtp_2 _1082_ (.CLK(clknet_4_2_0_clk),
    .D(_0092_),
    .RESET_B(net36),
    .Q(\u8.op1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1083_ (.CLK(clknet_4_2_0_clk),
    .D(_0093_),
    .RESET_B(net36),
    .Q(\u8.op1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1084_ (.CLK(clknet_4_0_0_clk),
    .D(_0094_),
    .RESET_B(net29),
    .Q(\u8.op1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1085_ (.CLK(clknet_4_2_0_clk),
    .D(_0095_),
    .RESET_B(net36),
    .Q(\u8.op1[7] ));
 sky130_fd_sc_hd__dfrtp_4 _1086_ (.CLK(clknet_4_2_0_clk),
    .D(_0096_),
    .RESET_B(net36),
    .Q(\u8.new_op1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1087_ (.CLK(clknet_4_7_0_clk),
    .D(_0097_),
    .RESET_B(net36),
    .Q(\u5.reg4[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1088_ (.CLK(clknet_4_6_0_clk),
    .D(_0098_),
    .RESET_B(net34),
    .Q(\u5.reg4[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1089_ (.CLK(clknet_4_6_0_clk),
    .D(_0099_),
    .RESET_B(net34),
    .Q(\u5.reg4[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1090_ (.CLK(clknet_4_6_0_clk),
    .D(_0100_),
    .RESET_B(net36),
    .Q(\u5.reg4[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1091_ (.CLK(clknet_4_3_0_clk),
    .D(_0101_),
    .RESET_B(net30),
    .Q(\u5.reg4[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1092_ (.CLK(clknet_4_4_0_clk),
    .D(_0102_),
    .RESET_B(net30),
    .Q(\u5.reg4[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1093_ (.CLK(clknet_4_5_0_clk),
    .D(_0103_),
    .RESET_B(net30),
    .Q(\u5.reg4[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1094_ (.CLK(clknet_4_5_0_clk),
    .D(_0104_),
    .RESET_B(net36),
    .Q(\u5.reg4[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1095_ (.CLK(clknet_4_7_0_clk),
    .D(_0105_),
    .RESET_B(net31),
    .Q(\u5.reg4[8] ));
 sky130_fd_sc_hd__dfrtp_4 _1096_ (.CLK(clknet_4_8_0_clk),
    .D(net48),
    .RESET_B(net33),
    .Q(\u8.b_assign_op1 ));
 sky130_fd_sc_hd__dfrtp_4 _1097_ (.CLK(clknet_4_10_0_clk),
    .D(net47),
    .RESET_B(net32),
    .Q(\u8.b_assign_op2 ));
 sky130_fd_sc_hd__dfrtp_1 _1098_ (.CLK(clknet_4_15_0_clk),
    .D(_0106_),
    .RESET_B(net35),
    .Q(\u1.state[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1099_ (.CLK(clknet_4_15_0_clk),
    .D(_0107_),
    .RESET_B(net35),
    .Q(\u1.state[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1100_ (.CLK(clknet_4_15_0_clk),
    .D(_0108_),
    .RESET_B(net35),
    .Q(\u1.state[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1101_ (.CLK(clknet_4_13_0_clk),
    .D(_0109_),
    .RESET_B(net35),
    .Q(\u1.state[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1102_ (.CLK(clknet_4_15_0_clk),
    .D(_0110_),
    .RESET_B(net35),
    .Q(\u1.state[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1103_ (.CLK(clknet_4_15_0_clk),
    .D(_0111_),
    .RESET_B(net36),
    .Q(\u1.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1104_ (.CLK(clknet_4_13_0_clk),
    .D(_0112_),
    .RESET_B(net36),
    .Q(\u1.state[1] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__buf_6 fanout29 (.A(net36),
    .X(net29));
 sky130_fd_sc_hd__buf_6 fanout30 (.A(net31),
    .X(net30));
 sky130_fd_sc_hd__buf_6 fanout31 (.A(net36),
    .X(net31));
 sky130_fd_sc_hd__buf_6 fanout32 (.A(net33),
    .X(net32));
 sky130_fd_sc_hd__buf_6 fanout33 (.A(net36),
    .X(net33));
 sky130_fd_sc_hd__buf_6 fanout34 (.A(net36),
    .X(net34));
 sky130_fd_sc_hd__buf_6 fanout35 (.A(net36),
    .X(net35));
 sky130_fd_sc_hd__buf_8 fanout36 (.A(net1),
    .X(net36));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\u3.keypad_async[1] ),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\u1.s_e_detect_w.s_signal ),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\u5.reg_val[1] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\u7.assign_op2 ),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\u7.assign_op1 ),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\u6.reg_async[3] ),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\u7.s_e_detect.s_signal ),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\u3.keypad_sync[1] ),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\u3.keypad_sync[0] ),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\u1.keypad_sync[0] ),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\u6.reg_sync[2] ),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\u6.reg_sync[0] ),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\u6.reg_async[1] ),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\u1.keypad_sync[1] ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\u6.reg_sync[3] ),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\u6.reg_sync[1] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\u7.state[5] ),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\u7.state[6] ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\u1.state[11] ),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0009_),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net12),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\u7.state[4] ),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\u1.state[9] ),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\u3.keypad_async[0] ),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\u1.state[8] ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\u7.state[0] ),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0011_),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\u1.state[0] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0006_),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\u1.state[13] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net13),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\u4.op1[0] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\u4.op1[6] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\u3.keypad_13[0] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\u1.s_e_detect_w.i_signal ),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0129_),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\u4.op1[5] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\u5.reg4[1] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\u5.reg1[7] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\u5.reg2[1] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\u4.op1[2] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\u5.reg2[4] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\u5.reg1[0] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\u4.op1[4] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\u5.reg2[6] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\u6.reg_async[0] ),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\u5.reg1[3] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\u4.op1[7] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\u5.reg2[7] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\u5.reg3[0] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\u5.reg4[0] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\u4.op1[3] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\u5.reg1[6] ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\u5.reg3[8] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\u5.reg3[3] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\u5.reg_val[0] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\u7.s_e_detect.i_signal ),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\u4.op1[1] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\u5.reg2[2] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\u5.reg1[4] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\u5.reg3[6] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\u5.reg4[5] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\u5.reg2[8] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\u5.reg1[2] ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\u5.reg2[5] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\u5.reg2[3] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\u5.reg3[5] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\u1.keypad_async[0] ),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\u5.reg1[8] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\u5.reg3[1] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\u5.reg4[2] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\u5.reg1[1] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\u5.reg3[7] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\u5.reg4[8] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\u5.reg3[2] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\u5.reg1[5] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\u4.ssdec[6] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\u5.reg3[4] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\u1.keypad_async[1] ),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\u5.reg4[7] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\u5.reg4[3] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\u1.state[1] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_0465_),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\u5.reg4[4] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\u4.ssdec[2] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\u5.reg2[0] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\u1.state[14] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\u4.ssdec[5] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\u5.reg4[6] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\u6.reg_async[2] ),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\u1.state[4] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\u5.reg_val[3] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\u1.state[6] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_0466_),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\u5.reg_val[1] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\u1.state[12] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\u4.op1[8] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\u1.state[2] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\u5.reg_val[3] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\u5.reg_val[1] ),
    .X(net135));
 sky130_fd_sc_hd__buf_1 input1 (.A(nrst),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(pb[8]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(pb[9]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(pb[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(pb[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(pb[2]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(pb[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(pb[4]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(pb[5]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(pb[6]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(pb[7]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 max_cap28 (.A(_0337_),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 output12 (.A(net12),
    .X(blue));
 sky130_fd_sc_hd__clkbuf_4 output13 (.A(net13),
    .X(red));
 sky130_fd_sc_hd__clkbuf_4 output14 (.A(net14),
    .X(ss[0]));
 sky130_fd_sc_hd__clkbuf_4 output15 (.A(net15),
    .X(ss[10]));
 sky130_fd_sc_hd__clkbuf_4 output16 (.A(net16),
    .X(ss[11]));
 sky130_fd_sc_hd__clkbuf_4 output17 (.A(net17),
    .X(ss[12]));
 sky130_fd_sc_hd__clkbuf_4 output18 (.A(net18),
    .X(ss[13]));
 sky130_fd_sc_hd__clkbuf_4 output19 (.A(net19),
    .X(ss[1]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(ss[2]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(ss[3]));
 sky130_fd_sc_hd__clkbuf_4 output22 (.A(net22),
    .X(ss[4]));
 sky130_fd_sc_hd__clkbuf_4 output23 (.A(net23),
    .X(ss[5]));
 sky130_fd_sc_hd__clkbuf_4 output24 (.A(net24),
    .X(ss[6]));
 sky130_fd_sc_hd__clkbuf_4 output25 (.A(net25),
    .X(ss[7]));
 sky130_fd_sc_hd__clkbuf_4 output26 (.A(net26),
    .X(ss[8]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(ss[9]));
endmodule

