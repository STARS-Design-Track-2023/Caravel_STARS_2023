magic
tech sky130A
magscale 1 2
timestamp 1694454429
<< obsli1 >>
rect 1104 2159 44620 45713
<< obsm1 >>
rect 14 2128 44698 45744
<< metal2 >>
rect 6458 47077 6514 47877
rect 14830 47077 14886 47877
rect 23846 47077 23902 47877
rect 32218 47077 32274 47877
rect 41234 47077 41290 47877
rect 18 0 74 800
rect 8390 0 8446 800
rect 17406 0 17462 800
rect 25778 0 25834 800
rect 34794 0 34850 800
rect 43166 0 43222 800
<< obsm2 >>
rect 20 47021 6402 47077
rect 6570 47021 14774 47077
rect 14942 47021 23790 47077
rect 23958 47021 32162 47077
rect 32330 47021 41178 47077
rect 41346 47021 44694 47077
rect 20 856 44694 47021
rect 130 734 8334 856
rect 8502 734 17350 856
rect 17518 734 25722 856
rect 25890 734 34738 856
rect 34906 734 43110 856
rect 43278 734 44694 856
<< metal3 >>
rect 0 45568 800 45688
rect 44933 43528 45733 43648
rect 0 36728 800 36848
rect 44933 34008 45733 34128
rect 0 27208 800 27328
rect 44933 25168 45733 25288
rect 0 18368 800 18488
rect 44933 15648 45733 15768
rect 0 8848 800 8968
rect 44933 6808 45733 6928
<< obsm3 >>
rect 880 45488 44933 45729
rect 800 43728 44933 45488
rect 800 43448 44853 43728
rect 800 36928 44933 43448
rect 880 36648 44933 36928
rect 800 34208 44933 36648
rect 800 33928 44853 34208
rect 800 27408 44933 33928
rect 880 27128 44933 27408
rect 800 25368 44933 27128
rect 800 25088 44853 25368
rect 800 18568 44933 25088
rect 880 18288 44933 18568
rect 800 15848 44933 18288
rect 800 15568 44853 15848
rect 800 9048 44933 15568
rect 880 8768 44933 9048
rect 800 7008 44933 8768
rect 800 6728 44853 7008
rect 800 2143 44933 6728
<< metal4 >>
rect 4208 2128 4528 45744
rect 19568 2128 19888 45744
rect 34928 2128 35248 45744
<< obsm4 >>
rect 10547 5339 19488 30837
rect 19968 5339 31221 30837
<< labels >>
rlabel metal2 s 34794 0 34850 800 6 clk
port 1 nsew signal input
rlabel metal3 s 44933 43528 45733 43648 6 cs
port 2 nsew signal input
rlabel metal2 s 41234 47077 41290 47877 6 gpio[0]
port 3 nsew signal input
rlabel metal2 s 23846 47077 23902 47877 6 gpio[10]
port 4 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 gpio[11]
port 5 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 gpio[12]
port 6 nsew signal input
rlabel metal3 s 44933 6808 45733 6928 6 gpio[13]
port 7 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 gpio[14]
port 8 nsew signal input
rlabel metal3 s 44933 34008 45733 34128 6 gpio[15]
port 9 nsew signal input
rlabel metal2 s 18 0 74 800 6 gpio[16]
port 10 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 gpio[1]
port 11 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 gpio[2]
port 12 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 gpio[3]
port 13 nsew signal input
rlabel metal2 s 14830 47077 14886 47877 6 gpio[4]
port 14 nsew signal input
rlabel metal3 s 44933 25168 45733 25288 6 gpio[5]
port 15 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 gpio[6]
port 16 nsew signal input
rlabel metal2 s 32218 47077 32274 47877 6 gpio[7]
port 17 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 gpio[8]
port 18 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 gpio[9]
port 19 nsew signal input
rlabel metal2 s 6458 47077 6514 47877 6 nrst
port 20 nsew signal input
rlabel metal3 s 44933 15648 45733 15768 6 pwm
port 21 nsew signal output
rlabel metal4 s 4208 2128 4528 45744 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 45744 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 45744 6 vssd1
port 23 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 45733 47877
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5157914
string GDS_FILE /home/designer-05/Caravel_STARS_2023/openlane/silly-sythensizer/runs/23_09_11_10_43/results/signoff/silly_synthesizer.magic.gds
string GDS_START 763434
<< end >>

